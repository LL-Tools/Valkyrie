

module b20_C_SARLock_k_64_7 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10184;

  NAND2_X1 U4814 ( .A1(n7264), .A2(n9009), .ZN(n7507) );
  NAND2_X2 U4815 ( .A1(n5221), .A2(n5220), .ZN(n7632) );
  INV_X1 U4816 ( .A(n5824), .ZN(n7732) );
  NAND4_X2 U4818 ( .A1(n5035), .A2(n5034), .A3(n5033), .A4(n5032), .ZN(n9252)
         );
  INV_X1 U4819 ( .A(n4980), .ZN(n5692) );
  CLKBUF_X1 U4820 ( .A(n9216), .Z(n4315) );
  NAND2_X2 U4821 ( .A1(n7695), .A2(n4940), .ZN(n5059) );
  OR3_X1 U4822 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5771) );
  CLKBUF_X1 U4823 ( .A(n10184), .Z(P2_U3893) );
  NOR2_X1 U4824 ( .A1(n6452), .A2(P2_U3151), .ZN(n10184) );
  INV_X1 U4825 ( .A(n9564), .ZN(n4308) );
  INV_X2 U4826 ( .A(n4308), .ZN(n4309) );
  AND4_X1 U4827 ( .A1(n5760), .A2(n5948), .A3(n5788), .A4(n5794), .ZN(n5745)
         );
  INV_X1 U4828 ( .A(n8789), .ZN(n5805) );
  AOI21_X1 U4829 ( .B1(n10008), .B2(n10006), .A(n10007), .ZN(n10005) );
  CLKBUF_X2 U4830 ( .A(n5050), .Z(n5615) );
  INV_X1 U4831 ( .A(n4985), .ZN(n5628) );
  OR2_X1 U4832 ( .A1(n9252), .A2(n4523), .ZN(n8982) );
  NAND2_X1 U4833 ( .A1(n7521), .A2(n7523), .ZN(n7522) );
  INV_X2 U4834 ( .A(n6086), .ZN(n8018) );
  AND2_X1 U4835 ( .A1(n4669), .A2(n4668), .ZN(n8075) );
  AND2_X1 U4836 ( .A1(n4877), .A2(n4874), .ZN(n7712) );
  INV_X2 U4838 ( .A(n4313), .ZN(n5701) );
  NAND2_X1 U4839 ( .A1(n4346), .A2(n4438), .ZN(n9851) );
  OR2_X1 U4840 ( .A1(n4936), .A2(n9756), .ZN(n4481) );
  INV_X1 U4841 ( .A(n5839), .ZN(n6309) );
  XNOR2_X1 U4842 ( .A(n6360), .B(n7671), .ZN(n7659) );
  NAND2_X1 U4843 ( .A1(n6373), .A2(n5845), .ZN(n5860) );
  AND2_X1 U4844 ( .A1(n7709), .A2(n9347), .ZN(n9125) );
  CLKBUF_X3 U4845 ( .A(n5059), .Z(n5651) );
  XNOR2_X1 U4846 ( .A(n5555), .B(n5554), .ZN(n7637) );
  XNOR2_X1 U4847 ( .A(n5415), .B(n5414), .ZN(n7196) );
  NAND4_X2 U4849 ( .A1(n5063), .A2(n5062), .A3(n5061), .A4(n5060), .ZN(n9251)
         );
  OR2_X1 U4850 ( .A1(n4357), .A2(n9360), .ZN(n9622) );
  AND2_X1 U4851 ( .A1(n4583), .A2(n6488), .ZN(n4310) );
  AND2_X1 U4852 ( .A1(n4483), .A2(n4409), .ZN(n4311) );
  NOR2_X4 U4853 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5217) );
  INV_X2 U4854 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4949) );
  OR2_X2 U4855 ( .A1(n9321), .A2(n9857), .ZN(n4346) );
  NAND2_X4 U4856 ( .A1(n4713), .A2(n5860), .ZN(n6602) );
  NAND2_X1 U4857 ( .A1(n6613), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5035) );
  AND2_X1 U4858 ( .A1(n9212), .A2(n5716), .ZN(n9564) );
  OAI21_X2 U4859 ( .B1(n7458), .B2(n7457), .A(n7798), .ZN(n7475) );
  NAND2_X2 U4860 ( .A1(n7352), .A2(n7779), .ZN(n7458) );
  NAND2_X2 U4861 ( .A1(n5385), .A2(n5384), .ZN(n5415) );
  CLKBUF_X1 U4862 ( .A(n5011), .Z(n4312) );
  CLKBUF_X1 U4863 ( .A(n5011), .Z(n4313) );
  INV_X2 U4864 ( .A(n7675), .ZN(n9109) );
  XNOR2_X2 U4865 ( .A(n7712), .B(n7958), .ZN(n8450) );
  INV_X4 U4866 ( .A(n7978), .ZN(n6892) );
  XNOR2_X2 U4867 ( .A(n9255), .B(n4617), .ZN(n9093) );
  NAND2_X2 U4868 ( .A1(n4342), .A2(n4942), .ZN(n9255) );
  BUF_X4 U4869 ( .A(n5161), .Z(n6613) );
  NAND2_X2 U4870 ( .A1(n5190), .A2(n5189), .ZN(n9610) );
  AOI21_X2 U4871 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n6788), .A(n7592), .ZN(
        n6360) );
  XNOR2_X1 U4872 ( .A(n5795), .B(n5794), .ZN(n6072) );
  INV_X2 U4873 ( .A(n7705), .ZN(n4940) );
  XNOR2_X2 U4874 ( .A(n5072), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9278) );
  XNOR2_X2 U4875 ( .A(n6381), .B(n6422), .ZN(n7069) );
  OAI21_X2 U4876 ( .B1(n6955), .B2(n6416), .A(n6946), .ZN(n6381) );
  NAND2_X1 U4878 ( .A1(n9426), .A2(n9139), .ZN(n9409) );
  AND2_X1 U4879 ( .A1(n9622), .A2(n9621), .ZN(n9708) );
  NAND2_X1 U4880 ( .A1(n9522), .A2(n9523), .ZN(n9521) );
  OR2_X1 U4881 ( .A1(n9481), .A2(n9462), .ZN(n9460) );
  OAI211_X1 U4882 ( .C1(n4849), .C2(n4844), .A(n4842), .B(n4847), .ZN(n7107)
         );
  NAND2_X1 U4883 ( .A1(n9155), .A2(n8990), .ZN(n6909) );
  INV_X4 U4884 ( .A(n5628), .ZN(n5710) );
  INV_X2 U4885 ( .A(n5657), .ZN(n5036) );
  INV_X2 U4886 ( .A(n7101), .ZN(n9940) );
  NAND2_X1 U4887 ( .A1(n4319), .A2(n4317), .ZN(n5879) );
  NAND2_X2 U4888 ( .A1(n5716), .A2(n9763), .ZN(n6608) );
  OAI21_X1 U4889 ( .B1(n4317), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n5016), .ZN(
        n5043) );
  MUX2_X1 U4890 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n6334), .S(n10124), .Z(n6324) );
  MUX2_X1 U4891 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n6334), .S(n10110), .Z(n6335) );
  NAND2_X1 U4892 ( .A1(n8011), .A2(n8308), .ZN(n8311) );
  AND2_X1 U4893 ( .A1(n4630), .A2(n4624), .ZN(n9089) );
  AOI21_X1 U4894 ( .B1(n4629), .B2(n4625), .A(n9189), .ZN(n4624) );
  AOI21_X1 U4895 ( .B1(n9380), .B2(n9592), .A(n9379), .ZN(n9626) );
  OR2_X1 U4896 ( .A1(n8470), .A2(n6304), .ZN(n4879) );
  NAND2_X1 U4897 ( .A1(n9400), .A2(n9399), .ZN(n4773) );
  AOI21_X1 U4898 ( .B1(n7893), .B2(n7892), .A(n7891), .ZN(n7902) );
  NOR2_X1 U4899 ( .A1(n8436), .A2(n4418), .ZN(n4417) );
  XNOR2_X1 U4900 ( .A(n8458), .B(n8335), .ZN(n8019) );
  OR2_X1 U4901 ( .A1(n8408), .A2(n8592), .ZN(n4741) );
  AOI21_X1 U4902 ( .B1(n4891), .B2(n4889), .A(n4888), .ZN(n4887) );
  OAI22_X1 U4903 ( .A1(n9569), .A2(n6521), .B1(n9545), .B2(n9748), .ZN(n9538)
         );
  INV_X1 U4904 ( .A(n4891), .ZN(n4890) );
  OAI21_X1 U4905 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n9870), .A(n9867), .ZN(
        n9879) );
  NAND2_X1 U4906 ( .A1(n5512), .A2(n5511), .ZN(n9484) );
  OR2_X1 U4907 ( .A1(n7666), .A2(n7665), .ZN(n4738) );
  CLKBUF_X1 U4908 ( .A(n7414), .Z(n4441) );
  NAND2_X1 U4909 ( .A1(n6102), .A2(n6101), .ZN(n8738) );
  NOR2_X1 U4910 ( .A1(n7677), .A2(n9687), .ZN(n9570) );
  NAND2_X1 U4911 ( .A1(n7078), .A2(n4685), .ZN(n7152) );
  NAND2_X1 U4912 ( .A1(n5395), .A2(n5394), .ZN(n9574) );
  NAND2_X2 U4913 ( .A1(n5367), .A2(n5366), .ZN(n9687) );
  XNOR2_X1 U4914 ( .A(n5382), .B(n5381), .ZN(n7176) );
  AND2_X1 U4915 ( .A1(n4635), .A2(n4634), .ZN(n7548) );
  NAND2_X1 U4916 ( .A1(n6007), .A2(n6006), .ZN(n8682) );
  OR2_X1 U4917 ( .A1(n7307), .A2(n6356), .ZN(n4635) );
  NAND2_X1 U4918 ( .A1(n5309), .A2(n5308), .ZN(n5334) );
  OAI21_X1 U4919 ( .B1(n5234), .B2(n5211), .A(n5210), .ZN(n5259) );
  OAI21_X1 U4920 ( .B1(n5234), .B2(n4836), .A(n4833), .ZN(n5306) );
  OAI211_X1 U4921 ( .C1(n5830), .C2(n7311), .A(n5951), .B(n5950), .ZN(n7453)
         );
  NAND2_X1 U4922 ( .A1(n5206), .A2(n5205), .ZN(n5234) );
  AND2_X1 U4923 ( .A1(n4746), .A2(n4742), .ZN(n6383) );
  XNOR2_X1 U4924 ( .A(n5204), .B(n4915), .ZN(n6694) );
  NAND2_X1 U4925 ( .A1(n5178), .A2(n5177), .ZN(n5204) );
  OR2_X1 U4926 ( .A1(n5176), .A2(n5175), .ZN(n5178) );
  NAND2_X1 U4927 ( .A1(n5152), .A2(n5151), .ZN(n5176) );
  NOR2_X1 U4928 ( .A1(n6924), .A2(n7408), .ZN(n6944) );
  AND2_X1 U4929 ( .A1(n4354), .A2(n6947), .ZN(n6922) );
  NAND2_X1 U4930 ( .A1(n5793), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5795) );
  OR2_X1 U4931 ( .A1(n8349), .A2(n6975), .ZN(n7753) );
  INV_X1 U4932 ( .A(n9924), .ZN(n4523) );
  AND3_X1 U4933 ( .A1(n5848), .A2(n5847), .A3(n5846), .ZN(n10055) );
  AND4_X1 U4934 ( .A1(n5858), .A2(n5857), .A3(n5856), .A4(n5855), .ZN(n6268)
         );
  NAND4_X1 U4935 ( .A1(n5818), .A2(n5817), .A3(n5816), .A4(n5815), .ZN(n8349)
         );
  NAND2_X1 U4936 ( .A1(n6843), .A2(n4423), .ZN(n5657) );
  NAND4_X1 U4937 ( .A1(n5015), .A2(n5014), .A3(n5013), .A4(n5012), .ZN(n9253)
         );
  NAND2_X2 U4938 ( .A1(n6572), .A2(n9126), .ZN(n9548) );
  NAND2_X1 U4939 ( .A1(n5046), .A2(n5045), .ZN(n5065) );
  AND2_X1 U4940 ( .A1(n6347), .A2(n6826), .ZN(n6863) );
  XNOR2_X1 U4941 ( .A(n4953), .B(n4952), .ZN(n4980) );
  NAND2_X1 U4942 ( .A1(n6180), .A2(n6181), .ZN(n5830) );
  OR2_X1 U4943 ( .A1(n6346), .A2(n6861), .ZN(n6347) );
  XNOR2_X1 U4944 ( .A(n5803), .B(n5802), .ZN(n8789) );
  NOR2_X1 U4945 ( .A1(n5787), .A2(n5786), .ZN(n6031) );
  NAND2_X1 U4946 ( .A1(n4951), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4953) );
  NAND2_X1 U4947 ( .A1(n5756), .A2(n5755), .ZN(n6181) );
  NAND2_X1 U4948 ( .A1(n4951), .A2(n4948), .ZN(n9126) );
  XNOR2_X1 U4949 ( .A(n4950), .B(n4949), .ZN(n9216) );
  NAND2_X1 U4950 ( .A1(n9757), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4935) );
  MUX2_X1 U4951 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5754), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5756) );
  NAND2_X1 U4952 ( .A1(n4445), .A2(n4442), .ZN(n9763) );
  XNOR2_X1 U4953 ( .A(n4962), .B(n4873), .ZN(n9770) );
  NAND2_X2 U4954 ( .A1(n4518), .A2(P1_U3086), .ZN(n9769) );
  OR2_X1 U4955 ( .A1(n4970), .A2(n4933), .ZN(n4445) );
  NAND2_X1 U4956 ( .A1(n4971), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4968) );
  INV_X1 U4957 ( .A(n5757), .ZN(n5747) );
  XNOR2_X1 U4958 ( .A(n5878), .B(n5877), .ZN(n6841) );
  NAND4_X1 U4959 ( .A1(n6373), .A2(n4901), .A3(n5741), .A4(n4550), .ZN(n5757)
         );
  INV_X4 U4960 ( .A(n7727), .ZN(n4317) );
  NAND2_X1 U4961 ( .A1(n4715), .A2(n4714), .ZN(n4713) );
  AND2_X1 U4962 ( .A1(n5877), .A2(n5901), .ZN(n4901) );
  AND2_X1 U4963 ( .A1(n5887), .A2(n5742), .ZN(n4550) );
  INV_X1 U4964 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5758) );
  INV_X1 U4965 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5794) );
  INV_X1 U4966 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5948) );
  INV_X1 U4967 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5788) );
  INV_X1 U4968 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5759) );
  INV_X1 U4969 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5992) );
  INV_X1 U4970 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5669) );
  INV_X4 U4971 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U4972 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n4919) );
  NOR2_X1 U4973 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4920) );
  INV_X1 U4974 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n4944) );
  OR2_X1 U4975 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n4899) );
  INV_X1 U4976 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4946) );
  INV_X1 U4977 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4952) );
  INV_X1 U4978 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4955) );
  NOR2_X1 U4979 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5744) );
  NOR2_X1 U4980 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5070) );
  NOR2_X1 U4981 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5022) );
  INV_X4 U4982 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  AND2_X2 U4983 ( .A1(n4794), .A2(n4793), .ZN(n7727) );
  NAND2_X1 U4984 ( .A1(n7705), .A2(n4939), .ZN(n5011) );
  AND2_X4 U4985 ( .A1(n5810), .A2(n5805), .ZN(n6087) );
  INV_X1 U4987 ( .A(n7718), .ZN(n4318) );
  AOI21_X2 U4988 ( .B1(n6571), .B2(n9592), .A(n6570), .ZN(n9376) );
  NAND2_X1 U4989 ( .A1(n6180), .A2(n6181), .ZN(n4319) );
  NAND2_X4 U4990 ( .A1(n4939), .A2(n4940), .ZN(n5010) );
  AND2_X1 U4991 ( .A1(n6608), .A2(n4701), .ZN(n4320) );
  AND2_X4 U4992 ( .A1(n6608), .A2(n4701), .ZN(n5037) );
  AOI21_X1 U4993 ( .B1(n4575), .B2(n4576), .A(n6294), .ZN(n4573) );
  NAND2_X1 U4994 ( .A1(n5657), .A2(n4985), .ZN(n5050) );
  NAND2_X1 U4995 ( .A1(n5608), .A2(n5607), .ZN(n5636) );
  NOR2_X2 U4996 ( .A1(n4926), .A2(n4925), .ZN(n4929) );
  OAI21_X1 U4997 ( .B1(n5772), .B2(n5753), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5754) );
  INV_X1 U4998 ( .A(n5749), .ZN(n5753) );
  NAND2_X1 U4999 ( .A1(n5755), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5752) );
  CLKBUF_X1 U5000 ( .A(n5777), .Z(n5778) );
  OR2_X1 U5001 ( .A1(n6947), .A2(n6948), .ZN(n4641) );
  XNOR2_X1 U5002 ( .A(n5800), .B(n5799), .ZN(n5804) );
  NAND2_X1 U5003 ( .A1(n4581), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5800) );
  AOI21_X1 U5004 ( .B1(n9414), .B2(n6531), .A(n4771), .ZN(n9400) );
  NAND2_X1 U5005 ( .A1(n9445), .A2(n9064), .ZN(n4597) );
  OR2_X1 U5006 ( .A1(n8566), .A2(n8300), .ZN(n7746) );
  INV_X1 U5007 ( .A(n5502), .ZN(n5503) );
  NAND2_X1 U5008 ( .A1(n7717), .A2(n7716), .ZN(n7736) );
  NAND2_X1 U5009 ( .A1(n4877), .A2(n4365), .ZN(n7717) );
  NAND2_X1 U5010 ( .A1(n5810), .A2(n8789), .ZN(n5854) );
  NOR2_X1 U5011 ( .A1(n6948), .A2(n4643), .ZN(n4642) );
  OR2_X1 U5012 ( .A1(n6491), .A2(n8024), .ZN(n7903) );
  OR2_X1 U5013 ( .A1(n8751), .A2(n8590), .ZN(n7948) );
  NAND2_X1 U5014 ( .A1(n8340), .A2(n10095), .ZN(n7779) );
  AND2_X1 U5015 ( .A1(n6158), .A2(n5774), .ZN(n4670) );
  INV_X1 U5016 ( .A(n4557), .ZN(n4556) );
  AND2_X1 U5017 ( .A1(n6226), .A2(n8336), .ZN(n7925) );
  INV_X1 U5018 ( .A(n5838), .ZN(n6106) );
  OR2_X1 U5019 ( .A1(n8533), .A2(n8062), .ZN(n7741) );
  OR2_X1 U5020 ( .A1(n8744), .A2(n8063), .ZN(n7863) );
  OR2_X1 U5021 ( .A1(n8674), .A2(n8101), .ZN(n7947) );
  INV_X1 U5022 ( .A(n8632), .ZN(n4544) );
  NAND2_X1 U5023 ( .A1(n7339), .A2(n7773), .ZN(n4897) );
  OR2_X1 U5024 ( .A1(n6142), .A2(n6319), .ZN(n6965) );
  NOR2_X1 U5025 ( .A1(n4899), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n4688) );
  AOI21_X1 U5026 ( .B1(n7107), .B2(n4506), .A(n4503), .ZN(n5172) );
  NOR2_X1 U5027 ( .A1(n4323), .A2(n5123), .ZN(n4506) );
  OAI21_X1 U5028 ( .B1(n4504), .B2(n4323), .A(n4350), .ZN(n4503) );
  INV_X1 U5029 ( .A(n8883), .ZN(n4502) );
  AOI21_X1 U5030 ( .B1(n4612), .B2(n4610), .A(n4376), .ZN(n9079) );
  AOI21_X1 U5031 ( .B1(n9141), .B2(n4628), .A(n4611), .ZN(n4610) );
  INV_X1 U5032 ( .A(n4772), .ZN(n4770) );
  INV_X1 U5033 ( .A(n4477), .ZN(n4476) );
  NAND2_X1 U5034 ( .A1(n9521), .A2(n4709), .ZN(n4708) );
  NOR2_X1 U5035 ( .A1(n9508), .A2(n4710), .ZN(n4709) );
  NOR2_X1 U5036 ( .A1(n9512), .A2(n9531), .ZN(n4537) );
  AND2_X1 U5037 ( .A1(n4758), .A2(n4465), .ZN(n4464) );
  NAND2_X1 U5038 ( .A1(n4466), .A2(n7496), .ZN(n4465) );
  NOR2_X1 U5039 ( .A1(n4761), .A2(n4759), .ZN(n4758) );
  INV_X1 U5040 ( .A(n6518), .ZN(n4759) );
  NAND2_X1 U5041 ( .A1(n7415), .A2(n9104), .ZN(n7414) );
  INV_X1 U5042 ( .A(n4701), .ZN(n4518) );
  NAND3_X1 U5043 ( .A1(n4965), .A2(P1_STATE_REG_SCAN_IN), .A3(n6610), .ZN(
        n6611) );
  XNOR2_X1 U5044 ( .A(n7698), .B(n7697), .ZN(n7701) );
  NAND2_X1 U5045 ( .A1(n4804), .A2(n4805), .ZN(n5582) );
  AND2_X1 U5046 ( .A1(n4806), .A2(n4809), .ZN(n4805) );
  AOI21_X1 U5047 ( .B1(n5554), .B2(n4811), .A(n4810), .ZN(n4809) );
  INV_X1 U5048 ( .A(n5416), .ZN(n4832) );
  AOI21_X1 U5049 ( .B1(n4818), .B2(n4819), .A(n5381), .ZN(n4817) );
  AOI21_X1 U5050 ( .B1(n4681), .B2(n4680), .A(n4337), .ZN(n4678) );
  BUF_X1 U5051 ( .A(n5844), .Z(n6086) );
  INV_X1 U5052 ( .A(n8625), .ZN(n6289) );
  NOR2_X1 U5053 ( .A1(n8298), .A2(n4676), .ZN(n4675) );
  INV_X1 U5054 ( .A(n4906), .ZN(n4676) );
  AOI22_X1 U5055 ( .A1(n7737), .A2(n8637), .B1(n7736), .B2(n7959), .ZN(n7974)
         );
  NAND2_X1 U5056 ( .A1(n4421), .A2(n4420), .ZN(n7737) );
  NOR2_X1 U5057 ( .A1(n8699), .A2(n8439), .ZN(n4420) );
  INV_X1 U5058 ( .A(n7736), .ZN(n4421) );
  INV_X2 U5059 ( .A(n6087), .ZN(n6078) );
  NAND2_X1 U5060 ( .A1(n4641), .A2(n4375), .ZN(n4639) );
  AOI21_X1 U5061 ( .B1(n4749), .B2(n4747), .A(n4351), .ZN(n4746) );
  INV_X1 U5062 ( .A(n7549), .ZN(n4634) );
  OR2_X1 U5063 ( .A1(n7606), .A2(n7605), .ZN(n4720) );
  AND2_X1 U5064 ( .A1(n6256), .A2(n6255), .ZN(n8445) );
  NAND2_X1 U5065 ( .A1(n8465), .A2(n6305), .ZN(n6468) );
  AOI21_X1 U5066 ( .B1(n4573), .B2(n4574), .A(n4390), .ZN(n4570) );
  NAND2_X1 U5067 ( .A1(n8477), .A2(n6302), .ZN(n4566) );
  AOI21_X1 U5068 ( .B1(n8498), .B2(n6299), .A(n4908), .ZN(n8490) );
  AND2_X1 U5069 ( .A1(n5746), .A2(n4687), .ZN(n4686) );
  INV_X1 U5070 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4687) );
  INV_X1 U5071 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5901) );
  INV_X1 U5072 ( .A(n4954), .ZN(n4956) );
  AND2_X1 U5073 ( .A1(n5250), .A2(n5249), .ZN(n7558) );
  INV_X1 U5074 ( .A(n4424), .ZN(n4423) );
  OAI21_X1 U5075 ( .B1(n9088), .B2(n9194), .A(n4965), .ZN(n4424) );
  AOI22_X1 U5076 ( .A1(n9255), .A2(n5036), .B1(n4987), .B2(n4617), .ZN(n5009)
         );
  NAND2_X1 U5077 ( .A1(n4507), .A2(n5083), .ZN(n4843) );
  INV_X1 U5078 ( .A(n5102), .ZN(n4507) );
  NOR2_X1 U5079 ( .A1(n5726), .A2(n6611), .ZN(n5724) );
  INV_X1 U5080 ( .A(n7709), .ZN(n9088) );
  AND2_X1 U5081 ( .A1(n7705), .A2(n7695), .ZN(n5161) );
  AND2_X1 U5082 ( .A1(n9184), .A2(n9186), .ZN(n9120) );
  AOI21_X1 U5083 ( .B1(n9432), .B2(n6530), .A(n6529), .ZN(n9414) );
  NAND2_X1 U5084 ( .A1(n6805), .A2(n6505), .ZN(n6902) );
  NAND2_X1 U5085 ( .A1(n6806), .A2(n8988), .ZN(n6805) );
  NAND2_X1 U5086 ( .A1(n6709), .A2(n6543), .ZN(n7091) );
  AND2_X1 U5087 ( .A1(n5677), .A2(n9754), .ZN(n6751) );
  INV_X1 U5088 ( .A(n5184), .ZN(n9080) );
  NAND2_X1 U5089 ( .A1(n6608), .A2(n4317), .ZN(n5184) );
  NAND2_X1 U5090 ( .A1(n9087), .A2(n6564), .ZN(n9592) );
  AND2_X1 U5091 ( .A1(n4932), .A2(n4871), .ZN(n4870) );
  NOR2_X1 U5092 ( .A1(n4872), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n4871) );
  NAND2_X1 U5093 ( .A1(n5638), .A2(n5637), .ZN(n5696) );
  NAND2_X1 U5094 ( .A1(n5129), .A2(n5128), .ZN(n5148) );
  NAND3_X1 U5095 ( .A1(n4972), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4793) );
  INV_X1 U5096 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4972) );
  INV_X1 U5097 ( .A(n8491), .ZN(n8462) );
  OAI21_X1 U5098 ( .B1(n8898), .B2(n4489), .A(n4488), .ZN(n8807) );
  NAND2_X1 U5099 ( .A1(n5666), .A2(n4491), .ZN(n4488) );
  NAND2_X1 U5100 ( .A1(n5666), .A2(n8874), .ZN(n4489) );
  INV_X1 U5101 ( .A(n6544), .ZN(n4608) );
  OR2_X1 U5102 ( .A1(n7818), .A2(n7817), .ZN(n7823) );
  AOI21_X1 U5103 ( .B1(n8987), .B2(n4620), .A(n7161), .ZN(n4619) );
  NOR2_X1 U5104 ( .A1(n4621), .A2(n9125), .ZN(n4620) );
  NAND2_X1 U5105 ( .A1(n8567), .A2(n7838), .ZN(n4429) );
  AND2_X1 U5106 ( .A1(n7835), .A2(n7894), .ZN(n4430) );
  OR2_X1 U5107 ( .A1(n4601), .A2(n4599), .ZN(n4596) );
  OR2_X1 U5108 ( .A1(n9051), .A2(n9050), .ZN(n4601) );
  INV_X1 U5109 ( .A(n4595), .ZN(n4594) );
  OAI211_X1 U5110 ( .C1(n4599), .C2(n4600), .A(n9063), .B(n9064), .ZN(n4595)
         );
  INV_X1 U5111 ( .A(n9056), .ZN(n4600) );
  OAI21_X1 U5112 ( .B1(n9045), .B2(n9172), .A(n4586), .ZN(n9038) );
  NAND2_X1 U5113 ( .A1(n4336), .A2(n4597), .ZN(n4593) );
  INV_X1 U5114 ( .A(n9050), .ZN(n4598) );
  AOI21_X1 U5115 ( .B1(n9071), .B2(n9125), .A(n9377), .ZN(n4615) );
  OR2_X1 U5116 ( .A1(n4730), .A2(n6832), .ZN(n4729) );
  NAND2_X1 U5117 ( .A1(n4762), .A2(n4371), .ZN(n4761) );
  NAND2_X1 U5118 ( .A1(n6520), .A2(n7675), .ZN(n4762) );
  NAND2_X1 U5119 ( .A1(n4799), .A2(n4798), .ZN(n7698) );
  AOI21_X1 U5120 ( .B1(n4801), .B2(n4803), .A(n4412), .ZN(n4798) );
  NAND2_X1 U5121 ( .A1(n5696), .A2(n4801), .ZN(n4799) );
  INV_X1 U5122 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U5123 ( .A1(n5333), .A2(n5335), .ZN(n4821) );
  INV_X1 U5124 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5212) );
  NOR2_X1 U5125 ( .A1(n6126), .A2(n6125), .ZN(n8004) );
  AND2_X1 U5126 ( .A1(n8273), .A2(n6122), .ZN(n6126) );
  OAI21_X1 U5127 ( .B1(n6072), .B2(n7752), .A(n7441), .ZN(n5796) );
  NAND2_X1 U5128 ( .A1(n6015), .A2(n8266), .ZN(n4665) );
  NAND2_X1 U5129 ( .A1(n6379), .A2(n4727), .ZN(n4726) );
  NAND2_X1 U5130 ( .A1(n4729), .A2(n4723), .ZN(n4722) );
  AND2_X1 U5131 ( .A1(n4730), .A2(n6620), .ZN(n4723) );
  INV_X1 U5132 ( .A(n6379), .ZN(n4730) );
  AND2_X1 U5133 ( .A1(n4729), .A2(n6620), .ZN(n4728) );
  NOR2_X1 U5134 ( .A1(n8360), .A2(n4447), .ZN(n6363) );
  AND2_X1 U5135 ( .A1(n6996), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4447) );
  NAND2_X1 U5136 ( .A1(n6441), .A2(n6442), .ZN(n8427) );
  NAND2_X1 U5137 ( .A1(n7885), .A2(n7882), .ZN(n4876) );
  NAND2_X1 U5138 ( .A1(n8019), .A2(n4881), .ZN(n4880) );
  INV_X1 U5139 ( .A(n6252), .ZN(n4881) );
  NAND2_X1 U5140 ( .A1(n8019), .A2(n8469), .ZN(n4882) );
  NOR2_X1 U5141 ( .A1(n6022), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6036) );
  AND2_X1 U5142 ( .A1(n5923), .A2(n5807), .ZN(n5937) );
  INV_X1 U5143 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5807) );
  NOR2_X1 U5144 ( .A1(n5924), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5923) );
  INV_X1 U5145 ( .A(n6271), .ZN(n4552) );
  OR2_X1 U5146 ( .A1(n8717), .A2(n8500), .ZN(n7878) );
  NAND2_X1 U5147 ( .A1(n4355), .A2(n4558), .ZN(n4557) );
  NAND2_X1 U5148 ( .A1(n6297), .A2(n4559), .ZN(n4558) );
  INV_X1 U5149 ( .A(n6295), .ZN(n4559) );
  AOI21_X1 U5150 ( .B1(n4563), .B2(n8539), .A(n4561), .ZN(n4560) );
  INV_X1 U5151 ( .A(n4564), .ZN(n4563) );
  OAI21_X1 U5152 ( .B1(n8539), .B2(n8538), .A(n4565), .ZN(n4564) );
  INV_X1 U5153 ( .A(n8524), .ZN(n4565) );
  OR2_X1 U5154 ( .A1(n8738), .A2(n8528), .ZN(n7864) );
  AOI21_X1 U5155 ( .B1(n8586), .B2(n4580), .A(n4578), .ZN(n4575) );
  AND2_X1 U5156 ( .A1(n7948), .A2(n7831), .ZN(n6294) );
  INV_X1 U5157 ( .A(n8586), .ZN(n6221) );
  OR2_X1 U5158 ( .A1(n8691), .A2(n6289), .ZN(n7807) );
  AND2_X1 U5159 ( .A1(n6214), .A2(n7791), .ZN(n4896) );
  INV_X1 U5160 ( .A(n6963), .ZN(n6164) );
  AND2_X1 U5161 ( .A1(n5743), .A2(n5744), .ZN(n4452) );
  INV_X1 U5162 ( .A(n8852), .ZN(n4858) );
  NOR2_X1 U5163 ( .A1(n4500), .A2(n4499), .ZN(n4498) );
  INV_X1 U5164 ( .A(n8961), .ZN(n4499) );
  INV_X1 U5165 ( .A(n5409), .ZN(n4867) );
  INV_X1 U5166 ( .A(n4475), .ZN(n4474) );
  OAI21_X1 U5167 ( .B1(n4347), .B2(n4476), .A(n4479), .ZN(n4475) );
  NAND2_X1 U5168 ( .A1(n4480), .A2(n6556), .ZN(n4479) );
  AND2_X1 U5169 ( .A1(n6553), .A2(n4693), .ZN(n4692) );
  OR2_X1 U5170 ( .A1(n9677), .A2(n8845), .ZN(n9175) );
  INV_X1 U5171 ( .A(n4761), .ZN(n4756) );
  OR2_X1 U5172 ( .A1(n9687), .A2(n8965), .ZN(n9031) );
  INV_X1 U5173 ( .A(n6517), .ZN(n4467) );
  AND2_X1 U5174 ( .A1(n7496), .A2(n9017), .ZN(n4324) );
  NAND2_X1 U5175 ( .A1(n5692), .A2(n9126), .ZN(n4966) );
  NAND2_X1 U5176 ( .A1(n5584), .A2(n5583), .ZN(n5606) );
  NAND2_X1 U5177 ( .A1(n4830), .A2(n4829), .ZN(n4828) );
  AOI21_X1 U5178 ( .B1(n4827), .B2(n4830), .A(n4826), .ZN(n4825) );
  INV_X1 U5179 ( .A(n5453), .ZN(n4829) );
  AOI21_X1 U5180 ( .B1(n4835), .B2(n4834), .A(n4386), .ZN(n4833) );
  INV_X1 U5181 ( .A(n4840), .ZN(n4834) );
  INV_X1 U5182 ( .A(n5088), .ZN(n4791) );
  INV_X1 U5183 ( .A(n8058), .ZN(n4683) );
  NAND2_X1 U5184 ( .A1(n6028), .A2(n6029), .ZN(n6030) );
  INV_X1 U5185 ( .A(n8322), .ZN(n4656) );
  AND2_X1 U5187 ( .A1(n8251), .A2(n8252), .ZN(n6099) );
  NAND2_X1 U5188 ( .A1(n5976), .A2(n8338), .ZN(n4668) );
  OR2_X1 U5189 ( .A1(n8102), .A2(n8599), .ZN(n6058) );
  OR2_X1 U5190 ( .A1(n4662), .A2(n4660), .ZN(n4657) );
  INV_X1 U5191 ( .A(n4665), .ZN(n4660) );
  AND2_X1 U5192 ( .A1(n8038), .A2(n4663), .ZN(n4662) );
  AND2_X1 U5193 ( .A1(n6120), .A2(n6119), .ZN(n8062) );
  AND4_X1 U5194 ( .A1(n6095), .A2(n6094), .A3(n6093), .A4(n6092), .ZN(n8063)
         );
  AND4_X1 U5195 ( .A1(n5912), .A2(n5911), .A3(n5910), .A4(n5909), .ZN(n6274)
         );
  OR2_X1 U5196 ( .A1(n4318), .A2(n5853), .ZN(n5858) );
  AND2_X1 U5197 ( .A1(n4716), .A2(n6833), .ZN(n6866) );
  NAND2_X1 U5198 ( .A1(n4718), .A2(n4717), .ZN(n4716) );
  NAND2_X1 U5199 ( .A1(n6865), .A2(n6833), .ZN(n6378) );
  NAND2_X1 U5200 ( .A1(n6866), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6865) );
  NAND2_X1 U5201 ( .A1(n6922), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6949) );
  NAND2_X1 U5202 ( .A1(n6922), .A2(n4363), .ZN(n4636) );
  NAND2_X1 U5203 ( .A1(n6922), .A2(n4642), .ZN(n4640) );
  AND2_X1 U5204 ( .A1(n6381), .A2(n7072), .ZN(n4749) );
  INV_X1 U5205 ( .A(n10022), .ZN(n4747) );
  NAND2_X1 U5206 ( .A1(n4744), .A2(n5926), .ZN(n4743) );
  INV_X1 U5207 ( .A(n4749), .ZN(n4744) );
  NOR2_X1 U5208 ( .A1(n10120), .A2(n6355), .ZN(n7307) );
  NOR2_X1 U5209 ( .A1(n7541), .A2(n7355), .ZN(n4733) );
  NOR2_X1 U5210 ( .A1(n6385), .A2(n4370), .ZN(n6384) );
  AOI21_X1 U5211 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n6701), .A(n7540), .ZN(
        n6386) );
  NOR2_X1 U5212 ( .A1(n7554), .A2(n6404), .ZN(n4633) );
  AND2_X1 U5213 ( .A1(n8427), .A2(n8426), .ZN(n8429) );
  NAND2_X1 U5214 ( .A1(n4652), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4649) );
  INV_X1 U5215 ( .A(n8423), .ZN(n4652) );
  OR2_X1 U5216 ( .A1(n8408), .A2(n4414), .ZN(n4740) );
  OR2_X1 U5217 ( .A1(n4341), .A2(n8421), .ZN(n4739) );
  INV_X1 U5218 ( .A(n4573), .ZN(n4571) );
  AND4_X1 U5219 ( .A1(n6069), .A2(n6068), .A3(n6067), .A4(n6066), .ZN(n8590)
         );
  OR2_X1 U5220 ( .A1(n5962), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U5221 ( .A1(n7330), .A2(n6270), .ZN(n4553) );
  NAND2_X1 U5222 ( .A1(n7329), .A2(n7783), .ZN(n4895) );
  NAND2_X1 U5223 ( .A1(n6967), .A2(n6966), .ZN(n7038) );
  AND3_X1 U5224 ( .A1(n6965), .A2(n6964), .A3(n6963), .ZN(n6966) );
  OR2_X1 U5225 ( .A1(n10104), .A2(n7752), .ZN(n6321) );
  NAND2_X1 U5226 ( .A1(n6243), .A2(n6242), .ZN(n8028) );
  OR2_X1 U5227 ( .A1(n7925), .A2(n7924), .ZN(n8513) );
  INV_X1 U5228 ( .A(n8513), .ZN(n8511) );
  NAND2_X1 U5229 ( .A1(n4562), .A2(n4560), .ZN(n8521) );
  NAND2_X1 U5230 ( .A1(n8537), .A2(n4563), .ZN(n4562) );
  NOR2_X1 U5231 ( .A1(n6224), .A2(n7856), .ZN(n4894) );
  AND2_X1 U5232 ( .A1(n4892), .A2(n7864), .ZN(n4891) );
  OR2_X1 U5233 ( .A1(n6224), .A2(n4893), .ZN(n4892) );
  NAND2_X1 U5234 ( .A1(n6223), .A2(n7847), .ZN(n4893) );
  CLKBUF_X1 U5235 ( .A(n8548), .Z(n8550) );
  NAND2_X1 U5236 ( .A1(n4577), .A2(n8586), .ZN(n4576) );
  INV_X1 U5237 ( .A(n8597), .ZN(n4577) );
  INV_X1 U5238 ( .A(n4575), .ZN(n4574) );
  INV_X1 U5239 ( .A(n6294), .ZN(n8575) );
  OR2_X1 U5240 ( .A1(n8761), .A2(n8589), .ZN(n7835) );
  AND2_X1 U5241 ( .A1(n6293), .A2(n6292), .ZN(n8598) );
  AND2_X1 U5242 ( .A1(n7835), .A2(n7827), .ZN(n8597) );
  AOI21_X1 U5243 ( .B1(n4542), .B2(n6290), .A(n7815), .ZN(n4541) );
  INV_X1 U5244 ( .A(n8624), .ZN(n10037) );
  NAND2_X1 U5245 ( .A1(n6312), .A2(n7910), .ZN(n10039) );
  INV_X1 U5246 ( .A(n7945), .ZN(n8610) );
  INV_X1 U5247 ( .A(n6083), .ZN(n6073) );
  INV_X1 U5248 ( .A(n4549), .ZN(n4548) );
  OAI21_X1 U5249 ( .B1(n6290), .B2(n6287), .A(n4381), .ZN(n4549) );
  AND2_X1 U5250 ( .A1(n7807), .A2(n7808), .ZN(n7942) );
  NAND2_X1 U5251 ( .A1(n6306), .A2(n7971), .ZN(n8627) );
  INV_X1 U5252 ( .A(n10039), .ZN(n8622) );
  NOR2_X1 U5253 ( .A1(n6965), .A2(n6164), .ZN(n6329) );
  INV_X1 U5254 ( .A(n8627), .ZN(n10050) );
  AND2_X1 U5255 ( .A1(n6339), .A2(n6693), .ZN(n6658) );
  INV_X1 U5256 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5798) );
  INV_X1 U5257 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U5258 ( .A1(n5764), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5766) );
  INV_X1 U5259 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5765) );
  XNOR2_X1 U5260 ( .A(n6162), .B(n6163), .ZN(n7638) );
  NAND2_X1 U5261 ( .A1(n5791), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U5262 ( .A1(n4862), .A2(n4861), .ZN(n4859) );
  INV_X1 U5263 ( .A(n5171), .ZN(n4861) );
  OR2_X1 U5264 ( .A1(n5268), .A2(n7255), .ZN(n5289) );
  OR2_X1 U5265 ( .A1(n7626), .A2(n7558), .ZN(n5251) );
  AND2_X1 U5266 ( .A1(n8891), .A2(n8892), .ZN(n5409) );
  AND3_X1 U5267 ( .A1(n4859), .A2(n5173), .A3(n4858), .ZN(n8850) );
  NOR2_X1 U5268 ( .A1(n5003), .A2(n5001), .ZN(n6719) );
  XNOR2_X1 U5269 ( .A(n4508), .B(n5710), .ZN(n5102) );
  INV_X1 U5270 ( .A(n5101), .ZN(n4508) );
  INV_X1 U5271 ( .A(n5083), .ZN(n4848) );
  NAND2_X1 U5272 ( .A1(n8874), .A2(n4493), .ZN(n4492) );
  INV_X1 U5273 ( .A(n5580), .ZN(n4493) );
  NAND2_X1 U5274 ( .A1(n5351), .A2(n5350), .ZN(n4864) );
  OAI21_X1 U5275 ( .B1(n9620), .B2(n4628), .A(n4627), .ZN(n4626) );
  NAND2_X1 U5276 ( .A1(n9084), .A2(n9620), .ZN(n4629) );
  AND2_X1 U5277 ( .A1(n9706), .A2(n9355), .ZN(n9213) );
  NAND2_X1 U5278 ( .A1(n9089), .A2(n4623), .ZN(n9222) );
  NOR2_X1 U5279 ( .A1(n4316), .A2(n4340), .ZN(n4623) );
  OR2_X1 U5280 ( .A1(n5011), .A2(n6626), .ZN(n4991) );
  NOR3_X1 U5281 ( .A1(n9258), .A2(n6626), .A3(n9271), .ZN(n9257) );
  OR2_X1 U5282 ( .A1(n5022), .A2(n9756), .ZN(n5072) );
  NOR2_X1 U5283 ( .A1(n6670), .A2(n4360), .ZN(n9295) );
  AOI21_X1 U5284 ( .B1(n9831), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9823), .ZN(
        n9840) );
  OR2_X1 U5285 ( .A1(n9840), .A2(n9839), .ZN(n9842) );
  AND2_X1 U5286 ( .A1(n9321), .A2(n9857), .ZN(n9322) );
  NOR2_X1 U5287 ( .A1(n4528), .A2(n8978), .ZN(n4527) );
  INV_X1 U5288 ( .A(n4328), .ZN(n4528) );
  NOR2_X1 U5289 ( .A1(n4770), .A2(n4768), .ZN(n4767) );
  INV_X1 U5290 ( .A(n6531), .ZN(n4768) );
  OAI21_X1 U5291 ( .B1(n4770), .B2(n4775), .A(n4769), .ZN(n4766) );
  AOI21_X1 U5292 ( .B1(n4772), .B2(n9393), .A(n4380), .ZN(n4769) );
  AND2_X1 U5293 ( .A1(n9127), .A2(n9066), .ZN(n9413) );
  AOI21_X1 U5294 ( .B1(n9443), .B2(n6528), .A(n6527), .ZN(n9432) );
  AND2_X1 U5295 ( .A1(n9059), .A2(n9060), .ZN(n9466) );
  NAND2_X1 U5296 ( .A1(n4329), .A2(n4377), .ZN(n4477) );
  NAND2_X1 U5297 ( .A1(n6525), .A2(n4343), .ZN(n4478) );
  NOR2_X1 U5298 ( .A1(n9484), .A2(n4535), .ZN(n4533) );
  NOR2_X1 U5299 ( .A1(n9512), .A2(n9525), .ZN(n6523) );
  NAND2_X1 U5300 ( .A1(n4708), .A2(n4366), .ZN(n9491) );
  OR2_X1 U5301 ( .A1(n8981), .A2(n9240), .ZN(n6519) );
  NAND2_X1 U5302 ( .A1(n6552), .A2(n9108), .ZN(n7568) );
  AND2_X1 U5303 ( .A1(n9021), .A2(n9166), .ZN(n9108) );
  OAI21_X1 U5304 ( .B1(n7420), .B2(n7496), .A(n4466), .ZN(n9588) );
  OR2_X1 U5305 ( .A1(n7434), .A2(n7586), .ZN(n9017) );
  INV_X1 U5306 ( .A(n4441), .ZN(n4699) );
  NAND2_X1 U5307 ( .A1(n4441), .A2(n4324), .ZN(n7494) );
  OR2_X1 U5308 ( .A1(n7434), .A2(n9243), .ZN(n6517) );
  AOI21_X1 U5309 ( .B1(n7506), .B2(n4780), .A(n4379), .ZN(n4779) );
  NAND2_X1 U5310 ( .A1(n7270), .A2(n6514), .ZN(n7505) );
  NAND2_X1 U5311 ( .A1(n7263), .A2(n9091), .ZN(n7262) );
  INV_X1 U5312 ( .A(n4753), .ZN(n4752) );
  OAI21_X1 U5313 ( .B1(n6909), .B2(n4754), .A(n7056), .ZN(n4753) );
  INV_X1 U5314 ( .A(n6507), .ZN(n4754) );
  NAND2_X1 U5315 ( .A1(n6902), .A2(n6909), .ZN(n6901) );
  NAND2_X1 U5316 ( .A1(n6763), .A2(n6502), .ZN(n6806) );
  AND2_X1 U5317 ( .A1(n9212), .A2(n6649), .ZN(n9563) );
  NAND2_X1 U5318 ( .A1(n5537), .A2(n5536), .ZN(n9462) );
  INV_X1 U5319 ( .A(n9944), .ZN(n9953) );
  INV_X1 U5320 ( .A(n6596), .ZN(n4519) );
  NAND2_X1 U5321 ( .A1(n5675), .A2(n5674), .ZN(n9753) );
  AOI21_X1 U5322 ( .B1(n5673), .B2(n8222), .A(n9770), .ZN(n5674) );
  XNOR2_X1 U5323 ( .A(n7731), .B(n7730), .ZN(n8975) );
  OAI21_X1 U5324 ( .B1(n7726), .B2(n7725), .A(n7724), .ZN(n7731) );
  NAND4_X1 U5325 ( .A1(n4929), .A2(n4932), .A3(n4928), .A4(n4712), .ZN(n4971)
         );
  INV_X1 U5326 ( .A(n4872), .ZN(n4712) );
  INV_X1 U5327 ( .A(n4971), .ZN(n4444) );
  NOR2_X1 U5328 ( .A1(n5529), .A2(n4808), .ZN(n4807) );
  INV_X1 U5329 ( .A(n5504), .ZN(n4808) );
  NAND2_X1 U5330 ( .A1(n4815), .A2(n4814), .ZN(n4813) );
  NOR2_X1 U5331 ( .A1(n4378), .A2(n4514), .ZN(n4513) );
  NAND2_X1 U5332 ( .A1(n4515), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4947) );
  NAND2_X1 U5333 ( .A1(n5418), .A2(n4512), .ZN(n4515) );
  INV_X1 U5334 ( .A(n4514), .ZN(n4512) );
  NAND2_X1 U5335 ( .A1(n4947), .A2(n4946), .ZN(n4951) );
  NAND2_X1 U5336 ( .A1(n4824), .A2(n4830), .ZN(n5454) );
  NAND2_X1 U5337 ( .A1(n5415), .A2(n4831), .ZN(n4824) );
  NAND2_X1 U5338 ( .A1(n4944), .A2(n5418), .ZN(n5422) );
  NAND2_X1 U5339 ( .A1(n4816), .A2(n4819), .ZN(n5382) );
  NAND2_X1 U5340 ( .A1(n5334), .A2(n4822), .ZN(n4816) );
  OAI21_X1 U5341 ( .B1(n5334), .B2(n5333), .A(n5335), .ZN(n5359) );
  AND2_X1 U5342 ( .A1(n5265), .A2(n5284), .ZN(n9331) );
  NAND2_X1 U5343 ( .A1(n4837), .A2(n4838), .ZN(n5283) );
  NAND2_X1 U5344 ( .A1(n5234), .A2(n4840), .ZN(n4837) );
  OR2_X1 U5345 ( .A1(n5235), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5261) );
  XNOR2_X1 U5346 ( .A(n5234), .B(n5233), .ZN(n6698) );
  NOR2_X1 U5347 ( .A1(n5133), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5218) );
  XNOR2_X1 U5348 ( .A(n5105), .B(SI_5_), .ZN(n5103) );
  INV_X1 U5349 ( .A(n5830), .ZN(n6342) );
  NOR2_X1 U5350 ( .A1(n8045), .A2(n8336), .ZN(n8044) );
  AND4_X1 U5351 ( .A1(n5814), .A2(n5813), .A3(n5812), .A4(n5811), .ZN(n7535)
         );
  NAND2_X1 U5352 ( .A1(n4674), .A2(n4672), .ZN(n8253) );
  AND2_X1 U5353 ( .A1(n4673), .A2(n8051), .ZN(n4672) );
  INV_X1 U5354 ( .A(n6071), .ZN(n4673) );
  INV_X1 U5355 ( .A(n8337), .ZN(n8612) );
  AND3_X1 U5356 ( .A1(n6137), .A2(n6136), .A3(n6135), .ZN(n8088) );
  INV_X1 U5357 ( .A(n7013), .ZN(n5885) );
  AND4_X1 U5358 ( .A1(n6082), .A2(n6081), .A3(n6080), .A4(n6079), .ZN(n8300)
         );
  INV_X1 U5359 ( .A(n8317), .ZN(n8326) );
  INV_X1 U5360 ( .A(n8305), .ZN(n8320) );
  NAND2_X1 U5361 ( .A1(n7920), .A2(n7918), .ZN(n7921) );
  NAND2_X1 U5362 ( .A1(n7976), .A2(n7975), .ZN(n4786) );
  OR2_X1 U5363 ( .A1(n7974), .A2(n7739), .ZN(n7976) );
  NAND2_X1 U5364 ( .A1(n7967), .A2(n7738), .ZN(n7739) );
  INV_X1 U5365 ( .A(n6181), .ZN(n7978) );
  CLKBUF_X1 U5366 ( .A(n6180), .Z(n7977) );
  XNOR2_X1 U5367 ( .A(n6157), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7980) );
  AND2_X1 U5368 ( .A1(n7723), .A2(n6311), .ZN(n8024) );
  NAND2_X1 U5369 ( .A1(n6262), .A2(n6261), .ZN(n8335) );
  NAND2_X1 U5370 ( .A1(n6241), .A2(n6240), .ZN(n8491) );
  INV_X1 U5371 ( .A(n8088), .ZN(n8514) );
  INV_X1 U5372 ( .A(n8062), .ZN(n8542) );
  INV_X1 U5373 ( .A(n8300), .ZN(n8577) );
  INV_X1 U5374 ( .A(n8590), .ZN(n8560) );
  INV_X1 U5375 ( .A(n8101), .ZN(n8599) );
  INV_X1 U5376 ( .A(n6274), .ZN(n8343) );
  NOR2_X1 U5377 ( .A1(n6383), .A2(n6427), .ZN(n6385) );
  NAND2_X1 U5378 ( .A1(n4738), .A2(n4349), .ZN(n4737) );
  AND2_X1 U5379 ( .A1(n4737), .A2(n4736), .ZN(n8350) );
  INV_X1 U5380 ( .A(n8351), .ZN(n4736) );
  INV_X1 U5381 ( .A(n4651), .ZN(n8406) );
  NAND2_X1 U5382 ( .A1(n8408), .A2(n8592), .ZN(n4457) );
  OR2_X1 U5383 ( .A1(n4435), .A2(n8411), .ZN(n4434) );
  INV_X1 U5384 ( .A(n4436), .ZN(n4435) );
  NAND2_X1 U5385 ( .A1(n6254), .A2(n6253), .ZN(n8458) );
  NAND2_X1 U5386 ( .A1(n6116), .A2(n6115), .ZN(n8533) );
  AND3_X1 U5387 ( .A1(n5905), .A2(n5904), .A3(n5903), .ZN(n10042) );
  AOI21_X1 U5388 ( .B1(n7685), .B2(n7732), .A(n6132), .ZN(n8722) );
  NAND2_X1 U5389 ( .A1(n5644), .A2(n5643), .ZN(n9402) );
  OR2_X1 U5390 ( .A1(n5734), .A2(n8946), .ZN(n5735) );
  NOR2_X1 U5391 ( .A1(n6725), .A2(n6726), .ZN(n6724) );
  NOR2_X1 U5392 ( .A1(n4487), .A2(n8933), .ZN(n4485) );
  AOI21_X1 U5393 ( .B1(n6781), .B2(n6780), .A(n4916), .ZN(n8911) );
  AND2_X1 U5394 ( .A1(n5724), .A2(n5694), .ZN(n9806) );
  OR2_X1 U5395 ( .A1(n4313), .A2(n5054), .ZN(n5063) );
  OR2_X1 U5396 ( .A1(n5059), .A2(n6637), .ZN(n4942) );
  NAND2_X1 U5397 ( .A1(n4331), .A2(n4940), .ZN(n4852) );
  XNOR2_X1 U5398 ( .A(n4976), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9261) );
  NAND2_X1 U5399 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4976) );
  AOI21_X1 U5400 ( .B1(n9792), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9787), .ZN(
        n6737) );
  NOR2_X1 U5401 ( .A1(n9851), .A2(n9852), .ZN(n9850) );
  NAND2_X1 U5402 ( .A1(n6535), .A2(n6534), .ZN(n9370) );
  NAND2_X1 U5403 ( .A1(n9381), .A2(n4468), .ZN(n9627) );
  NAND2_X1 U5404 ( .A1(n4773), .A2(n4772), .ZN(n9381) );
  NAND2_X1 U5405 ( .A1(n4470), .A2(n4469), .ZN(n4468) );
  NAND2_X1 U5406 ( .A1(n4773), .A2(n4774), .ZN(n4470) );
  XNOR2_X1 U5407 ( .A(n4700), .B(n4469), .ZN(n9380) );
  AND2_X1 U5408 ( .A1(n9374), .A2(n9944), .ZN(n4433) );
  NAND2_X1 U5409 ( .A1(n5137), .A2(n5136), .ZN(n7208) );
  NAND2_X1 U5410 ( .A1(n4936), .A2(n4937), .ZN(n9757) );
  AND2_X1 U5411 ( .A1(n7791), .A2(n7790), .ZN(n4427) );
  NAND2_X1 U5412 ( .A1(n4606), .A2(n4605), .ZN(n8989) );
  NOR2_X1 U5413 ( .A1(n4608), .A2(n9125), .ZN(n4607) );
  NAND2_X1 U5414 ( .A1(n8982), .A2(n9098), .ZN(n4604) );
  NAND2_X1 U5415 ( .A1(n4622), .A2(n4619), .ZN(n4618) );
  AOI21_X1 U5416 ( .B1(n7836), .B2(n4430), .A(n4429), .ZN(n7839) );
  NAND2_X1 U5417 ( .A1(n7868), .A2(n4368), .ZN(n4455) );
  AOI22_X1 U5418 ( .A1(n9034), .A2(n4628), .B1(n9036), .B2(n9035), .ZN(n4588)
         );
  NAND2_X1 U5419 ( .A1(n9033), .A2(n9125), .ZN(n4589) );
  NOR2_X1 U5420 ( .A1(n4710), .A2(n4587), .ZN(n4586) );
  INV_X1 U5421 ( .A(n9042), .ZN(n4587) );
  NAND2_X1 U5422 ( .A1(n4591), .A2(n4597), .ZN(n4590) );
  NAND2_X1 U5423 ( .A1(n4596), .A2(n4594), .ZN(n4591) );
  NAND2_X1 U5424 ( .A1(n7959), .A2(n7903), .ZN(n4454) );
  INV_X1 U5425 ( .A(n4802), .ZN(n4801) );
  OAI21_X1 U5426 ( .B1(n5695), .B2(n4803), .A(n6458), .ZN(n4802) );
  INV_X1 U5427 ( .A(n5697), .ZN(n4803) );
  NAND2_X1 U5428 ( .A1(n4505), .A2(n7108), .ZN(n4504) );
  INV_X1 U5429 ( .A(n5123), .ZN(n4505) );
  INV_X1 U5430 ( .A(n9183), .ZN(n4611) );
  NAND2_X1 U5431 ( .A1(n4614), .A2(n4613), .ZN(n4612) );
  INV_X1 U5432 ( .A(n9141), .ZN(n4613) );
  NAND2_X1 U5433 ( .A1(n4616), .A2(n4615), .ZN(n4614) );
  NAND2_X1 U5434 ( .A1(n9072), .A2(n4628), .ZN(n4616) );
  OR2_X1 U5435 ( .A1(n9387), .A2(n6569), .ZN(n9183) );
  INV_X1 U5436 ( .A(n5528), .ZN(n4811) );
  INV_X1 U5437 ( .A(n5556), .ZN(n4810) );
  NOR2_X1 U5438 ( .A1(n4831), .A2(n5453), .ZN(n4827) );
  INV_X1 U5439 ( .A(n5452), .ZN(n4826) );
  INV_X1 U5440 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4923) );
  INV_X1 U5441 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4924) );
  INV_X1 U5442 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5387) );
  INV_X1 U5443 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5386) );
  INV_X1 U5444 ( .A(n4822), .ZN(n4818) );
  INV_X1 U5445 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n5336) );
  NOR2_X1 U5446 ( .A1(n5261), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5315) );
  INV_X1 U5447 ( .A(SI_11_), .ZN(n5213) );
  INV_X1 U5448 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U5449 ( .A1(n7448), .A2(n5961), .ZN(n5973) );
  NAND2_X1 U5450 ( .A1(n4788), .A2(n4787), .ZN(n7959) );
  AND2_X1 U5451 ( .A1(n8334), .A2(n7715), .ZN(n4787) );
  NAND2_X1 U5452 ( .A1(n4898), .A2(n5777), .ZN(n5755) );
  AOI21_X1 U5453 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n6660), .A(n10005), .ZN(
        n6354) );
  NOR2_X1 U5454 ( .A1(n10022), .A2(n5926), .ZN(n4745) );
  NOR2_X1 U5455 ( .A1(n6133), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6185) );
  AND2_X1 U5456 ( .A1(n6089), .A2(n6088), .ZN(n6103) );
  NOR2_X1 U5457 ( .A1(n6076), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6089) );
  NOR2_X1 U5458 ( .A1(n5982), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5996) );
  INV_X1 U5459 ( .A(n7457), .ZN(n7799) );
  OR2_X1 U5460 ( .A1(n6298), .A2(n8088), .ZN(n7923) );
  INV_X1 U5461 ( .A(n7740), .ZN(n4888) );
  INV_X1 U5462 ( .A(n4894), .ZN(n4889) );
  AND2_X1 U5463 ( .A1(n7998), .A2(n8613), .ZN(n7824) );
  OR2_X1 U5464 ( .A1(n7998), .A2(n8613), .ZN(n7826) );
  OR2_X1 U5465 ( .A1(n7535), .A2(n8294), .ZN(n7803) );
  INV_X1 U5466 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6163) );
  INV_X1 U5467 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5785) );
  INV_X1 U5468 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5742) );
  NOR2_X1 U5469 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n4511) );
  AND2_X1 U5470 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5094) );
  AND2_X1 U5471 ( .A1(n4860), .A2(n4858), .ZN(n4857) );
  INV_X1 U5472 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5288) );
  NOR2_X1 U5473 ( .A1(n9370), .A2(n9387), .ZN(n4530) );
  INV_X1 U5474 ( .A(n9233), .ZN(n6532) );
  OR2_X1 U5475 ( .A1(n9402), .A2(n6532), .ZN(n9075) );
  INV_X1 U5476 ( .A(n7506), .ZN(n4781) );
  NOR2_X1 U5477 ( .A1(n4781), .A2(n4778), .ZN(n4777) );
  INV_X1 U5478 ( .A(n6515), .ZN(n4780) );
  OR2_X1 U5479 ( .A1(n9610), .A2(n6511), .ZN(n9008) );
  NAND2_X1 U5480 ( .A1(n4751), .A2(n4750), .ZN(n7162) );
  AOI21_X1 U5481 ( .B1(n4752), .B2(n4754), .A(n4382), .ZN(n4750) );
  NAND2_X1 U5482 ( .A1(n4752), .A2(n6902), .ZN(n4751) );
  NAND2_X1 U5483 ( .A1(n7162), .A2(n7161), .ZN(n7160) );
  NOR2_X2 U5484 ( .A1(n9256), .A2(n6684), .ZN(n6706) );
  OAI21_X1 U5485 ( .B1(n7701), .B2(n7700), .A(n7699), .ZN(n7726) );
  NAND2_X1 U5486 ( .A1(n4933), .A2(n4873), .ZN(n4872) );
  AND2_X1 U5487 ( .A1(n5637), .A2(n5612), .ZN(n5635) );
  AND2_X1 U5488 ( .A1(n5607), .A2(n5588), .ZN(n5605) );
  AND2_X1 U5489 ( .A1(n5583), .A2(n5560), .ZN(n5581) );
  NAND2_X1 U5490 ( .A1(n4944), .A2(n4949), .ZN(n4514) );
  INV_X1 U5491 ( .A(SI_20_), .ZN(n5480) );
  AOI21_X1 U5492 ( .B1(n4831), .B2(n5414), .A(n4403), .ZN(n4830) );
  NAND2_X1 U5493 ( .A1(n5389), .A2(n5388), .ZN(n5416) );
  INV_X1 U5494 ( .A(SI_17_), .ZN(n5388) );
  NOR2_X1 U5495 ( .A1(n5358), .A2(n4823), .ZN(n4822) );
  INV_X1 U5496 ( .A(n5335), .ZN(n4823) );
  NAND2_X1 U5497 ( .A1(n5311), .A2(n5310), .ZN(n5335) );
  INV_X1 U5498 ( .A(SI_14_), .ZN(n5310) );
  AOI21_X1 U5499 ( .B1(n4840), .B2(n5211), .A(n4839), .ZN(n4838) );
  INV_X1 U5500 ( .A(n5260), .ZN(n4839) );
  NOR2_X1 U5501 ( .A1(n5258), .A2(n4841), .ZN(n4840) );
  INV_X1 U5502 ( .A(n5210), .ZN(n4841) );
  OAI21_X1 U5503 ( .B1(n4317), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n5047), .ZN(
        n5066) );
  INV_X1 U5504 ( .A(n8263), .ZN(n4663) );
  AND2_X1 U5505 ( .A1(n6070), .A2(n8590), .ZN(n6071) );
  AND2_X1 U5506 ( .A1(n8307), .A2(n8009), .ZN(n8082) );
  NAND2_X1 U5507 ( .A1(n4677), .A2(n4681), .ZN(n8273) );
  NAND2_X1 U5508 ( .A1(n4666), .A2(n7522), .ZN(n4669) );
  AND2_X1 U5509 ( .A1(n5974), .A2(n4667), .ZN(n4666) );
  INV_X1 U5510 ( .A(n8291), .ZN(n4667) );
  OR2_X1 U5511 ( .A1(n6059), .A2(n8101), .ZN(n4906) );
  INV_X1 U5512 ( .A(n7919), .ZN(n4784) );
  NAND2_X1 U5513 ( .A1(n4425), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9971) );
  OR2_X1 U5514 ( .A1(n9963), .A2(n9962), .ZN(n9965) );
  NAND2_X1 U5515 ( .A1(n9971), .A2(n6375), .ZN(n9991) );
  OAI22_X1 U5516 ( .A1(n9999), .A2(n10000), .B1(n9989), .B2(n6410), .ZN(n6873)
         );
  NAND2_X1 U5517 ( .A1(n6863), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6862) );
  AND2_X1 U5518 ( .A1(n4722), .A2(n4725), .ZN(n4721) );
  OR2_X1 U5519 ( .A1(n6832), .A2(n4726), .ZN(n4725) );
  OAI21_X1 U5520 ( .B1(n6378), .B2(n4730), .A(n4728), .ZN(n6380) );
  OAI21_X1 U5521 ( .B1(n6944), .B2(n6942), .A(n6943), .ZN(n6946) );
  NOR2_X1 U5522 ( .A1(n5947), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5969) );
  NOR2_X1 U5523 ( .A1(n6431), .A2(n7542), .ZN(n7645) );
  INV_X1 U5524 ( .A(n4738), .ZN(n7664) );
  AND2_X1 U5525 ( .A1(n4720), .A2(n4719), .ZN(n6389) );
  NAND2_X1 U5526 ( .A1(n6788), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4719) );
  NAND2_X1 U5527 ( .A1(n4646), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4645) );
  INV_X1 U5528 ( .A(n8361), .ZN(n4646) );
  AND2_X1 U5529 ( .A1(n6996), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4735) );
  INV_X1 U5530 ( .A(n8409), .ZN(n4437) );
  INV_X1 U5531 ( .A(n8427), .ZN(n8425) );
  NAND2_X1 U5532 ( .A1(n6466), .A2(n6465), .ZN(n6470) );
  NOR2_X1 U5533 ( .A1(n4875), .A2(n4335), .ZN(n4874) );
  NOR2_X1 U5534 ( .A1(n4882), .A2(n4876), .ZN(n4875) );
  NOR2_X1 U5535 ( .A1(n4882), .A2(n7886), .ZN(n4878) );
  OR2_X1 U5536 ( .A1(n8445), .A2(n6257), .ZN(n8452) );
  NOR2_X1 U5537 ( .A1(n6244), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6256) );
  OR2_X1 U5538 ( .A1(n6235), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6244) );
  OR2_X1 U5539 ( .A1(n6117), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U5540 ( .A1(n6103), .A2(n8061), .ZN(n6117) );
  NAND2_X1 U5541 ( .A1(n6051), .A2(n6050), .ZN(n6064) );
  OR2_X1 U5542 ( .A1(n5964), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5982) );
  INV_X1 U5543 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5808) );
  CLKBUF_X1 U5544 ( .A(n7339), .Z(n7364) );
  AND4_X1 U5545 ( .A1(n5930), .A2(n5929), .A3(n5928), .A4(n5927), .ZN(n10038)
         );
  NOR2_X1 U5546 ( .A1(n4345), .A2(n4552), .ZN(n4551) );
  OR2_X1 U5547 ( .A1(n5907), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5924) );
  INV_X1 U5548 ( .A(n7376), .ZN(n7929) );
  INV_X1 U5549 ( .A(n6264), .ZN(n7927) );
  NAND2_X1 U5550 ( .A1(n6207), .A2(n7926), .ZN(n6879) );
  OR2_X1 U5551 ( .A1(n6143), .A2(n6155), .ZN(n6963) );
  NAND2_X1 U5552 ( .A1(n7713), .A2(n7732), .ZN(n4788) );
  NAND2_X1 U5553 ( .A1(n6464), .A2(n6463), .ZN(n6491) );
  OR2_X1 U5554 ( .A1(n7885), .A2(n7886), .ZN(n8476) );
  AND2_X1 U5555 ( .A1(n7878), .A2(n7879), .ZN(n8488) );
  AND2_X1 U5556 ( .A1(n7923), .A2(n7922), .ZN(n8505) );
  OR2_X1 U5557 ( .A1(n4392), .A2(n4557), .ZN(n4555) );
  AND4_X1 U5558 ( .A1(n6110), .A2(n6109), .A3(n6108), .A4(n6107), .ZN(n8528)
         );
  AOI21_X1 U5559 ( .B1(n8537), .B2(n8538), .A(n8539), .ZN(n8522) );
  AOI21_X1 U5560 ( .B1(n4569), .B2(n4568), .A(n4567), .ZN(n8552) );
  NOR2_X1 U5561 ( .A1(n4571), .A2(n8567), .ZN(n4568) );
  OAI21_X1 U5562 ( .B1(n4570), .B2(n8567), .A(n4384), .ZN(n4567) );
  NAND2_X1 U5563 ( .A1(n8552), .A2(n8551), .ZN(n8537) );
  NOR2_X1 U5564 ( .A1(n4543), .A2(n4348), .ZN(n4540) );
  OAI21_X1 U5565 ( .B1(n4541), .B2(n4348), .A(n4322), .ZN(n4539) );
  NAND2_X1 U5566 ( .A1(n4897), .A2(n7791), .ZN(n7354) );
  AND3_X1 U5567 ( .A1(n5921), .A2(n5920), .A3(n5919), .ZN(n10083) );
  OR2_X1 U5568 ( .A1(n7919), .A2(n7980), .ZN(n10104) );
  XNOR2_X1 U5569 ( .A(n5773), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U5570 ( .A1(n4353), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5773) );
  XNOR2_X1 U5571 ( .A(n5780), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7752) );
  OR2_X1 U5572 ( .A1(n6004), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U5573 ( .A1(n5747), .A2(n5758), .ZN(n5947) );
  CLKBUF_X1 U5574 ( .A(n5757), .Z(n5917) );
  NAND2_X1 U5575 ( .A1(n5829), .A2(n5828), .ZN(n9960) );
  NAND2_X1 U5576 ( .A1(n4956), .A2(n4511), .ZN(n5667) );
  AND2_X1 U5577 ( .A1(n4511), .A2(n5671), .ZN(n4510) );
  OR2_X1 U5578 ( .A1(n5289), .A2(n5288), .ZN(n5321) );
  AND2_X1 U5579 ( .A1(n5329), .A2(n5303), .ZN(n4516) );
  AND2_X1 U5580 ( .A1(n8901), .A2(n5553), .ZN(n8826) );
  INV_X1 U5581 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7255) );
  INV_X1 U5582 ( .A(n4846), .ZN(n4845) );
  INV_X1 U5583 ( .A(n4843), .ZN(n4851) );
  NAND2_X1 U5584 ( .A1(n4865), .A2(n8960), .ZN(n8882) );
  INV_X1 U5585 ( .A(n8826), .ZN(n4487) );
  NAND2_X1 U5586 ( .A1(n4486), .A2(n8826), .ZN(n8828) );
  NAND2_X1 U5587 ( .A1(n8824), .A2(n8825), .ZN(n4486) );
  AND2_X1 U5588 ( .A1(n5474), .A2(n5473), .ZN(n8924) );
  AOI21_X1 U5589 ( .B1(n4868), .B2(n4867), .A(n4388), .ZN(n4866) );
  NAND2_X1 U5590 ( .A1(n5459), .A2(n5458), .ZN(n5487) );
  INV_X1 U5591 ( .A(n5461), .ZN(n5459) );
  NAND2_X1 U5592 ( .A1(n7583), .A2(n7584), .ZN(n7582) );
  OR2_X1 U5593 ( .A1(n5241), .A2(n5224), .ZN(n5268) );
  XNOR2_X1 U5594 ( .A(n4986), .B(n4985), .ZN(n5007) );
  NAND2_X1 U5595 ( .A1(n9255), .A2(n4987), .ZN(n4984) );
  AND2_X1 U5596 ( .A1(n8890), .A2(n5413), .ZN(n8837) );
  AND2_X1 U5597 ( .A1(n5692), .A2(n9088), .ZN(n9212) );
  NAND2_X1 U5598 ( .A1(n5320), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5342) );
  INV_X1 U5599 ( .A(n5321), .ZN(n5320) );
  INV_X1 U5600 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5341) );
  INV_X1 U5601 ( .A(n4966), .ZN(n6538) );
  NOR2_X1 U5602 ( .A1(n9257), .A2(n4344), .ZN(n9284) );
  NOR2_X1 U5603 ( .A1(n9295), .A2(n9294), .ZN(n9293) );
  AOI21_X1 U5604 ( .B1(n9311), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9304), .ZN(
        n6674) );
  NOR2_X1 U5605 ( .A1(n6789), .A2(n4439), .ZN(n6792) );
  NOR2_X1 U5606 ( .A1(n4440), .A2(n6735), .ZN(n4439) );
  INV_X1 U5607 ( .A(n6798), .ZN(n4440) );
  NAND2_X1 U5608 ( .A1(n6792), .A2(n6791), .ZN(n7248) );
  AOI21_X1 U5609 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n9780), .A(n9775), .ZN(
        n9816) );
  AOI21_X1 U5610 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9819), .A(n9814), .ZN(
        n7253) );
  OR2_X1 U5611 ( .A1(n5360), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U5612 ( .A1(n9874), .A2(n4415), .ZN(n9892) );
  OR2_X1 U5613 ( .A1(n9882), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4415) );
  OR2_X1 U5614 ( .A1(n9891), .A2(n9892), .ZN(n9888) );
  INV_X1 U5615 ( .A(n9232), .ZN(n6569) );
  INV_X1 U5616 ( .A(n9120), .ZN(n9078) );
  AND2_X1 U5617 ( .A1(n9382), .A2(n4774), .ZN(n4772) );
  NAND2_X1 U5618 ( .A1(n9715), .A2(n6532), .ZN(n4774) );
  OR2_X1 U5619 ( .A1(n5538), .A2(n8833), .ZN(n5594) );
  AOI21_X1 U5620 ( .B1(n4474), .B2(n4476), .A(n4374), .ZN(n4472) );
  NAND2_X1 U5621 ( .A1(n5513), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5538) );
  INV_X1 U5622 ( .A(n5515), .ZN(n5513) );
  NAND2_X1 U5623 ( .A1(n4708), .A2(n9047), .ZN(n9489) );
  NAND2_X1 U5624 ( .A1(n9521), .A2(n9181), .ZN(n9503) );
  NAND2_X1 U5625 ( .A1(n9528), .A2(n9742), .ZN(n9529) );
  NAND2_X1 U5626 ( .A1(n9528), .A2(n4537), .ZN(n9510) );
  INV_X1 U5627 ( .A(n9238), .ZN(n9546) );
  AOI21_X1 U5628 ( .B1(n4692), .B2(n7675), .A(n4690), .ZN(n4689) );
  INV_X1 U5629 ( .A(n9037), .ZN(n4690) );
  NAND2_X1 U5630 ( .A1(n4756), .A2(n4372), .ZN(n4755) );
  NAND2_X1 U5631 ( .A1(n7568), .A2(n9166), .ZN(n7680) );
  NAND2_X1 U5632 ( .A1(n7680), .A2(n9109), .ZN(n9558) );
  OAI21_X1 U5633 ( .B1(n4324), .B2(n4697), .A(n9026), .ZN(n4696) );
  NAND2_X1 U5634 ( .A1(n7494), .A2(n9163), .ZN(n9582) );
  NAND2_X1 U5635 ( .A1(n7504), .A2(n4325), .ZN(n9595) );
  NAND2_X1 U5636 ( .A1(n7504), .A2(n9804), .ZN(n7491) );
  NAND2_X1 U5637 ( .A1(n7123), .A2(n6510), .ZN(n7225) );
  NOR2_X1 U5638 ( .A1(n7226), .A2(n9610), .ZN(n7270) );
  NAND2_X1 U5639 ( .A1(n4521), .A2(n4520), .ZN(n7226) );
  NAND2_X1 U5640 ( .A1(n7160), .A2(n4461), .ZN(n7125) );
  NAND2_X1 U5641 ( .A1(n4462), .A2(n7111), .ZN(n4461) );
  NOR2_X1 U5642 ( .A1(n6807), .A2(n8914), .ZN(n6903) );
  NAND2_X1 U5643 ( .A1(n6499), .A2(n9940), .ZN(n6500) );
  NAND2_X1 U5644 ( .A1(n4523), .A2(n4522), .ZN(n6807) );
  NAND2_X1 U5645 ( .A1(n5590), .A2(n5589), .ZN(n9436) );
  NAND2_X1 U5646 ( .A1(n5562), .A2(n5561), .ZN(n9645) );
  AOI211_X1 U5647 ( .C1(n9495), .C2(n9510), .A(n9548), .B(n4401), .ZN(n9661)
         );
  AND2_X1 U5648 ( .A1(n6572), .A2(n9194), .ZN(n9949) );
  NOR2_X1 U5649 ( .A1(n6751), .A2(n6576), .ZN(n6580) );
  XNOR2_X1 U5650 ( .A(n7726), .B(n7725), .ZN(n7713) );
  NAND2_X1 U5651 ( .A1(n5667), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5672) );
  NAND2_X1 U5652 ( .A1(n4813), .A2(n5504), .ZN(n5530) );
  AOI21_X1 U5653 ( .B1(n5103), .B2(n4791), .A(n4385), .ZN(n4790) );
  XNOR2_X1 U5654 ( .A(n5040), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6671) );
  NAND2_X1 U5655 ( .A1(n4996), .A2(n5821), .ZN(n4782) );
  INV_X1 U5656 ( .A(n4317), .ZN(n4701) );
  NAND2_X1 U5658 ( .A1(n8311), .A2(n8013), .ZN(n8030) );
  NAND2_X1 U5659 ( .A1(n6127), .A2(n8002), .ZN(n8045) );
  NAND2_X1 U5660 ( .A1(n8250), .A2(n8059), .ZN(n4684) );
  INV_X1 U5661 ( .A(n4653), .ZN(n8094) );
  NOR2_X1 U5662 ( .A1(n4656), .A2(n4661), .ZN(n4654) );
  INV_X1 U5663 ( .A(n6988), .ZN(n5866) );
  INV_X1 U5665 ( .A(n4674), .ZN(n8297) );
  NAND2_X1 U5666 ( .A1(n6060), .A2(n4906), .ZN(n8296) );
  INV_X1 U5667 ( .A(n10042), .ZN(n10080) );
  AND2_X1 U5668 ( .A1(n7153), .A2(n5899), .ZN(n4685) );
  NAND2_X1 U5669 ( .A1(n6178), .A2(n6177), .ZN(n8317) );
  AND2_X1 U5670 ( .A1(n6021), .A2(n6020), .ZN(n8333) );
  OR2_X1 U5671 ( .A1(n6195), .A2(n6313), .ZN(n8324) );
  NAND2_X1 U5672 ( .A1(n4658), .A2(n4657), .ZN(n8323) );
  NAND2_X1 U5673 ( .A1(n8323), .A2(n8322), .ZN(n8321) );
  AND2_X1 U5674 ( .A1(n6194), .A2(n6313), .ZN(n8329) );
  INV_X1 U5675 ( .A(n8500), .ZN(n8479) );
  INV_X1 U5676 ( .A(n8528), .ZN(n8553) );
  INV_X1 U5677 ( .A(n10038), .ZN(n8342) );
  NAND2_X1 U5678 ( .A1(n5839), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5840) );
  CLKBUF_X1 U5679 ( .A(n6206), .Z(n8348) );
  INV_X1 U5680 ( .A(P2_U3893), .ZN(n8347) );
  NAND2_X1 U5681 ( .A1(n6378), .A2(n6832), .ZN(n6836) );
  NAND2_X1 U5682 ( .A1(n4640), .A2(n4641), .ZN(n6951) );
  NOR2_X1 U5683 ( .A1(n4638), .A2(n4639), .ZN(n6351) );
  NOR2_X1 U5684 ( .A1(n6939), .A2(n6419), .ZN(n7067) );
  AOI21_X1 U5685 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n7069), .A(n4749), .ZN(
        n10023) );
  OAI211_X1 U5686 ( .C1(n4749), .C2(n7069), .A(n4743), .B(n4747), .ZN(n4748)
         );
  AND2_X1 U5687 ( .A1(n6384), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7313) );
  INV_X1 U5688 ( .A(n4635), .ZN(n7550) );
  NAND2_X1 U5689 ( .A1(n4731), .A2(n4732), .ZN(n7540) );
  NAND2_X1 U5690 ( .A1(n6385), .A2(n4734), .ZN(n4732) );
  NAND2_X1 U5691 ( .A1(n6384), .A2(n4733), .ZN(n4731) );
  INV_X1 U5692 ( .A(n4720), .ZN(n7604) );
  NOR2_X1 U5693 ( .A1(n7649), .A2(n6358), .ZN(n7594) );
  NOR2_X1 U5694 ( .A1(n7659), .A2(n8685), .ZN(n7658) );
  MUX2_X1 U5695 ( .A(n8432), .B(n8431), .S(n8430), .Z(n8434) );
  AND2_X1 U5696 ( .A1(n4650), .A2(n8423), .ZN(n4446) );
  INV_X1 U5697 ( .A(n6366), .ZN(n4650) );
  NAND2_X1 U5698 ( .A1(n4740), .A2(n4739), .ZN(n8420) );
  AND3_X1 U5699 ( .A1(n4740), .A2(n4739), .A3(n6395), .ZN(n6396) );
  INV_X1 U5700 ( .A(n4584), .ZN(n4583) );
  OAI21_X1 U5701 ( .B1(n6486), .B2(n6485), .A(n6481), .ZN(n4584) );
  AOI21_X1 U5702 ( .B1(n6315), .B2(n8627), .A(n6314), .ZN(n8460) );
  NAND2_X1 U5703 ( .A1(n4879), .A2(n6252), .ZN(n6483) );
  NAND2_X1 U5704 ( .A1(n6234), .A2(n6233), .ZN(n8483) );
  NAND2_X1 U5705 ( .A1(n6075), .A2(n6074), .ZN(n8566) );
  OAI21_X1 U5706 ( .B1(n8598), .B2(n4571), .A(n4570), .ZN(n8559) );
  OAI21_X1 U5707 ( .B1(n8598), .B2(n8597), .A(n4579), .ZN(n8587) );
  NAND2_X1 U5708 ( .A1(n6049), .A2(n6048), .ZN(n8674) );
  AND2_X1 U5709 ( .A1(n7471), .A2(n6287), .ZN(n4917) );
  NAND2_X1 U5710 ( .A1(n5981), .A2(n5980), .ZN(n8691) );
  NAND2_X1 U5711 ( .A1(n5972), .A2(n5971), .ZN(n7466) );
  NAND2_X1 U5712 ( .A1(n4553), .A2(n6271), .ZN(n7404) );
  NAND2_X1 U5713 ( .A1(n4895), .A2(n7768), .ZN(n7407) );
  OR2_X1 U5714 ( .A1(n5830), .A2(n6602), .ZN(n5846) );
  INV_X1 U5715 ( .A(n10053), .ZN(n6975) );
  NAND2_X1 U5716 ( .A1(n6968), .A2(n8630), .ZN(n10043) );
  NOR2_X2 U5717 ( .A1(n6321), .A2(n6327), .ZN(n8604) );
  AND2_X1 U5718 ( .A1(n7734), .A2(n7733), .ZN(n8637) );
  INV_X1 U5719 ( .A(n8656), .ZN(n8686) );
  AND2_X1 U5720 ( .A1(n10124), .A2(n10074), .ZN(n8687) );
  INV_X1 U5721 ( .A(n8637), .ZN(n8695) );
  NAND2_X1 U5722 ( .A1(n4788), .A2(n7715), .ZN(n8699) );
  NAND2_X1 U5723 ( .A1(n4566), .A2(n6303), .ZN(n8461) );
  INV_X1 U5724 ( .A(n8028), .ZN(n8708) );
  NAND2_X1 U5725 ( .A1(n6231), .A2(n6230), .ZN(n8717) );
  NAND2_X1 U5726 ( .A1(n8521), .A2(n6295), .ZN(n8512) );
  CLKBUF_X1 U5727 ( .A(n8509), .Z(n8510) );
  NAND2_X1 U5728 ( .A1(n4886), .A2(n4891), .ZN(n8520) );
  NAND2_X1 U5729 ( .A1(n8550), .A2(n4894), .ZN(n4886) );
  OAI21_X1 U5730 ( .B1(n8550), .B2(n6223), .A(n7847), .ZN(n8536) );
  NAND2_X1 U5731 ( .A1(n6085), .A2(n6084), .ZN(n8744) );
  NAND2_X1 U5732 ( .A1(n6063), .A2(n6062), .ZN(n8751) );
  NOR2_X1 U5733 ( .A1(n4572), .A2(n4574), .ZN(n8576) );
  NOR2_X1 U5734 ( .A1(n8598), .A2(n4576), .ZN(n4572) );
  NAND2_X1 U5735 ( .A1(n4883), .A2(n7835), .ZN(n8585) );
  NAND2_X1 U5736 ( .A1(n6034), .A2(n6033), .ZN(n8761) );
  INV_X1 U5737 ( .A(n8333), .ZN(n7998) );
  NAND2_X1 U5738 ( .A1(n4538), .A2(n4541), .ZN(n8609) );
  NAND2_X1 U5739 ( .A1(n7471), .A2(n4542), .ZN(n4538) );
  NAND2_X1 U5740 ( .A1(n5994), .A2(n5993), .ZN(n8773) );
  NAND2_X1 U5741 ( .A1(n4545), .A2(n4548), .ZN(n8621) );
  NAND2_X1 U5742 ( .A1(n4547), .A2(n4546), .ZN(n4545) );
  INV_X1 U5743 ( .A(n8766), .ZN(n8774) );
  OR2_X1 U5744 ( .A1(n10108), .A2(n10102), .ZN(n8766) );
  AND2_X1 U5745 ( .A1(n7638), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6693) );
  AND2_X1 U5746 ( .A1(n5802), .A2(n5798), .ZN(n4431) );
  INV_X1 U5747 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U5748 ( .A1(n5767), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5769) );
  INV_X1 U5749 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7688) );
  INV_X1 U5750 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8239) );
  INV_X1 U5751 ( .A(n7752), .ZN(n7749) );
  INV_X1 U5752 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7391) );
  INV_X1 U5753 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7294) );
  INV_X1 U5754 ( .A(n8393), .ZN(n7178) );
  INV_X1 U5755 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7031) );
  INV_X1 U5756 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6787) );
  INV_X1 U5757 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6732) );
  INV_X1 U5758 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6700) );
  INV_X1 U5759 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6696) );
  INV_X1 U5760 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6662) );
  INV_X1 U5761 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6657) );
  INV_X1 U5762 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6635) );
  AND3_X1 U5763 ( .A1(n4900), .A2(n6373), .A3(n5741), .ZN(n5900) );
  AND2_X1 U5764 ( .A1(n5887), .A2(n5877), .ZN(n4900) );
  INV_X1 U5765 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6622) );
  AND3_X1 U5766 ( .A1(n6373), .A2(n5741), .A3(n5877), .ZN(n5886) );
  CLKBUF_X1 U5767 ( .A(n9960), .Z(n4426) );
  NAND2_X1 U5768 ( .A1(n4956), .A2(n4955), .ZN(n5689) );
  NAND2_X1 U5769 ( .A1(n4859), .A2(n5173), .ZN(n8851) );
  NAND2_X1 U5770 ( .A1(n5004), .A2(n5628), .ZN(n5005) );
  INV_X1 U5771 ( .A(n5003), .ZN(n5004) );
  INV_X1 U5772 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8868) );
  AND2_X1 U5773 ( .A1(n5255), .A2(n5254), .ZN(n5256) );
  NAND2_X1 U5774 ( .A1(n8873), .A2(n8874), .ZN(n8872) );
  NAND2_X1 U5775 ( .A1(n8881), .A2(n5409), .ZN(n8890) );
  INV_X1 U5776 ( .A(n8850), .ZN(n4855) );
  NAND2_X1 U5777 ( .A1(n5457), .A2(n5456), .ZN(n9512) );
  NAND2_X1 U5778 ( .A1(n5527), .A2(n8825), .ZN(n8932) );
  INV_X1 U5779 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8942) );
  NAND2_X1 U5780 ( .A1(n4843), .A2(n4850), .ZN(n4842) );
  NOR2_X1 U5781 ( .A1(n7107), .A2(n7108), .ZN(n7106) );
  OAI21_X1 U5782 ( .B1(n8898), .B2(n4494), .A(n4490), .ZN(n8951) );
  NAND2_X1 U5783 ( .A1(n5614), .A2(n5613), .ZN(n9417) );
  NAND2_X1 U5784 ( .A1(n5715), .A2(n9920), .ZN(n8957) );
  AND2_X1 U5785 ( .A1(n4864), .A2(n4865), .ZN(n8962) );
  NAND2_X1 U5786 ( .A1(n9085), .A2(n9086), .ZN(n4630) );
  NOR2_X1 U5787 ( .A1(n4626), .A2(n9706), .ZN(n4625) );
  AND2_X1 U5788 ( .A1(n8978), .A2(n9203), .ZN(n9189) );
  INV_X1 U5789 ( .A(n9213), .ZN(n9190) );
  INV_X1 U5790 ( .A(n9322), .ZN(n4438) );
  NOR2_X1 U5791 ( .A1(n9850), .A2(n9322), .ZN(n9868) );
  NAND2_X1 U5792 ( .A1(n9876), .A2(n9875), .ZN(n9874) );
  INV_X1 U5793 ( .A(n9889), .ZN(n9883) );
  INV_X1 U5794 ( .A(n9343), .ZN(n9901) );
  AOI21_X1 U5795 ( .B1(n9346), .B2(n9880), .A(n4315), .ZN(n4449) );
  INV_X1 U5796 ( .A(n9345), .ZN(n4450) );
  NOR2_X1 U5797 ( .A1(n9352), .A2(n9548), .ZN(n9617) );
  NAND2_X1 U5798 ( .A1(n4528), .A2(n8978), .ZN(n4524) );
  INV_X1 U5799 ( .A(n4766), .ZN(n4765) );
  OR2_X1 U5800 ( .A1(n9396), .A2(n9395), .ZN(n9398) );
  NAND2_X1 U5801 ( .A1(n4473), .A2(n4477), .ZN(n9459) );
  NAND2_X1 U5802 ( .A1(n9487), .A2(n4347), .ZN(n4473) );
  OAI21_X1 U5803 ( .B1(n9487), .B2(n6525), .A(n4343), .ZN(n9476) );
  NAND2_X1 U5804 ( .A1(n5424), .A2(n5423), .ZN(n9677) );
  INV_X1 U5805 ( .A(n4760), .ZN(n7676) );
  AOI21_X1 U5806 ( .B1(n4763), .B2(n4321), .A(n6520), .ZN(n4760) );
  AND2_X1 U5807 ( .A1(n4763), .A2(n4327), .ZN(n7567) );
  NOR2_X1 U5808 ( .A1(n4699), .A2(n4698), .ZN(n7495) );
  INV_X1 U5809 ( .A(n9017), .ZN(n4698) );
  NAND2_X1 U5810 ( .A1(n7488), .A2(n9106), .ZN(n7487) );
  NAND2_X1 U5811 ( .A1(n7420), .A2(n6517), .ZN(n7488) );
  NAND2_X1 U5812 ( .A1(n7503), .A2(n7506), .ZN(n7502) );
  NAND2_X1 U5813 ( .A1(n7262), .A2(n6515), .ZN(n7503) );
  OAI21_X1 U5814 ( .B1(n6902), .B2(n4754), .A(n4752), .ZN(n7052) );
  NAND2_X1 U5815 ( .A1(n6901), .A2(n6507), .ZN(n7053) );
  OR2_X1 U5816 ( .A1(n9934), .A2(n9347), .ZN(n9928) );
  NOR2_X1 U5817 ( .A1(n9934), .A2(n6754), .ZN(n9925) );
  NAND2_X1 U5818 ( .A1(n9957), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n4705) );
  OR2_X1 U5819 ( .A1(n9627), .A2(n9953), .ZN(n4707) );
  NAND2_X1 U5820 ( .A1(n5267), .A2(n5266), .ZN(n7434) );
  NAND2_X1 U5821 ( .A1(n5239), .A2(n5238), .ZN(n7301) );
  INV_X1 U5822 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n4482) );
  NAND2_X1 U5823 ( .A1(n9710), .A2(n9946), .ZN(n4483) );
  INV_X1 U5824 ( .A(n9402), .ZN(n9715) );
  INV_X1 U5825 ( .A(n9417), .ZN(n9719) );
  INV_X1 U5826 ( .A(n9436), .ZN(n9723) );
  INV_X1 U5827 ( .A(n9512), .ZN(n9738) );
  INV_X1 U5828 ( .A(n7434), .ZN(n9804) );
  AND2_X1 U5829 ( .A1(n4978), .A2(n4517), .ZN(n4702) );
  NAND2_X1 U5830 ( .A1(n9946), .A2(n9949), .ZN(n9747) );
  INV_X1 U5831 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4934) );
  INV_X1 U5832 ( .A(n4939), .ZN(n7695) );
  XNOR2_X1 U5833 ( .A(n6459), .B(n6458), .ZN(n8791) );
  NAND2_X1 U5834 ( .A1(n4800), .A2(n5697), .ZN(n6459) );
  XNOR2_X1 U5835 ( .A(n5696), .B(n5695), .ZN(n9762) );
  NOR2_X1 U5836 ( .A1(n4444), .A2(n4443), .ZN(n4442) );
  NOR2_X1 U5837 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4443) );
  NAND2_X1 U5838 ( .A1(n4932), .A2(n5418), .ZN(n4961) );
  NAND2_X1 U5839 ( .A1(n4812), .A2(n5528), .ZN(n5555) );
  NAND2_X1 U5840 ( .A1(n4813), .A2(n4807), .ZN(n4812) );
  INV_X1 U5841 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7711) );
  XNOR2_X1 U5842 ( .A(n4945), .B(n4955), .ZN(n7709) );
  INV_X1 U5843 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8221) );
  OR2_X1 U5844 ( .A1(n4947), .A2(n4946), .ZN(n4948) );
  INV_X1 U5845 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7393) );
  XNOR2_X1 U5846 ( .A(n5285), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9831) );
  INV_X1 U5847 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6814) );
  AND2_X1 U5848 ( .A1(n5135), .A2(n5134), .ZN(n9792) );
  NAND2_X1 U5849 ( .A1(n4792), .A2(n5088), .ZN(n5104) );
  XNOR2_X1 U5850 ( .A(n4782), .B(n5017), .ZN(n6596) );
  OAI21_X1 U5851 ( .B1(n6169), .B2(n6168), .A(n8320), .ZN(n6201) );
  NOR2_X1 U5852 ( .A1(n4786), .A2(n4419), .ZN(n7984) );
  INV_X1 U5853 ( .A(n4737), .ZN(n8352) );
  AOI21_X1 U5854 ( .B1(n4387), .B2(n6928), .A(n4434), .ZN(n8418) );
  NOR2_X1 U5855 ( .A1(n4904), .A2(n5733), .ZN(n5739) );
  OR2_X1 U5856 ( .A1(n8807), .A2(n5737), .ZN(n5738) );
  OR2_X1 U5857 ( .A1(n6583), .A2(n9685), .ZN(n4902) );
  NAND2_X1 U5858 ( .A1(n4706), .A2(n4703), .ZN(P1_U3550) );
  INV_X1 U5859 ( .A(n4704), .ZN(n4703) );
  NAND2_X1 U5860 ( .A1(n9710), .A2(n9959), .ZN(n4706) );
  OAI21_X1 U5861 ( .B1(n9711), .B2(n9685), .A(n4705), .ZN(n4704) );
  NOR2_X1 U5862 ( .A1(n4459), .A2(n4402), .ZN(n4458) );
  NOR2_X1 U5863 ( .A1(n9946), .A2(n6582), .ZN(n4459) );
  AND2_X2 U5864 ( .A1(n4965), .A2(n6538), .ZN(n4987) );
  AND2_X1 U5865 ( .A1(n4327), .A2(n6519), .ZN(n4321) );
  OR2_X1 U5866 ( .A1(n8623), .A2(n8682), .ZN(n4322) );
  AND2_X1 U5867 ( .A1(n7864), .A2(n7869), .ZN(n8539) );
  INV_X1 U5868 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8784) );
  AND2_X1 U5869 ( .A1(n5145), .A2(n7200), .ZN(n4323) );
  NAND2_X1 U5870 ( .A1(n4548), .A2(n4544), .ZN(n4543) );
  AND2_X1 U5871 ( .A1(n9804), .A2(n4531), .ZN(n4325) );
  AND2_X1 U5872 ( .A1(n4631), .A2(n6827), .ZN(n4326) );
  AND2_X1 U5873 ( .A1(n8695), .A2(n7914), .ZN(n7966) );
  NAND2_X1 U5874 ( .A1(n9599), .A2(n8966), .ZN(n4327) );
  AND2_X1 U5875 ( .A1(n4530), .A2(n4529), .ZN(n4328) );
  OR2_X1 U5876 ( .A1(n9484), .A2(n9236), .ZN(n4329) );
  AND2_X1 U5877 ( .A1(n4310), .A2(n10124), .ZN(n4330) );
  INV_X1 U5878 ( .A(n6290), .ZN(n4546) );
  NAND2_X1 U5879 ( .A1(n6373), .A2(n5741), .ZN(n5862) );
  INV_X1 U5880 ( .A(n7541), .ZN(n4734) );
  AND2_X1 U5881 ( .A1(n4939), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4331) );
  AND2_X1 U5882 ( .A1(n4325), .A2(n9599), .ZN(n4332) );
  OR2_X1 U5883 ( .A1(n7967), .A2(n4314), .ZN(n4333) );
  INV_X1 U5884 ( .A(n9484), .ZN(n9731) );
  INV_X1 U5885 ( .A(n9462), .ZN(n4480) );
  XNOR2_X1 U5886 ( .A(n6446), .B(n6396), .ZN(n4334) );
  INV_X1 U5887 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5748) );
  NAND2_X1 U5888 ( .A1(n4880), .A2(n4391), .ZN(n4335) );
  AND2_X1 U5889 ( .A1(n4603), .A2(n4598), .ZN(n4336) );
  NAND2_X1 U5890 ( .A1(n6125), .A2(n6122), .ZN(n4337) );
  AND2_X1 U5891 ( .A1(n4865), .A2(n8961), .ZN(n4338) );
  INV_X1 U5892 ( .A(n9097), .ZN(n4621) );
  AND2_X1 U5893 ( .A1(n5556), .A2(n5535), .ZN(n5554) );
  OR2_X1 U5894 ( .A1(n9959), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n4339) );
  OR2_X1 U5895 ( .A1(n9126), .A2(n4315), .ZN(n4340) );
  OR2_X1 U5896 ( .A1(n8412), .A2(n6394), .ZN(n4341) );
  AND3_X1 U5897 ( .A1(n4941), .A2(n4852), .A3(n4943), .ZN(n4342) );
  XNOR2_X1 U5898 ( .A(n5766), .B(n5765), .ZN(n5775) );
  OR2_X1 U5899 ( .A1(n9495), .A2(n9237), .ZN(n4343) );
  NAND2_X1 U5900 ( .A1(n8882), .A2(n8883), .ZN(n8881) );
  INV_X1 U5901 ( .A(n6268), .ZN(n6209) );
  AND2_X1 U5902 ( .A1(n9261), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4344) );
  INV_X1 U5903 ( .A(n7496), .ZN(n9106) );
  AND2_X1 U5904 ( .A1(n9025), .A2(n9163), .ZN(n7496) );
  NOR2_X1 U5905 ( .A1(n8344), .A2(n7084), .ZN(n4345) );
  AND2_X1 U5906 ( .A1(n4329), .A2(n4343), .ZN(n4347) );
  AND2_X1 U5907 ( .A1(n8682), .A2(n8623), .ZN(n4348) );
  INV_X1 U5908 ( .A(n9488), .ZN(n4711) );
  OR2_X1 U5909 ( .A1(n7671), .A2(n6389), .ZN(n4349) );
  NAND2_X1 U5910 ( .A1(n7201), .A2(n5146), .ZN(n4350) );
  AND2_X1 U5911 ( .A1(n6660), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4351) );
  INV_X1 U5912 ( .A(n8857), .ZN(n4520) );
  AND3_X1 U5913 ( .A1(n4991), .A2(n4990), .A3(n4989), .ZN(n4352) );
  OR2_X1 U5914 ( .A1(n5772), .A2(n5771), .ZN(n4353) );
  OR2_X1 U5915 ( .A1(n6350), .A2(n6620), .ZN(n4354) );
  INV_X1 U5916 ( .A(n9181), .ZN(n4710) );
  INV_X1 U5917 ( .A(n9163), .ZN(n4697) );
  OR2_X1 U5918 ( .A1(n6296), .A2(n8336), .ZN(n4355) );
  INV_X1 U5919 ( .A(n9382), .ZN(n4469) );
  NAND2_X1 U5920 ( .A1(n5442), .A2(n5441), .ZN(n9531) );
  NAND2_X2 U5921 ( .A1(n4982), .A2(n4965), .ZN(n4985) );
  AND2_X1 U5922 ( .A1(n8838), .A2(n8941), .ZN(n4356) );
  NAND2_X1 U5923 ( .A1(n5318), .A2(n5317), .ZN(n9691) );
  INV_X1 U5924 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4937) );
  AND2_X1 U5925 ( .A1(n9383), .A2(n4328), .ZN(n4357) );
  OR2_X1 U5926 ( .A1(n7869), .A2(n7894), .ZN(n4358) );
  AND3_X1 U5927 ( .A1(n7902), .A2(n7901), .A3(n8335), .ZN(n4359) );
  XNOR2_X1 U5928 ( .A(n8028), .B(n8478), .ZN(n8469) );
  OAI21_X1 U5929 ( .B1(n6142), .B2(n7968), .A(n5796), .ZN(n5797) );
  INV_X1 U5930 ( .A(n8523), .ZN(n4561) );
  AND2_X1 U5931 ( .A1(n6671), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4360) );
  AND2_X1 U5932 ( .A1(n4684), .A2(n4683), .ZN(n4361) );
  XNOR2_X1 U5933 ( .A(n5844), .B(n7323), .ZN(n5836) );
  AND2_X1 U5934 ( .A1(n5103), .A2(n5084), .ZN(n4362) );
  NAND2_X1 U5935 ( .A1(n5778), .A2(n5748), .ZN(n6156) );
  AND2_X1 U5936 ( .A1(n4642), .A2(n7072), .ZN(n4363) );
  NOR2_X1 U5937 ( .A1(n7658), .A2(n6361), .ZN(n4364) );
  AND2_X1 U5938 ( .A1(n4874), .A2(n7903), .ZN(n4365) );
  INV_X1 U5939 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9756) );
  INV_X1 U5940 ( .A(n4580), .ZN(n4579) );
  NOR2_X1 U5941 ( .A1(n8099), .A2(n8589), .ZN(n4580) );
  INV_X1 U5942 ( .A(n9387), .ZN(n9711) );
  NAND2_X1 U5943 ( .A1(n5699), .A2(n5698), .ZN(n9387) );
  AND2_X1 U5944 ( .A1(n4711), .A2(n9047), .ZN(n4366) );
  AND2_X1 U5945 ( .A1(n5008), .A2(n5009), .ZN(n4367) );
  AND2_X1 U5946 ( .A1(n4561), .A2(n4358), .ZN(n4368) );
  AND2_X1 U5947 ( .A1(n5885), .A2(n5870), .ZN(n4369) );
  AND2_X1 U5948 ( .A1(n6383), .A2(n6427), .ZN(n4370) );
  INV_X1 U5949 ( .A(n4869), .ZN(n4868) );
  OAI21_X1 U5950 ( .B1(n8838), .B2(n8941), .A(n5413), .ZN(n4869) );
  NAND2_X1 U5951 ( .A1(n9687), .A2(n9562), .ZN(n4371) );
  NAND2_X1 U5952 ( .A1(n4321), .A2(n7675), .ZN(n4372) );
  INV_X1 U5953 ( .A(n4491), .ZN(n4490) );
  NAND2_X1 U5954 ( .A1(n5634), .A2(n4492), .ZN(n4491) );
  NOR2_X1 U5955 ( .A1(n9697), .A2(n9242), .ZN(n4373) );
  NOR2_X1 U5956 ( .A1(n4480), .A2(n6556), .ZN(n4374) );
  NAND2_X1 U5957 ( .A1(n6633), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4375) );
  AND2_X1 U5958 ( .A1(n9076), .A2(n4628), .ZN(n4376) );
  NAND2_X1 U5959 ( .A1(n6526), .A2(n4478), .ZN(n4377) );
  OR2_X1 U5960 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4378) );
  NOR2_X1 U5961 ( .A1(n7632), .A2(n9244), .ZN(n4379) );
  XNOR2_X1 U5962 ( .A(n7701), .B(SI_29_), .ZN(n6533) );
  NOR2_X1 U5963 ( .A1(n9711), .A2(n6569), .ZN(n4380) );
  OR2_X1 U5964 ( .A1(n6288), .A2(n6289), .ZN(n4381) );
  AND2_X1 U5965 ( .A1(n6508), .A2(n7205), .ZN(n4382) );
  AND2_X1 U5966 ( .A1(n6470), .A2(n6469), .ZN(n4383) );
  INV_X1 U5967 ( .A(n4535), .ZN(n4534) );
  NAND2_X1 U5968 ( .A1(n4537), .A2(n4536), .ZN(n4535) );
  INV_X1 U5969 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5690) );
  INV_X1 U5970 ( .A(n4661), .ZN(n4659) );
  NAND2_X1 U5971 ( .A1(n4665), .A2(n8261), .ZN(n4661) );
  INV_X1 U5972 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4967) );
  NAND2_X1 U5973 ( .A1(n8566), .A2(n8577), .ZN(n4384) );
  AND2_X1 U5974 ( .A1(n5106), .A2(SI_5_), .ZN(n4385) );
  AND2_X1 U5975 ( .A1(n5282), .A2(SI_12_), .ZN(n4386) );
  INV_X1 U5976 ( .A(n4836), .ZN(n4835) );
  NAND2_X1 U5977 ( .A1(n4838), .A2(n5280), .ZN(n4836) );
  NAND2_X1 U5978 ( .A1(n4741), .A2(n4457), .ZN(n4387) );
  OR2_X1 U5979 ( .A1(n8839), .A2(n4356), .ZN(n4388) );
  NOR3_X1 U5980 ( .A1(n9382), .A2(n9399), .A3(n9118), .ZN(n4389) );
  NOR2_X1 U5981 ( .A1(n7849), .A2(n8590), .ZN(n4390) );
  INV_X1 U5982 ( .A(n4603), .ZN(n4599) );
  AND2_X1 U5983 ( .A1(n9466), .A2(n9478), .ZN(n4603) );
  OR2_X1 U5984 ( .A1(n8458), .A2(n8463), .ZN(n4391) );
  INV_X1 U5985 ( .A(n7958), .ZN(n6484) );
  AND2_X1 U5986 ( .A1(n7903), .A2(n7901), .ZN(n7958) );
  AND2_X1 U5987 ( .A1(n4560), .A2(n6297), .ZN(n4392) );
  AND2_X1 U5988 ( .A1(n4979), .A2(n4702), .ZN(n9145) );
  INV_X1 U5989 ( .A(n9145), .ZN(n4617) );
  AND2_X1 U5990 ( .A1(n7768), .A2(n6211), .ZN(n4393) );
  AOI21_X1 U5991 ( .B1(n9106), .B2(n4467), .A(n4373), .ZN(n4466) );
  AND2_X1 U5992 ( .A1(n6304), .A2(n6303), .ZN(n4394) );
  AND2_X1 U5993 ( .A1(n7214), .A2(n5914), .ZN(n4395) );
  INV_X1 U5994 ( .A(n4820), .ZN(n4819) );
  OAI21_X1 U5995 ( .B1(n5358), .B2(n4821), .A(n5357), .ZN(n4820) );
  INV_X1 U5996 ( .A(n4682), .ZN(n4681) );
  OAI21_X1 U5997 ( .B1(n8275), .B2(n4683), .A(n8274), .ZN(n4682) );
  AND2_X1 U5998 ( .A1(n5958), .A2(n5946), .ZN(n4396) );
  INV_X1 U5999 ( .A(n4501), .ZN(n4500) );
  NOR2_X1 U6000 ( .A1(n4869), .A2(n4502), .ZN(n4501) );
  AND2_X1 U6001 ( .A1(n4741), .A2(n4341), .ZN(n4397) );
  AND2_X1 U6002 ( .A1(n6221), .A2(n7835), .ZN(n4398) );
  AND2_X1 U6003 ( .A1(n4556), .A2(n4563), .ZN(n4399) );
  OAI21_X1 U6004 ( .B1(n4657), .B2(n4656), .A(n6030), .ZN(n4655) );
  INV_X1 U6005 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4933) );
  AND2_X1 U6006 ( .A1(n8977), .A2(n8976), .ZN(n9706) );
  INV_X1 U6007 ( .A(n8981), .ZN(n8974) );
  NAND2_X1 U6008 ( .A1(n5340), .A2(n5339), .ZN(n8981) );
  AND3_X1 U6009 ( .A1(n7970), .A2(n4333), .A3(n4912), .ZN(n4400) );
  INV_X1 U6010 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4873) );
  INV_X1 U6011 ( .A(n6620), .ZN(n4727) );
  NAND2_X1 U6012 ( .A1(n9588), .A2(n6518), .ZN(n4763) );
  NAND2_X1 U6013 ( .A1(n9082), .A2(n9081), .ZN(n9620) );
  INV_X1 U6014 ( .A(n9620), .ZN(n4529) );
  INV_X1 U6015 ( .A(n8623), .ZN(n8266) );
  AND2_X1 U6016 ( .A1(n9528), .A2(n4534), .ZN(n4401) );
  NOR2_X1 U6017 ( .A1(n5434), .A2(n4832), .ZN(n4831) );
  AND4_X1 U6018 ( .A1(n6027), .A2(n6026), .A3(n6025), .A4(n6024), .ZN(n8613)
         );
  INV_X1 U6019 ( .A(n7554), .ZN(n6701) );
  INV_X1 U6020 ( .A(n9091), .ZN(n4778) );
  INV_X1 U6021 ( .A(n9166), .ZN(n4694) );
  OAI21_X1 U6022 ( .B1(n7987), .B2(n7824), .A(n7826), .ZN(n8596) );
  NAND2_X1 U6023 ( .A1(n4885), .A2(n6218), .ZN(n8608) );
  INV_X1 U6024 ( .A(n8874), .ZN(n4494) );
  INV_X1 U6025 ( .A(n9445), .ZN(n4602) );
  XNOR2_X1 U6026 ( .A(n5769), .B(n5768), .ZN(n6144) );
  NAND2_X1 U6027 ( .A1(n7522), .A2(n5974), .ZN(n8289) );
  NOR2_X1 U6028 ( .A1(n9571), .A2(n9677), .ZN(n9528) );
  INV_X1 U6029 ( .A(n8933), .ZN(n4863) );
  NAND2_X1 U6030 ( .A1(n4671), .A2(n6158), .ZN(n6143) );
  NOR2_X1 U6031 ( .A1(n6583), .A2(n9747), .ZN(n4402) );
  INV_X1 U6032 ( .A(n4680), .ZN(n4679) );
  OR2_X1 U6033 ( .A1(n8275), .A2(n6100), .ZN(n4680) );
  INV_X1 U6034 ( .A(n4543), .ZN(n4542) );
  INV_X1 U6035 ( .A(n4775), .ZN(n4771) );
  NAND2_X1 U6036 ( .A1(n9417), .A2(n9234), .ZN(n4775) );
  AND2_X1 U6037 ( .A1(n5433), .A2(SI_18_), .ZN(n4403) );
  AND2_X1 U6038 ( .A1(n4664), .A2(n4663), .ZN(n4404) );
  AND2_X1 U6039 ( .A1(n5554), .A2(n4807), .ZN(n4405) );
  AND2_X1 U6040 ( .A1(n8014), .A2(n8013), .ZN(n4406) );
  INV_X1 U6041 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U6042 ( .A1(n5486), .A2(n5485), .ZN(n9495) );
  INV_X1 U6043 ( .A(n9495), .ZN(n4536) );
  AND2_X2 U6044 ( .A1(n6962), .A2(n6323), .ZN(n10124) );
  NAND2_X1 U6045 ( .A1(n5287), .A2(n5286), .ZN(n9697) );
  INV_X1 U6046 ( .A(n9697), .ZN(n4531) );
  NAND2_X1 U6047 ( .A1(n6986), .A2(n4369), .ZN(n7011) );
  AND4_X1 U6048 ( .A1(n6042), .A2(n6041), .A3(n6040), .A4(n6039), .ZN(n8589)
         );
  OAI21_X1 U6049 ( .B1(n7369), .B2(n6281), .A(n6280), .ZN(n7357) );
  OAI21_X1 U6050 ( .B1(n7475), .B2(n6215), .A(n7803), .ZN(n7533) );
  NOR2_X1 U6051 ( .A1(n7106), .A2(n5123), .ZN(n4407) );
  AND2_X1 U6052 ( .A1(n4855), .A2(n5173), .ZN(n4408) );
  OR2_X1 U6053 ( .A1(n9946), .A2(n4482), .ZN(n4409) );
  INV_X1 U6054 ( .A(n7471), .ZN(n4547) );
  NAND2_X1 U6055 ( .A1(n7279), .A2(n5946), .ZN(n7447) );
  AND2_X1 U6056 ( .A1(n7152), .A2(n5914), .ZN(n7211) );
  NOR2_X1 U6057 ( .A1(n7313), .A2(n6385), .ZN(n4410) );
  INV_X1 U6058 ( .A(n4521), .ZN(n7168) );
  NOR2_X1 U6059 ( .A1(n7169), .A2(n7208), .ZN(n4521) );
  NAND2_X1 U6060 ( .A1(n7504), .A2(n4332), .ZN(n4532) );
  NAND2_X1 U6061 ( .A1(n5772), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U6062 ( .A1(n8909), .A2(n4851), .ZN(n4411) );
  AND2_X1 U6063 ( .A1(n6461), .A2(n6460), .ZN(n4412) );
  INV_X1 U6064 ( .A(n7655), .ZN(n6730) );
  AND2_X1 U6065 ( .A1(n5977), .A2(n5761), .ZN(n7655) );
  AND2_X1 U6066 ( .A1(n7078), .A2(n5899), .ZN(n4413) );
  INV_X1 U6067 ( .A(n9125), .ZN(n4628) );
  AND2_X2 U6068 ( .A1(n6580), .A2(n6579), .ZN(n9959) );
  OR2_X1 U6069 ( .A1(n4966), .A2(n4315), .ZN(n6843) );
  NAND2_X1 U6070 ( .A1(n6891), .A2(n7978), .ZN(n10024) );
  INV_X1 U6071 ( .A(n7208), .ZN(n4462) );
  NAND2_X1 U6072 ( .A1(n6986), .A2(n5870), .ZN(n7010) );
  INV_X1 U6073 ( .A(n9119), .ZN(n4627) );
  NAND2_X1 U6074 ( .A1(n9940), .A2(n7098), .ZN(n7097) );
  INV_X1 U6075 ( .A(n7097), .ZN(n4522) );
  OR2_X1 U6076 ( .A1(n8421), .A2(n8592), .ZN(n4414) );
  INV_X1 U6077 ( .A(n6861), .ZN(n4717) );
  NAND2_X1 U6078 ( .A1(n6346), .A2(n6861), .ZN(n6826) );
  INV_X1 U6079 ( .A(n6826), .ZN(n4632) );
  INV_X1 U6080 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n4643) );
  AOI21_X1 U6081 ( .B1(n10011), .B2(n8412), .A(n4437), .ZN(n4436) );
  XNOR2_X1 U6082 ( .A(n6394), .B(n8412), .ZN(n8408) );
  NAND2_X1 U6083 ( .A1(n9990), .A2(n6376), .ZN(n6377) );
  NOR2_X1 U6084 ( .A1(n7641), .A2(n6387), .ZN(n7606) );
  NOR2_X1 U6085 ( .A1(n6392), .A2(n8368), .ZN(n8389) );
  NOR2_X1 U6086 ( .A1(n8350), .A2(n4735), .ZN(n6391) );
  NAND2_X1 U6087 ( .A1(n9888), .A2(n9339), .ZN(n9341) );
  NOR2_X1 U6088 ( .A1(n5344), .A2(n9854), .ZN(n9853) );
  NAND2_X1 U6089 ( .A1(n9348), .A2(n4315), .ZN(n4451) );
  NOR2_X1 U6090 ( .A1(n9863), .A2(n9862), .ZN(n9861) );
  AOI21_X1 U6091 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9831), .A(n9826), .ZN(
        n9837) );
  AOI21_X1 U6092 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9780), .A(n9772), .ZN(
        n9813) );
  AOI21_X1 U6093 ( .B1(n9843), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9835), .ZN(
        n9334) );
  AOI21_X1 U6094 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6739), .A(n6738), .ZN(
        n9786) );
  AOI21_X1 U6095 ( .B1(n6798), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6797), .ZN(
        n6801) );
  NAND2_X1 U6096 ( .A1(n8982), .A2(n9149), .ZN(n6764) );
  OAI21_X2 U6097 ( .B1(n7117), .B2(n9101), .A(n6550), .ZN(n7266) );
  NOR2_X1 U6098 ( .A1(n9395), .A2(n9377), .ZN(n4700) );
  NAND2_X1 U6099 ( .A1(n6766), .A2(n8982), .ZN(n6810) );
  NAND3_X1 U6100 ( .A1(n4707), .A2(n9625), .A3(n9626), .ZN(n9710) );
  AOI21_X1 U6101 ( .B1(n8429), .B2(P2_U3893), .A(n10011), .ZN(n8431) );
  NOR2_X1 U6102 ( .A1(n7306), .A2(n7305), .ZN(n7304) );
  OAI21_X1 U6103 ( .B1(n7595), .B2(n7599), .A(n7597), .ZN(n7662) );
  AOI21_X1 U6104 ( .B1(n6412), .B2(n6841), .A(n6821), .ZN(n6934) );
  NAND2_X1 U6105 ( .A1(n8414), .A2(n8415), .ZN(n8413) );
  NAND2_X1 U6106 ( .A1(n8372), .A2(n8373), .ZN(n8371) );
  NAND2_X1 U6107 ( .A1(n4417), .A2(n4416), .ZN(P2_U3200) );
  INV_X1 U6108 ( .A(n8435), .ZN(n4416) );
  NOR2_X1 U6109 ( .A1(n8437), .A2(n10024), .ZN(n4418) );
  NOR2_X1 U6110 ( .A1(n6434), .A2(n7644), .ZN(n7599) );
  NOR3_X1 U6111 ( .A1(n6872), .A2(n6823), .A3(n6822), .ZN(n6821) );
  NAND3_X1 U6112 ( .A1(n5747), .A2(n4688), .A3(n5746), .ZN(n5772) );
  NAND3_X1 U6113 ( .A1(n4783), .A2(n7921), .A3(n4400), .ZN(n4419) );
  NAND2_X2 U6114 ( .A1(n6232), .A2(n7878), .ZN(n8475) );
  NAND2_X1 U6115 ( .A1(n5750), .A2(n5749), .ZN(n5751) );
  OAI21_X2 U6116 ( .B1(n6863), .B2(n4632), .A(n4326), .ZN(n6828) );
  OAI211_X1 U6117 ( .C1(n6371), .C2(n9967), .A(n4422), .B(n6457), .ZN(P2_U3201) );
  NAND2_X1 U6118 ( .A1(n4334), .A2(n6928), .ZN(n4422) );
  NOR2_X2 U6119 ( .A1(n6364), .A2(n8378), .ZN(n8399) );
  OAI21_X1 U6120 ( .B1(n7659), .B2(n4645), .A(n4644), .ZN(n8360) );
  XNOR2_X1 U6121 ( .A(n6363), .B(n8374), .ZN(n8379) );
  NOR2_X1 U6122 ( .A1(n7548), .A2(n4633), .ZN(n6357) );
  NOR2_X1 U6123 ( .A1(n7594), .A2(n7593), .ZN(n7592) );
  NOR2_X1 U6124 ( .A1(n7650), .A2(n7651), .ZN(n7649) );
  INV_X1 U6125 ( .A(n9969), .ZN(n4425) );
  NOR3_X2 U6126 ( .A1(n9395), .A2(n9377), .A3(n9382), .ZN(n6562) );
  NAND2_X1 U6127 ( .A1(n6581), .A2(n9959), .ZN(n4432) );
  NAND2_X1 U6128 ( .A1(n4432), .A2(n4339), .ZN(n6578) );
  OAI21_X1 U6129 ( .B1(n7881), .B2(n6300), .A(n7880), .ZN(n7884) );
  NAND2_X1 U6130 ( .A1(n4455), .A2(n7870), .ZN(n7875) );
  NAND2_X1 U6131 ( .A1(n4428), .A2(n4427), .ZN(n7795) );
  NAND3_X1 U6132 ( .A1(n7789), .A2(n7788), .A3(n7934), .ZN(n4428) );
  NAND2_X1 U6133 ( .A1(n7916), .A2(n7915), .ZN(n7920) );
  MUX2_X1 U6134 ( .A(n7797), .B(n7796), .S(n7910), .Z(n7806) );
  NAND3_X1 U6135 ( .A1(n4898), .A2(n5777), .A3(n4431), .ZN(n4581) );
  NAND2_X1 U6136 ( .A1(n4785), .A2(n4784), .ZN(n4783) );
  NAND2_X1 U6137 ( .A1(n5069), .A2(n5068), .ZN(n5085) );
  NAND2_X1 U6138 ( .A1(n5021), .A2(n5020), .ZN(n5042) );
  NAND2_X1 U6139 ( .A1(n7907), .A2(n7906), .ZN(n7909) );
  OAI21_X1 U6140 ( .B1(n7904), .B2(n8458), .A(n4453), .ZN(n7905) );
  NOR2_X2 U6141 ( .A1(n6574), .A2(n4433), .ZN(n6581) );
  NAND2_X1 U6142 ( .A1(n6826), .A2(n5853), .ZN(n4631) );
  NAND2_X1 U6143 ( .A1(n7068), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10008) );
  NAND2_X1 U6144 ( .A1(n6361), .A2(n4646), .ZN(n4644) );
  XNOR2_X1 U6145 ( .A(n6357), .B(n7655), .ZN(n7650) );
  AOI21_X1 U6146 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n7178), .A(n8397), .ZN(
        n6365) );
  NOR2_X1 U6147 ( .A1(n9284), .A2(n9283), .ZN(n9282) );
  AOI21_X1 U6148 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(n9278), .A(n9282), .ZN(
        n6648) );
  NAND2_X1 U6149 ( .A1(n4450), .A2(n4449), .ZN(n4448) );
  NAND2_X1 U6150 ( .A1(n4451), .A2(n4448), .ZN(n9350) );
  NAND2_X2 U6151 ( .A1(n7091), .A2(n9148), .ZN(n6545) );
  NAND2_X1 U6152 ( .A1(n4456), .A2(n9097), .ZN(n7117) );
  OR2_X1 U6153 ( .A1(n9253), .A2(n9940), .ZN(n6544) );
  INV_X1 U6154 ( .A(n7055), .ZN(n4456) );
  INV_X1 U6155 ( .A(n4696), .ZN(n4695) );
  AOI21_X1 U6156 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n7178), .A(n8387), .ZN(
        n6394) );
  NAND2_X1 U6157 ( .A1(n4639), .A2(n7072), .ZN(n4637) );
  AOI21_X1 U6158 ( .B1(n4651), .B2(n4446), .A(n8422), .ZN(n8424) );
  NOR2_X1 U6159 ( .A1(n6354), .A2(n6427), .ZN(n6356) );
  NAND2_X2 U6160 ( .A1(n9446), .A2(n6559), .ZN(n9426) );
  AND3_X2 U6161 ( .A1(n4903), .A2(n5745), .A3(n4452), .ZN(n5746) );
  NAND2_X1 U6162 ( .A1(n4883), .A2(n4398), .ZN(n8571) );
  INV_X1 U6163 ( .A(n6377), .ZN(n4718) );
  NAND2_X1 U6164 ( .A1(n7909), .A2(n7959), .ZN(n7911) );
  INV_X1 U6165 ( .A(n7920), .ZN(n4785) );
  MUX2_X1 U6166 ( .A(n7877), .B(n7876), .S(n7910), .Z(n7881) );
  NOR2_X1 U6167 ( .A1(n4359), .A2(n4454), .ZN(n4453) );
  AOI21_X2 U6168 ( .B1(n9409), .B2(n9413), .A(n9197), .ZN(n9394) );
  OR2_X2 U6169 ( .A1(n9541), .A2(n9542), .ZN(n9539) );
  NAND2_X1 U6170 ( .A1(n6547), .A2(n8990), .ZN(n7055) );
  NAND2_X1 U6171 ( .A1(n6555), .A2(n9057), .ZN(n9465) );
  NOR2_X1 U6172 ( .A1(n7642), .A2(n7643), .ZN(n7641) );
  NAND2_X1 U6173 ( .A1(n8596), .A2(n7827), .ZN(n4883) );
  NAND2_X1 U6174 ( .A1(n8631), .A2(n6217), .ZN(n4885) );
  XNOR2_X1 U6175 ( .A(n5752), .B(n5798), .ZN(n6180) );
  NAND2_X1 U6176 ( .A1(n4310), .A2(n4582), .ZN(n6493) );
  NOR2_X2 U6177 ( .A1(n5771), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n5749) );
  AND3_X2 U6178 ( .A1(n5825), .A2(n5826), .A3(n5831), .ZN(n7323) );
  NAND2_X1 U6179 ( .A1(n4460), .A2(n4458), .ZN(P1_U3519) );
  OR2_X1 U6180 ( .A1(n6581), .A2(n9955), .ZN(n4460) );
  NAND2_X1 U6181 ( .A1(n9109), .A2(n4694), .ZN(n4693) );
  NAND2_X1 U6182 ( .A1(n4691), .A2(n4689), .ZN(n9541) );
  NAND2_X1 U6183 ( .A1(n7125), .A2(n7124), .ZN(n7123) );
  NAND2_X1 U6184 ( .A1(n7420), .A2(n4466), .ZN(n4463) );
  NAND2_X1 U6185 ( .A1(n4464), .A2(n4463), .ZN(n4757) );
  NAND2_X1 U6186 ( .A1(n9487), .A2(n4474), .ZN(n4471) );
  NAND2_X1 U6187 ( .A1(n4471), .A2(n4472), .ZN(n9443) );
  XNOR2_X2 U6188 ( .A(n4481), .B(P1_IR_REG_29__SCAN_IN), .ZN(n4939) );
  AND2_X2 U6189 ( .A1(n4870), .A2(n5418), .ZN(n4936) );
  OAI211_X1 U6190 ( .C1(n8825), .C2(n4487), .A(n4484), .B(n8901), .ZN(n5579)
         );
  NAND3_X1 U6191 ( .A1(n5527), .A2(n8825), .A3(n4485), .ZN(n4484) );
  NAND3_X1 U6192 ( .A1(n5527), .A2(n8825), .A3(n4863), .ZN(n8824) );
  NAND2_X1 U6193 ( .A1(n8898), .A2(n5580), .ZN(n8873) );
  INV_X1 U6194 ( .A(n4865), .ZN(n4495) );
  NAND2_X1 U6195 ( .A1(n4495), .A2(n4501), .ZN(n4496) );
  NAND3_X1 U6196 ( .A1(n4497), .A2(n4496), .A3(n4866), .ZN(n8922) );
  NAND3_X1 U6197 ( .A1(n4864), .A2(n4498), .A3(n4865), .ZN(n4497) );
  NAND2_X1 U6198 ( .A1(n4864), .A2(n4338), .ZN(n8960) );
  NAND3_X1 U6199 ( .A1(n4964), .A2(n4963), .A3(n4509), .ZN(n4965) );
  NAND2_X1 U6200 ( .A1(n4956), .A2(n4510), .ZN(n4509) );
  AND2_X2 U6201 ( .A1(n4929), .A2(n4928), .ZN(n5418) );
  NAND3_X1 U6202 ( .A1(n4929), .A2(n4928), .A3(n4513), .ZN(n4954) );
  NAND2_X1 U6203 ( .A1(n7582), .A2(n5303), .ZN(n5331) );
  NAND2_X1 U6204 ( .A1(n7582), .A2(n4516), .ZN(n8816) );
  NAND2_X1 U6205 ( .A1(n8816), .A2(n8817), .ZN(n5332) );
  NAND3_X1 U6206 ( .A1(n4519), .A2(n6608), .A3(n4317), .ZN(n4517) );
  AND2_X1 U6207 ( .A1(n9145), .A2(n6684), .ZN(n7098) );
  OR2_X1 U6208 ( .A1(n9383), .A2(n9706), .ZN(n4525) );
  NAND2_X1 U6209 ( .A1(n9383), .A2(n4530), .ZN(n9358) );
  NAND2_X1 U6210 ( .A1(n9383), .A2(n9711), .ZN(n9384) );
  NAND3_X1 U6211 ( .A1(n4526), .A2(n4525), .A3(n4524), .ZN(n9352) );
  NAND2_X1 U6212 ( .A1(n9383), .A2(n4527), .ZN(n4526) );
  NAND3_X1 U6213 ( .A1(n8974), .A2(n4332), .A3(n7504), .ZN(n7677) );
  INV_X1 U6214 ( .A(n4532), .ZN(n9594) );
  NAND2_X1 U6215 ( .A1(n9528), .A2(n4533), .ZN(n9481) );
  NAND2_X1 U6216 ( .A1(n6882), .A2(n6883), .ZN(n6881) );
  NAND2_X1 U6217 ( .A1(n6208), .A2(n7754), .ZN(n6882) );
  INV_X1 U6218 ( .A(n6882), .ZN(n7926) );
  AOI21_X1 U6219 ( .B1(n7471), .B2(n4540), .A(n4539), .ZN(n7989) );
  NAND4_X1 U6220 ( .A1(n4901), .A2(n6373), .A3(n5741), .A4(n5887), .ZN(n5915)
         );
  NAND2_X1 U6221 ( .A1(n4553), .A2(n4551), .ZN(n6273) );
  NAND2_X1 U6222 ( .A1(n8537), .A2(n4399), .ZN(n4554) );
  NAND2_X1 U6223 ( .A1(n4554), .A2(n4555), .ZN(n8498) );
  NAND2_X1 U6224 ( .A1(n4566), .A2(n4394), .ZN(n8465) );
  INV_X1 U6225 ( .A(n8598), .ZN(n4569) );
  AND2_X1 U6226 ( .A1(n8674), .A2(n8599), .ZN(n4578) );
  NAND3_X1 U6227 ( .A1(n5777), .A2(n4898), .A3(n5798), .ZN(n5801) );
  NAND2_X1 U6228 ( .A1(n4383), .A2(n4585), .ZN(n4582) );
  NAND2_X1 U6229 ( .A1(n4582), .A2(n4330), .ZN(n6495) );
  AND2_X1 U6230 ( .A1(n4582), .A2(n4583), .ZN(n8444) );
  INV_X1 U6231 ( .A(n6482), .ZN(n4585) );
  AOI21_X1 U6232 ( .B1(n4589), .B2(n4588), .A(n9568), .ZN(n9045) );
  NAND2_X1 U6233 ( .A1(n4592), .A2(n4590), .ZN(n9069) );
  OR2_X1 U6234 ( .A1(n9052), .A2(n4593), .ZN(n4592) );
  NAND2_X1 U6235 ( .A1(n8983), .A2(n9125), .ZN(n4606) );
  NAND2_X2 U6236 ( .A1(n6545), .A2(n6544), .ZN(n8983) );
  AOI21_X1 U6237 ( .B1(n8989), .B2(n9149), .A(n4604), .ZN(n8992) );
  NAND3_X1 U6238 ( .A1(n8982), .A2(n4607), .A3(n6545), .ZN(n4605) );
  NAND3_X1 U6239 ( .A1(n8982), .A2(n6545), .A3(n6544), .ZN(n4609) );
  INV_X1 U6240 ( .A(n9093), .ZN(n6707) );
  NAND2_X1 U6241 ( .A1(n6706), .A2(n9093), .ZN(n6709) );
  NAND2_X2 U6242 ( .A1(n4352), .A2(n4993), .ZN(n9256) );
  AOI21_X1 U6243 ( .B1(n4618), .B2(n9004), .A(n9003), .ZN(n9011) );
  NAND3_X1 U6244 ( .A1(n8994), .A2(n9125), .A3(n8993), .ZN(n4622) );
  NAND2_X1 U6245 ( .A1(n4637), .A2(n4636), .ZN(n6352) );
  INV_X1 U6246 ( .A(n4640), .ZN(n4638) );
  OAI21_X1 U6247 ( .B1(n8407), .B2(n4649), .A(n4647), .ZN(n8422) );
  NAND2_X1 U6248 ( .A1(n6366), .A2(n4652), .ZN(n4647) );
  XNOR2_X1 U6249 ( .A(n6365), .B(n8412), .ZN(n8407) );
  NAND2_X1 U6250 ( .A1(n4648), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4651) );
  INV_X1 U6251 ( .A(n8407), .ZN(n4648) );
  NAND2_X1 U6252 ( .A1(n8265), .A2(n4659), .ZN(n4658) );
  AOI21_X1 U6253 ( .B1(n8265), .B2(n4654), .A(n4655), .ZN(n4653) );
  NAND2_X1 U6254 ( .A1(n8265), .A2(n8261), .ZN(n4664) );
  INV_X1 U6255 ( .A(n4669), .ZN(n8290) );
  NAND2_X1 U6256 ( .A1(n4671), .A2(n4670), .ZN(n5776) );
  NAND2_X1 U6257 ( .A1(n5770), .A2(n6144), .ZN(n4671) );
  NAND2_X1 U6258 ( .A1(n5867), .A2(n5866), .ZN(n6986) );
  NAND2_X1 U6259 ( .A1(n6060), .A2(n4675), .ZN(n4674) );
  NOR2_X1 U6260 ( .A1(n8297), .A2(n6071), .ZN(n8052) );
  NAND2_X1 U6261 ( .A1(n8250), .A2(n4679), .ZN(n4677) );
  OAI21_X1 U6262 ( .B1(n8250), .B2(n4682), .A(n4678), .ZN(n8002) );
  NAND2_X1 U6263 ( .A1(n8311), .A2(n4406), .ZN(n8031) );
  NAND2_X1 U6264 ( .A1(n7279), .A2(n4396), .ZN(n7448) );
  NAND2_X1 U6265 ( .A1(n7152), .A2(n4395), .ZN(n7212) );
  AND2_X1 U6266 ( .A1(n5747), .A2(n4686), .ZN(n5777) );
  NAND2_X1 U6267 ( .A1(n5747), .A2(n5746), .ZN(n5781) );
  NAND2_X1 U6268 ( .A1(n7568), .A2(n4692), .ZN(n4691) );
  OAI21_X2 U6269 ( .B1(n7414), .B2(n4697), .A(n4695), .ZN(n7570) );
  AND2_X2 U6270 ( .A1(n9394), .A2(n9393), .ZN(n9395) );
  MUX2_X1 U6271 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6372), .S(n6602), .Z(n9992)
         );
  NAND2_X1 U6272 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5845), .ZN(n4714) );
  OAI21_X1 U6273 ( .B1(n6373), .B2(n8784), .A(P2_IR_REG_2__SCAN_IN), .ZN(n4715) );
  NAND2_X1 U6274 ( .A1(n6378), .A2(n4728), .ZN(n4724) );
  OAI211_X1 U6275 ( .C1(n6378), .C2(n4726), .A(n4724), .B(n4721), .ZN(n6924)
         );
  INV_X1 U6276 ( .A(n6384), .ZN(n7314) );
  NAND2_X1 U6277 ( .A1(n7069), .A2(n4745), .ZN(n4742) );
  INV_X1 U6278 ( .A(n4748), .ZN(n10021) );
  NAND2_X1 U6279 ( .A1(n4757), .A2(n4755), .ZN(n9569) );
  NAND2_X1 U6280 ( .A1(n4764), .A2(n4765), .ZN(n6537) );
  NAND2_X1 U6281 ( .A1(n9414), .A2(n4767), .ZN(n4764) );
  NAND2_X1 U6282 ( .A1(n7263), .A2(n4777), .ZN(n4776) );
  NAND2_X1 U6283 ( .A1(n4776), .A2(n4779), .ZN(n7422) );
  NAND2_X1 U6284 ( .A1(n6707), .A2(n6703), .ZN(n6705) );
  NAND4_X1 U6285 ( .A1(n4932), .A2(n4929), .A3(n4873), .A4(n4928), .ZN(n4969)
         );
  NAND2_X1 U6286 ( .A1(n4782), .A2(n5017), .ZN(n5021) );
  NAND2_X1 U6287 ( .A1(n5085), .A2(n4362), .ZN(n4789) );
  NAND2_X1 U6288 ( .A1(n4789), .A2(n4790), .ZN(n5125) );
  NAND2_X1 U6289 ( .A1(n5085), .A2(n5084), .ZN(n4792) );
  INV_X1 U6290 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4797) );
  INV_X1 U6291 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4796) );
  INV_X1 U6292 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4795) );
  NAND3_X1 U6293 ( .A1(n4797), .A2(n4796), .A3(n4795), .ZN(n4794) );
  NAND2_X1 U6294 ( .A1(n5696), .A2(n5695), .ZN(n4800) );
  INV_X1 U6295 ( .A(n5506), .ZN(n4815) );
  NAND2_X1 U6296 ( .A1(n5506), .A2(n4405), .ZN(n4804) );
  NAND3_X1 U6297 ( .A1(n5554), .A2(n4807), .A3(n5505), .ZN(n4806) );
  INV_X1 U6298 ( .A(n5505), .ZN(n4814) );
  OAI21_X1 U6299 ( .B1(n5334), .B2(n4820), .A(n4817), .ZN(n5385) );
  OAI21_X1 U6300 ( .B1(n5415), .B2(n5414), .A(n5416), .ZN(n5435) );
  OAI21_X1 U6301 ( .B1(n5415), .B2(n4828), .A(n4825), .ZN(n5481) );
  INV_X1 U6302 ( .A(n8911), .ZN(n4844) );
  OAI21_X1 U6303 ( .B1(n8911), .B2(n4848), .A(n4845), .ZN(n6585) );
  OAI21_X1 U6304 ( .B1(n8910), .B2(n4848), .A(n5102), .ZN(n4846) );
  NAND2_X1 U6305 ( .A1(n8911), .A2(n8910), .ZN(n8909) );
  NAND2_X1 U6306 ( .A1(n5102), .A2(n4848), .ZN(n4847) );
  OAI21_X1 U6307 ( .B1(n5102), .B2(n4850), .A(n8910), .ZN(n4849) );
  INV_X1 U6308 ( .A(n6586), .ZN(n4850) );
  NOR2_X1 U6309 ( .A1(n6724), .A2(n4367), .ZN(n6771) );
  XNOR2_X1 U6310 ( .A(n5007), .B(n5006), .ZN(n6726) );
  NAND2_X1 U6311 ( .A1(n4853), .A2(n5005), .ZN(n6725) );
  OR2_X1 U6312 ( .A1(n6719), .A2(n6718), .ZN(n4853) );
  NAND2_X1 U6313 ( .A1(n5174), .A2(n4860), .ZN(n4854) );
  NAND3_X1 U6314 ( .A1(n4854), .A2(n4856), .A3(n7394), .ZN(n7557) );
  NAND3_X1 U6315 ( .A1(n4859), .A2(n5173), .A3(n4857), .ZN(n4856) );
  INV_X1 U6316 ( .A(n7396), .ZN(n4860) );
  INV_X1 U6317 ( .A(n5172), .ZN(n4862) );
  NAND2_X1 U6318 ( .A1(n5353), .A2(n5352), .ZN(n4865) );
  OAI21_X1 U6319 ( .B1(n8475), .B2(n7885), .A(n7882), .ZN(n8470) );
  NAND2_X1 U6320 ( .A1(n8475), .A2(n4878), .ZN(n4877) );
  NAND2_X1 U6321 ( .A1(n4885), .A2(n4884), .ZN(n6220) );
  AND2_X1 U6322 ( .A1(n6219), .A2(n6218), .ZN(n4884) );
  OAI21_X1 U6323 ( .B1(n8548), .B2(n4890), .A(n4887), .ZN(n6225) );
  NAND2_X1 U6324 ( .A1(n4895), .A2(n4393), .ZN(n10031) );
  NAND2_X1 U6325 ( .A1(n4897), .A2(n4896), .ZN(n7352) );
  NOR2_X2 U6326 ( .A1(n5751), .A2(n4899), .ZN(n4898) );
  OR2_X1 U6327 ( .A1(n7727), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5016) );
  OAI21_X1 U6328 ( .B1(n7727), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n4973), .ZN(
        n5018) );
  NAND2_X1 U6329 ( .A1(n7727), .A2(n6595), .ZN(n4973) );
  AND2_X1 U6330 ( .A1(n9495), .A2(n9237), .ZN(n6525) );
  NAND2_X1 U6331 ( .A1(n7718), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5842) );
  OR2_X2 U6332 ( .A1(n7266), .A2(n9091), .ZN(n7264) );
  XNOR2_X1 U6333 ( .A(n6537), .B(n9120), .ZN(n9374) );
  AOI21_X2 U6334 ( .B1(n7507), .B2(n4781), .A(n6551), .ZN(n7415) );
  OR2_X1 U6335 ( .A1(n5973), .A2(n8339), .ZN(n5974) );
  CLKBUF_X1 U6337 ( .A(n7035), .Z(n7377) );
  NAND2_X1 U6338 ( .A1(n5526), .A2(n5525), .ZN(n8825) );
  NOR2_X4 U6339 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6373) );
  OAI22_X1 U6340 ( .A1(n8075), .A2(n8074), .B1(n6289), .B2(n5988), .ZN(n8265)
         );
  AND2_X2 U6341 ( .A1(n6580), .A2(n6752), .ZN(n9946) );
  AND2_X1 U6342 ( .A1(n6753), .A2(n9920), .ZN(n9934) );
  INV_X2 U6343 ( .A(n8634), .ZN(n8616) );
  INV_X1 U6344 ( .A(n9531), .ZN(n9742) );
  AND4_X1 U6345 ( .A1(n5992), .A2(n5759), .A3(n6016), .A4(n5758), .ZN(n4903)
         );
  AND3_X1 U6346 ( .A1(n5734), .A2(n9806), .A3(n5736), .ZN(n4904) );
  AND2_X1 U6347 ( .A1(n5476), .A2(n5475), .ZN(n4905) );
  OR2_X1 U6348 ( .A1(n9738), .A2(n8844), .ZN(n4907) );
  AND2_X1 U6349 ( .A1(n6298), .A2(n8514), .ZN(n4908) );
  OR2_X1 U6350 ( .A1(n6336), .A2(n8656), .ZN(n4909) );
  OR2_X1 U6351 ( .A1(n8447), .A2(n8656), .ZN(n4910) );
  OR2_X1 U6352 ( .A1(n8447), .A2(n8766), .ZN(n4911) );
  OR3_X1 U6353 ( .A1(n7969), .A2(n4314), .A3(n7968), .ZN(n4912) );
  OR2_X1 U6354 ( .A1(n6336), .A2(n8766), .ZN(n4913) );
  AND2_X1 U6355 ( .A1(n8003), .A2(n8529), .ZN(n4914) );
  INV_X1 U6356 ( .A(n9948), .ZN(n6508) );
  AND2_X1 U6357 ( .A1(n5205), .A2(n5183), .ZN(n4915) );
  INV_X1 U6358 ( .A(n9251), .ZN(n6504) );
  INV_X1 U6359 ( .A(n7925), .ZN(n6227) );
  INV_X1 U6360 ( .A(n9253), .ZN(n6499) );
  INV_X1 U6361 ( .A(n4987), .ZN(n5200) );
  INV_X1 U6362 ( .A(n7301), .ZN(n6514) );
  INV_X1 U6363 ( .A(n5330), .ZN(n5329) );
  NAND2_X1 U6364 ( .A1(n6284), .A2(n6283), .ZN(n7459) );
  AND2_X1 U6365 ( .A1(n5053), .A2(n5052), .ZN(n4916) );
  AND2_X1 U6366 ( .A1(n7622), .A2(n5251), .ZN(n4918) );
  INV_X1 U6367 ( .A(n8469), .ZN(n6304) );
  INV_X1 U6368 ( .A(n9383), .ZN(n9401) );
  NAND2_X1 U6369 ( .A1(n7905), .A2(n7910), .ZN(n7906) );
  NOR2_X1 U6370 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5743) );
  NAND2_X1 U6371 ( .A1(n7911), .A2(n7894), .ZN(n7912) );
  NAND2_X1 U6372 ( .A1(n6043), .A2(n6044), .ZN(n6045) );
  OR2_X1 U6373 ( .A1(n8533), .A2(n8542), .ZN(n6295) );
  AND2_X1 U6374 ( .A1(n6036), .A2(n6035), .ZN(n6051) );
  INV_X1 U6375 ( .A(n8488), .ZN(n6300) );
  OR2_X1 U6376 ( .A1(n5302), .A2(n5301), .ZN(n5303) );
  OR2_X1 U6377 ( .A1(n5252), .A2(n7624), .ZN(n5255) );
  NAND2_X1 U6378 ( .A1(n5081), .A2(n5082), .ZN(n5083) );
  INV_X1 U6379 ( .A(n5370), .ZN(n5368) );
  INV_X1 U6380 ( .A(n6905), .ZN(n6506) );
  INV_X1 U6381 ( .A(n9245), .ZN(n6513) );
  INV_X1 U6382 ( .A(n9247), .ZN(n6509) );
  INV_X1 U6383 ( .A(n8914), .ZN(n6503) );
  OR2_X1 U6384 ( .A1(n7698), .A2(n7697), .ZN(n7699) );
  INV_X1 U6385 ( .A(SI_22_), .ZN(n5507) );
  INV_X1 U6386 ( .A(n5131), .ZN(n4928) );
  NOR2_X1 U6387 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4927) );
  INV_X1 U6388 ( .A(n10100), .ZN(n6485) );
  OR2_X1 U6389 ( .A1(n6064), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6076) );
  OR2_X1 U6390 ( .A1(n6009), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6022) );
  INV_X1 U6391 ( .A(n7767), .ZN(n6211) );
  NAND2_X1 U6392 ( .A1(n8489), .A2(n6301), .ZN(n8477) );
  NAND2_X1 U6393 ( .A1(n7973), .A2(n7441), .ZN(n7919) );
  OR2_X1 U6394 ( .A1(n6306), .A2(n7968), .ZN(n6326) );
  INV_X1 U6395 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5760) );
  AND2_X1 U6396 ( .A1(n5122), .A2(n5121), .ZN(n5123) );
  INV_X1 U6397 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5163) );
  AND2_X1 U6398 ( .A1(n5094), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5112) );
  AND2_X1 U6399 ( .A1(n5580), .A2(n5578), .ZN(n8899) );
  AND2_X1 U6400 ( .A1(n5000), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5001) );
  OR2_X1 U6401 ( .A1(n5594), .A2(n5591), .ZN(n5618) );
  NAND2_X1 U6402 ( .A1(n5368), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5398) );
  INV_X1 U6403 ( .A(n9075), .ZN(n9377) );
  AND2_X1 U6404 ( .A1(n9645), .A2(n9235), .ZN(n6527) );
  NAND2_X1 U6405 ( .A1(n5396), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5425) );
  NOR2_X1 U6406 ( .A1(n9586), .A2(n8974), .ZN(n6520) );
  AND2_X1 U6407 ( .A1(n5112), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5138) );
  OR2_X1 U6408 ( .A1(n9610), .A2(n9246), .ZN(n6512) );
  NAND2_X1 U6409 ( .A1(n6497), .A2(n9145), .ZN(n6498) );
  OR2_X1 U6410 ( .A1(n5337), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U6411 ( .A1(n4317), .A2(n6599), .ZN(n5047) );
  AND2_X1 U6412 ( .A1(n6159), .A2(n6158), .ZN(n6160) );
  INV_X1 U6413 ( .A(n4314), .ZN(n7973) );
  INV_X1 U6414 ( .A(n7311), .ZN(n6427) );
  AOI21_X1 U6415 ( .B1(n6456), .B2(n10001), .A(n6455), .ZN(n6457) );
  INV_X1 U6416 ( .A(n8478), .ZN(n8315) );
  OR2_X1 U6417 ( .A1(n6128), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6133) );
  INV_X1 U6418 ( .A(n7952), .ZN(n8567) );
  INV_X1 U6419 ( .A(n6658), .ZN(n6327) );
  AND2_X1 U6420 ( .A1(n6313), .A2(n7910), .ZN(n8624) );
  NOR2_X1 U6421 ( .A1(n6322), .A2(n6164), .ZN(n6331) );
  NOR2_X1 U6422 ( .A1(n5164), .A2(n5163), .ZN(n5191) );
  OR2_X1 U6423 ( .A1(n5487), .A2(n8868), .ZN(n5515) );
  OR2_X1 U6424 ( .A1(n5342), .A2(n5341), .ZN(n5370) );
  OR2_X1 U6425 ( .A1(n5425), .A2(n8942), .ZN(n5461) );
  INV_X1 U6426 ( .A(n5010), .ZN(n5700) );
  NAND2_X1 U6427 ( .A1(n9183), .A2(n9074), .ZN(n9382) );
  AND2_X1 U6428 ( .A1(n9058), .A2(n9057), .ZN(n9478) );
  AND2_X1 U6429 ( .A1(n9174), .A2(n9181), .ZN(n9523) );
  AND2_X1 U6430 ( .A1(n9589), .A2(n6843), .ZN(n6844) );
  OR2_X1 U6431 ( .A1(n9753), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5676) );
  AND2_X1 U6432 ( .A1(n4316), .A2(n7709), .ZN(n6572) );
  INV_X1 U6433 ( .A(n9241), .ZN(n8966) );
  INV_X1 U6434 ( .A(n9548), .ZN(n9698) );
  INV_X1 U6435 ( .A(n9592), .ZN(n9544) );
  AND2_X1 U6436 ( .A1(n5697), .A2(n5642), .ZN(n5695) );
  NAND2_X1 U6437 ( .A1(n6161), .A2(n6160), .ZN(n6339) );
  INV_X1 U6438 ( .A(n8324), .ZN(n8283) );
  NAND2_X1 U6439 ( .A1(n6170), .A2(n10040), .ZN(n8303) );
  AND2_X1 U6440 ( .A1(n6193), .A2(n6192), .ZN(n8500) );
  AND4_X1 U6441 ( .A1(n6057), .A2(n6056), .A3(n6055), .A4(n6054), .ZN(n8101)
         );
  INV_X1 U6442 ( .A(n9982), .ZN(n10013) );
  AND2_X1 U6443 ( .A1(P2_U3893), .A2(n7977), .ZN(n10001) );
  INV_X1 U6444 ( .A(n10083), .ZN(n7344) );
  INV_X1 U6445 ( .A(n8604), .ZN(n10040) );
  INV_X1 U6446 ( .A(n10043), .ZN(n8605) );
  OR2_X1 U6447 ( .A1(n10124), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6494) );
  AND4_X1 U6448 ( .A1(n6322), .A2(n6964), .A3(n6963), .A4(n6321), .ZN(n6323)
         );
  AND2_X1 U6449 ( .A1(n7833), .A2(n7826), .ZN(n7988) );
  AND2_X1 U6450 ( .A1(n6485), .A2(n10104), .ZN(n10090) );
  AND2_X1 U6451 ( .A1(n6205), .A2(n6204), .ZN(n10100) );
  INV_X1 U6452 ( .A(n10090), .ZN(n10074) );
  INV_X1 U6453 ( .A(n10102), .ZN(n10081) );
  INV_X1 U6454 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5887) );
  OR2_X1 U6455 ( .A1(n5736), .A2(n5735), .ZN(n5737) );
  OR2_X1 U6456 ( .A1(n8810), .A2(n5010), .ZN(n5655) );
  OR2_X1 U6457 ( .A1(n6650), .A2(n6649), .ZN(n9343) );
  OR2_X1 U6458 ( .A1(n6650), .A2(n6641), .ZN(n9889) );
  OR2_X1 U6459 ( .A1(n6650), .A2(n6646), .ZN(n9895) );
  INV_X1 U6460 ( .A(n9895), .ZN(n9880) );
  INV_X1 U6461 ( .A(n4315), .ZN(n9347) );
  INV_X1 U6462 ( .A(n9928), .ZN(n9905) );
  AND2_X1 U6463 ( .A1(n5676), .A2(n9755), .ZN(n6579) );
  NAND2_X1 U6464 ( .A1(n9589), .A2(n9695), .ZN(n9944) );
  AND2_X1 U6465 ( .A1(n9125), .A2(n9126), .ZN(n7514) );
  AND2_X1 U6466 ( .A1(n5365), .A2(n5392), .ZN(n9870) );
  AND2_X1 U6467 ( .A1(n5237), .A2(n5261), .ZN(n9780) );
  INV_X1 U6468 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7149) );
  OR2_X1 U6469 ( .A1(n6339), .A2(n6338), .ZN(n6452) );
  INV_X1 U6470 ( .A(n6199), .ZN(n6200) );
  OR2_X1 U6471 ( .A1(n6167), .A2(n6166), .ZN(n8305) );
  INV_X1 U6472 ( .A(n8303), .ZN(n8332) );
  NAND2_X1 U6473 ( .A1(n6251), .A2(n6250), .ZN(n8478) );
  INV_X1 U6474 ( .A(n8063), .ZN(n8561) );
  OR2_X1 U6475 ( .A1(P2_U3150), .A2(n6453), .ZN(n9982) );
  INV_X1 U6476 ( .A(n10001), .ZN(n10019) );
  NAND2_X1 U6477 ( .A1(n6891), .A2(n6892), .ZN(n9967) );
  AND2_X1 U6478 ( .A1(n7038), .A2(n10040), .ZN(n8634) );
  NAND2_X1 U6479 ( .A1(n7321), .A2(n8616), .ZN(n10047) );
  NAND2_X1 U6480 ( .A1(n10124), .A2(n10081), .ZN(n8656) );
  INV_X1 U6481 ( .A(n8687), .ZN(n8694) );
  INV_X1 U6482 ( .A(n10124), .ZN(n10122) );
  INV_X1 U6483 ( .A(n8483), .ZN(n8714) );
  OR2_X1 U6484 ( .A1(n10108), .A2(n10090), .ZN(n8782) );
  AND2_X1 U6485 ( .A1(n6333), .A2(n6332), .ZN(n10108) );
  INV_X2 U6486 ( .A(n10108), .ZN(n10110) );
  AND2_X1 U6487 ( .A1(n6658), .A2(n6143), .ZN(n6687) );
  INV_X1 U6488 ( .A(n6687), .ZN(n6682) );
  INV_X1 U6489 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8794) );
  INV_X1 U6490 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7581) );
  INV_X1 U6491 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6998) );
  XNOR2_X1 U6492 ( .A(n5691), .B(n5690), .ZN(n6610) );
  NAND2_X1 U6493 ( .A1(n5729), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9810) );
  INV_X1 U6494 ( .A(n9806), .ZN(n8946) );
  INV_X1 U6495 ( .A(n8957), .ZN(n9803) );
  NAND2_X1 U6496 ( .A1(n5601), .A2(n5600), .ZN(n9449) );
  INV_X1 U6497 ( .A(n9866), .ZN(n9904) );
  INV_X1 U6498 ( .A(n9925), .ZN(n9913) );
  INV_X1 U6499 ( .A(n9931), .ZN(n9556) );
  INV_X1 U6500 ( .A(n9922), .ZN(n9910) );
  NAND2_X1 U6501 ( .A1(n9959), .A2(n9949), .ZN(n9685) );
  INV_X1 U6502 ( .A(n9959), .ZN(n9957) );
  INV_X1 U6503 ( .A(n9574), .ZN(n9748) );
  INV_X1 U6504 ( .A(n9936), .ZN(n9937) );
  INV_X1 U6505 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7692) );
  INV_X1 U6506 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6995) );
  NOR2_X1 U6507 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4922) );
  NOR2_X1 U6508 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4921) );
  NAND4_X1 U6509 ( .A1(n4922), .A2(n4921), .A3(n4920), .A4(n4919), .ZN(n4926)
         );
  NAND3_X1 U6510 ( .A1(n5217), .A2(n4924), .A3(n4923), .ZN(n4925) );
  NAND3_X1 U6511 ( .A1(n5022), .A2(n5070), .A3(n4927), .ZN(n5131) );
  NAND4_X1 U6512 ( .A1(n4944), .A2(n4946), .A3(n5671), .A4(n5669), .ZN(n4931)
         );
  NAND4_X1 U6513 ( .A1(n4955), .A2(n4949), .A3(n4952), .A4(n5690), .ZN(n4930)
         );
  NOR2_X2 U6514 ( .A1(n4931), .A2(n4930), .ZN(n4932) );
  XNOR2_X2 U6515 ( .A(n4935), .B(n4934), .ZN(n7705) );
  NAND2_X1 U6516 ( .A1(n5161), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4943) );
  INV_X1 U6517 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6637) );
  INV_X1 U6518 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n4938) );
  OR2_X1 U6519 ( .A1(n5011), .A2(n4938), .ZN(n4941) );
  NAND2_X1 U6520 ( .A1(n4954), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4945) );
  NAND2_X1 U6521 ( .A1(n5422), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4950) );
  NAND2_X1 U6522 ( .A1(n9126), .A2(n9216), .ZN(n9194) );
  AND2_X1 U6523 ( .A1(n5669), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4960) );
  NAND3_X1 U6524 ( .A1(n9756), .A2(P1_IR_REG_25__SCAN_IN), .A3(
        P1_IR_REG_24__SCAN_IN), .ZN(n4958) );
  NAND2_X1 U6525 ( .A1(n5669), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4957) );
  AND2_X1 U6526 ( .A1(n4958), .A2(n4957), .ZN(n4959) );
  AOI21_X1 U6527 ( .B1(n5667), .B2(n4960), .A(n4959), .ZN(n4964) );
  NAND2_X1 U6528 ( .A1(n4961), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4962) );
  INV_X1 U6529 ( .A(n9770), .ZN(n4963) );
  XNOR2_X2 U6530 ( .A(n4968), .B(n4967), .ZN(n5716) );
  NAND2_X1 U6531 ( .A1(n4969), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4970) );
  INV_X1 U6532 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6597) );
  INV_X1 U6533 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6595) );
  XNOR2_X1 U6534 ( .A(n5018), .B(SI_1_), .ZN(n5017) );
  AND2_X1 U6535 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4974) );
  NAND2_X1 U6536 ( .A1(n4317), .A2(n4974), .ZN(n4996) );
  AND2_X1 U6537 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4975) );
  NAND2_X1 U6538 ( .A1(n7727), .A2(n4975), .ZN(n5821) );
  NAND2_X1 U6539 ( .A1(n4320), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4979) );
  INV_X1 U6540 ( .A(n6608), .ZN(n4977) );
  NAND2_X1 U6541 ( .A1(n4977), .A2(n9261), .ZN(n4978) );
  NAND2_X1 U6542 ( .A1(n9088), .A2(n4315), .ZN(n6540) );
  NAND2_X1 U6543 ( .A1(n6540), .A2(n4316), .ZN(n4981) );
  INV_X1 U6544 ( .A(n9126), .ZN(n9217) );
  NAND2_X1 U6545 ( .A1(n5692), .A2(n9217), .ZN(n9087) );
  NAND2_X1 U6546 ( .A1(n4981), .A2(n9087), .ZN(n4982) );
  NAND2_X1 U6547 ( .A1(n5050), .A2(n4617), .ZN(n4983) );
  NAND2_X1 U6548 ( .A1(n4984), .A2(n4983), .ZN(n4986) );
  INV_X1 U6549 ( .A(n5007), .ZN(n5008) );
  INV_X1 U6550 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6626) );
  INV_X1 U6551 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n4988) );
  OR2_X1 U6552 ( .A1(n5010), .A2(n4988), .ZN(n4990) );
  NAND2_X1 U6553 ( .A1(n5161), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n4989) );
  INV_X1 U6554 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n4992) );
  OR2_X1 U6555 ( .A1(n5059), .A2(n4992), .ZN(n4993) );
  NAND2_X1 U6556 ( .A1(n4987), .A2(n9256), .ZN(n4999) );
  INV_X1 U6557 ( .A(SI_0_), .ZN(n4995) );
  INV_X1 U6558 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4994) );
  OAI21_X1 U6559 ( .B1(n4701), .B2(n4995), .A(n4994), .ZN(n4997) );
  AND2_X1 U6560 ( .A1(n4997), .A2(n4996), .ZN(n9771) );
  MUX2_X1 U6561 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9771), .S(n6608), .Z(n6755) );
  NAND2_X1 U6562 ( .A1(n5050), .A2(n6755), .ZN(n4998) );
  NAND2_X1 U6563 ( .A1(n4999), .A2(n4998), .ZN(n5003) );
  INV_X1 U6564 ( .A(n4965), .ZN(n5000) );
  INV_X1 U6565 ( .A(n6755), .ZN(n6684) );
  INV_X1 U6566 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9271) );
  OAI22_X1 U6567 ( .A1(n6684), .A2(n5200), .B1(n9271), .B2(n4965), .ZN(n5002)
         );
  AOI21_X1 U6568 ( .B1(n9256), .B2(n5036), .A(n5002), .ZN(n6718) );
  INV_X1 U6569 ( .A(n5009), .ZN(n5006) );
  NAND2_X1 U6570 ( .A1(n6613), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5015) );
  INV_X1 U6571 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9275) );
  OR2_X1 U6572 ( .A1(n5010), .A2(n9275), .ZN(n5014) );
  INV_X1 U6573 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6640) );
  OR2_X1 U6574 ( .A1(n5059), .A2(n6640), .ZN(n5013) );
  INV_X1 U6575 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6645) );
  OR2_X1 U6576 ( .A1(n4312), .A2(n6645), .ZN(n5012) );
  INV_X1 U6577 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6604) );
  XNOR2_X1 U6578 ( .A(n5043), .B(SI_2_), .ZN(n5041) );
  INV_X1 U6579 ( .A(n5018), .ZN(n5019) );
  NAND2_X1 U6580 ( .A1(n5019), .A2(SI_1_), .ZN(n5020) );
  XNOR2_X1 U6581 ( .A(n5042), .B(n5041), .ZN(n6603) );
  NAND2_X1 U6582 ( .A1(n5037), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5024) );
  INV_X2 U6583 ( .A(n6608), .ZN(n5440) );
  NAND2_X1 U6584 ( .A1(n5440), .A2(n9278), .ZN(n5023) );
  OAI211_X1 U6585 ( .C1(n5184), .C2(n6603), .A(n5024), .B(n5023), .ZN(n7101)
         );
  AOI22_X1 U6586 ( .A1(n9253), .A2(n4987), .B1(n7101), .B2(n5050), .ZN(n5025)
         );
  XNOR2_X1 U6587 ( .A(n5025), .B(n5710), .ZN(n5027) );
  AND2_X1 U6588 ( .A1(n7101), .A2(n4987), .ZN(n5026) );
  AOI21_X1 U6589 ( .B1(n9253), .B2(n5036), .A(n5026), .ZN(n5028) );
  XNOR2_X1 U6590 ( .A(n5027), .B(n5028), .ZN(n6772) );
  INV_X1 U6591 ( .A(n5027), .ZN(n5030) );
  INV_X1 U6592 ( .A(n5028), .ZN(n5029) );
  OAI22_X1 U6593 ( .A1(n6771), .A2(n6772), .B1(n5030), .B2(n5029), .ZN(n6781)
         );
  INV_X1 U6594 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5031) );
  OR2_X1 U6595 ( .A1(n4313), .A2(n5031), .ZN(n5034) );
  INV_X1 U6596 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9921) );
  OR2_X1 U6597 ( .A1(n5059), .A2(n9921), .ZN(n5033) );
  OR2_X1 U6598 ( .A1(n5010), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5032) );
  INV_X1 U6599 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5038) );
  NAND2_X1 U6600 ( .A1(n5072), .A2(n5038), .ZN(n5039) );
  NAND2_X1 U6601 ( .A1(n5039), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5040) );
  AOI22_X1 U6602 ( .A1(n5037), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n5440), .B2(
        n6671), .ZN(n5049) );
  NAND2_X1 U6603 ( .A1(n5042), .A2(n5041), .ZN(n5046) );
  INV_X1 U6604 ( .A(n5043), .ZN(n5044) );
  NAND2_X1 U6605 ( .A1(n5044), .A2(SI_2_), .ZN(n5045) );
  INV_X1 U6606 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6601) );
  INV_X1 U6607 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6599) );
  XNOR2_X1 U6608 ( .A(n5066), .B(SI_3_), .ZN(n5064) );
  XNOR2_X1 U6609 ( .A(n5065), .B(n5064), .ZN(n6600) );
  OR2_X1 U6610 ( .A1(n6600), .A2(n5184), .ZN(n5048) );
  NAND2_X1 U6611 ( .A1(n5049), .A2(n5048), .ZN(n9924) );
  AOI22_X1 U6612 ( .A1(n9252), .A2(n5036), .B1(n5569), .B2(n9924), .ZN(n5052)
         );
  AOI22_X1 U6613 ( .A1(n9252), .A2(n5569), .B1(n9924), .B2(n5615), .ZN(n5051)
         );
  XNOR2_X1 U6614 ( .A(n5051), .B(n5710), .ZN(n5053) );
  XOR2_X1 U6615 ( .A(n5053), .B(n5052), .Z(n6780) );
  INV_X1 U6616 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5054) );
  INV_X1 U6617 ( .A(n5161), .ZN(n5373) );
  INV_X1 U6618 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5055) );
  OR2_X1 U6619 ( .A1(n5373), .A2(n5055), .ZN(n5062) );
  INV_X1 U6620 ( .A(n5094), .ZN(n5095) );
  INV_X1 U6621 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5057) );
  INV_X1 U6622 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5056) );
  NAND2_X1 U6623 ( .A1(n5057), .A2(n5056), .ZN(n5058) );
  NAND2_X1 U6624 ( .A1(n5095), .A2(n5058), .ZN(n8912) );
  OR2_X1 U6625 ( .A1(n5010), .A2(n8912), .ZN(n5061) );
  INV_X1 U6626 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6847) );
  OR2_X1 U6627 ( .A1(n5651), .A2(n6847), .ZN(n5060) );
  NAND2_X1 U6628 ( .A1(n9251), .A2(n5036), .ZN(n5077) );
  NAND2_X1 U6629 ( .A1(n5065), .A2(n5064), .ZN(n5069) );
  INV_X1 U6630 ( .A(n5066), .ZN(n5067) );
  NAND2_X1 U6631 ( .A1(n5067), .A2(SI_3_), .ZN(n5068) );
  INV_X1 U6632 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6605) );
  INV_X1 U6633 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6607) );
  MUX2_X1 U6634 ( .A(n6605), .B(n6607), .S(n4317), .Z(n5086) );
  XNOR2_X1 U6635 ( .A(n5086), .B(SI_4_), .ZN(n5084) );
  XNOR2_X1 U6636 ( .A(n5085), .B(n5084), .ZN(n6606) );
  OR2_X1 U6637 ( .A1(n6606), .A2(n5184), .ZN(n5075) );
  OR2_X1 U6638 ( .A1(n5070), .A2(n9756), .ZN(n5071) );
  NAND2_X1 U6639 ( .A1(n5072), .A2(n5071), .ZN(n5089) );
  INV_X1 U6640 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5073) );
  XNOR2_X1 U6641 ( .A(n5089), .B(n5073), .ZN(n9292) );
  AOI22_X1 U6642 ( .A1(n5037), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n5440), .B2(
        n9292), .ZN(n5074) );
  NAND2_X1 U6643 ( .A1(n5075), .A2(n5074), .ZN(n8914) );
  NAND2_X1 U6644 ( .A1(n8914), .A2(n4987), .ZN(n5076) );
  NAND2_X1 U6645 ( .A1(n5077), .A2(n5076), .ZN(n5082) );
  NAND2_X1 U6646 ( .A1(n9251), .A2(n4987), .ZN(n5079) );
  NAND2_X1 U6647 ( .A1(n8914), .A2(n5615), .ZN(n5078) );
  NAND2_X1 U6648 ( .A1(n5079), .A2(n5078), .ZN(n5080) );
  XNOR2_X1 U6649 ( .A(n5080), .B(n5710), .ZN(n5081) );
  XOR2_X1 U6650 ( .A(n5082), .B(n5081), .Z(n8910) );
  INV_X1 U6651 ( .A(n5086), .ZN(n5087) );
  NAND2_X1 U6652 ( .A1(n5087), .A2(SI_4_), .ZN(n5088) );
  INV_X1 U6653 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6619) );
  MUX2_X1 U6654 ( .A(n6622), .B(n6619), .S(n4317), .Z(n5105) );
  XNOR2_X1 U6655 ( .A(n5104), .B(n5103), .ZN(n6621) );
  OR2_X1 U6656 ( .A1(n6621), .A2(n5184), .ZN(n5092) );
  OAI21_X1 U6657 ( .B1(n5089), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5090) );
  XNOR2_X1 U6658 ( .A(n5090), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9311) );
  AOI22_X1 U6659 ( .A1(n5037), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5440), .B2(
        n9311), .ZN(n5091) );
  NAND2_X1 U6660 ( .A1(n5092), .A2(n5091), .ZN(n6905) );
  NAND2_X1 U6661 ( .A1(n5701), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5100) );
  INV_X1 U6662 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5093) );
  OR2_X1 U6663 ( .A1(n5373), .A2(n5093), .ZN(n5099) );
  INV_X1 U6664 ( .A(n5112), .ZN(n5113) );
  INV_X1 U6665 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8141) );
  NAND2_X1 U6666 ( .A1(n5095), .A2(n8141), .ZN(n5096) );
  NAND2_X1 U6667 ( .A1(n5113), .A2(n5096), .ZN(n6906) );
  OR2_X1 U6668 ( .A1(n5010), .A2(n6906), .ZN(n5098) );
  INV_X1 U6669 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6666) );
  OR2_X1 U6670 ( .A1(n5651), .A2(n6666), .ZN(n5097) );
  NAND4_X1 U6671 ( .A1(n5100), .A2(n5099), .A3(n5098), .A4(n5097), .ZN(n9250)
         );
  AOI22_X1 U6672 ( .A1(n6905), .A2(n5615), .B1(n5569), .B2(n9250), .ZN(n5101)
         );
  AOI22_X1 U6673 ( .A1(n6905), .A2(n5569), .B1(n5036), .B2(n9250), .ZN(n6586)
         );
  INV_X1 U6674 ( .A(n5105), .ZN(n5106) );
  INV_X1 U6675 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5107) );
  MUX2_X1 U6676 ( .A(n6635), .B(n5107), .S(n4317), .Z(n5126) );
  XNOR2_X1 U6677 ( .A(n5126), .B(SI_6_), .ZN(n5124) );
  XNOR2_X1 U6678 ( .A(n5125), .B(n5124), .ZN(n6634) );
  OR2_X1 U6679 ( .A1(n6634), .A2(n5184), .ZN(n5110) );
  NAND2_X1 U6680 ( .A1(n5131), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5108) );
  XNOR2_X1 U6681 ( .A(n5108), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6739) );
  AOI22_X1 U6682 ( .A1(n5037), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5440), .B2(
        n6739), .ZN(n5109) );
  NAND2_X1 U6683 ( .A1(n5110), .A2(n5109), .ZN(n9948) );
  NAND2_X1 U6684 ( .A1(n5701), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5119) );
  INV_X1 U6685 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5111) );
  OR2_X1 U6686 ( .A1(n5373), .A2(n5111), .ZN(n5118) );
  INV_X1 U6687 ( .A(n5138), .ZN(n5115) );
  INV_X1 U6688 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7109) );
  NAND2_X1 U6689 ( .A1(n5113), .A2(n7109), .ZN(n5114) );
  NAND2_X1 U6690 ( .A1(n5115), .A2(n5114), .ZN(n7110) );
  OR2_X1 U6691 ( .A1(n5010), .A2(n7110), .ZN(n5117) );
  INV_X1 U6692 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7058) );
  OR2_X1 U6693 ( .A1(n5651), .A2(n7058), .ZN(n5116) );
  NAND4_X1 U6694 ( .A1(n5119), .A2(n5118), .A3(n5117), .A4(n5116), .ZN(n9249)
         );
  AOI22_X1 U6695 ( .A1(n9948), .A2(n5615), .B1(n5569), .B2(n9249), .ZN(n5120)
         );
  XNOR2_X1 U6696 ( .A(n5120), .B(n5710), .ZN(n5122) );
  AOI22_X1 U6697 ( .A1(n9948), .A2(n5569), .B1(n5036), .B2(n9249), .ZN(n5121)
         );
  XNOR2_X1 U6698 ( .A(n5122), .B(n5121), .ZN(n7108) );
  NAND2_X1 U6699 ( .A1(n5125), .A2(n5124), .ZN(n5129) );
  INV_X1 U6700 ( .A(n5126), .ZN(n5127) );
  NAND2_X1 U6701 ( .A1(n5127), .A2(SI_6_), .ZN(n5128) );
  INV_X1 U6702 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5130) );
  MUX2_X1 U6703 ( .A(n6657), .B(n5130), .S(n4317), .Z(n5149) );
  XNOR2_X1 U6704 ( .A(n5149), .B(SI_7_), .ZN(n5147) );
  XNOR2_X1 U6705 ( .A(n5148), .B(n5147), .ZN(n6656) );
  OR2_X1 U6706 ( .A1(n6656), .A2(n5184), .ZN(n5137) );
  OR2_X1 U6707 ( .A1(n5131), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5133) );
  NAND2_X1 U6708 ( .A1(n5133), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5132) );
  MUX2_X1 U6709 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5132), .S(
        P1_IR_REG_7__SCAN_IN), .Z(n5135) );
  INV_X1 U6710 ( .A(n5218), .ZN(n5134) );
  AOI22_X1 U6711 ( .A1(n5037), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5440), .B2(
        n9792), .ZN(n5136) );
  NAND2_X1 U6712 ( .A1(n6613), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5142) );
  INV_X1 U6713 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6734) );
  OR2_X1 U6714 ( .A1(n4312), .A2(n6734), .ZN(n5141) );
  NAND2_X1 U6715 ( .A1(n5138), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5164) );
  OAI21_X1 U6716 ( .B1(n5138), .B2(P1_REG3_REG_7__SCAN_IN), .A(n5164), .ZN(
        n7204) );
  OR2_X1 U6717 ( .A1(n5010), .A2(n7204), .ZN(n5140) );
  INV_X1 U6718 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7170) );
  OR2_X1 U6719 ( .A1(n5651), .A2(n7170), .ZN(n5139) );
  NAND4_X1 U6720 ( .A1(n5142), .A2(n5141), .A3(n5140), .A4(n5139), .ZN(n9248)
         );
  AOI22_X1 U6721 ( .A1(n7208), .A2(n5615), .B1(n5569), .B2(n9248), .ZN(n5143)
         );
  XOR2_X1 U6722 ( .A(n5710), .B(n5143), .Z(n7201) );
  INV_X1 U6723 ( .A(n7201), .ZN(n5145) );
  AND2_X1 U6724 ( .A1(n9248), .A2(n5036), .ZN(n5144) );
  AOI21_X1 U6725 ( .B1(n7208), .B2(n5569), .A(n5144), .ZN(n7200) );
  INV_X1 U6726 ( .A(n7200), .ZN(n5146) );
  NAND2_X1 U6727 ( .A1(n5148), .A2(n5147), .ZN(n5152) );
  INV_X1 U6728 ( .A(n5149), .ZN(n5150) );
  NAND2_X1 U6729 ( .A1(n5150), .A2(SI_7_), .ZN(n5151) );
  INV_X1 U6730 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5153) );
  MUX2_X1 U6731 ( .A(n6662), .B(n5153), .S(n4317), .Z(n5155) );
  INV_X1 U6732 ( .A(SI_8_), .ZN(n5154) );
  NAND2_X1 U6733 ( .A1(n5155), .A2(n5154), .ZN(n5177) );
  INV_X1 U6734 ( .A(n5155), .ZN(n5156) );
  NAND2_X1 U6735 ( .A1(n5156), .A2(SI_8_), .ZN(n5157) );
  NAND2_X1 U6736 ( .A1(n5177), .A2(n5157), .ZN(n5175) );
  INV_X1 U6737 ( .A(n5175), .ZN(n5158) );
  XNOR2_X1 U6738 ( .A(n5176), .B(n5158), .ZN(n6661) );
  OR2_X1 U6739 ( .A1(n6661), .A2(n5184), .ZN(n5160) );
  OR2_X1 U6740 ( .A1(n5218), .A2(n9756), .ZN(n5186) );
  XNOR2_X1 U6741 ( .A(n5186), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6798) );
  AOI22_X1 U6742 ( .A1(n5037), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5440), .B2(
        n6798), .ZN(n5159) );
  NAND2_X1 U6743 ( .A1(n5160), .A2(n5159), .ZN(n8857) );
  NAND2_X1 U6744 ( .A1(n6613), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5169) );
  INV_X1 U6745 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5162) );
  OR2_X1 U6746 ( .A1(n5059), .A2(n5162), .ZN(n5168) );
  AND2_X1 U6747 ( .A1(n5164), .A2(n5163), .ZN(n5165) );
  OR2_X1 U6748 ( .A1(n5165), .A2(n5191), .ZN(n8858) );
  OR2_X1 U6749 ( .A1(n5010), .A2(n8858), .ZN(n5167) );
  INV_X1 U6750 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6735) );
  OR2_X1 U6751 ( .A1(n4313), .A2(n6735), .ZN(n5166) );
  NAND4_X1 U6752 ( .A1(n5169), .A2(n5168), .A3(n5167), .A4(n5166), .ZN(n9247)
         );
  AOI22_X1 U6753 ( .A1(n8857), .A2(n5615), .B1(n5569), .B2(n9247), .ZN(n5170)
         );
  XNOR2_X1 U6754 ( .A(n5170), .B(n5710), .ZN(n5171) );
  NAND2_X1 U6755 ( .A1(n5172), .A2(n5171), .ZN(n5173) );
  OAI22_X1 U6756 ( .A1(n4520), .A2(n5200), .B1(n6509), .B2(n5657), .ZN(n8852)
         );
  INV_X1 U6757 ( .A(n5173), .ZN(n5174) );
  INV_X1 U6758 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5179) );
  MUX2_X1 U6759 ( .A(n6696), .B(n5179), .S(n4317), .Z(n5181) );
  INV_X1 U6760 ( .A(SI_9_), .ZN(n5180) );
  NAND2_X1 U6761 ( .A1(n5181), .A2(n5180), .ZN(n5205) );
  INV_X1 U6762 ( .A(n5181), .ZN(n5182) );
  NAND2_X1 U6763 ( .A1(n5182), .A2(SI_9_), .ZN(n5183) );
  NAND2_X1 U6764 ( .A1(n6694), .A2(n9080), .ZN(n5190) );
  INV_X1 U6765 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6766 ( .A1(n5186), .A2(n5185), .ZN(n5187) );
  NAND2_X1 U6767 ( .A1(n5187), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5188) );
  XNOR2_X1 U6768 ( .A(n5188), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7249) );
  AOI22_X1 U6769 ( .A1(n5037), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5440), .B2(
        n7249), .ZN(n5189) );
  NAND2_X1 U6770 ( .A1(n9610), .A2(n5615), .ZN(n5198) );
  NAND2_X1 U6771 ( .A1(n6613), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5196) );
  INV_X1 U6772 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6790) );
  OR2_X1 U6773 ( .A1(n4313), .A2(n6790), .ZN(n5195) );
  NAND2_X1 U6774 ( .A1(n5191), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5241) );
  OR2_X1 U6775 ( .A1(n5191), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6776 ( .A1(n5241), .A2(n5192), .ZN(n9608) );
  OR2_X1 U6777 ( .A1(n5010), .A2(n9608), .ZN(n5194) );
  INV_X1 U6778 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6799) );
  OR2_X1 U6779 ( .A1(n5651), .A2(n6799), .ZN(n5193) );
  NAND4_X1 U6780 ( .A1(n5196), .A2(n5195), .A3(n5194), .A4(n5193), .ZN(n9246)
         );
  CLKBUF_X3 U6781 ( .A(n4987), .Z(n5569) );
  NAND2_X1 U6782 ( .A1(n9246), .A2(n5569), .ZN(n5197) );
  NAND2_X1 U6783 ( .A1(n5198), .A2(n5197), .ZN(n5199) );
  XNOR2_X1 U6784 ( .A(n5199), .B(n5628), .ZN(n5203) );
  AND2_X1 U6785 ( .A1(n9246), .A2(n5036), .ZN(n5201) );
  AOI21_X1 U6786 ( .B1(n9610), .B2(n5569), .A(n5201), .ZN(n5202) );
  NOR2_X1 U6787 ( .A1(n5203), .A2(n5202), .ZN(n7396) );
  NAND2_X1 U6788 ( .A1(n5203), .A2(n5202), .ZN(n7394) );
  NAND2_X1 U6789 ( .A1(n5204), .A2(n4915), .ZN(n5206) );
  MUX2_X1 U6790 ( .A(n6700), .B(n5207), .S(n4317), .Z(n5208) );
  XNOR2_X1 U6791 ( .A(n5208), .B(SI_10_), .ZN(n5233) );
  INV_X1 U6792 ( .A(n5233), .ZN(n5211) );
  INV_X1 U6793 ( .A(n5208), .ZN(n5209) );
  NAND2_X1 U6794 ( .A1(n5209), .A2(SI_10_), .ZN(n5210) );
  MUX2_X1 U6795 ( .A(n6732), .B(n5212), .S(n4317), .Z(n5214) );
  NAND2_X1 U6796 ( .A1(n5214), .A2(n5213), .ZN(n5260) );
  INV_X1 U6797 ( .A(n5214), .ZN(n5215) );
  NAND2_X1 U6798 ( .A1(n5215), .A2(SI_11_), .ZN(n5216) );
  NAND2_X1 U6799 ( .A1(n5260), .A2(n5216), .ZN(n5258) );
  XNOR2_X1 U6800 ( .A(n5259), .B(n5258), .ZN(n6722) );
  NAND2_X1 U6801 ( .A1(n6722), .A2(n9080), .ZN(n5221) );
  NAND2_X1 U6802 ( .A1(n5218), .A2(n5217), .ZN(n5235) );
  NAND2_X1 U6803 ( .A1(n5261), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5219) );
  XNOR2_X1 U6804 ( .A(n5219), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9819) );
  AOI22_X1 U6805 ( .A1(n5037), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5440), .B2(
        n9819), .ZN(n5220) );
  NAND2_X1 U6806 ( .A1(n7632), .A2(n5615), .ZN(n5231) );
  NAND2_X1 U6807 ( .A1(n6613), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5229) );
  INV_X1 U6808 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5222) );
  OR2_X1 U6809 ( .A1(n5651), .A2(n5222), .ZN(n5228) );
  INV_X1 U6810 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7561) );
  INV_X1 U6811 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5223) );
  OAI21_X1 U6812 ( .B1(n5241), .B2(n7561), .A(n5223), .ZN(n5225) );
  NAND2_X1 U6813 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n5224) );
  NAND2_X1 U6814 ( .A1(n5225), .A2(n5268), .ZN(n9907) );
  OR2_X1 U6815 ( .A1(n5010), .A2(n9907), .ZN(n5227) );
  INV_X1 U6816 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7251) );
  OR2_X1 U6817 ( .A1(n4312), .A2(n7251), .ZN(n5226) );
  NAND4_X1 U6818 ( .A1(n5229), .A2(n5228), .A3(n5227), .A4(n5226), .ZN(n9244)
         );
  NAND2_X1 U6819 ( .A1(n9244), .A2(n4987), .ZN(n5230) );
  NAND2_X1 U6820 ( .A1(n5231), .A2(n5230), .ZN(n5232) );
  XNOR2_X1 U6821 ( .A(n5232), .B(n4985), .ZN(n7624) );
  INV_X1 U6822 ( .A(n7632), .ZN(n9914) );
  INV_X1 U6823 ( .A(n9244), .ZN(n6516) );
  OAI22_X1 U6824 ( .A1(n9914), .A2(n5200), .B1(n6516), .B2(n5657), .ZN(n7623)
         );
  NAND2_X1 U6825 ( .A1(n7624), .A2(n7623), .ZN(n7622) );
  NAND2_X1 U6826 ( .A1(n6698), .A2(n9080), .ZN(n5239) );
  NAND2_X1 U6827 ( .A1(n5235), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5236) );
  MUX2_X1 U6828 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5236), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5237) );
  AOI22_X1 U6829 ( .A1(n5037), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5440), .B2(
        n9780), .ZN(n5238) );
  NAND2_X1 U6830 ( .A1(n7301), .A2(n5615), .ZN(n5247) );
  NAND2_X1 U6831 ( .A1(n6613), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5245) );
  INV_X1 U6832 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5240) );
  OR2_X1 U6833 ( .A1(n5651), .A2(n5240), .ZN(n5244) );
  XNOR2_X1 U6834 ( .A(n5241), .B(n7561), .ZN(n7273) );
  OR2_X1 U6835 ( .A1(n5010), .A2(n7273), .ZN(n5243) );
  INV_X1 U6836 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7250) );
  OR2_X1 U6837 ( .A1(n4313), .A2(n7250), .ZN(n5242) );
  NAND4_X1 U6838 ( .A1(n5245), .A2(n5244), .A3(n5243), .A4(n5242), .ZN(n9245)
         );
  NAND2_X1 U6839 ( .A1(n9245), .A2(n4987), .ZN(n5246) );
  NAND2_X1 U6840 ( .A1(n5247), .A2(n5246), .ZN(n5248) );
  XNOR2_X1 U6841 ( .A(n5248), .B(n5628), .ZN(n7626) );
  NAND2_X1 U6842 ( .A1(n7301), .A2(n4987), .ZN(n5250) );
  NAND2_X1 U6843 ( .A1(n9245), .A2(n5036), .ZN(n5249) );
  NAND2_X1 U6844 ( .A1(n7557), .A2(n4918), .ZN(n5257) );
  INV_X1 U6845 ( .A(n7623), .ZN(n5253) );
  AOI21_X1 U6846 ( .B1(n7626), .B2(n7558), .A(n5253), .ZN(n5252) );
  NAND3_X1 U6847 ( .A1(n5253), .A2(n7558), .A3(n7626), .ZN(n5254) );
  NAND2_X1 U6848 ( .A1(n5257), .A2(n5256), .ZN(n9797) );
  MUX2_X1 U6849 ( .A(n6787), .B(n6814), .S(n4317), .Z(n5281) );
  XNOR2_X1 U6850 ( .A(n5281), .B(SI_12_), .ZN(n5280) );
  XNOR2_X1 U6851 ( .A(n5283), .B(n5280), .ZN(n6786) );
  NAND2_X1 U6852 ( .A1(n6786), .A2(n9080), .ZN(n5267) );
  OR2_X1 U6853 ( .A1(n5315), .A2(n9756), .ZN(n5264) );
  INV_X1 U6854 ( .A(n5264), .ZN(n5262) );
  NAND2_X1 U6855 ( .A1(n5262), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5265) );
  INV_X1 U6856 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5263) );
  NAND2_X1 U6857 ( .A1(n5264), .A2(n5263), .ZN(n5284) );
  AOI22_X1 U6858 ( .A1(n5037), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9331), .B2(
        n5440), .ZN(n5266) );
  NAND2_X1 U6859 ( .A1(n6613), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5274) );
  NAND2_X1 U6860 ( .A1(n5268), .A2(n7255), .ZN(n5269) );
  NAND2_X1 U6861 ( .A1(n5289), .A2(n5269), .ZN(n9809) );
  OR2_X1 U6862 ( .A1(n5010), .A2(n9809), .ZN(n5273) );
  INV_X1 U6863 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7425) );
  OR2_X1 U6864 ( .A1(n5059), .A2(n7425), .ZN(n5272) );
  INV_X1 U6865 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5270) );
  OR2_X1 U6866 ( .A1(n4312), .A2(n5270), .ZN(n5271) );
  NAND4_X1 U6867 ( .A1(n5274), .A2(n5273), .A3(n5272), .A4(n5271), .ZN(n9243)
         );
  AOI22_X1 U6868 ( .A1(n7434), .A2(n5615), .B1(n5569), .B2(n9243), .ZN(n5275)
         );
  XOR2_X1 U6869 ( .A(n4985), .B(n5275), .Z(n5277) );
  INV_X1 U6870 ( .A(n9243), .ZN(n7586) );
  OAI22_X1 U6871 ( .A1(n9804), .A2(n5200), .B1(n7586), .B2(n5657), .ZN(n5276)
         );
  NOR2_X1 U6872 ( .A1(n5277), .A2(n5276), .ZN(n5278) );
  AOI21_X1 U6873 ( .B1(n5277), .B2(n5276), .A(n5278), .ZN(n9798) );
  NAND2_X1 U6874 ( .A1(n9797), .A2(n9798), .ZN(n9796) );
  INV_X1 U6875 ( .A(n5278), .ZN(n5279) );
  NAND2_X1 U6876 ( .A1(n9796), .A2(n5279), .ZN(n7583) );
  INV_X1 U6877 ( .A(n5281), .ZN(n5282) );
  MUX2_X1 U6878 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4518), .Z(n5307) );
  XNOR2_X1 U6879 ( .A(n5307), .B(SI_13_), .ZN(n5304) );
  XNOR2_X1 U6880 ( .A(n5306), .B(n5304), .ZN(n6815) );
  NAND2_X1 U6881 ( .A1(n6815), .A2(n9080), .ZN(n5287) );
  NAND2_X1 U6882 ( .A1(n5284), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5285) );
  AOI22_X1 U6883 ( .A1(n9831), .A2(n5440), .B1(n5037), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6884 ( .A1(n9697), .A2(n5615), .ZN(n5298) );
  NAND2_X1 U6885 ( .A1(n6613), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5296) );
  NAND2_X1 U6886 ( .A1(n5289), .A2(n5288), .ZN(n5290) );
  NAND2_X1 U6887 ( .A1(n5321), .A2(n5290), .ZN(n7492) );
  OR2_X1 U6888 ( .A1(n5010), .A2(n7492), .ZN(n5295) );
  INV_X1 U6889 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n5291) );
  OR2_X1 U6890 ( .A1(n5651), .A2(n5291), .ZN(n5294) );
  INV_X1 U6891 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n5292) );
  OR2_X1 U6892 ( .A1(n4312), .A2(n5292), .ZN(n5293) );
  NAND4_X1 U6893 ( .A1(n5296), .A2(n5295), .A3(n5294), .A4(n5293), .ZN(n9242)
         );
  NAND2_X1 U6894 ( .A1(n9242), .A2(n5569), .ZN(n5297) );
  NAND2_X1 U6895 ( .A1(n5298), .A2(n5297), .ZN(n5299) );
  XNOR2_X1 U6896 ( .A(n5299), .B(n4985), .ZN(n5302) );
  AOI22_X1 U6897 ( .A1(n9697), .A2(n5569), .B1(n5036), .B2(n9242), .ZN(n5300)
         );
  XNOR2_X1 U6898 ( .A(n5302), .B(n5300), .ZN(n7584) );
  INV_X1 U6899 ( .A(n5300), .ZN(n5301) );
  INV_X1 U6900 ( .A(n5304), .ZN(n5305) );
  NAND2_X1 U6901 ( .A1(n5306), .A2(n5305), .ZN(n5309) );
  NAND2_X1 U6902 ( .A1(n5307), .A2(SI_13_), .ZN(n5308) );
  MUX2_X1 U6903 ( .A(n6998), .B(n6995), .S(n4317), .Z(n5311) );
  INV_X1 U6904 ( .A(n5311), .ZN(n5312) );
  NAND2_X1 U6905 ( .A1(n5312), .A2(SI_14_), .ZN(n5313) );
  NAND2_X1 U6906 ( .A1(n5335), .A2(n5313), .ZN(n5333) );
  XNOR2_X1 U6907 ( .A(n5334), .B(n5333), .ZN(n6994) );
  NAND2_X1 U6908 ( .A1(n6994), .A2(n9080), .ZN(n5318) );
  NOR2_X1 U6909 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5314) );
  NAND2_X1 U6910 ( .A1(n5315), .A2(n5314), .ZN(n5337) );
  NAND2_X1 U6911 ( .A1(n5337), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5316) );
  XNOR2_X1 U6912 ( .A(n5316), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9843) );
  AOI22_X1 U6913 ( .A1(n5440), .A2(n9843), .B1(n5037), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6914 ( .A1(n5701), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5327) );
  INV_X1 U6915 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5319) );
  OR2_X1 U6916 ( .A1(n5373), .A2(n5319), .ZN(n5326) );
  INV_X1 U6917 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8819) );
  NAND2_X1 U6918 ( .A1(n5321), .A2(n8819), .ZN(n5322) );
  NAND2_X1 U6919 ( .A1(n5342), .A2(n5322), .ZN(n9596) );
  OR2_X1 U6920 ( .A1(n5010), .A2(n9596), .ZN(n5325) );
  INV_X1 U6921 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n5323) );
  OR2_X1 U6922 ( .A1(n5059), .A2(n5323), .ZN(n5324) );
  NAND4_X1 U6923 ( .A1(n5327), .A2(n5326), .A3(n5325), .A4(n5324), .ZN(n9241)
         );
  AOI22_X1 U6924 ( .A1(n9691), .A2(n5615), .B1(n5569), .B2(n9241), .ZN(n5328)
         );
  XNOR2_X1 U6925 ( .A(n5328), .B(n4985), .ZN(n5330) );
  AOI22_X1 U6926 ( .A1(n9691), .A2(n5569), .B1(n5036), .B2(n9241), .ZN(n8817)
         );
  NAND2_X1 U6927 ( .A1(n5331), .A2(n5330), .ZN(n8815) );
  NAND2_X1 U6928 ( .A1(n5332), .A2(n8815), .ZN(n5353) );
  INV_X1 U6929 ( .A(n5353), .ZN(n5351) );
  MUX2_X1 U6930 ( .A(n7031), .B(n5336), .S(n4317), .Z(n5355) );
  XNOR2_X1 U6931 ( .A(n5355), .B(SI_15_), .ZN(n5354) );
  XNOR2_X1 U6932 ( .A(n5359), .B(n5354), .ZN(n7008) );
  NAND2_X1 U6933 ( .A1(n7008), .A2(n9080), .ZN(n5340) );
  NAND2_X1 U6934 ( .A1(n5360), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5338) );
  XNOR2_X1 U6935 ( .A(n5338), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9857) );
  AOI22_X1 U6936 ( .A1(n9857), .A2(n5440), .B1(n5037), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6937 ( .A1(n5342), .A2(n5341), .ZN(n5343) );
  AND2_X1 U6938 ( .A1(n5370), .A2(n5343), .ZN(n8970) );
  NAND2_X1 U6939 ( .A1(n5700), .A2(n8970), .ZN(n5348) );
  NAND2_X1 U6940 ( .A1(n6613), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5347) );
  INV_X1 U6941 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9852) );
  OR2_X1 U6942 ( .A1(n4312), .A2(n9852), .ZN(n5346) );
  INV_X1 U6943 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n5344) );
  OR2_X1 U6944 ( .A1(n5059), .A2(n5344), .ZN(n5345) );
  NAND4_X1 U6945 ( .A1(n5348), .A2(n5347), .A3(n5346), .A4(n5345), .ZN(n9240)
         );
  AOI22_X1 U6946 ( .A1(n8981), .A2(n5615), .B1(n5569), .B2(n9240), .ZN(n5349)
         );
  XNOR2_X1 U6947 ( .A(n5349), .B(n4985), .ZN(n5352) );
  INV_X1 U6948 ( .A(n5352), .ZN(n5350) );
  AOI22_X1 U6949 ( .A1(n8981), .A2(n5569), .B1(n5036), .B2(n9240), .ZN(n8961)
         );
  INV_X1 U6950 ( .A(n5354), .ZN(n5358) );
  INV_X1 U6951 ( .A(n5355), .ZN(n5356) );
  NAND2_X1 U6952 ( .A1(n5356), .A2(SI_15_), .ZN(n5357) );
  MUX2_X1 U6953 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n4518), .Z(n5383) );
  XNOR2_X1 U6954 ( .A(n5383), .B(SI_16_), .ZN(n5381) );
  NAND2_X1 U6955 ( .A1(n7176), .A2(n9080), .ZN(n5367) );
  NAND2_X1 U6956 ( .A1(n5361), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5364) );
  INV_X1 U6957 ( .A(n5364), .ZN(n5362) );
  NAND2_X1 U6958 ( .A1(n5362), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n5365) );
  INV_X1 U6959 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5363) );
  NAND2_X1 U6960 ( .A1(n5364), .A2(n5363), .ZN(n5392) );
  AOI22_X1 U6961 ( .A1(n9870), .A2(n5440), .B1(n5037), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U6962 ( .A1(n9687), .A2(n5615), .ZN(n5379) );
  INV_X1 U6963 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9338) );
  INV_X1 U6964 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5369) );
  NAND2_X1 U6965 ( .A1(n5370), .A2(n5369), .ZN(n5371) );
  NAND2_X1 U6966 ( .A1(n5398), .A2(n5371), .ZN(n7678) );
  OR2_X1 U6967 ( .A1(n7678), .A2(n5010), .ZN(n5377) );
  INV_X1 U6968 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9318) );
  OR2_X1 U6969 ( .A1(n4313), .A2(n9318), .ZN(n5375) );
  INV_X1 U6970 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n5372) );
  OR2_X1 U6971 ( .A1(n5373), .A2(n5372), .ZN(n5374) );
  AND2_X1 U6972 ( .A1(n5375), .A2(n5374), .ZN(n5376) );
  OAI211_X1 U6973 ( .C1(n5651), .C2(n9338), .A(n5377), .B(n5376), .ZN(n9562)
         );
  NAND2_X1 U6974 ( .A1(n9562), .A2(n5569), .ZN(n5378) );
  NAND2_X1 U6975 ( .A1(n5379), .A2(n5378), .ZN(n5380) );
  XNOR2_X1 U6976 ( .A(n5380), .B(n4985), .ZN(n5406) );
  AOI22_X1 U6977 ( .A1(n9687), .A2(n5569), .B1(n5036), .B2(n9562), .ZN(n5407)
         );
  XNOR2_X1 U6978 ( .A(n5406), .B(n5407), .ZN(n8883) );
  NAND2_X1 U6979 ( .A1(n5383), .A2(SI_16_), .ZN(n5384) );
  MUX2_X1 U6980 ( .A(n5387), .B(n5386), .S(n4518), .Z(n5389) );
  INV_X1 U6981 ( .A(n5389), .ZN(n5390) );
  NAND2_X1 U6982 ( .A1(n5390), .A2(SI_17_), .ZN(n5391) );
  NAND2_X1 U6983 ( .A1(n5416), .A2(n5391), .ZN(n5414) );
  NAND2_X1 U6984 ( .A1(n7196), .A2(n9080), .ZN(n5395) );
  NAND2_X1 U6985 ( .A1(n5392), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5393) );
  XNOR2_X1 U6986 ( .A(n5393), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9882) );
  AOI22_X1 U6987 ( .A1(n9882), .A2(n5440), .B1(n5037), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n5394) );
  NAND2_X1 U6988 ( .A1(n9574), .A2(n5615), .ZN(n5403) );
  INV_X1 U6989 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9683) );
  INV_X1 U6990 ( .A(n5398), .ZN(n5396) );
  INV_X1 U6991 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6992 ( .A1(n5398), .A2(n5397), .ZN(n5399) );
  NAND2_X1 U6993 ( .A1(n5425), .A2(n5399), .ZN(n9575) );
  OR2_X1 U6994 ( .A1(n9575), .A2(n5010), .ZN(n5401) );
  INV_X1 U6995 ( .A(n5059), .ZN(n5427) );
  AOI22_X1 U6996 ( .A1(n5427), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n6613), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n5400) );
  OAI211_X1 U6997 ( .C1(n4313), .C2(n9683), .A(n5401), .B(n5400), .ZN(n9239)
         );
  NAND2_X1 U6998 ( .A1(n9239), .A2(n5569), .ZN(n5402) );
  NAND2_X1 U6999 ( .A1(n5403), .A2(n5402), .ZN(n5404) );
  XNOR2_X1 U7000 ( .A(n5404), .B(n5710), .ZN(n5412) );
  AND2_X1 U7001 ( .A1(n9239), .A2(n5036), .ZN(n5405) );
  AOI21_X1 U7002 ( .B1(n9574), .B2(n5569), .A(n5405), .ZN(n5410) );
  XNOR2_X1 U7003 ( .A(n5412), .B(n5410), .ZN(n8891) );
  INV_X1 U7004 ( .A(n5406), .ZN(n5408) );
  NAND2_X1 U7005 ( .A1(n5408), .A2(n5407), .ZN(n8892) );
  INV_X1 U7006 ( .A(n5410), .ZN(n5411) );
  NAND2_X1 U7007 ( .A1(n5412), .A2(n5411), .ZN(n5413) );
  MUX2_X1 U7008 ( .A(n7294), .B(n5417), .S(n4518), .Z(n5432) );
  XNOR2_X1 U7009 ( .A(n5432), .B(SI_18_), .ZN(n5431) );
  XNOR2_X1 U7010 ( .A(n5435), .B(n5431), .ZN(n7222) );
  NAND2_X1 U7011 ( .A1(n7222), .A2(n9080), .ZN(n5424) );
  INV_X1 U7012 ( .A(n5418), .ZN(n5419) );
  NAND2_X1 U7013 ( .A1(n5419), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5420) );
  MUX2_X1 U7014 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5420), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n5421) );
  AND2_X1 U7015 ( .A1(n5422), .A2(n5421), .ZN(n9900) );
  AOI22_X1 U7016 ( .A1(n5037), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5440), .B2(
        n9900), .ZN(n5423) );
  NAND2_X1 U7017 ( .A1(n5425), .A2(n8942), .ZN(n5426) );
  NAND2_X1 U7018 ( .A1(n5461), .A2(n5426), .ZN(n9549) );
  AOI22_X1 U7019 ( .A1(n5701), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n6613), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U7020 ( .A1(n5427), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5428) );
  OAI211_X1 U7021 ( .C1(n9549), .C2(n5010), .A(n5429), .B(n5428), .ZN(n9565)
         );
  AOI22_X1 U7022 ( .A1(n9677), .A2(n5569), .B1(n5036), .B2(n9565), .ZN(n8941)
         );
  AOI22_X1 U7023 ( .A1(n9677), .A2(n5615), .B1(n5569), .B2(n9565), .ZN(n5430)
         );
  XNOR2_X1 U7024 ( .A(n5430), .B(n5710), .ZN(n8838) );
  INV_X1 U7025 ( .A(n5431), .ZN(n5434) );
  INV_X1 U7026 ( .A(n5432), .ZN(n5433) );
  MUX2_X1 U7027 ( .A(n7391), .B(n7393), .S(n4518), .Z(n5437) );
  INV_X1 U7028 ( .A(SI_19_), .ZN(n5436) );
  NAND2_X1 U7029 ( .A1(n5437), .A2(n5436), .ZN(n5452) );
  INV_X1 U7030 ( .A(n5437), .ZN(n5438) );
  NAND2_X1 U7031 ( .A1(n5438), .A2(SI_19_), .ZN(n5439) );
  NAND2_X1 U7032 ( .A1(n5452), .A2(n5439), .ZN(n5453) );
  XNOR2_X1 U7033 ( .A(n5454), .B(n5453), .ZN(n7390) );
  NAND2_X1 U7034 ( .A1(n7390), .A2(n9080), .ZN(n5442) );
  AOI22_X1 U7035 ( .A1(n5037), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9347), .B2(
        n5440), .ZN(n5441) );
  NAND2_X1 U7036 ( .A1(n9531), .A2(n5615), .ZN(n5449) );
  XNOR2_X1 U7037 ( .A(n5461), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n9532) );
  NAND2_X1 U7038 ( .A1(n9532), .A2(n5700), .ZN(n5447) );
  INV_X1 U7039 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9340) );
  NAND2_X1 U7040 ( .A1(n6613), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U7041 ( .A1(n5701), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5443) );
  OAI211_X1 U7042 ( .C1(n5651), .C2(n9340), .A(n5444), .B(n5443), .ZN(n5445)
         );
  INV_X1 U7043 ( .A(n5445), .ZN(n5446) );
  NAND2_X1 U7044 ( .A1(n5447), .A2(n5446), .ZN(n9238) );
  NAND2_X1 U7045 ( .A1(n9238), .A2(n5569), .ZN(n5448) );
  NAND2_X1 U7046 ( .A1(n5449), .A2(n5448), .ZN(n5450) );
  XNOR2_X1 U7047 ( .A(n5450), .B(n5628), .ZN(n5471) );
  AND2_X1 U7048 ( .A1(n9238), .A2(n5036), .ZN(n5451) );
  AOI21_X1 U7049 ( .B1(n9531), .B2(n5569), .A(n5451), .ZN(n5472) );
  AND2_X1 U7050 ( .A1(n5471), .A2(n5472), .ZN(n8839) );
  MUX2_X1 U7051 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n4518), .Z(n5478) );
  XNOR2_X1 U7052 ( .A(n5478), .B(n5480), .ZN(n5455) );
  XNOR2_X1 U7053 ( .A(n5481), .B(n5455), .ZN(n7440) );
  NAND2_X1 U7054 ( .A1(n7440), .A2(n9080), .ZN(n5457) );
  NAND2_X1 U7055 ( .A1(n5037), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5456) );
  AND2_X1 U7056 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5458) );
  INV_X1 U7057 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8842) );
  INV_X1 U7058 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5460) );
  OAI21_X1 U7059 ( .B1(n5461), .B2(n8842), .A(n5460), .ZN(n5462) );
  NAND2_X1 U7060 ( .A1(n5487), .A2(n5462), .ZN(n9513) );
  OR2_X1 U7061 ( .A1(n9513), .A2(n5010), .ZN(n5467) );
  INV_X1 U7062 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9514) );
  NAND2_X1 U7063 ( .A1(n5701), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U7064 ( .A1(n6613), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5463) );
  OAI211_X1 U7065 ( .C1(n9514), .C2(n5059), .A(n5464), .B(n5463), .ZN(n5465)
         );
  INV_X1 U7066 ( .A(n5465), .ZN(n5466) );
  NAND2_X1 U7067 ( .A1(n5467), .A2(n5466), .ZN(n9525) );
  AOI22_X1 U7068 ( .A1(n9512), .A2(n5615), .B1(n5569), .B2(n9525), .ZN(n5468)
         );
  XNOR2_X1 U7069 ( .A(n5468), .B(n5710), .ZN(n5470) );
  AOI22_X1 U7070 ( .A1(n9512), .A2(n5569), .B1(n5036), .B2(n9525), .ZN(n5469)
         );
  NAND2_X1 U7071 ( .A1(n5470), .A2(n5469), .ZN(n5477) );
  OAI21_X1 U7072 ( .B1(n5470), .B2(n5469), .A(n5477), .ZN(n8923) );
  INV_X1 U7073 ( .A(n8923), .ZN(n5476) );
  INV_X1 U7074 ( .A(n5471), .ZN(n5474) );
  INV_X1 U7075 ( .A(n5472), .ZN(n5473) );
  INV_X1 U7076 ( .A(n8924), .ZN(n5475) );
  NAND2_X1 U7077 ( .A1(n8922), .A2(n4905), .ZN(n8926) );
  NAND2_X1 U7078 ( .A1(n8926), .A2(n5477), .ZN(n8863) );
  INV_X1 U7079 ( .A(n5478), .ZN(n5479) );
  OAI21_X1 U7080 ( .B1(n5481), .B2(n5480), .A(n5479), .ZN(n5483) );
  NAND2_X1 U7081 ( .A1(n5481), .A2(n5480), .ZN(n5482) );
  NAND2_X1 U7082 ( .A1(n5483), .A2(n5482), .ZN(n5506) );
  MUX2_X1 U7083 ( .A(n8239), .B(n8221), .S(n4518), .Z(n5502) );
  XNOR2_X1 U7084 ( .A(n5502), .B(SI_21_), .ZN(n5484) );
  XNOR2_X1 U7085 ( .A(n5506), .B(n5484), .ZN(n7501) );
  NAND2_X1 U7086 ( .A1(n7501), .A2(n9080), .ZN(n5486) );
  NAND2_X1 U7087 ( .A1(n5037), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U7088 ( .A1(n9495), .A2(n5615), .ZN(n5496) );
  NAND2_X1 U7089 ( .A1(n5487), .A2(n8868), .ZN(n5488) );
  AND2_X1 U7090 ( .A1(n5515), .A2(n5488), .ZN(n9496) );
  NAND2_X1 U7091 ( .A1(n9496), .A2(n5700), .ZN(n5494) );
  INV_X1 U7092 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U7093 ( .A1(n5701), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U7094 ( .A1(n6613), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5489) );
  OAI211_X1 U7095 ( .C1(n5491), .C2(n5059), .A(n5490), .B(n5489), .ZN(n5492)
         );
  INV_X1 U7096 ( .A(n5492), .ZN(n5493) );
  NAND2_X1 U7097 ( .A1(n5494), .A2(n5493), .ZN(n9237) );
  NAND2_X1 U7098 ( .A1(n9237), .A2(n5569), .ZN(n5495) );
  NAND2_X1 U7099 ( .A1(n5496), .A2(n5495), .ZN(n5497) );
  XNOR2_X1 U7100 ( .A(n5497), .B(n5710), .ZN(n5498) );
  AOI22_X1 U7101 ( .A1(n9495), .A2(n5569), .B1(n5036), .B2(n9237), .ZN(n5499)
         );
  XNOR2_X1 U7102 ( .A(n5498), .B(n5499), .ZN(n8865) );
  NAND2_X1 U7103 ( .A1(n8863), .A2(n8865), .ZN(n8864) );
  INV_X1 U7104 ( .A(n5498), .ZN(n5500) );
  NAND2_X1 U7105 ( .A1(n5500), .A2(n5499), .ZN(n5501) );
  NAND2_X1 U7106 ( .A1(n8864), .A2(n5501), .ZN(n5526) );
  INV_X1 U7107 ( .A(n5526), .ZN(n5524) );
  NOR2_X1 U7108 ( .A1(n5503), .A2(SI_21_), .ZN(n5505) );
  NAND2_X1 U7109 ( .A1(n5503), .A2(SI_21_), .ZN(n5504) );
  MUX2_X1 U7110 ( .A(n7581), .B(n7711), .S(n4518), .Z(n5508) );
  NAND2_X1 U7111 ( .A1(n5508), .A2(n5507), .ZN(n5528) );
  INV_X1 U7112 ( .A(n5508), .ZN(n5509) );
  NAND2_X1 U7113 ( .A1(n5509), .A2(SI_22_), .ZN(n5510) );
  NAND2_X1 U7114 ( .A1(n5528), .A2(n5510), .ZN(n5529) );
  XNOR2_X1 U7115 ( .A(n5530), .B(n5529), .ZN(n7579) );
  NAND2_X1 U7116 ( .A1(n7579), .A2(n9080), .ZN(n5512) );
  NAND2_X1 U7117 ( .A1(n5037), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5511) );
  INV_X1 U7118 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U7119 ( .A1(n5515), .A2(n5514), .ZN(n5516) );
  NAND2_X1 U7120 ( .A1(n5538), .A2(n5516), .ZN(n9479) );
  OR2_X1 U7121 ( .A1(n9479), .A2(n5010), .ZN(n5521) );
  INV_X1 U7122 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9480) );
  NAND2_X1 U7123 ( .A1(n5701), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5518) );
  NAND2_X1 U7124 ( .A1(n6613), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5517) );
  OAI211_X1 U7125 ( .C1(n9480), .C2(n5651), .A(n5518), .B(n5517), .ZN(n5519)
         );
  INV_X1 U7126 ( .A(n5519), .ZN(n5520) );
  NAND2_X1 U7127 ( .A1(n5521), .A2(n5520), .ZN(n9236) );
  AOI22_X1 U7128 ( .A1(n9484), .A2(n5615), .B1(n5569), .B2(n9236), .ZN(n5522)
         );
  XNOR2_X1 U7129 ( .A(n5522), .B(n5710), .ZN(n5525) );
  INV_X1 U7130 ( .A(n5525), .ZN(n5523) );
  NAND2_X1 U7131 ( .A1(n5524), .A2(n5523), .ZN(n5527) );
  INV_X1 U7132 ( .A(n9236), .ZN(n6554) );
  OAI22_X1 U7133 ( .A1(n9731), .A2(n5200), .B1(n6554), .B2(n5657), .ZN(n8933)
         );
  INV_X1 U7134 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7640) );
  INV_X1 U7135 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5531) );
  MUX2_X1 U7136 ( .A(n7640), .B(n5531), .S(n4518), .Z(n5533) );
  INV_X1 U7137 ( .A(SI_23_), .ZN(n5532) );
  NAND2_X1 U7138 ( .A1(n5533), .A2(n5532), .ZN(n5556) );
  INV_X1 U7139 ( .A(n5533), .ZN(n5534) );
  NAND2_X1 U7140 ( .A1(n5534), .A2(SI_23_), .ZN(n5535) );
  NAND2_X1 U7141 ( .A1(n7637), .A2(n9080), .ZN(n5537) );
  NAND2_X1 U7142 ( .A1(n5037), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U7143 ( .A1(n9462), .A2(n5615), .ZN(n5546) );
  INV_X1 U7144 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8833) );
  NAND2_X1 U7145 ( .A1(n5538), .A2(n8833), .ZN(n5539) );
  NAND2_X1 U7146 ( .A1(n5594), .A2(n5539), .ZN(n9464) );
  OR2_X1 U7147 ( .A1(n9464), .A2(n5010), .ZN(n5544) );
  INV_X1 U7148 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9463) );
  NAND2_X1 U7149 ( .A1(n6613), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7150 ( .A1(n5701), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5540) );
  OAI211_X1 U7151 ( .C1(n9463), .C2(n5651), .A(n5541), .B(n5540), .ZN(n5542)
         );
  INV_X1 U7152 ( .A(n5542), .ZN(n5543) );
  NAND2_X1 U7153 ( .A1(n5544), .A2(n5543), .ZN(n9448) );
  NAND2_X1 U7154 ( .A1(n9448), .A2(n5569), .ZN(n5545) );
  NAND2_X1 U7155 ( .A1(n5546), .A2(n5545), .ZN(n5547) );
  XNOR2_X1 U7156 ( .A(n5547), .B(n5628), .ZN(n5549) );
  AND2_X1 U7157 ( .A1(n9448), .A2(n5036), .ZN(n5548) );
  AOI21_X1 U7158 ( .B1(n9462), .B2(n5569), .A(n5548), .ZN(n5550) );
  NAND2_X1 U7159 ( .A1(n5549), .A2(n5550), .ZN(n8901) );
  INV_X1 U7160 ( .A(n5549), .ZN(n5552) );
  INV_X1 U7161 ( .A(n5550), .ZN(n5551) );
  NAND2_X1 U7162 ( .A1(n5552), .A2(n5551), .ZN(n5553) );
  INV_X1 U7163 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7686) );
  MUX2_X1 U7164 ( .A(n7688), .B(n7686), .S(n4518), .Z(n5558) );
  INV_X1 U7165 ( .A(SI_24_), .ZN(n5557) );
  NAND2_X1 U7166 ( .A1(n5558), .A2(n5557), .ZN(n5583) );
  INV_X1 U7167 ( .A(n5558), .ZN(n5559) );
  NAND2_X1 U7168 ( .A1(n5559), .A2(SI_24_), .ZN(n5560) );
  XNOR2_X1 U7169 ( .A(n5582), .B(n5581), .ZN(n7685) );
  NAND2_X1 U7170 ( .A1(n7685), .A2(n9080), .ZN(n5562) );
  NAND2_X1 U7171 ( .A1(n5037), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U7172 ( .A1(n9645), .A2(n5615), .ZN(n5571) );
  XNOR2_X1 U7173 ( .A(n5594), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n9453) );
  NAND2_X1 U7174 ( .A1(n9453), .A2(n5700), .ZN(n5568) );
  INV_X1 U7175 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U7176 ( .A1(n6613), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7177 ( .A1(n5701), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5563) );
  OAI211_X1 U7178 ( .C1(n5059), .C2(n5565), .A(n5564), .B(n5563), .ZN(n5566)
         );
  INV_X1 U7179 ( .A(n5566), .ZN(n5567) );
  NAND2_X1 U7180 ( .A1(n5568), .A2(n5567), .ZN(n9235) );
  NAND2_X1 U7181 ( .A1(n9235), .A2(n5569), .ZN(n5570) );
  NAND2_X1 U7182 ( .A1(n5571), .A2(n5570), .ZN(n5572) );
  XNOR2_X1 U7183 ( .A(n5572), .B(n5628), .ZN(n5574) );
  AND2_X1 U7184 ( .A1(n9235), .A2(n5036), .ZN(n5573) );
  AOI21_X1 U7185 ( .B1(n9645), .B2(n5569), .A(n5573), .ZN(n5575) );
  NAND2_X1 U7186 ( .A1(n5574), .A2(n5575), .ZN(n5580) );
  INV_X1 U7187 ( .A(n5574), .ZN(n5577) );
  INV_X1 U7188 ( .A(n5575), .ZN(n5576) );
  NAND2_X1 U7189 ( .A1(n5577), .A2(n5576), .ZN(n5578) );
  NAND2_X1 U7190 ( .A1(n5579), .A2(n8899), .ZN(n8898) );
  NAND2_X1 U7191 ( .A1(n5582), .A2(n5581), .ZN(n5584) );
  INV_X1 U7192 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7691) );
  MUX2_X1 U7193 ( .A(n7691), .B(n7692), .S(n4518), .Z(n5586) );
  INV_X1 U7194 ( .A(SI_25_), .ZN(n5585) );
  NAND2_X1 U7195 ( .A1(n5586), .A2(n5585), .ZN(n5607) );
  INV_X1 U7196 ( .A(n5586), .ZN(n5587) );
  NAND2_X1 U7197 ( .A1(n5587), .A2(SI_25_), .ZN(n5588) );
  XNOR2_X1 U7198 ( .A(n5606), .B(n5605), .ZN(n7690) );
  NAND2_X1 U7199 ( .A1(n7690), .A2(n9080), .ZN(n5590) );
  NAND2_X1 U7200 ( .A1(n5037), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U7201 ( .A1(n9436), .A2(n5615), .ZN(n5603) );
  NAND2_X1 U7202 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n5591) );
  INV_X1 U7203 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5593) );
  INV_X1 U7204 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5592) );
  OAI21_X1 U7205 ( .B1(n5594), .B2(n5593), .A(n5592), .ZN(n5595) );
  AND2_X1 U7206 ( .A1(n5618), .A2(n5595), .ZN(n9437) );
  NAND2_X1 U7207 ( .A1(n9437), .A2(n5700), .ZN(n5601) );
  INV_X1 U7208 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U7209 ( .A1(n6613), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U7210 ( .A1(n5701), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5596) );
  OAI211_X1 U7211 ( .C1(n5598), .C2(n5059), .A(n5597), .B(n5596), .ZN(n5599)
         );
  INV_X1 U7212 ( .A(n5599), .ZN(n5600) );
  NAND2_X1 U7213 ( .A1(n9449), .A2(n4987), .ZN(n5602) );
  NAND2_X1 U7214 ( .A1(n5603), .A2(n5602), .ZN(n5604) );
  XNOR2_X1 U7215 ( .A(n5604), .B(n5710), .ZN(n5633) );
  AOI22_X1 U7216 ( .A1(n9436), .A2(n5569), .B1(n5036), .B2(n9449), .ZN(n5631)
         );
  XNOR2_X1 U7217 ( .A(n5633), .B(n5631), .ZN(n8874) );
  NAND2_X1 U7218 ( .A1(n5606), .A2(n5605), .ZN(n5608) );
  INV_X1 U7219 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8801) );
  INV_X1 U7220 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9767) );
  MUX2_X1 U7221 ( .A(n8801), .B(n9767), .S(n4518), .Z(n5610) );
  INV_X1 U7222 ( .A(SI_26_), .ZN(n5609) );
  NAND2_X1 U7223 ( .A1(n5610), .A2(n5609), .ZN(n5637) );
  INV_X1 U7224 ( .A(n5610), .ZN(n5611) );
  NAND2_X1 U7225 ( .A1(n5611), .A2(SI_26_), .ZN(n5612) );
  XNOR2_X1 U7226 ( .A(n5636), .B(n5635), .ZN(n8799) );
  NAND2_X1 U7227 ( .A1(n8799), .A2(n9080), .ZN(n5614) );
  NAND2_X1 U7228 ( .A1(n5037), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7229 ( .A1(n9417), .A2(n5615), .ZN(n5627) );
  INV_X1 U7230 ( .A(n5618), .ZN(n5616) );
  NAND2_X1 U7231 ( .A1(n5616), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5647) );
  INV_X1 U7232 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U7233 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  AND2_X1 U7234 ( .A1(n5647), .A2(n5619), .ZN(n9418) );
  NAND2_X1 U7235 ( .A1(n9418), .A2(n5700), .ZN(n5625) );
  INV_X1 U7236 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U7237 ( .A1(n6613), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U7238 ( .A1(n5701), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5620) );
  OAI211_X1 U7239 ( .C1(n5622), .C2(n5651), .A(n5621), .B(n5620), .ZN(n5623)
         );
  INV_X1 U7240 ( .A(n5623), .ZN(n5624) );
  NAND2_X1 U7241 ( .A1(n5625), .A2(n5624), .ZN(n9234) );
  NAND2_X1 U7242 ( .A1(n9234), .A2(n4987), .ZN(n5626) );
  NAND2_X1 U7243 ( .A1(n5627), .A2(n5626), .ZN(n5629) );
  XNOR2_X1 U7244 ( .A(n5629), .B(n5628), .ZN(n5660) );
  AND2_X1 U7245 ( .A1(n9234), .A2(n5036), .ZN(n5630) );
  AOI21_X1 U7246 ( .B1(n9417), .B2(n5569), .A(n5630), .ZN(n5661) );
  XNOR2_X1 U7247 ( .A(n5660), .B(n5661), .ZN(n8948) );
  INV_X1 U7248 ( .A(n5631), .ZN(n5632) );
  NOR2_X1 U7249 ( .A1(n5633), .A2(n5632), .ZN(n8949) );
  NOR2_X1 U7250 ( .A1(n8948), .A2(n8949), .ZN(n5634) );
  NAND2_X1 U7251 ( .A1(n5636), .A2(n5635), .ZN(n5638) );
  INV_X1 U7252 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8798) );
  INV_X1 U7253 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9765) );
  MUX2_X1 U7254 ( .A(n8798), .B(n9765), .S(n4518), .Z(n5640) );
  INV_X1 U7255 ( .A(SI_27_), .ZN(n5639) );
  NAND2_X1 U7256 ( .A1(n5640), .A2(n5639), .ZN(n5697) );
  INV_X1 U7257 ( .A(n5640), .ZN(n5641) );
  NAND2_X1 U7258 ( .A1(n5641), .A2(SI_27_), .ZN(n5642) );
  NAND2_X1 U7259 ( .A1(n9762), .A2(n9080), .ZN(n5644) );
  NAND2_X1 U7260 ( .A1(n5037), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5643) );
  INV_X1 U7261 ( .A(n5647), .ZN(n5645) );
  NAND2_X1 U7262 ( .A1(n5645), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9368) );
  INV_X1 U7263 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U7264 ( .A1(n5647), .A2(n5646), .ZN(n5648) );
  NAND2_X1 U7265 ( .A1(n9368), .A2(n5648), .ZN(n8810) );
  INV_X1 U7266 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U7267 ( .A1(n6613), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U7268 ( .A1(n5701), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5649) );
  OAI211_X1 U7269 ( .C1(n5652), .C2(n5651), .A(n5650), .B(n5649), .ZN(n5653)
         );
  INV_X1 U7270 ( .A(n5653), .ZN(n5654) );
  NAND2_X1 U7271 ( .A1(n5655), .A2(n5654), .ZN(n9233) );
  AOI22_X1 U7272 ( .A1(n9402), .A2(n5615), .B1(n5569), .B2(n9233), .ZN(n5656)
         );
  XOR2_X1 U7273 ( .A(n5710), .B(n5656), .Z(n5659) );
  OAI22_X1 U7274 ( .A1(n9715), .A2(n5200), .B1(n6532), .B2(n5657), .ZN(n5658)
         );
  NOR2_X1 U7275 ( .A1(n5659), .A2(n5658), .ZN(n5734) );
  AOI21_X1 U7276 ( .B1(n5659), .B2(n5658), .A(n5734), .ZN(n8805) );
  INV_X1 U7277 ( .A(n8805), .ZN(n5665) );
  INV_X1 U7278 ( .A(n5660), .ZN(n5663) );
  INV_X1 U7279 ( .A(n5661), .ZN(n5662) );
  NAND2_X1 U7280 ( .A1(n5663), .A2(n5662), .ZN(n8806) );
  INV_X1 U7281 ( .A(n8806), .ZN(n5664) );
  NOR2_X1 U7282 ( .A1(n5665), .A2(n5664), .ZN(n5666) );
  NAND2_X1 U7283 ( .A1(n5672), .A2(n5671), .ZN(n5668) );
  NAND2_X1 U7284 ( .A1(n5668), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5670) );
  XNOR2_X1 U7285 ( .A(n5670), .B(n5669), .ZN(n7694) );
  XNOR2_X1 U7286 ( .A(n5672), .B(n5671), .ZN(n7687) );
  NAND3_X1 U7287 ( .A1(n7694), .A2(P1_B_REG_SCAN_IN), .A3(n7687), .ZN(n5675)
         );
  INV_X1 U7288 ( .A(n7687), .ZN(n5673) );
  INV_X1 U7289 ( .A(P1_B_REG_SCAN_IN), .ZN(n8222) );
  NAND2_X1 U7290 ( .A1(n7687), .A2(n9770), .ZN(n9755) );
  OR2_X1 U7291 ( .A1(n9753), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U7292 ( .A1(n7694), .A2(n9770), .ZN(n9754) );
  NOR2_X1 U7293 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n5681) );
  NOR4_X1 U7294 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5680) );
  NOR4_X1 U7295 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5679) );
  NOR4_X1 U7296 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5678) );
  NAND4_X1 U7297 ( .A1(n5681), .A2(n5680), .A3(n5679), .A4(n5678), .ZN(n5687)
         );
  NOR4_X1 U7298 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5685) );
  NOR4_X1 U7299 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5684) );
  NOR4_X1 U7300 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5683) );
  NOR4_X1 U7301 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5682) );
  NAND4_X1 U7302 ( .A1(n5685), .A2(n5684), .A3(n5683), .A4(n5682), .ZN(n5686)
         );
  NOR2_X1 U7303 ( .A1(n5687), .A2(n5686), .ZN(n5688) );
  OR2_X1 U7304 ( .A1(n9753), .A2(n5688), .ZN(n6749) );
  NAND3_X1 U7305 ( .A1(n6579), .A2(n6751), .A3(n6749), .ZN(n5726) );
  NAND2_X1 U7306 ( .A1(n5689), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5691) );
  INV_X1 U7307 ( .A(n9949), .ZN(n9939) );
  INV_X1 U7308 ( .A(n9212), .ZN(n5693) );
  AND2_X1 U7309 ( .A1(n9939), .A2(n5693), .ZN(n5694) );
  INV_X1 U7310 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7986) );
  MUX2_X1 U7311 ( .A(n8794), .B(n7986), .S(n4518), .Z(n6461) );
  XNOR2_X1 U7312 ( .A(n6461), .B(SI_28_), .ZN(n6458) );
  NAND2_X1 U7313 ( .A1(n8791), .A2(n9080), .ZN(n5699) );
  NAND2_X1 U7314 ( .A1(n5037), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5698) );
  NAND2_X1 U7315 ( .A1(n9387), .A2(n4987), .ZN(n5709) );
  XNOR2_X1 U7316 ( .A(n9368), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U7317 ( .A1(n9386), .A2(n5700), .ZN(n5707) );
  INV_X1 U7318 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U7319 ( .A1(n6613), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U7320 ( .A1(n5701), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5702) );
  OAI211_X1 U7321 ( .C1(n5704), .C2(n5059), .A(n5703), .B(n5702), .ZN(n5705)
         );
  INV_X1 U7322 ( .A(n5705), .ZN(n5706) );
  NAND2_X1 U7323 ( .A1(n5707), .A2(n5706), .ZN(n9232) );
  NAND2_X1 U7324 ( .A1(n9232), .A2(n5036), .ZN(n5708) );
  NAND2_X1 U7325 ( .A1(n5709), .A2(n5708), .ZN(n5711) );
  XNOR2_X1 U7326 ( .A(n5711), .B(n5710), .ZN(n5713) );
  AOI22_X1 U7327 ( .A1(n9387), .A2(n5615), .B1(n5569), .B2(n9232), .ZN(n5712)
         );
  XNOR2_X1 U7328 ( .A(n5713), .B(n5712), .ZN(n5736) );
  NAND3_X1 U7329 ( .A1(n8807), .A2(n9806), .A3(n5736), .ZN(n5740) );
  INV_X1 U7330 ( .A(n6572), .ZN(n6685) );
  OR2_X1 U7331 ( .A1(n6685), .A2(n9126), .ZN(n6754) );
  INV_X1 U7332 ( .A(n6754), .ZN(n5714) );
  NAND2_X1 U7333 ( .A1(n5724), .A2(n5714), .ZN(n5715) );
  INV_X1 U7334 ( .A(n6611), .ZN(n9752) );
  NAND3_X1 U7335 ( .A1(n9752), .A2(n7514), .A3(n4316), .ZN(n9920) );
  INV_X1 U7336 ( .A(n5716), .ZN(n6649) );
  INV_X1 U7337 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9365) );
  OR2_X1 U7338 ( .A1(n5010), .A2(n9365), .ZN(n5717) );
  OR2_X1 U7339 ( .A1(n9368), .A2(n5717), .ZN(n5722) );
  INV_X1 U7340 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9366) );
  NAND2_X1 U7341 ( .A1(n6613), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5719) );
  INV_X1 U7342 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6577) );
  OR2_X1 U7343 ( .A1(n4313), .A2(n6577), .ZN(n5718) );
  OAI211_X1 U7344 ( .C1(n9366), .C2(n5059), .A(n5719), .B(n5718), .ZN(n5720)
         );
  INV_X1 U7345 ( .A(n5720), .ZN(n5721) );
  NAND2_X1 U7346 ( .A1(n5722), .A2(n5721), .ZN(n6819) );
  AOI22_X1 U7347 ( .A1(n9233), .A2(n9563), .B1(n4309), .B2(n6819), .ZN(n9378)
         );
  INV_X1 U7348 ( .A(n9194), .ZN(n5723) );
  NAND2_X1 U7349 ( .A1(n5724), .A2(n5723), .ZN(n8955) );
  NAND2_X1 U7350 ( .A1(n9949), .A2(n6754), .ZN(n5725) );
  NAND2_X1 U7351 ( .A1(n5726), .A2(n5725), .ZN(n5728) );
  NAND2_X1 U7352 ( .A1(n9212), .A2(n9194), .ZN(n5727) );
  AND3_X1 U7353 ( .A1(n5727), .A2(n6610), .A3(n4965), .ZN(n6748) );
  NAND2_X1 U7354 ( .A1(n5728), .A2(n6748), .ZN(n5729) );
  INV_X1 U7355 ( .A(n9810), .ZN(n8971) );
  AOI22_X1 U7356 ( .A1(n9386), .A2(n8971), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n5730) );
  OAI21_X1 U7357 ( .B1(n9378), .B2(n8955), .A(n5730), .ZN(n5731) );
  AOI21_X1 U7358 ( .B1(n9387), .B2(n8957), .A(n5731), .ZN(n5732) );
  INV_X1 U7359 ( .A(n5732), .ZN(n5733) );
  NAND3_X1 U7360 ( .A1(n5740), .A2(n5739), .A3(n5738), .ZN(P1_U3220) );
  NOR2_X2 U7361 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5741) );
  INV_X2 U7362 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7363 ( .A1(n4319), .A2(n4701), .ZN(n5824) );
  NAND2_X1 U7364 ( .A1(n6722), .A2(n7732), .ZN(n5763) );
  NAND2_X1 U7365 ( .A1(n5969), .A2(n5759), .ZN(n5787) );
  NAND2_X1 U7366 ( .A1(n5787), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7367 ( .A1(n5991), .A2(n5760), .ZN(n5977) );
  OR2_X1 U7368 ( .A1(n5991), .A2(n5760), .ZN(n5761) );
  AOI22_X1 U7369 ( .A1(n6073), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6342), .B2(
        n7655), .ZN(n5762) );
  NAND2_X1 U7370 ( .A1(n5763), .A2(n5762), .ZN(n8294) );
  NAND2_X1 U7371 ( .A1(n6162), .A2(n6163), .ZN(n5764) );
  XNOR2_X1 U7372 ( .A(n5775), .B(P2_B_REG_SCAN_IN), .ZN(n5770) );
  NAND2_X1 U7373 ( .A1(n5766), .A2(n5765), .ZN(n5767) );
  INV_X1 U7374 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5774) );
  INV_X1 U7375 ( .A(n6158), .ZN(n8802) );
  NAND2_X1 U7376 ( .A1(n5775), .A2(n8802), .ZN(n6691) );
  NAND2_X1 U7377 ( .A1(n5776), .A2(n6691), .ZN(n6142) );
  INV_X1 U7378 ( .A(n5778), .ZN(n5779) );
  NAND2_X1 U7379 ( .A1(n5779), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U7380 ( .A1(n5781), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5782) );
  MUX2_X1 U7381 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5782), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5783) );
  INV_X1 U7382 ( .A(n5783), .ZN(n5784) );
  NOR2_X1 U7383 ( .A1(n5784), .A2(n5778), .ZN(n6316) );
  NAND2_X1 U7384 ( .A1(n7749), .A2(n6316), .ZN(n7968) );
  NOR2_X1 U7385 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5989) );
  NAND4_X1 U7386 ( .A1(n5989), .A2(n5992), .A3(n6016), .A4(n5785), .ZN(n5786)
         );
  NAND2_X1 U7387 ( .A1(n6031), .A2(n5788), .ZN(n6046) );
  INV_X1 U7388 ( .A(n6046), .ZN(n5790) );
  INV_X1 U7389 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U7390 ( .A1(n5790), .A2(n5789), .ZN(n5791) );
  INV_X1 U7391 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U7392 ( .A1(n6061), .A2(n5792), .ZN(n5793) );
  INV_X1 U7393 ( .A(n6316), .ZN(n7441) );
  INV_X1 U7394 ( .A(n5797), .ZN(n5844) );
  XNOR2_X1 U7395 ( .A(n8294), .B(n8018), .ZN(n5975) );
  INV_X1 U7396 ( .A(n5975), .ZN(n5976) );
  INV_X1 U7397 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U7398 ( .A1(n5801), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5803) );
  INV_X1 U7399 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5802) );
  AND2_X2 U7400 ( .A1(n7707), .A2(n8789), .ZN(n5838) );
  INV_X2 U7401 ( .A(n6106), .ZN(n6475) );
  NAND2_X1 U7402 ( .A1(n6475), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5814) );
  AND2_X4 U7403 ( .A1(n5804), .A2(n5805), .ZN(n7718) );
  INV_X1 U7404 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7651) );
  OR2_X1 U7405 ( .A1(n5906), .A2(n7651), .ZN(n5813) );
  INV_X1 U7406 ( .A(n5804), .ZN(n5810) );
  NOR2_X1 U7407 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5871) );
  INV_X1 U7408 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5806) );
  NAND2_X1 U7409 ( .A1(n5871), .A2(n5806), .ZN(n5907) );
  NAND2_X1 U7410 ( .A1(n5937), .A2(n5808), .ZN(n5962) );
  NAND2_X1 U7411 ( .A1(n5964), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5809) );
  AND2_X1 U7412 ( .A1(n5982), .A2(n5809), .ZN(n7483) );
  OR2_X1 U7413 ( .A1(n6078), .A2(n7483), .ZN(n5812) );
  INV_X2 U7414 ( .A(n5854), .ZN(n5839) );
  INV_X1 U7415 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7643) );
  OR2_X1 U7416 ( .A1(n6309), .A2(n7643), .ZN(n5811) );
  INV_X1 U7417 ( .A(n7535), .ZN(n8338) );
  NAND2_X1 U7418 ( .A1(n5839), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U7419 ( .A1(n6087), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5817) );
  NAND2_X1 U7420 ( .A1(n7718), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U7421 ( .A1(n5838), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U7422 ( .A1(n4701), .A2(SI_0_), .ZN(n5820) );
  INV_X1 U7423 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U7424 ( .A1(n5820), .A2(n5819), .ZN(n5822) );
  AND2_X1 U7425 ( .A1(n5822), .A2(n5821), .ZN(n8804) );
  MUX2_X1 U7426 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8804), .S(n5830), .Z(n10053)
         );
  NAND2_X1 U7427 ( .A1(n6086), .A2(n6975), .ZN(n5823) );
  NAND2_X1 U7428 ( .A1(n7753), .A2(n5823), .ZN(n7003) );
  OR2_X1 U7429 ( .A1(n5879), .A2(n6595), .ZN(n5826) );
  OR2_X1 U7430 ( .A1(n5824), .A2(n6596), .ZN(n5825) );
  NAND2_X1 U7431 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5827) );
  MUX2_X1 U7432 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5827), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5829) );
  INV_X1 U7433 ( .A(n6373), .ZN(n5828) );
  OR2_X1 U7434 ( .A1(n4319), .A2(n4426), .ZN(n5831) );
  NAND2_X1 U7435 ( .A1(n5839), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5835) );
  NAND2_X1 U7436 ( .A1(n6087), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U7437 ( .A1(n7718), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U7438 ( .A1(n5838), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5832) );
  NAND4_X2 U7439 ( .A1(n5835), .A2(n5834), .A3(n5833), .A4(n5832), .ZN(n6206)
         );
  XNOR2_X1 U7440 ( .A(n5836), .B(n6206), .ZN(n7001) );
  NAND2_X1 U7441 ( .A1(n7003), .A2(n7001), .ZN(n7002) );
  INV_X1 U7442 ( .A(n8348), .ZN(n6981) );
  NAND2_X1 U7443 ( .A1(n5836), .A2(n6981), .ZN(n5837) );
  NAND2_X1 U7444 ( .A1(n7002), .A2(n5837), .ZN(n6976) );
  NAND2_X1 U7445 ( .A1(n5838), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U7446 ( .A1(n6087), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5841) );
  NAND4_X2 U7447 ( .A1(n5843), .A2(n5842), .A3(n5841), .A4(n5840), .ZN(n8346)
         );
  INV_X1 U7448 ( .A(n8346), .ZN(n5850) );
  INV_X1 U7449 ( .A(n5844), .ZN(n5859) );
  OR2_X1 U7450 ( .A1(n5879), .A2(n6604), .ZN(n5848) );
  OR2_X1 U7451 ( .A1(n5824), .A2(n6603), .ZN(n5847) );
  INV_X1 U7452 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5845) );
  XNOR2_X1 U7453 ( .A(n5859), .B(n10055), .ZN(n5849) );
  XNOR2_X1 U7454 ( .A(n5850), .B(n5849), .ZN(n6979) );
  NAND2_X1 U7455 ( .A1(n6976), .A2(n6979), .ZN(n6977) );
  INV_X1 U7456 ( .A(n5849), .ZN(n5851) );
  NAND2_X1 U7457 ( .A1(n5851), .A2(n5850), .ZN(n5852) );
  NAND2_X1 U7458 ( .A1(n6977), .A2(n5852), .ZN(n6985) );
  INV_X1 U7459 ( .A(n6985), .ZN(n5867) );
  INV_X1 U7460 ( .A(n7718), .ZN(n5906) );
  INV_X1 U7461 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5853) );
  NAND2_X1 U7462 ( .A1(n5838), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5857) );
  OR2_X1 U7463 ( .A1(n6078), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5856) );
  INV_X1 U7464 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7385) );
  OR2_X1 U7465 ( .A1(n5854), .A2(n7385), .ZN(n5855) );
  NAND2_X1 U7466 ( .A1(n5860), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5861) );
  MUX2_X1 U7467 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5861), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5863) );
  NAND2_X1 U7468 ( .A1(n5863), .A2(n5862), .ZN(n6861) );
  OR2_X1 U7469 ( .A1(n5879), .A2(n6601), .ZN(n5865) );
  OR2_X1 U7470 ( .A1(n5824), .A2(n6600), .ZN(n5864) );
  OAI211_X1 U7471 ( .C1(n5830), .C2(n6861), .A(n5865), .B(n5864), .ZN(n7387)
         );
  XNOR2_X1 U7472 ( .A(n5859), .B(n7387), .ZN(n5868) );
  XNOR2_X1 U7473 ( .A(n6268), .B(n5868), .ZN(n6988) );
  INV_X1 U7474 ( .A(n5868), .ZN(n5869) );
  NAND2_X1 U7475 ( .A1(n6209), .A2(n5869), .ZN(n5870) );
  NAND2_X1 U7476 ( .A1(n7718), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5876) );
  INV_X1 U7477 ( .A(n5871), .ZN(n5891) );
  NAND2_X1 U7478 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5872) );
  AND2_X1 U7479 ( .A1(n5891), .A2(n5872), .ZN(n7333) );
  OR2_X1 U7480 ( .A1(n6078), .A2(n7333), .ZN(n5875) );
  NAND2_X1 U7481 ( .A1(n5839), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7482 ( .A1(n5838), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5873) );
  NAND4_X1 U7483 ( .A1(n5876), .A2(n5875), .A3(n5874), .A4(n5873), .ZN(n8345)
         );
  INV_X1 U7484 ( .A(n8345), .ZN(n6991) );
  NAND2_X1 U7485 ( .A1(n5862), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5878) );
  INV_X1 U7486 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5877) );
  OR2_X1 U7487 ( .A1(n5824), .A2(n6606), .ZN(n5881) );
  OR2_X1 U7488 ( .A1(n5879), .A2(n6605), .ZN(n5880) );
  OAI211_X1 U7489 ( .C1(n5830), .C2(n6841), .A(n5881), .B(n5880), .ZN(n7335)
         );
  XNOR2_X1 U7490 ( .A(n5797), .B(n7335), .ZN(n5882) );
  NAND2_X1 U7491 ( .A1(n6991), .A2(n5882), .ZN(n7080) );
  INV_X1 U7492 ( .A(n5882), .ZN(n5883) );
  NAND2_X1 U7493 ( .A1(n5883), .A2(n8345), .ZN(n5884) );
  NAND2_X1 U7494 ( .A1(n7080), .A2(n5884), .ZN(n7013) );
  NAND2_X1 U7495 ( .A1(n7011), .A2(n7080), .ZN(n5897) );
  OR2_X1 U7496 ( .A1(n5886), .A2(n8784), .ZN(n5888) );
  XNOR2_X1 U7497 ( .A(n5888), .B(n5887), .ZN(n6620) );
  OR2_X1 U7498 ( .A1(n5824), .A2(n6621), .ZN(n5890) );
  OR2_X1 U7499 ( .A1(n6083), .A2(n6622), .ZN(n5889) );
  OAI211_X1 U7500 ( .C1(n5830), .C2(n6620), .A(n5890), .B(n5889), .ZN(n7084)
         );
  XNOR2_X1 U7501 ( .A(n8018), .B(n7084), .ZN(n5898) );
  NAND2_X1 U7502 ( .A1(n6475), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U7503 ( .A1(n5891), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5892) );
  AND2_X1 U7504 ( .A1(n5907), .A2(n5892), .ZN(n7409) );
  OR2_X1 U7505 ( .A1(n6078), .A2(n7409), .ZN(n5895) );
  NAND2_X1 U7506 ( .A1(n7718), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U7507 ( .A1(n5839), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5893) );
  NAND4_X1 U7508 ( .A1(n5896), .A2(n5895), .A3(n5894), .A4(n5893), .ZN(n8344)
         );
  XNOR2_X1 U7509 ( .A(n5898), .B(n8344), .ZN(n7079) );
  NAND2_X1 U7510 ( .A1(n5897), .A2(n7079), .ZN(n7078) );
  INV_X1 U7511 ( .A(n8344), .ZN(n10036) );
  NAND2_X1 U7512 ( .A1(n10036), .A2(n5898), .ZN(n5899) );
  OR2_X1 U7513 ( .A1(n5824), .A2(n6634), .ZN(n5905) );
  OR2_X1 U7514 ( .A1(n6083), .A2(n6635), .ZN(n5904) );
  OR2_X1 U7515 ( .A1(n5900), .A2(n8784), .ZN(n5902) );
  XNOR2_X1 U7516 ( .A(n5902), .B(n5901), .ZN(n6633) );
  OR2_X1 U7517 ( .A1(n5830), .A2(n6633), .ZN(n5903) );
  XNOR2_X1 U7518 ( .A(n8018), .B(n10042), .ZN(n5913) );
  NAND2_X1 U7519 ( .A1(n5838), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5912) );
  INV_X1 U7520 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6415) );
  OR2_X1 U7521 ( .A1(n5906), .A2(n6415), .ZN(n5911) );
  NAND2_X1 U7522 ( .A1(n5907), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5908) );
  AND2_X1 U7523 ( .A1(n5924), .A2(n5908), .ZN(n10041) );
  OR2_X1 U7524 ( .A1(n6078), .A2(n10041), .ZN(n5910) );
  INV_X1 U7525 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6416) );
  OR2_X1 U7526 ( .A1(n6309), .A2(n6416), .ZN(n5909) );
  XNOR2_X1 U7527 ( .A(n5913), .B(n6274), .ZN(n7153) );
  NAND2_X1 U7528 ( .A1(n8343), .A2(n5913), .ZN(n5914) );
  OR2_X1 U7529 ( .A1(n5824), .A2(n6656), .ZN(n5921) );
  OR2_X1 U7530 ( .A1(n6083), .A2(n6657), .ZN(n5920) );
  NAND2_X1 U7531 ( .A1(n5915), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5916) );
  MUX2_X1 U7532 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5916), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5918) );
  NAND2_X1 U7533 ( .A1(n5918), .A2(n5917), .ZN(n7072) );
  OR2_X1 U7534 ( .A1(n5830), .A2(n7072), .ZN(n5919) );
  XNOR2_X1 U7535 ( .A(n7344), .B(n8018), .ZN(n5931) );
  NAND2_X1 U7536 ( .A1(n6475), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5930) );
  INV_X1 U7537 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5922) );
  OR2_X1 U7538 ( .A1(n5906), .A2(n5922), .ZN(n5929) );
  INV_X1 U7539 ( .A(n5923), .ZN(n5938) );
  NAND2_X1 U7540 ( .A1(n5924), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5925) );
  AND2_X1 U7541 ( .A1(n5938), .A2(n5925), .ZN(n7342) );
  OR2_X1 U7542 ( .A1(n6078), .A2(n7342), .ZN(n5928) );
  INV_X1 U7543 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5926) );
  OR2_X1 U7544 ( .A1(n6309), .A2(n5926), .ZN(n5927) );
  NAND2_X1 U7545 ( .A1(n5931), .A2(n10038), .ZN(n7281) );
  INV_X1 U7546 ( .A(n5931), .ZN(n5932) );
  NAND2_X1 U7547 ( .A1(n8342), .A2(n5932), .ZN(n5933) );
  AND2_X1 U7548 ( .A1(n7281), .A2(n5933), .ZN(n7214) );
  NAND2_X1 U7549 ( .A1(n7212), .A2(n7281), .ZN(n5944) );
  NAND2_X1 U7550 ( .A1(n5917), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5934) );
  XNOR2_X1 U7551 ( .A(n5934), .B(n5758), .ZN(n6660) );
  OR2_X1 U7552 ( .A1(n5824), .A2(n6661), .ZN(n5936) );
  OR2_X1 U7553 ( .A1(n6083), .A2(n6662), .ZN(n5935) );
  OAI211_X1 U7554 ( .C1(n5830), .C2(n6660), .A(n5936), .B(n5935), .ZN(n7368)
         );
  XNOR2_X1 U7555 ( .A(n8018), .B(n7368), .ZN(n5945) );
  NAND2_X1 U7556 ( .A1(n6475), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5943) );
  INV_X1 U7557 ( .A(n5937), .ZN(n5952) );
  NAND2_X1 U7558 ( .A1(n5938), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5939) );
  AND2_X1 U7559 ( .A1(n5952), .A2(n5939), .ZN(n7366) );
  OR2_X1 U7560 ( .A1(n6078), .A2(n7366), .ZN(n5942) );
  NAND2_X1 U7561 ( .A1(n7718), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U7562 ( .A1(n5839), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5940) );
  NAND4_X1 U7563 ( .A1(n5943), .A2(n5942), .A3(n5941), .A4(n5940), .ZN(n8341)
         );
  XNOR2_X1 U7564 ( .A(n5945), .B(n8341), .ZN(n7280) );
  NAND2_X1 U7565 ( .A1(n5944), .A2(n7280), .ZN(n7279) );
  INV_X1 U7566 ( .A(n8341), .ZN(n6279) );
  NAND2_X1 U7567 ( .A1(n6279), .A2(n5945), .ZN(n5946) );
  NAND2_X1 U7568 ( .A1(n5947), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5949) );
  XNOR2_X1 U7569 ( .A(n5949), .B(n5948), .ZN(n7311) );
  NAND2_X1 U7570 ( .A1(n6694), .A2(n7732), .ZN(n5951) );
  OR2_X1 U7571 ( .A1(n6083), .A2(n6696), .ZN(n5950) );
  XNOR2_X1 U7572 ( .A(n7453), .B(n8018), .ZN(n5959) );
  NAND2_X1 U7573 ( .A1(n6475), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U7574 ( .A1(n5952), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5953) );
  AND2_X1 U7575 ( .A1(n5962), .A2(n5953), .ZN(n7442) );
  OR2_X1 U7576 ( .A1(n6078), .A2(n7442), .ZN(n5956) );
  NAND2_X1 U7577 ( .A1(n7718), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7578 ( .A1(n5839), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5954) );
  NAND4_X1 U7579 ( .A1(n5957), .A2(n5956), .A3(n5955), .A4(n5954), .ZN(n8340)
         );
  INV_X1 U7580 ( .A(n8340), .ZN(n7460) );
  XNOR2_X1 U7581 ( .A(n5959), .B(n7460), .ZN(n7450) );
  INV_X1 U7582 ( .A(n7450), .ZN(n5958) );
  INV_X1 U7583 ( .A(n5959), .ZN(n5960) );
  NAND2_X1 U7584 ( .A1(n5960), .A2(n8340), .ZN(n5961) );
  INV_X1 U7585 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6404) );
  OR2_X1 U7586 ( .A1(n5906), .A2(n6404), .ZN(n5968) );
  NAND2_X1 U7587 ( .A1(n5962), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5963) );
  AND2_X1 U7588 ( .A1(n5964), .A2(n5963), .ZN(n7525) );
  OR2_X1 U7589 ( .A1(n6078), .A2(n7525), .ZN(n5967) );
  INV_X1 U7590 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7464) );
  OR2_X1 U7591 ( .A1(n6309), .A2(n7464), .ZN(n5966) );
  NAND2_X1 U7592 ( .A1(n6475), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5965) );
  NAND4_X1 U7593 ( .A1(n5968), .A2(n5967), .A3(n5966), .A4(n5965), .ZN(n8339)
         );
  INV_X1 U7594 ( .A(n8339), .ZN(n8287) );
  XNOR2_X1 U7595 ( .A(n5973), .B(n8287), .ZN(n7521) );
  NAND2_X1 U7596 ( .A1(n6698), .A2(n7732), .ZN(n5972) );
  OR2_X1 U7597 ( .A1(n5969), .A2(n8784), .ZN(n5970) );
  XNOR2_X1 U7598 ( .A(n5970), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7554) );
  AOI22_X1 U7599 ( .A1(n6073), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6342), .B2(
        n7554), .ZN(n5971) );
  XNOR2_X1 U7600 ( .A(n7466), .B(n8018), .ZN(n7523) );
  XNOR2_X1 U7601 ( .A(n5975), .B(n7535), .ZN(n8291) );
  NAND2_X1 U7602 ( .A1(n6786), .A2(n7732), .ZN(n5981) );
  NAND2_X1 U7603 ( .A1(n5977), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5979) );
  INV_X1 U7604 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5978) );
  XNOR2_X1 U7605 ( .A(n5979), .B(n5978), .ZN(n6788) );
  INV_X1 U7606 ( .A(n6788), .ZN(n7610) );
  AOI22_X1 U7607 ( .A1(n6073), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6342), .B2(
        n7610), .ZN(n5980) );
  XNOR2_X1 U7608 ( .A(n8691), .B(n8018), .ZN(n5988) );
  NAND2_X1 U7609 ( .A1(n7718), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5987) );
  INV_X1 U7610 ( .A(n5996), .ZN(n5997) );
  NAND2_X1 U7611 ( .A1(n5982), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5983) );
  AND2_X1 U7612 ( .A1(n5997), .A2(n5983), .ZN(n8069) );
  OR2_X1 U7613 ( .A1(n6078), .A2(n8069), .ZN(n5986) );
  NAND2_X1 U7614 ( .A1(n6475), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U7615 ( .A1(n5839), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5984) );
  NAND4_X1 U7616 ( .A1(n5987), .A2(n5986), .A3(n5985), .A4(n5984), .ZN(n8625)
         );
  XNOR2_X1 U7617 ( .A(n5988), .B(n6289), .ZN(n8074) );
  NAND2_X1 U7618 ( .A1(n6815), .A2(n7732), .ZN(n5994) );
  OR2_X1 U7619 ( .A1(n5989), .A2(n8784), .ZN(n5990) );
  NAND2_X1 U7620 ( .A1(n5991), .A2(n5990), .ZN(n6004) );
  XNOR2_X1 U7621 ( .A(n6004), .B(n5992), .ZN(n7671) );
  AOI22_X1 U7622 ( .A1(n6073), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6342), .B2(
        n7671), .ZN(n5993) );
  XNOR2_X1 U7623 ( .A(n8773), .B(n8018), .ZN(n6003) );
  INV_X1 U7624 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8685) );
  OR2_X1 U7625 ( .A1(n5906), .A2(n8685), .ZN(n6002) );
  INV_X1 U7626 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7627 ( .A1(n5996), .A2(n5995), .ZN(n6009) );
  NAND2_X1 U7628 ( .A1(n5997), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5998) );
  AND2_X1 U7629 ( .A1(n6009), .A2(n5998), .ZN(n8620) );
  OR2_X1 U7630 ( .A1(n6078), .A2(n8620), .ZN(n6001) );
  INV_X1 U7631 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7665) );
  OR2_X1 U7632 ( .A1(n6309), .A2(n7665), .ZN(n6000) );
  NAND2_X1 U7633 ( .A1(n6475), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5999) );
  NAND4_X1 U7634 ( .A1(n6002), .A2(n6001), .A3(n6000), .A4(n5999), .ZN(n8337)
         );
  NAND2_X1 U7635 ( .A1(n6003), .A2(n8612), .ZN(n8261) );
  NOR2_X1 U7636 ( .A1(n6003), .A2(n8612), .ZN(n8263) );
  NAND2_X1 U7637 ( .A1(n6994), .A2(n7732), .ZN(n6007) );
  NAND2_X1 U7638 ( .A1(n6005), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6017) );
  XNOR2_X1 U7639 ( .A(n6016), .B(n6017), .ZN(n6996) );
  INV_X1 U7640 ( .A(n6996), .ZN(n8356) );
  AOI22_X1 U7641 ( .A1(n6073), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6342), .B2(
        n8356), .ZN(n6006) );
  XNOR2_X1 U7642 ( .A(n8682), .B(n8018), .ZN(n6015) );
  INV_X1 U7643 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8681) );
  OR2_X1 U7644 ( .A1(n5906), .A2(n8681), .ZN(n6014) );
  INV_X1 U7645 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6008) );
  OR2_X1 U7646 ( .A1(n6309), .A2(n6008), .ZN(n6013) );
  NAND2_X1 U7647 ( .A1(n6009), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6010) );
  AND2_X1 U7648 ( .A1(n6022), .A2(n6010), .ZN(n8614) );
  OR2_X1 U7649 ( .A1(n6078), .A2(n8614), .ZN(n6012) );
  NAND2_X1 U7650 ( .A1(n6475), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6011) );
  NAND4_X1 U7651 ( .A1(n6014), .A2(n6013), .A3(n6012), .A4(n6011), .ZN(n8623)
         );
  XNOR2_X1 U7652 ( .A(n6015), .B(n8623), .ZN(n8038) );
  NAND2_X1 U7653 ( .A1(n7008), .A2(n7732), .ZN(n6021) );
  NAND2_X1 U7654 ( .A1(n6017), .A2(n6016), .ZN(n6018) );
  NAND2_X1 U7655 ( .A1(n6018), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6019) );
  XNOR2_X1 U7656 ( .A(n6019), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8374) );
  AOI22_X1 U7657 ( .A1(n6073), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6342), .B2(
        n8374), .ZN(n6020) );
  XNOR2_X1 U7658 ( .A(n8333), .B(n8018), .ZN(n6028) );
  NAND2_X1 U7659 ( .A1(n6475), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6027) );
  INV_X1 U7660 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8380) );
  OR2_X1 U7661 ( .A1(n5906), .A2(n8380), .ZN(n6026) );
  INV_X1 U7662 ( .A(n6036), .ZN(n6037) );
  NAND2_X1 U7663 ( .A1(n6022), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6023) );
  AND2_X1 U7664 ( .A1(n6037), .A2(n6023), .ZN(n8325) );
  OR2_X1 U7665 ( .A1(n6078), .A2(n8325), .ZN(n6025) );
  INV_X1 U7666 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8369) );
  OR2_X1 U7667 ( .A1(n6309), .A2(n8369), .ZN(n6024) );
  XNOR2_X1 U7668 ( .A(n6028), .B(n8613), .ZN(n8322) );
  INV_X1 U7669 ( .A(n8613), .ZN(n6029) );
  NAND2_X1 U7670 ( .A1(n7176), .A2(n7732), .ZN(n6034) );
  OR2_X1 U7671 ( .A1(n6031), .A2(n8784), .ZN(n6032) );
  XNOR2_X1 U7672 ( .A(n6032), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8393) );
  AOI22_X1 U7673 ( .A1(n6073), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6342), .B2(
        n8393), .ZN(n6033) );
  INV_X1 U7674 ( .A(n8761), .ZN(n8099) );
  XNOR2_X1 U7675 ( .A(n8099), .B(n8018), .ZN(n6043) );
  NAND2_X1 U7676 ( .A1(n6475), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6042) );
  INV_X1 U7677 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8677) );
  OR2_X1 U7678 ( .A1(n5906), .A2(n8677), .ZN(n6041) );
  INV_X1 U7679 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8601) );
  OR2_X1 U7680 ( .A1(n6309), .A2(n8601), .ZN(n6040) );
  INV_X1 U7681 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6035) );
  INV_X1 U7682 ( .A(n6051), .ZN(n6052) );
  NAND2_X1 U7683 ( .A1(n6037), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6038) );
  AND2_X1 U7684 ( .A1(n6052), .A2(n6038), .ZN(n8602) );
  OR2_X1 U7685 ( .A1(n6078), .A2(n8602), .ZN(n6039) );
  XNOR2_X1 U7686 ( .A(n6043), .B(n8589), .ZN(n8093) );
  NAND2_X1 U7687 ( .A1(n8094), .A2(n8093), .ZN(n8092) );
  INV_X1 U7688 ( .A(n8589), .ZN(n6044) );
  NAND2_X1 U7689 ( .A1(n8092), .A2(n6045), .ZN(n8100) );
  NAND2_X1 U7690 ( .A1(n7196), .A2(n7732), .ZN(n6049) );
  NAND2_X1 U7691 ( .A1(n6046), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6047) );
  XNOR2_X1 U7692 ( .A(n6047), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8412) );
  AOI22_X1 U7693 ( .A1(n6073), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6342), .B2(
        n8412), .ZN(n6048) );
  XNOR2_X1 U7694 ( .A(n6086), .B(n8674), .ZN(n8102) );
  NAND2_X1 U7695 ( .A1(n6475), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6057) );
  INV_X1 U7696 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8675) );
  OR2_X1 U7697 ( .A1(n5906), .A2(n8675), .ZN(n6056) );
  INV_X1 U7698 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8592) );
  OR2_X1 U7699 ( .A1(n6309), .A2(n8592), .ZN(n6055) );
  INV_X1 U7700 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7701 ( .A1(n6052), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6053) );
  AND2_X1 U7702 ( .A1(n6064), .A2(n6053), .ZN(n8591) );
  OR2_X1 U7703 ( .A1(n6078), .A2(n8591), .ZN(n6054) );
  NAND2_X1 U7704 ( .A1(n8100), .A2(n6058), .ZN(n6060) );
  INV_X1 U7705 ( .A(n8102), .ZN(n6059) );
  NAND2_X1 U7706 ( .A1(n7222), .A2(n7732), .ZN(n6063) );
  XNOR2_X1 U7707 ( .A(n6061), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8430) );
  AOI22_X1 U7708 ( .A1(n6073), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6342), .B2(
        n8430), .ZN(n6062) );
  XNOR2_X1 U7709 ( .A(n8751), .B(n8018), .ZN(n6070) );
  NAND2_X1 U7710 ( .A1(n6475), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6069) );
  INV_X1 U7711 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8670) );
  OR2_X1 U7712 ( .A1(n5906), .A2(n8670), .ZN(n6068) );
  NAND2_X1 U7713 ( .A1(n6064), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6065) );
  AND2_X1 U7714 ( .A1(n6076), .A2(n6065), .ZN(n8580) );
  OR2_X1 U7715 ( .A1(n6078), .A2(n8580), .ZN(n6067) );
  INV_X1 U7716 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8579) );
  OR2_X1 U7717 ( .A1(n6309), .A2(n8579), .ZN(n6066) );
  XNOR2_X1 U7718 ( .A(n6070), .B(n8590), .ZN(n8298) );
  NAND2_X1 U7719 ( .A1(n7390), .A2(n7732), .ZN(n6075) );
  AOI22_X1 U7720 ( .A1(n6073), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7973), .B2(
        n6342), .ZN(n6074) );
  XNOR2_X1 U7721 ( .A(n8566), .B(n8018), .ZN(n6097) );
  NAND2_X1 U7722 ( .A1(n6475), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6082) );
  INV_X1 U7723 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n6369) );
  OR2_X1 U7724 ( .A1(n5906), .A2(n6369), .ZN(n6081) );
  INV_X1 U7725 ( .A(n6089), .ZN(n6090) );
  NAND2_X1 U7726 ( .A1(n6076), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6077) );
  AND2_X1 U7727 ( .A1(n6090), .A2(n6077), .ZN(n8563) );
  OR2_X1 U7728 ( .A1(n6078), .A2(n8563), .ZN(n6080) );
  INV_X1 U7729 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8564) );
  OR2_X1 U7730 ( .A1(n6309), .A2(n8564), .ZN(n6079) );
  XNOR2_X1 U7731 ( .A(n6097), .B(n8577), .ZN(n8051) );
  NAND2_X1 U7732 ( .A1(n7440), .A2(n7732), .ZN(n6085) );
  INV_X1 U7733 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8164) );
  OR2_X1 U7734 ( .A1(n6083), .A2(n8164), .ZN(n6084) );
  XNOR2_X1 U7735 ( .A(n6086), .B(n8744), .ZN(n6096) );
  INV_X1 U7736 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6088) );
  INV_X1 U7737 ( .A(n6103), .ZN(n6104) );
  NAND2_X1 U7738 ( .A1(n6090), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7739 ( .A1(n6104), .A2(n6091), .ZN(n8556) );
  NAND2_X1 U7740 ( .A1(n6087), .A2(n8556), .ZN(n6095) );
  INV_X1 U7741 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8743) );
  OR2_X1 U7742 ( .A1(n6106), .A2(n8743), .ZN(n6094) );
  INV_X1 U7743 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8662) );
  OR2_X1 U7744 ( .A1(n5906), .A2(n8662), .ZN(n6093) );
  INV_X1 U7745 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8555) );
  OR2_X1 U7746 ( .A1(n6309), .A2(n8555), .ZN(n6092) );
  NOR2_X1 U7747 ( .A1(n6096), .A2(n8561), .ZN(n6100) );
  AOI21_X1 U7748 ( .B1(n6096), .B2(n8561), .A(n6100), .ZN(n8251) );
  INV_X1 U7749 ( .A(n6097), .ZN(n6098) );
  NAND2_X1 U7750 ( .A1(n6098), .A2(n8577), .ZN(n8252) );
  NAND2_X1 U7751 ( .A1(n8253), .A2(n6099), .ZN(n8250) );
  INV_X1 U7752 ( .A(n6100), .ZN(n8059) );
  NAND2_X1 U7753 ( .A1(n7501), .A2(n7732), .ZN(n6102) );
  OR2_X1 U7754 ( .A1(n6083), .A2(n8239), .ZN(n6101) );
  XNOR2_X1 U7755 ( .A(n8738), .B(n8018), .ZN(n6111) );
  INV_X1 U7756 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8061) );
  NAND2_X1 U7757 ( .A1(n6104), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7758 ( .A1(n6117), .A2(n6105), .ZN(n8545) );
  NAND2_X1 U7759 ( .A1(n6087), .A2(n8545), .ZN(n6110) );
  INV_X1 U7760 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8737) );
  OR2_X1 U7761 ( .A1(n6106), .A2(n8737), .ZN(n6109) );
  INV_X1 U7762 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8659) );
  OR2_X1 U7763 ( .A1(n5906), .A2(n8659), .ZN(n6108) );
  INV_X1 U7764 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8544) );
  OR2_X1 U7765 ( .A1(n6309), .A2(n8544), .ZN(n6107) );
  NAND2_X1 U7766 ( .A1(n6111), .A2(n8528), .ZN(n6114) );
  INV_X1 U7767 ( .A(n6111), .ZN(n6112) );
  NAND2_X1 U7768 ( .A1(n6112), .A2(n8553), .ZN(n6113) );
  NAND2_X1 U7769 ( .A1(n6114), .A2(n6113), .ZN(n8058) );
  INV_X1 U7770 ( .A(n6114), .ZN(n8275) );
  NAND2_X1 U7771 ( .A1(n7579), .A2(n7732), .ZN(n6116) );
  OR2_X1 U7772 ( .A1(n6083), .A2(n7581), .ZN(n6115) );
  XNOR2_X1 U7773 ( .A(n8533), .B(n8018), .ZN(n6121) );
  NAND2_X1 U7774 ( .A1(n6117), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U7775 ( .A1(n6128), .A2(n6118), .ZN(n8532) );
  AOI22_X1 U7776 ( .A1(n8532), .A2(n6087), .B1(n5839), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n6120) );
  AOI22_X1 U7777 ( .A1(n5838), .A2(P2_REG0_REG_22__SCAN_IN), .B1(n7718), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n6119) );
  XNOR2_X1 U7778 ( .A(n6121), .B(n8542), .ZN(n8274) );
  NAND2_X1 U7779 ( .A1(n6121), .A2(n8062), .ZN(n6122) );
  NAND2_X1 U7780 ( .A1(n7637), .A2(n7732), .ZN(n6124) );
  OR2_X1 U7781 ( .A1(n6083), .A2(n7640), .ZN(n6123) );
  NAND2_X1 U7782 ( .A1(n6124), .A2(n6123), .ZN(n6296) );
  INV_X1 U7783 ( .A(n6296), .ZN(n6226) );
  XNOR2_X1 U7784 ( .A(n6226), .B(n8018), .ZN(n6125) );
  INV_X1 U7785 ( .A(n6141), .ZN(n6127) );
  INV_X1 U7786 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8516) );
  NAND2_X1 U7787 ( .A1(n6128), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7788 ( .A1(n6133), .A2(n6129), .ZN(n8517) );
  NAND2_X1 U7789 ( .A1(n8517), .A2(n6087), .ZN(n6131) );
  AOI22_X1 U7790 ( .A1(n6475), .A2(P2_REG0_REG_23__SCAN_IN), .B1(n7718), .B2(
        P2_REG1_REG_23__SCAN_IN), .ZN(n6130) );
  OAI211_X1 U7791 ( .C1(n6309), .C2(n8516), .A(n6131), .B(n6130), .ZN(n8336)
         );
  NOR2_X1 U7792 ( .A1(n6083), .A2(n7688), .ZN(n6132) );
  XNOR2_X1 U7793 ( .A(n8722), .B(n8018), .ZN(n6138) );
  INV_X1 U7794 ( .A(n6185), .ZN(n6186) );
  NAND2_X1 U7795 ( .A1(n6133), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U7796 ( .A1(n6186), .A2(n6134), .ZN(n8502) );
  NAND2_X1 U7797 ( .A1(n8502), .A2(n6087), .ZN(n6137) );
  AOI22_X1 U7798 ( .A1(n6475), .A2(P2_REG0_REG_24__SCAN_IN), .B1(n7718), .B2(
        P2_REG1_REG_24__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7799 ( .A1(n5839), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7800 ( .A1(n6138), .A2(n8514), .ZN(n8003) );
  INV_X1 U7801 ( .A(n6138), .ZN(n6139) );
  NAND2_X1 U7802 ( .A1(n6139), .A2(n8088), .ZN(n8080) );
  AND2_X1 U7803 ( .A1(n8003), .A2(n8080), .ZN(n6140) );
  OAI21_X1 U7804 ( .B1(n8044), .B2(n6141), .A(n6140), .ZN(n8085) );
  INV_X1 U7805 ( .A(n8085), .ZN(n6169) );
  NOR3_X1 U7806 ( .A1(n8044), .A2(n6141), .A3(n6140), .ZN(n6168) );
  OR2_X1 U7807 ( .A1(n6143), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7808 ( .A1(n6144), .A2(n8802), .ZN(n6688) );
  NAND2_X1 U7809 ( .A1(n6145), .A2(n6688), .ZN(n6319) );
  NAND2_X1 U7810 ( .A1(n6142), .A2(n6319), .ZN(n6322) );
  NOR4_X1 U7811 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6154) );
  INV_X1 U7812 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n8138) );
  INV_X1 U7813 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n8236) );
  INV_X1 U7814 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n8173) );
  INV_X1 U7815 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n8219) );
  NAND4_X1 U7816 ( .A1(n8138), .A2(n8236), .A3(n8173), .A4(n8219), .ZN(n6151)
         );
  NOR4_X1 U7817 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6149) );
  NOR4_X1 U7818 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6148) );
  NOR4_X1 U7819 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6147) );
  NOR4_X1 U7820 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6146) );
  NAND4_X1 U7821 ( .A1(n6149), .A2(n6148), .A3(n6147), .A4(n6146), .ZN(n6150)
         );
  NOR4_X1 U7822 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        n6151), .A4(n6150), .ZN(n6153) );
  NOR4_X1 U7823 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6152) );
  AND3_X1 U7824 ( .A1(n6154), .A2(n6153), .A3(n6152), .ZN(n6155) );
  NAND2_X1 U7825 ( .A1(n6156), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6157) );
  NAND2_X1 U7826 ( .A1(n7973), .A2(n7980), .ZN(n6306) );
  OR2_X1 U7827 ( .A1(n6331), .A2(n6326), .ZN(n6174) );
  INV_X1 U7828 ( .A(n6144), .ZN(n6161) );
  INV_X1 U7829 ( .A(n5775), .ZN(n6159) );
  NAND2_X1 U7830 ( .A1(n6174), .A2(n6658), .ZN(n6167) );
  NAND2_X2 U7831 ( .A1(n7980), .A2(n7752), .ZN(n7894) );
  INV_X1 U7832 ( .A(n7980), .ZN(n7580) );
  NAND2_X1 U7833 ( .A1(n7580), .A2(n7749), .ZN(n10102) );
  AND2_X1 U7834 ( .A1(n7894), .A2(n10102), .ZN(n6171) );
  INV_X1 U7835 ( .A(n6326), .ZN(n6165) );
  AOI21_X1 U7836 ( .B1(n6329), .B2(n6171), .A(n6165), .ZN(n6166) );
  NAND2_X1 U7837 ( .A1(n7919), .A2(n10081), .ZN(n8615) );
  INV_X1 U7838 ( .A(n8615), .ZN(n8630) );
  NAND3_X1 U7839 ( .A1(n6329), .A2(n6658), .A3(n8630), .ZN(n6170) );
  NAND2_X1 U7840 ( .A1(n6326), .A2(n6171), .ZN(n6172) );
  NAND2_X1 U7841 ( .A1(n6172), .A2(n8615), .ZN(n6330) );
  INV_X1 U7842 ( .A(n6330), .ZN(n6175) );
  NAND2_X1 U7843 ( .A1(n4314), .A2(n7441), .ZN(n7917) );
  NAND2_X1 U7844 ( .A1(n7917), .A2(n7910), .ZN(n6320) );
  AND3_X1 U7845 ( .A1(n6320), .A2(n6339), .A3(n7638), .ZN(n6173) );
  OAI211_X1 U7846 ( .C1(n6329), .C2(n6175), .A(n6174), .B(n6173), .ZN(n6176)
         );
  NAND2_X1 U7847 ( .A1(n6176), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6178) );
  OR3_X1 U7848 ( .A1(n7973), .A2(n6316), .A3(n7894), .ZN(n6204) );
  INV_X1 U7849 ( .A(n6204), .ZN(n6969) );
  NAND2_X1 U7850 ( .A1(n6969), .A2(n6658), .ZN(n7979) );
  OR2_X1 U7851 ( .A1(n6331), .A2(n7979), .ZN(n6177) );
  INV_X1 U7852 ( .A(n8336), .ZN(n8529) );
  INV_X1 U7853 ( .A(n7979), .ZN(n6179) );
  AND2_X1 U7854 ( .A1(n6331), .A2(n6179), .ZN(n6194) );
  INV_X1 U7855 ( .A(n7977), .ZN(n6182) );
  NAND2_X1 U7856 ( .A1(n6182), .A2(n7978), .ZN(n6183) );
  NAND2_X1 U7857 ( .A1(n5830), .A2(n6183), .ZN(n6312) );
  INV_X1 U7858 ( .A(n6312), .ZN(n6313) );
  INV_X1 U7859 ( .A(n8329), .ZN(n8288) );
  INV_X1 U7860 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7861 ( .A1(n6185), .A2(n6184), .ZN(n6235) );
  NAND2_X1 U7862 ( .A1(n6186), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U7863 ( .A1(n6235), .A2(n6187), .ZN(n8495) );
  NAND2_X1 U7864 ( .A1(n8495), .A2(n6087), .ZN(n6193) );
  INV_X1 U7865 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7866 ( .A1(n7718), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U7867 ( .A1(n6475), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6188) );
  OAI211_X1 U7868 ( .C1(n6309), .C2(n6190), .A(n6189), .B(n6188), .ZN(n6191)
         );
  INV_X1 U7869 ( .A(n6191), .ZN(n6192) );
  INV_X1 U7870 ( .A(n6194), .ZN(n6195) );
  AOI22_X1 U7871 ( .A1(n8479), .A2(n8283), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n6196) );
  OAI21_X1 U7872 ( .B1(n8529), .B2(n8288), .A(n6196), .ZN(n6197) );
  AOI21_X1 U7873 ( .B1(n8502), .B2(n8317), .A(n6197), .ZN(n6198) );
  OAI21_X1 U7874 ( .B1(n8722), .B2(n8332), .A(n6198), .ZN(n6199) );
  NAND2_X1 U7875 ( .A1(n6201), .A2(n6200), .ZN(P2_U3169) );
  NAND2_X1 U7876 ( .A1(n7580), .A2(n6316), .ZN(n6202) );
  AND2_X1 U7877 ( .A1(n10102), .A2(n6202), .ZN(n6203) );
  AND2_X1 U7878 ( .A1(n4314), .A2(n6203), .ZN(n6205) );
  OR2_X2 U7879 ( .A1(n6206), .A2(n7323), .ZN(n6208) );
  NAND2_X1 U7880 ( .A1(n6206), .A2(n7323), .ZN(n7754) );
  INV_X1 U7881 ( .A(n7753), .ZN(n6207) );
  NAND2_X1 U7882 ( .A1(n6879), .A2(n6208), .ZN(n7034) );
  OR2_X1 U7883 ( .A1(n8346), .A2(n10055), .ZN(n7758) );
  NAND2_X1 U7884 ( .A1(n8346), .A2(n10055), .ZN(n7760) );
  NAND2_X1 U7885 ( .A1(n7758), .A2(n7760), .ZN(n6264) );
  NAND2_X1 U7886 ( .A1(n7034), .A2(n7927), .ZN(n7035) );
  NAND2_X1 U7887 ( .A1(n7035), .A2(n7758), .ZN(n6210) );
  NAND2_X1 U7888 ( .A1(n6268), .A2(n7387), .ZN(n7782) );
  INV_X1 U7889 ( .A(n7387), .ZN(n10061) );
  NAND2_X1 U7890 ( .A1(n6209), .A2(n10061), .ZN(n7759) );
  NAND2_X1 U7891 ( .A1(n7782), .A2(n7759), .ZN(n7376) );
  NAND2_X1 U7892 ( .A1(n6210), .A2(n7929), .ZN(n7379) );
  NAND2_X1 U7893 ( .A1(n7379), .A2(n7782), .ZN(n7329) );
  INV_X1 U7894 ( .A(n7335), .ZN(n10067) );
  NAND2_X1 U7895 ( .A1(n8345), .A2(n10067), .ZN(n7783) );
  NAND2_X1 U7896 ( .A1(n6991), .A2(n7335), .ZN(n7768) );
  INV_X1 U7897 ( .A(n7084), .ZN(n10072) );
  NOR2_X1 U7898 ( .A1(n8344), .A2(n10072), .ZN(n7767) );
  NAND2_X1 U7899 ( .A1(n8344), .A2(n10072), .ZN(n10030) );
  NAND2_X1 U7900 ( .A1(n8343), .A2(n10042), .ZN(n7788) );
  AND2_X1 U7901 ( .A1(n10030), .A2(n7788), .ZN(n7770) );
  NAND2_X1 U7902 ( .A1(n10031), .A2(n7770), .ZN(n6212) );
  NAND2_X1 U7903 ( .A1(n6274), .A2(n10080), .ZN(n7786) );
  NAND2_X1 U7904 ( .A1(n6212), .A2(n7786), .ZN(n7341) );
  INV_X1 U7905 ( .A(n7341), .ZN(n6213) );
  NAND2_X1 U7906 ( .A1(n10038), .A2(n7344), .ZN(n7790) );
  NAND2_X1 U7907 ( .A1(n8342), .A2(n10083), .ZN(n7363) );
  NAND2_X1 U7908 ( .A1(n7790), .A2(n7363), .ZN(n7346) );
  NAND2_X1 U7909 ( .A1(n6213), .A2(n7934), .ZN(n7339) );
  INV_X1 U7910 ( .A(n7368), .ZN(n10089) );
  NAND2_X1 U7911 ( .A1(n8341), .A2(n10089), .ZN(n7775) );
  AND2_X1 U7912 ( .A1(n7775), .A2(n7363), .ZN(n7773) );
  NAND2_X1 U7913 ( .A1(n6279), .A2(n7368), .ZN(n7791) );
  NAND2_X1 U7914 ( .A1(n7460), .A2(n7453), .ZN(n7792) );
  INV_X1 U7915 ( .A(n7453), .ZN(n10095) );
  NAND2_X1 U7916 ( .A1(n7792), .A2(n7779), .ZN(n7938) );
  INV_X1 U7917 ( .A(n7938), .ZN(n6214) );
  INV_X1 U7918 ( .A(n7466), .ZN(n10103) );
  AND2_X1 U7919 ( .A1(n10103), .A2(n8339), .ZN(n7457) );
  NAND2_X1 U7920 ( .A1(n8287), .A2(n7466), .ZN(n7798) );
  NAND2_X1 U7921 ( .A1(n8294), .A2(n7535), .ZN(n7802) );
  INV_X1 U7922 ( .A(n7802), .ZN(n6215) );
  NAND2_X1 U7923 ( .A1(n8691), .A2(n6289), .ZN(n7808) );
  NAND2_X1 U7924 ( .A1(n7533), .A2(n7942), .ZN(n6216) );
  NAND2_X1 U7925 ( .A1(n6216), .A2(n7807), .ZN(n8631) );
  NAND2_X1 U7926 ( .A1(n8773), .A2(n8612), .ZN(n6217) );
  OR2_X1 U7927 ( .A1(n8773), .A2(n8612), .ZN(n6218) );
  NOR2_X1 U7928 ( .A1(n8682), .A2(n8266), .ZN(n7819) );
  INV_X1 U7929 ( .A(n7819), .ZN(n6219) );
  NAND2_X1 U7930 ( .A1(n8682), .A2(n8266), .ZN(n7811) );
  NAND2_X1 U7931 ( .A1(n6220), .A2(n7811), .ZN(n7987) );
  NAND2_X1 U7932 ( .A1(n8761), .A2(n8589), .ZN(n7827) );
  NAND2_X1 U7933 ( .A1(n8674), .A2(n8101), .ZN(n7830) );
  NAND2_X1 U7934 ( .A1(n7947), .A2(n7830), .ZN(n8586) );
  NAND2_X1 U7935 ( .A1(n8751), .A2(n8590), .ZN(n7831) );
  INV_X1 U7936 ( .A(n7830), .ZN(n8572) );
  NOR2_X1 U7937 ( .A1(n8575), .A2(n8572), .ZN(n6222) );
  NAND2_X1 U7938 ( .A1(n8571), .A2(n6222), .ZN(n8573) );
  NAND2_X1 U7939 ( .A1(n8573), .A2(n7948), .ZN(n8568) );
  NAND2_X1 U7940 ( .A1(n8566), .A2(n8300), .ZN(n7854) );
  NAND2_X1 U7941 ( .A1(n7746), .A2(n7854), .ZN(n7952) );
  NAND2_X1 U7942 ( .A1(n8568), .A2(n8567), .ZN(n8665) );
  NAND2_X1 U7943 ( .A1(n8665), .A2(n7746), .ZN(n8548) );
  INV_X1 U7944 ( .A(n7863), .ZN(n6223) );
  NAND2_X1 U7945 ( .A1(n8744), .A2(n8063), .ZN(n7847) );
  NAND2_X1 U7946 ( .A1(n8738), .A2(n8528), .ZN(n7869) );
  INV_X1 U7947 ( .A(n7869), .ZN(n6224) );
  NAND2_X1 U7948 ( .A1(n8533), .A2(n8062), .ZN(n7740) );
  NAND2_X1 U7949 ( .A1(n6225), .A2(n7741), .ZN(n8509) );
  INV_X1 U7950 ( .A(n8509), .ZN(n6228) );
  NAND2_X1 U7951 ( .A1(n6228), .A2(n6227), .ZN(n8504) );
  INV_X1 U7952 ( .A(n8722), .ZN(n6298) );
  NAND2_X1 U7953 ( .A1(n6298), .A2(n8088), .ZN(n7922) );
  NAND2_X1 U7954 ( .A1(n6296), .A2(n8529), .ZN(n8503) );
  AND2_X1 U7955 ( .A1(n7922), .A2(n8503), .ZN(n7874) );
  NAND2_X1 U7956 ( .A1(n8504), .A2(n7874), .ZN(n6229) );
  NAND2_X1 U7957 ( .A1(n6229), .A2(n7923), .ZN(n8487) );
  NAND2_X1 U7958 ( .A1(n7690), .A2(n7732), .ZN(n6231) );
  OR2_X1 U7959 ( .A1(n6083), .A2(n7691), .ZN(n6230) );
  NAND2_X1 U7960 ( .A1(n8717), .A2(n8500), .ZN(n7879) );
  NAND2_X1 U7961 ( .A1(n8487), .A2(n7879), .ZN(n6232) );
  NAND2_X1 U7962 ( .A1(n8799), .A2(n7732), .ZN(n6234) );
  OR2_X1 U7963 ( .A1(n6083), .A2(n8801), .ZN(n6233) );
  NAND2_X1 U7964 ( .A1(n6235), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7965 ( .A1(n6244), .A2(n6236), .ZN(n8482) );
  NAND2_X1 U7966 ( .A1(n8482), .A2(n6087), .ZN(n6241) );
  INV_X1 U7967 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8481) );
  NAND2_X1 U7968 ( .A1(n6475), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U7969 ( .A1(n7718), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6237) );
  OAI211_X1 U7970 ( .C1(n8481), .C2(n6309), .A(n6238), .B(n6237), .ZN(n6239)
         );
  INV_X1 U7971 ( .A(n6239), .ZN(n6240) );
  NOR2_X1 U7972 ( .A1(n8483), .A2(n8462), .ZN(n7885) );
  NAND2_X1 U7973 ( .A1(n8483), .A2(n8462), .ZN(n7882) );
  NAND2_X1 U7974 ( .A1(n9762), .A2(n7732), .ZN(n6243) );
  OR2_X1 U7975 ( .A1(n6083), .A2(n8798), .ZN(n6242) );
  INV_X1 U7976 ( .A(n6256), .ZN(n6246) );
  NAND2_X1 U7977 ( .A1(n6244), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7978 ( .A1(n6246), .A2(n6245), .ZN(n8468) );
  NAND2_X1 U7979 ( .A1(n8468), .A2(n6087), .ZN(n6251) );
  INV_X1 U7980 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8471) );
  NAND2_X1 U7981 ( .A1(n6475), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U7982 ( .A1(n7718), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6247) );
  OAI211_X1 U7983 ( .C1(n8471), .C2(n6309), .A(n6248), .B(n6247), .ZN(n6249)
         );
  INV_X1 U7984 ( .A(n6249), .ZN(n6250) );
  OR2_X1 U7985 ( .A1(n8028), .A2(n8315), .ZN(n6252) );
  NAND2_X1 U7986 ( .A1(n8791), .A2(n7732), .ZN(n6254) );
  OR2_X1 U7987 ( .A1(n6083), .A2(n8794), .ZN(n6253) );
  INV_X1 U7988 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6255) );
  NOR2_X1 U7989 ( .A1(n6256), .A2(n6255), .ZN(n6257) );
  NAND2_X1 U7990 ( .A1(n8452), .A2(n6087), .ZN(n6262) );
  INV_X1 U7991 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U7992 ( .A1(n6475), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U7993 ( .A1(n7718), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6258) );
  OAI211_X1 U7994 ( .C1(n8453), .C2(n6309), .A(n6259), .B(n6258), .ZN(n6260)
         );
  INV_X1 U7995 ( .A(n6260), .ZN(n6261) );
  XNOR2_X1 U7996 ( .A(n6483), .B(n8019), .ZN(n8455) );
  NAND2_X1 U7997 ( .A1(n8349), .A2(n10053), .ZN(n6883) );
  INV_X1 U7998 ( .A(n7323), .ZN(n6263) );
  OR2_X1 U7999 ( .A1(n8348), .A2(n6263), .ZN(n7039) );
  NAND2_X1 U8000 ( .A1(n6881), .A2(n7039), .ZN(n6265) );
  NAND2_X1 U8001 ( .A1(n6265), .A2(n6264), .ZN(n7381) );
  INV_X1 U8002 ( .A(n10055), .ZN(n6266) );
  OR2_X1 U8003 ( .A1(n8346), .A2(n6266), .ZN(n7380) );
  NAND2_X1 U8004 ( .A1(n7381), .A2(n7380), .ZN(n6267) );
  NAND2_X1 U8005 ( .A1(n6267), .A2(n7376), .ZN(n7383) );
  NAND2_X1 U8006 ( .A1(n6268), .A2(n10061), .ZN(n6269) );
  NAND2_X1 U8007 ( .A1(n7383), .A2(n6269), .ZN(n7330) );
  NAND2_X1 U8008 ( .A1(n8345), .A2(n7335), .ZN(n6270) );
  NAND2_X1 U8009 ( .A1(n6991), .A2(n10067), .ZN(n6271) );
  NAND2_X1 U8010 ( .A1(n8344), .A2(n7084), .ZN(n6272) );
  NAND2_X1 U8011 ( .A1(n6273), .A2(n6272), .ZN(n10033) );
  NAND2_X1 U8012 ( .A1(n6274), .A2(n10042), .ZN(n7932) );
  NAND2_X1 U8013 ( .A1(n10033), .A2(n7932), .ZN(n6275) );
  NAND2_X1 U8014 ( .A1(n8343), .A2(n10080), .ZN(n7931) );
  NAND2_X1 U8015 ( .A1(n6275), .A2(n7931), .ZN(n7345) );
  NAND2_X1 U8016 ( .A1(n10038), .A2(n10083), .ZN(n6276) );
  NAND2_X1 U8017 ( .A1(n7345), .A2(n6276), .ZN(n6278) );
  NAND2_X1 U8018 ( .A1(n8342), .A2(n7344), .ZN(n6277) );
  NAND2_X1 U8019 ( .A1(n6278), .A2(n6277), .ZN(n7369) );
  AND2_X1 U8020 ( .A1(n8341), .A2(n7368), .ZN(n6281) );
  NAND2_X1 U8021 ( .A1(n6279), .A2(n10089), .ZN(n6280) );
  NAND2_X1 U8022 ( .A1(n8340), .A2(n7453), .ZN(n6282) );
  NAND2_X1 U8023 ( .A1(n7357), .A2(n6282), .ZN(n6284) );
  NAND2_X1 U8024 ( .A1(n7460), .A2(n10095), .ZN(n6283) );
  NAND2_X1 U8025 ( .A1(n8339), .A2(n7466), .ZN(n6286) );
  NOR2_X1 U8026 ( .A1(n8339), .A2(n7466), .ZN(n6285) );
  AOI21_X1 U8027 ( .B1(n7459), .B2(n6286), .A(n6285), .ZN(n7470) );
  NAND2_X1 U8028 ( .A1(n7803), .A2(n7802), .ZN(n7940) );
  NAND2_X1 U8029 ( .A1(n7470), .A2(n7940), .ZN(n7471) );
  NAND2_X1 U8030 ( .A1(n8294), .A2(n8338), .ZN(n6287) );
  NOR2_X1 U8031 ( .A1(n8691), .A2(n8625), .ZN(n6290) );
  INV_X1 U8032 ( .A(n8691), .ZN(n6288) );
  OR2_X1 U8033 ( .A1(n8773), .A2(n8337), .ZN(n7813) );
  NAND2_X1 U8034 ( .A1(n8773), .A2(n8337), .ZN(n7812) );
  NAND2_X1 U8035 ( .A1(n7813), .A2(n7812), .ZN(n8632) );
  INV_X1 U8036 ( .A(n8682), .ZN(n8767) );
  NAND2_X1 U8037 ( .A1(n8333), .A2(n8613), .ZN(n6291) );
  NAND2_X1 U8038 ( .A1(n7989), .A2(n6291), .ZN(n6293) );
  NAND2_X1 U8039 ( .A1(n7998), .A2(n6029), .ZN(n6292) );
  INV_X1 U8040 ( .A(n8751), .ZN(n7849) );
  NAND2_X1 U8041 ( .A1(n7863), .A2(n7847), .ZN(n8551) );
  INV_X1 U8042 ( .A(n8744), .ZN(n8260) );
  NAND2_X1 U8043 ( .A1(n8260), .A2(n8063), .ZN(n8538) );
  NOR2_X1 U8044 ( .A1(n8738), .A2(n8553), .ZN(n8524) );
  NAND2_X1 U8045 ( .A1(n7741), .A2(n7740), .ZN(n8523) );
  NAND2_X1 U8046 ( .A1(n6296), .A2(n8336), .ZN(n6297) );
  NAND2_X1 U8047 ( .A1(n8722), .A2(n8088), .ZN(n6299) );
  NAND2_X1 U8048 ( .A1(n8490), .A2(n6300), .ZN(n8489) );
  INV_X1 U8049 ( .A(n8717), .ZN(n8493) );
  NAND2_X1 U8050 ( .A1(n8493), .A2(n8500), .ZN(n6301) );
  NAND2_X1 U8051 ( .A1(n8483), .A2(n8491), .ZN(n6302) );
  NAND2_X1 U8052 ( .A1(n8714), .A2(n8462), .ZN(n6303) );
  NAND2_X1 U8053 ( .A1(n8028), .A2(n8478), .ZN(n6305) );
  XNOR2_X1 U8054 ( .A(n6468), .B(n8019), .ZN(n6315) );
  NAND2_X1 U8055 ( .A1(n6316), .A2(n7752), .ZN(n7971) );
  NAND2_X1 U8056 ( .A1(n8445), .A2(n6087), .ZN(n7723) );
  INV_X1 U8057 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8233) );
  NAND2_X1 U8058 ( .A1(n7718), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6308) );
  NAND2_X1 U8059 ( .A1(n6475), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6307) );
  OAI211_X1 U8060 ( .C1(n8233), .C2(n6309), .A(n6308), .B(n6307), .ZN(n6310)
         );
  INV_X1 U8061 ( .A(n6310), .ZN(n6311) );
  OAI22_X1 U8062 ( .A1(n8024), .A2(n10039), .B1(n8315), .B2(n10037), .ZN(n6314) );
  OAI21_X1 U8063 ( .B1(n10090), .B2(n8455), .A(n8460), .ZN(n6334) );
  NAND3_X1 U8064 ( .A1(n4314), .A2(n6316), .A3(n7980), .ZN(n6317) );
  NAND2_X1 U8065 ( .A1(n6317), .A2(n7894), .ZN(n6318) );
  MUX2_X1 U8066 ( .A(n6319), .B(n6142), .S(n6318), .Z(n6962) );
  AND2_X1 U8067 ( .A1(n6320), .A2(n6658), .ZN(n6964) );
  INV_X1 U8068 ( .A(n6324), .ZN(n6325) );
  INV_X1 U8069 ( .A(n8458), .ZN(n6336) );
  NAND2_X1 U8070 ( .A1(n6325), .A2(n4909), .ZN(P2_U3487) );
  OAI21_X1 U8071 ( .B1(n6327), .B2(n6326), .A(n7979), .ZN(n6328) );
  NAND2_X1 U8072 ( .A1(n6329), .A2(n6328), .ZN(n6333) );
  NAND3_X1 U8073 ( .A1(n6331), .A2(n6658), .A3(n6330), .ZN(n6332) );
  INV_X1 U8074 ( .A(n6335), .ZN(n6337) );
  NAND2_X1 U8075 ( .A1(n6337), .A2(n4913), .ZN(P2_U3455) );
  INV_X1 U8076 ( .A(n7638), .ZN(n6338) );
  NAND2_X1 U8077 ( .A1(n7910), .A2(n7638), .ZN(n6341) );
  NAND2_X1 U8078 ( .A1(n6452), .A2(n6341), .ZN(n6450) );
  OAI21_X1 U8079 ( .B1(n6450), .B2(n6342), .A(P2_STATE_REG_SCAN_IN), .ZN(
        P2_U3150) );
  INV_X1 U8080 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10112) );
  MUX2_X1 U8081 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10112), .S(n6602), .Z(n9985)
         );
  INV_X1 U8082 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6893) );
  AND2_X1 U8083 ( .A1(n6893), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6343) );
  NAND2_X1 U8084 ( .A1(n6373), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6344) );
  OAI21_X1 U8085 ( .B1(n9960), .B2(n6343), .A(n6344), .ZN(n9963) );
  INV_X1 U8086 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9962) );
  NAND2_X1 U8087 ( .A1(n9965), .A2(n6344), .ZN(n9984) );
  NAND2_X1 U8088 ( .A1(n9985), .A2(n9984), .ZN(n9983) );
  NAND2_X1 U8089 ( .A1(n6602), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6345) );
  NAND2_X1 U8090 ( .A1(n9983), .A2(n6345), .ZN(n6346) );
  INV_X1 U8091 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6348) );
  XNOR2_X1 U8092 ( .A(n6841), .B(n6348), .ZN(n6827) );
  NAND2_X1 U8093 ( .A1(n6841), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6349) );
  NAND2_X1 U8094 ( .A1(n6828), .A2(n6349), .ZN(n6350) );
  NAND2_X1 U8095 ( .A1(n6350), .A2(n6620), .ZN(n6947) );
  MUX2_X1 U8096 ( .A(n6415), .B(P2_REG1_REG_6__SCAN_IN), .S(n6633), .Z(n6948)
         );
  INV_X1 U8097 ( .A(n7072), .ZN(n6422) );
  AOI21_X1 U8098 ( .B1(n6351), .B2(n6422), .A(n6352), .ZN(n7068) );
  INV_X1 U8099 ( .A(n6352), .ZN(n10006) );
  INV_X1 U8100 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6353) );
  MUX2_X1 U8101 ( .A(n6353), .B(P2_REG1_REG_8__SCAN_IN), .S(n6660), .Z(n10007)
         );
  INV_X1 U8102 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10120) );
  AOI21_X1 U8103 ( .B1(n6354), .B2(n6427), .A(n6356), .ZN(n7309) );
  INV_X1 U8104 ( .A(n7309), .ZN(n6355) );
  AOI22_X1 U8105 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7554), .B1(n6701), .B2(
        n6404), .ZN(n7549) );
  NOR2_X1 U8106 ( .A1(n7655), .A2(n6357), .ZN(n6358) );
  NAND2_X1 U8107 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n6788), .ZN(n6359) );
  OAI21_X1 U8108 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n6788), .A(n6359), .ZN(
        n7593) );
  NOR2_X1 U8109 ( .A1(n7671), .A2(n6360), .ZN(n6361) );
  NAND2_X1 U8110 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n6996), .ZN(n6362) );
  OAI21_X1 U8111 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n6996), .A(n6362), .ZN(
        n8361) );
  NOR2_X1 U8112 ( .A1(n8374), .A2(n6363), .ZN(n6364) );
  INV_X1 U8113 ( .A(n8374), .ZN(n7032) );
  NOR2_X1 U8114 ( .A1(n8380), .A2(n8379), .ZN(n8378) );
  AOI22_X1 U8115 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8393), .B1(n7178), .B2(
        n8677), .ZN(n8398) );
  NOR2_X1 U8116 ( .A1(n8399), .A2(n8398), .ZN(n8397) );
  NOR2_X1 U8117 ( .A1(n8412), .A2(n6365), .ZN(n6366) );
  INV_X1 U8118 ( .A(n8430), .ZN(n7293) );
  NAND2_X1 U8119 ( .A1(n7293), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6367) );
  OAI21_X1 U8120 ( .B1(n7293), .B2(P2_REG1_REG_18__SCAN_IN), .A(n6367), .ZN(
        n8423) );
  INV_X1 U8121 ( .A(n6367), .ZN(n6368) );
  NOR2_X1 U8122 ( .A1(n8422), .A2(n6368), .ZN(n6370) );
  XNOR2_X1 U8123 ( .A(n4314), .B(n6369), .ZN(n6445) );
  XNOR2_X1 U8124 ( .A(n6370), .B(n6445), .ZN(n6371) );
  OR2_X1 U8125 ( .A1(n7977), .A2(P2_U3151), .ZN(n8792) );
  NOR2_X1 U8126 ( .A1(n6450), .A2(n8792), .ZN(n6891) );
  MUX2_X1 U8127 ( .A(n8564), .B(P2_REG2_REG_19__SCAN_IN), .S(n4314), .Z(n6446)
         );
  INV_X1 U8128 ( .A(n6633), .ZN(n6955) );
  INV_X1 U8129 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6372) );
  AND2_X1 U8130 ( .A1(n6893), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U8131 ( .A1(n6373), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6375) );
  OAI21_X1 U8132 ( .B1(n9960), .B2(n6374), .A(n6375), .ZN(n9969) );
  INV_X1 U8133 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9968) );
  NAND2_X1 U8134 ( .A1(n9992), .A2(n9991), .ZN(n9990) );
  NAND2_X1 U8135 ( .A1(n6602), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U8136 ( .A1(n6377), .A2(n6861), .ZN(n6833) );
  INV_X1 U8137 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7332) );
  XNOR2_X1 U8138 ( .A(n6841), .B(n7332), .ZN(n6832) );
  NAND2_X1 U8139 ( .A1(n6841), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6379) );
  INV_X1 U8140 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7408) );
  INV_X1 U8141 ( .A(n6380), .ZN(n6942) );
  MUX2_X1 U8142 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6416), .S(n6633), .Z(n6943)
         );
  INV_X1 U8143 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6382) );
  MUX2_X1 U8144 ( .A(n6382), .B(P2_REG2_REG_8__SCAN_IN), .S(n6660), .Z(n10022)
         );
  INV_X1 U8145 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7355) );
  AOI22_X1 U8146 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7554), .B1(n6701), .B2(
        n7464), .ZN(n7541) );
  NOR2_X1 U8147 ( .A1(n7655), .A2(n6386), .ZN(n6387) );
  XOR2_X1 U8148 ( .A(n6730), .B(n6386), .Z(n7642) );
  NAND2_X1 U8149 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n6788), .ZN(n6388) );
  OAI21_X1 U8150 ( .B1(n6788), .B2(P2_REG2_REG_12__SCAN_IN), .A(n6388), .ZN(
        n7605) );
  XNOR2_X1 U8151 ( .A(n7671), .B(n6389), .ZN(n7666) );
  NAND2_X1 U8152 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n6996), .ZN(n6390) );
  OAI21_X1 U8153 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n6996), .A(n6390), .ZN(
        n8351) );
  NOR2_X1 U8154 ( .A1(n8374), .A2(n6391), .ZN(n6392) );
  XNOR2_X1 U8155 ( .A(n6391), .B(n8374), .ZN(n8370) );
  NOR2_X1 U8156 ( .A1(n8369), .A2(n8370), .ZN(n8368) );
  NAND2_X1 U8157 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n7178), .ZN(n6393) );
  OAI21_X1 U8158 ( .B1(n7178), .B2(P2_REG2_REG_16__SCAN_IN), .A(n6393), .ZN(
        n8388) );
  NOR2_X1 U8159 ( .A1(n8389), .A2(n8388), .ZN(n8387) );
  NAND2_X1 U8160 ( .A1(n7293), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6395) );
  OAI21_X1 U8161 ( .B1(n7293), .B2(P2_REG2_REG_18__SCAN_IN), .A(n6395), .ZN(
        n8421) );
  MUX2_X1 U8162 ( .A(n8592), .B(n8675), .S(n6892), .Z(n6397) );
  NAND2_X1 U8163 ( .A1(n6397), .A2(n8412), .ZN(n6440) );
  XOR2_X1 U8164 ( .A(n8412), .B(n6397), .Z(n8415) );
  MUX2_X1 U8165 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n6892), .Z(n6398) );
  OR2_X1 U8166 ( .A1(n6398), .A2(n7178), .ZN(n6439) );
  XNOR2_X1 U8167 ( .A(n6398), .B(n8393), .ZN(n8392) );
  MUX2_X1 U8168 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n6892), .Z(n6399) );
  OR2_X1 U8169 ( .A1(n6399), .A2(n7032), .ZN(n6438) );
  XNOR2_X1 U8170 ( .A(n6399), .B(n8374), .ZN(n8373) );
  MUX2_X1 U8171 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n6892), .Z(n6400) );
  OR2_X1 U8172 ( .A1(n6400), .A2(n6996), .ZN(n6437) );
  XNOR2_X1 U8173 ( .A(n6400), .B(n8356), .ZN(n8355) );
  MUX2_X1 U8174 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n6892), .Z(n6402) );
  INV_X1 U8175 ( .A(n6402), .ZN(n6401) );
  NAND2_X1 U8176 ( .A1(n7671), .A2(n6401), .ZN(n6436) );
  XNOR2_X1 U8177 ( .A(n6402), .B(n7671), .ZN(n7661) );
  MUX2_X1 U8178 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n6892), .Z(n6403) );
  AND2_X1 U8179 ( .A1(n6403), .A2(n6788), .ZN(n7595) );
  MUX2_X1 U8180 ( .A(n7643), .B(n7651), .S(n6892), .Z(n6433) );
  AND2_X1 U8181 ( .A1(n6433), .A2(n7655), .ZN(n6434) );
  MUX2_X1 U8182 ( .A(n7464), .B(n6404), .S(n6892), .Z(n6430) );
  AND2_X1 U8183 ( .A1(n6430), .A2(n7554), .ZN(n6431) );
  MUX2_X1 U8184 ( .A(n7355), .B(n10120), .S(n6892), .Z(n6426) );
  AND2_X1 U8185 ( .A1(n6426), .A2(n6427), .ZN(n6428) );
  INV_X1 U8186 ( .A(n6660), .ZN(n10012) );
  MUX2_X1 U8187 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n6892), .Z(n6423) );
  INV_X1 U8188 ( .A(n6423), .ZN(n6424) );
  MUX2_X1 U8189 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n6892), .Z(n6420) );
  INV_X1 U8190 ( .A(n6420), .ZN(n6421) );
  MUX2_X1 U8191 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n6892), .Z(n6412) );
  MUX2_X1 U8192 ( .A(n9968), .B(n9962), .S(n6181), .Z(n6407) );
  XNOR2_X1 U8193 ( .A(n6407), .B(n4426), .ZN(n9977) );
  INV_X1 U8194 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6971) );
  INV_X1 U8195 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6405) );
  MUX2_X1 U8196 ( .A(n6971), .B(n6405), .S(n6892), .Z(n6406) );
  NAND2_X1 U8197 ( .A1(n6406), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9978) );
  INV_X1 U8198 ( .A(n6407), .ZN(n6408) );
  AOI22_X1 U8199 ( .A1(n9977), .A2(n9978), .B1(n4426), .B2(n6408), .ZN(n9999)
         );
  MUX2_X1 U8200 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6892), .Z(n6409) );
  XNOR2_X1 U8201 ( .A(n6409), .B(n6602), .ZN(n10000) );
  INV_X1 U8202 ( .A(n6602), .ZN(n9989) );
  INV_X1 U8203 ( .A(n6409), .ZN(n6410) );
  MUX2_X1 U8204 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n6892), .Z(n6411) );
  XNOR2_X1 U8205 ( .A(n6411), .B(n6861), .ZN(n6874) );
  NOR2_X1 U8206 ( .A1(n6873), .A2(n6874), .ZN(n6872) );
  NOR2_X1 U8207 ( .A1(n6411), .A2(n6861), .ZN(n6823) );
  XNOR2_X1 U8208 ( .A(n6412), .B(n6841), .ZN(n6822) );
  MUX2_X1 U8209 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n6892), .Z(n6413) );
  XNOR2_X1 U8210 ( .A(n6413), .B(n6620), .ZN(n6933) );
  INV_X1 U8211 ( .A(n6413), .ZN(n6414) );
  OAI22_X1 U8212 ( .A1(n6934), .A2(n6933), .B1(n4727), .B2(n6414), .ZN(n6940)
         );
  MUX2_X1 U8213 ( .A(n6416), .B(n6415), .S(n6892), .Z(n6417) );
  NAND2_X1 U8214 ( .A1(n6417), .A2(n6955), .ZN(n6418) );
  OAI21_X1 U8215 ( .B1(n6955), .B2(n6417), .A(n6418), .ZN(n6941) );
  NOR2_X1 U8216 ( .A1(n6940), .A2(n6941), .ZN(n6939) );
  INV_X1 U8217 ( .A(n6418), .ZN(n6419) );
  XNOR2_X1 U8218 ( .A(n6420), .B(n7072), .ZN(n7066) );
  NOR2_X1 U8219 ( .A1(n7067), .A2(n7066), .ZN(n7065) );
  AOI21_X1 U8220 ( .B1(n6422), .B2(n6421), .A(n7065), .ZN(n10018) );
  XNOR2_X1 U8221 ( .A(n6423), .B(n6660), .ZN(n10017) );
  NOR2_X1 U8222 ( .A1(n10018), .A2(n10017), .ZN(n10016) );
  AOI21_X1 U8223 ( .B1(n10012), .B2(n6424), .A(n10016), .ZN(n7306) );
  INV_X1 U8224 ( .A(n6428), .ZN(n6425) );
  OAI21_X1 U8225 ( .B1(n6427), .B2(n6426), .A(n6425), .ZN(n7305) );
  NOR2_X1 U8226 ( .A1(n6428), .A2(n7304), .ZN(n7543) );
  INV_X1 U8227 ( .A(n6431), .ZN(n6429) );
  OAI21_X1 U8228 ( .B1(n7554), .B2(n6430), .A(n6429), .ZN(n7544) );
  NOR2_X1 U8229 ( .A1(n7543), .A2(n7544), .ZN(n7542) );
  INV_X1 U8230 ( .A(n6434), .ZN(n6432) );
  OAI21_X1 U8231 ( .B1(n7655), .B2(n6433), .A(n6432), .ZN(n7646) );
  NOR2_X1 U8232 ( .A1(n7645), .A2(n7646), .ZN(n7644) );
  INV_X1 U8233 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7536) );
  INV_X1 U8234 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8692) );
  MUX2_X1 U8235 ( .A(n7536), .B(n8692), .S(n6892), .Z(n6435) );
  NAND2_X1 U8236 ( .A1(n6435), .A2(n7610), .ZN(n7597) );
  NAND2_X1 U8237 ( .A1(n7661), .A2(n7662), .ZN(n7660) );
  NAND2_X1 U8238 ( .A1(n6436), .A2(n7660), .ZN(n8354) );
  NAND2_X1 U8239 ( .A1(n8355), .A2(n8354), .ZN(n8353) );
  NAND2_X1 U8240 ( .A1(n6437), .A2(n8353), .ZN(n8372) );
  NAND2_X1 U8241 ( .A1(n6438), .A2(n8371), .ZN(n8391) );
  NAND2_X1 U8242 ( .A1(n8392), .A2(n8391), .ZN(n8390) );
  NAND2_X1 U8243 ( .A1(n6439), .A2(n8390), .ZN(n8414) );
  NAND2_X1 U8244 ( .A1(n6440), .A2(n8413), .ZN(n6441) );
  MUX2_X1 U8245 ( .A(n8579), .B(n8670), .S(n6892), .Z(n6442) );
  INV_X1 U8246 ( .A(n6441), .ZN(n6444) );
  INV_X1 U8247 ( .A(n6442), .ZN(n6443) );
  NAND2_X1 U8248 ( .A1(n6444), .A2(n6443), .ZN(n8426) );
  OAI21_X1 U8249 ( .B1(n8425), .B2(n8430), .A(n8426), .ZN(n6449) );
  INV_X1 U8250 ( .A(n6445), .ZN(n6447) );
  MUX2_X1 U8251 ( .A(n6447), .B(n6446), .S(n7978), .Z(n6448) );
  XNOR2_X1 U8252 ( .A(n6449), .B(n6448), .ZN(n6456) );
  NAND2_X1 U8253 ( .A1(n7978), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8796) );
  NOR2_X1 U8254 ( .A1(n6450), .A2(n8796), .ZN(n6451) );
  MUX2_X1 U8255 ( .A(P2_U3893), .B(n6451), .S(n7977), .Z(n10011) );
  INV_X1 U8256 ( .A(n10011), .ZN(n7312) );
  NAND2_X1 U8257 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8053) );
  INV_X1 U8258 ( .A(n6452), .ZN(n6453) );
  NAND2_X1 U8259 ( .A1(n10013), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n6454) );
  OAI211_X1 U8260 ( .C1(n7312), .C2(n4314), .A(n8053), .B(n6454), .ZN(n6455)
         );
  INV_X1 U8261 ( .A(n6468), .ZN(n6466) );
  INV_X1 U8262 ( .A(SI_28_), .ZN(n6460) );
  INV_X1 U8263 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n6462) );
  INV_X1 U8264 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7696) );
  MUX2_X1 U8265 ( .A(n6462), .B(n7696), .S(n4518), .Z(n7697) );
  NAND2_X1 U8266 ( .A1(n6533), .A2(n7732), .ZN(n6464) );
  OR2_X1 U8267 ( .A1(n6083), .A2(n6462), .ZN(n6463) );
  NAND2_X1 U8268 ( .A1(n6491), .A2(n8024), .ZN(n7901) );
  AND2_X1 U8269 ( .A1(n8458), .A2(n8335), .ZN(n6472) );
  NOR2_X1 U8270 ( .A1(n6484), .A2(n6472), .ZN(n6465) );
  NOR2_X1 U8271 ( .A1(n8458), .A2(n8335), .ZN(n6471) );
  NOR2_X1 U8272 ( .A1(n7958), .A2(n6471), .ZN(n6467) );
  NAND2_X1 U8273 ( .A1(n6468), .A2(n6467), .ZN(n6469) );
  INV_X1 U8274 ( .A(n6471), .ZN(n6474) );
  NAND2_X1 U8275 ( .A1(n6484), .A2(n6472), .ZN(n6473) );
  OAI211_X1 U8276 ( .C1(n6484), .C2(n6474), .A(n6473), .B(n8627), .ZN(n6482)
         );
  INV_X1 U8277 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8224) );
  NAND2_X1 U8278 ( .A1(n6475), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U8279 ( .A1(n5839), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6476) );
  OAI211_X1 U8280 ( .C1(n5906), .C2(n8224), .A(n6477), .B(n6476), .ZN(n6478)
         );
  INV_X1 U8281 ( .A(n6478), .ZN(n6479) );
  NAND2_X1 U8282 ( .A1(n7723), .A2(n6479), .ZN(n8334) );
  AND2_X1 U8283 ( .A1(n5830), .A2(P2_B_REG_SCAN_IN), .ZN(n6480) );
  NOR2_X1 U8284 ( .A1(n10039), .A2(n6480), .ZN(n8438) );
  AOI22_X1 U8285 ( .A1(n8335), .A2(n8624), .B1(n8334), .B2(n8438), .ZN(n6481)
         );
  INV_X1 U8286 ( .A(n8335), .ZN(n8463) );
  INV_X1 U8287 ( .A(n8450), .ZN(n6486) );
  INV_X1 U8288 ( .A(n10104), .ZN(n6487) );
  NAND2_X1 U8289 ( .A1(n8450), .A2(n6487), .ZN(n6488) );
  OR2_X1 U8290 ( .A1(n6493), .A2(n10108), .ZN(n6490) );
  OR2_X1 U8291 ( .A1(n10110), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6489) );
  NAND2_X1 U8292 ( .A1(n6490), .A2(n6489), .ZN(n6492) );
  INV_X1 U8293 ( .A(n6491), .ZN(n8447) );
  NAND2_X1 U8294 ( .A1(n6492), .A2(n4911), .ZN(P2_U3456) );
  NAND2_X1 U8295 ( .A1(n6495), .A2(n6494), .ZN(n6496) );
  NAND2_X1 U8296 ( .A1(n6496), .A2(n4910), .ZN(P2_U3488) );
  NAND2_X1 U8297 ( .A1(n9253), .A2(n9940), .ZN(n9148) );
  NAND2_X1 U8298 ( .A1(n6544), .A2(n9148), .ZN(n7089) );
  NAND2_X1 U8299 ( .A1(n9256), .A2(n6755), .ZN(n6703) );
  INV_X1 U8300 ( .A(n9255), .ZN(n6497) );
  NAND2_X1 U8301 ( .A1(n6705), .A2(n6498), .ZN(n7096) );
  NAND2_X1 U8302 ( .A1(n7089), .A2(n7096), .ZN(n7095) );
  NAND2_X1 U8303 ( .A1(n7095), .A2(n6500), .ZN(n6765) );
  NAND2_X1 U8304 ( .A1(n9252), .A2(n4523), .ZN(n9149) );
  NAND2_X1 U8305 ( .A1(n6765), .A2(n6764), .ZN(n6763) );
  INV_X1 U8306 ( .A(n9252), .ZN(n6501) );
  NAND2_X1 U8307 ( .A1(n6501), .A2(n4523), .ZN(n6502) );
  XNOR2_X2 U8308 ( .A(n6503), .B(n9251), .ZN(n8988) );
  NAND2_X1 U8309 ( .A1(n6504), .A2(n6503), .ZN(n6505) );
  INV_X1 U8310 ( .A(n9250), .ZN(n7112) );
  OR2_X1 U8311 ( .A1(n6905), .A2(n7112), .ZN(n9155) );
  NAND2_X1 U8312 ( .A1(n6905), .A2(n7112), .ZN(n8990) );
  NAND2_X1 U8313 ( .A1(n7112), .A2(n6506), .ZN(n6507) );
  INV_X1 U8314 ( .A(n9249), .ZN(n7205) );
  OR2_X1 U8315 ( .A1(n9948), .A2(n7205), .ZN(n8993) );
  NAND2_X1 U8316 ( .A1(n9948), .A2(n7205), .ZN(n9097) );
  NAND2_X1 U8317 ( .A1(n8993), .A2(n9097), .ZN(n7056) );
  INV_X1 U8318 ( .A(n9248), .ZN(n7111) );
  OR2_X1 U8319 ( .A1(n7208), .A2(n7111), .ZN(n8996) );
  NAND2_X1 U8320 ( .A1(n7208), .A2(n7111), .ZN(n7118) );
  NAND2_X1 U8321 ( .A1(n8996), .A2(n7118), .ZN(n7161) );
  OR2_X1 U8322 ( .A1(n8857), .A2(n6509), .ZN(n8997) );
  NAND2_X1 U8323 ( .A1(n8857), .A2(n6509), .ZN(n9000) );
  NAND2_X1 U8324 ( .A1(n8997), .A2(n9000), .ZN(n7124) );
  NAND2_X1 U8325 ( .A1(n4520), .A2(n6509), .ZN(n6510) );
  INV_X1 U8326 ( .A(n9246), .ZN(n6511) );
  NAND2_X1 U8327 ( .A1(n9610), .A2(n6511), .ZN(n9005) );
  NAND2_X1 U8328 ( .A1(n9008), .A2(n9005), .ZN(n7235) );
  NAND2_X1 U8329 ( .A1(n7225), .A2(n7235), .ZN(n7224) );
  NAND2_X1 U8330 ( .A1(n7224), .A2(n6512), .ZN(n7263) );
  OR2_X1 U8331 ( .A1(n7301), .A2(n6513), .ZN(n9013) );
  NAND2_X1 U8332 ( .A1(n7301), .A2(n6513), .ZN(n9009) );
  NAND2_X1 U8333 ( .A1(n9013), .A2(n9009), .ZN(n9091) );
  NAND2_X1 U8334 ( .A1(n6514), .A2(n6513), .ZN(n6515) );
  OR2_X1 U8335 ( .A1(n7632), .A2(n6516), .ZN(n9012) );
  NAND2_X1 U8336 ( .A1(n7632), .A2(n6516), .ZN(n9015) );
  NAND2_X1 U8337 ( .A1(n9012), .A2(n9015), .ZN(n7506) );
  NAND2_X1 U8338 ( .A1(n7434), .A2(n7586), .ZN(n9162) );
  NAND2_X1 U8339 ( .A1(n9017), .A2(n9162), .ZN(n7421) );
  NAND2_X1 U8340 ( .A1(n7422), .A2(n7421), .ZN(n7420) );
  INV_X1 U8341 ( .A(n9242), .ZN(n9584) );
  OR2_X1 U8342 ( .A1(n9697), .A2(n9584), .ZN(n9025) );
  NAND2_X1 U8343 ( .A1(n9697), .A2(n9584), .ZN(n9163) );
  NAND2_X1 U8344 ( .A1(n9691), .A2(n9241), .ZN(n6518) );
  INV_X1 U8345 ( .A(n9691), .ZN(n9599) );
  INV_X1 U8346 ( .A(n9240), .ZN(n9586) );
  INV_X1 U8347 ( .A(n9562), .ZN(n8965) );
  NAND2_X1 U8348 ( .A1(n9687), .A2(n8965), .ZN(n9557) );
  NAND2_X1 U8349 ( .A1(n9031), .A2(n9557), .ZN(n7675) );
  NOR2_X1 U8350 ( .A1(n9574), .A2(n9239), .ZN(n6521) );
  INV_X1 U8351 ( .A(n9239), .ZN(n9545) );
  INV_X1 U8352 ( .A(n9565), .ZN(n8845) );
  NAND2_X1 U8353 ( .A1(n9677), .A2(n8845), .ZN(n9042) );
  NAND2_X1 U8354 ( .A1(n9175), .A2(n9042), .ZN(n9542) );
  AOI22_X1 U8355 ( .A1(n9538), .A2(n9542), .B1(n9677), .B2(n9565), .ZN(n9520)
         );
  NAND2_X1 U8356 ( .A1(n9531), .A2(n9238), .ZN(n6522) );
  AOI22_X1 U8357 ( .A1(n9520), .A2(n6522), .B1(n9546), .B2(n9742), .ZN(n9509)
         );
  INV_X1 U8358 ( .A(n9509), .ZN(n6524) );
  INV_X1 U8359 ( .A(n9525), .ZN(n8844) );
  OAI21_X2 U8360 ( .B1(n6524), .B2(n6523), .A(n4907), .ZN(n9487) );
  INV_X1 U8361 ( .A(n9237), .ZN(n9046) );
  NAND2_X1 U8362 ( .A1(n9484), .A2(n9236), .ZN(n6526) );
  INV_X1 U8363 ( .A(n9448), .ZN(n6556) );
  INV_X1 U8364 ( .A(n9645), .ZN(n9456) );
  INV_X1 U8365 ( .A(n9235), .ZN(n6558) );
  NAND2_X1 U8366 ( .A1(n9456), .A2(n6558), .ZN(n6528) );
  NAND2_X1 U8367 ( .A1(n9436), .A2(n9449), .ZN(n6530) );
  NOR2_X1 U8368 ( .A1(n9436), .A2(n9449), .ZN(n6529) );
  INV_X1 U8369 ( .A(n9234), .ZN(n6560) );
  NAND2_X1 U8370 ( .A1(n9719), .A2(n6560), .ZN(n6531) );
  NAND2_X1 U8371 ( .A1(n9402), .A2(n6532), .ZN(n9073) );
  NAND2_X1 U8372 ( .A1(n9075), .A2(n9073), .ZN(n9399) );
  NAND2_X1 U8373 ( .A1(n9387), .A2(n6569), .ZN(n9074) );
  NAND2_X1 U8374 ( .A1(n6533), .A2(n9080), .ZN(n6535) );
  NAND2_X1 U8375 ( .A1(n5037), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6534) );
  INV_X1 U8376 ( .A(n6819), .ZN(n6536) );
  OR2_X1 U8377 ( .A1(n9370), .A2(n6536), .ZN(n9184) );
  NAND2_X1 U8378 ( .A1(n9370), .A2(n6536), .ZN(n9186) );
  INV_X1 U8379 ( .A(n6540), .ZN(n6539) );
  NAND2_X1 U8380 ( .A1(n6539), .A2(n6538), .ZN(n9226) );
  NAND2_X1 U8381 ( .A1(n9226), .A2(n6685), .ZN(n6758) );
  AND2_X1 U8382 ( .A1(n6540), .A2(n9194), .ZN(n6541) );
  OR2_X1 U8383 ( .A1(n6758), .A2(n6541), .ZN(n9589) );
  INV_X1 U8384 ( .A(n7514), .ZN(n9695) );
  INV_X1 U8385 ( .A(n9449), .ZN(n6542) );
  OR2_X1 U8386 ( .A1(n9436), .A2(n6542), .ZN(n9137) );
  NAND2_X1 U8387 ( .A1(n9436), .A2(n6542), .ZN(n9139) );
  NAND2_X1 U8388 ( .A1(n9137), .A2(n9139), .ZN(n9431) );
  NOR2_X1 U8389 ( .A1(n9645), .A2(n6558), .ZN(n9136) );
  NOR2_X1 U8390 ( .A1(n9431), .A2(n9136), .ZN(n6559) );
  OR2_X1 U8391 ( .A1(n9255), .A2(n9145), .ZN(n6543) );
  INV_X1 U8392 ( .A(n6764), .ZN(n9094) );
  NAND2_X1 U8393 ( .A1(n8983), .A2(n9094), .ZN(n6766) );
  INV_X1 U8394 ( .A(n8988), .ZN(n9098) );
  NAND2_X1 U8395 ( .A1(n6810), .A2(n9098), .ZN(n6546) );
  NAND2_X1 U8396 ( .A1(n6504), .A2(n8914), .ZN(n8985) );
  NAND2_X1 U8397 ( .A1(n6546), .A2(n8985), .ZN(n6910) );
  INV_X1 U8398 ( .A(n6909), .ZN(n9095) );
  NAND2_X1 U8399 ( .A1(n6910), .A2(n9095), .ZN(n6547) );
  AND2_X1 U8400 ( .A1(n9000), .A2(n7118), .ZN(n8999) );
  NAND2_X1 U8401 ( .A1(n9005), .A2(n8999), .ZN(n9101) );
  NAND2_X1 U8402 ( .A1(n9008), .A2(n8997), .ZN(n9002) );
  NAND2_X1 U8403 ( .A1(n9002), .A2(n9005), .ZN(n6548) );
  NAND2_X1 U8404 ( .A1(n6548), .A2(n9101), .ZN(n9157) );
  NAND2_X1 U8405 ( .A1(n8996), .A2(n8993), .ZN(n6549) );
  OR2_X1 U8406 ( .A1(n9002), .A2(n6549), .ZN(n9159) );
  NAND2_X1 U8407 ( .A1(n9157), .A2(n9159), .ZN(n6550) );
  INV_X1 U8408 ( .A(n9015), .ZN(n6551) );
  INV_X1 U8409 ( .A(n7421), .ZN(n9104) );
  OR2_X1 U8410 ( .A1(n9691), .A2(n8966), .ZN(n9026) );
  NAND2_X1 U8411 ( .A1(n9691), .A2(n8966), .ZN(n9027) );
  NAND2_X1 U8412 ( .A1(n7570), .A2(n9027), .ZN(n6552) );
  OR2_X1 U8413 ( .A1(n8981), .A2(n9586), .ZN(n9021) );
  NAND2_X1 U8414 ( .A1(n8981), .A2(n9586), .ZN(n9166) );
  OR2_X1 U8415 ( .A1(n9574), .A2(n9545), .ZN(n9037) );
  NAND2_X1 U8416 ( .A1(n9574), .A2(n9545), .ZN(n9041) );
  NAND2_X1 U8417 ( .A1(n9037), .A2(n9041), .ZN(n9568) );
  INV_X1 U8418 ( .A(n9557), .ZN(n9030) );
  NOR2_X1 U8419 ( .A1(n9568), .A2(n9030), .ZN(n6553) );
  NAND2_X1 U8420 ( .A1(n9539), .A2(n9042), .ZN(n9522) );
  OR2_X1 U8421 ( .A1(n9531), .A2(n9546), .ZN(n9174) );
  NAND2_X1 U8422 ( .A1(n9531), .A2(n9546), .ZN(n9181) );
  XNOR2_X1 U8423 ( .A(n9512), .B(n8844), .ZN(n9508) );
  OR2_X1 U8424 ( .A1(n9512), .A2(n8844), .ZN(n9047) );
  XNOR2_X1 U8425 ( .A(n9495), .B(n9046), .ZN(n9488) );
  NAND2_X1 U8426 ( .A1(n9495), .A2(n9046), .ZN(n9053) );
  NAND2_X1 U8427 ( .A1(n9491), .A2(n9053), .ZN(n9473) );
  OR2_X1 U8428 ( .A1(n9484), .A2(n6554), .ZN(n9058) );
  NAND2_X1 U8429 ( .A1(n9484), .A2(n6554), .ZN(n9057) );
  NAND2_X1 U8430 ( .A1(n9473), .A2(n9478), .ZN(n6555) );
  OR2_X1 U8431 ( .A1(n9462), .A2(n6556), .ZN(n9059) );
  NAND2_X1 U8432 ( .A1(n9462), .A2(n6556), .ZN(n9060) );
  NAND2_X1 U8433 ( .A1(n9465), .A2(n9466), .ZN(n6557) );
  NAND2_X1 U8434 ( .A1(n6557), .A2(n9060), .ZN(n9444) );
  INV_X1 U8435 ( .A(n9136), .ZN(n9424) );
  NAND2_X1 U8436 ( .A1(n9645), .A2(n6558), .ZN(n9134) );
  NAND2_X1 U8437 ( .A1(n9424), .A2(n9134), .ZN(n9445) );
  OR2_X2 U8438 ( .A1(n9444), .A2(n9445), .ZN(n9446) );
  OR2_X1 U8439 ( .A1(n9417), .A2(n6560), .ZN(n9127) );
  NAND2_X1 U8440 ( .A1(n9417), .A2(n6560), .ZN(n9066) );
  INV_X1 U8441 ( .A(n9066), .ZN(n9197) );
  INV_X1 U8442 ( .A(n9399), .ZN(n9393) );
  INV_X1 U8443 ( .A(n9074), .ZN(n6561) );
  NOR2_X1 U8444 ( .A1(n6562), .A2(n6561), .ZN(n6563) );
  XNOR2_X1 U8445 ( .A(n6563), .B(n9078), .ZN(n6571) );
  OR2_X1 U8446 ( .A1(n7709), .A2(n4315), .ZN(n6564) );
  INV_X1 U8447 ( .A(n9563), .ZN(n9583) );
  NAND2_X1 U8448 ( .A1(n6613), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6567) );
  INV_X1 U8449 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9623) );
  OR2_X1 U8450 ( .A1(n4313), .A2(n9623), .ZN(n6566) );
  INV_X1 U8451 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9361) );
  OR2_X1 U8452 ( .A1(n5651), .A2(n9361), .ZN(n6565) );
  AND3_X1 U8453 ( .A1(n6567), .A2(n6566), .A3(n6565), .ZN(n9119) );
  INV_X1 U8454 ( .A(n9763), .ZN(n6646) );
  NAND2_X1 U8455 ( .A1(n6646), .A2(P1_B_REG_SCAN_IN), .ZN(n6568) );
  NAND2_X1 U8456 ( .A1(n4309), .A2(n6568), .ZN(n9353) );
  OAI22_X1 U8457 ( .A1(n6569), .A2(n9583), .B1(n9119), .B2(n9353), .ZN(n6570)
         );
  AND2_X1 U8458 ( .A1(n6903), .A2(n6506), .ZN(n7059) );
  NAND2_X1 U8459 ( .A1(n7059), .A2(n6508), .ZN(n7169) );
  NOR2_X2 U8460 ( .A1(n7505), .A2(n7632), .ZN(n7504) );
  NAND2_X1 U8461 ( .A1(n9748), .A2(n9570), .ZN(n9571) );
  NOR2_X2 U8462 ( .A1(n9645), .A2(n9460), .ZN(n9452) );
  NAND2_X1 U8463 ( .A1(n9723), .A2(n9452), .ZN(n9433) );
  OR2_X2 U8464 ( .A1(n9433), .A2(n9417), .ZN(n9415) );
  NOR2_X2 U8465 ( .A1(n9415), .A2(n9402), .ZN(n9383) );
  AOI21_X1 U8466 ( .B1(n9370), .B2(n9384), .A(n9548), .ZN(n6573) );
  NAND2_X1 U8467 ( .A1(n6573), .A2(n9358), .ZN(n9372) );
  NAND2_X1 U8468 ( .A1(n9376), .A2(n9372), .ZN(n6574) );
  AOI21_X1 U8469 ( .B1(n7514), .B2(n4316), .A(P1_U3086), .ZN(n6575) );
  NAND3_X1 U8470 ( .A1(n6749), .A2(n6748), .A3(n6575), .ZN(n6576) );
  INV_X1 U8471 ( .A(n9370), .ZN(n6583) );
  NAND2_X1 U8472 ( .A1(n6578), .A2(n4902), .ZN(P1_U3551) );
  INV_X1 U8473 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6582) );
  INV_X1 U8474 ( .A(n6579), .ZN(n6752) );
  NOR2_X1 U8475 ( .A1(n4965), .A2(P1_U3086), .ZN(n6584) );
  AND2_X2 U8476 ( .A1(n6584), .A2(n6610), .ZN(P1_U3973) );
  NAND2_X1 U8477 ( .A1(n4411), .A2(n6585), .ZN(n6587) );
  XNOR2_X1 U8478 ( .A(n6587), .B(n6586), .ZN(n6588) );
  NOR2_X1 U8479 ( .A1(n6588), .A2(n8946), .ZN(n6594) );
  AND2_X1 U8480 ( .A1(n8957), .A2(n6905), .ZN(n6593) );
  NOR2_X1 U8481 ( .A1(n9810), .A2(n6906), .ZN(n6592) );
  NAND2_X1 U8482 ( .A1(n9251), .A2(n9563), .ZN(n6590) );
  NAND2_X1 U8483 ( .A1(n9249), .A2(n4309), .ZN(n6589) );
  AND2_X1 U8484 ( .A1(n6590), .A2(n6589), .ZN(n6911) );
  OAI22_X1 U8485 ( .A1(n8955), .A2(n6911), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8141), .ZN(n6591) );
  OR4_X1 U8486 ( .A1(n6594), .A2(n6593), .A3(n6592), .A4(n6591), .ZN(P1_U3227)
         );
  NOR2_X1 U8487 ( .A1(n4701), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8786) );
  INV_X2 U8488 ( .A(n8786), .ZN(n8800) );
  NAND2_X1 U8489 ( .A1(n4701), .A2(P2_U3151), .ZN(n8788) );
  OAI222_X1 U8490 ( .A1(n8800), .A2(n6595), .B1(n8788), .B2(n6596), .C1(
        P2_U3151), .C2(n4426), .ZN(P2_U3294) );
  NAND2_X1 U8491 ( .A1(n4701), .A2(P1_U3086), .ZN(n9766) );
  INV_X1 U8492 ( .A(n9261), .ZN(n6638) );
  OAI222_X1 U8493 ( .A1(n9766), .A2(n6597), .B1(n9769), .B2(n6596), .C1(
        P1_U3086), .C2(n6638), .ZN(P1_U3354) );
  INV_X1 U8494 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6598) );
  INV_X1 U8495 ( .A(n9278), .ZN(n6639) );
  OAI222_X1 U8496 ( .A1(n9766), .A2(n6598), .B1(n9769), .B2(n6603), .C1(
        P1_U3086), .C2(n6639), .ZN(P1_U3353) );
  INV_X1 U8497 ( .A(n6671), .ZN(n6664) );
  OAI222_X1 U8498 ( .A1(n9766), .A2(n6599), .B1(n9769), .B2(n6600), .C1(
        P1_U3086), .C2(n6664), .ZN(P1_U3352) );
  INV_X1 U8499 ( .A(n8788), .ZN(n8795) );
  INV_X1 U8500 ( .A(n8795), .ZN(n8803) );
  OAI222_X1 U8501 ( .A1(n8800), .A2(n6601), .B1(n8803), .B2(n6600), .C1(
        P2_U3151), .C2(n6861), .ZN(P2_U3292) );
  OAI222_X1 U8502 ( .A1(n8800), .A2(n6604), .B1(n8803), .B2(n6603), .C1(
        P2_U3151), .C2(n6602), .ZN(P2_U3293) );
  OAI222_X1 U8503 ( .A1(n8800), .A2(n6605), .B1(n8803), .B2(n6606), .C1(
        P2_U3151), .C2(n6841), .ZN(P2_U3291) );
  INV_X1 U8504 ( .A(n9292), .ZN(n6665) );
  OAI222_X1 U8505 ( .A1(n6607), .A2(n9766), .B1(P1_U3086), .B2(n6665), .C1(
        n9769), .C2(n6606), .ZN(P1_U3351) );
  NAND2_X1 U8506 ( .A1(n9212), .A2(n6610), .ZN(n6609) );
  AND2_X1 U8507 ( .A1(n6609), .A2(n6608), .ZN(n6623) );
  INV_X1 U8508 ( .A(n6623), .ZN(n6612) );
  OR2_X1 U8509 ( .A1(n6610), .A2(P1_U3086), .ZN(n9123) );
  NAND2_X1 U8510 ( .A1(n6611), .A2(n9123), .ZN(n6624) );
  AND2_X1 U8511 ( .A1(n6612), .A2(n6624), .ZN(n9866) );
  NOR2_X1 U8512 ( .A1(n9866), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8513 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6618) );
  INV_X1 U8514 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6616) );
  NAND2_X1 U8515 ( .A1(n6613), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6615) );
  INV_X1 U8516 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9618) );
  OR2_X1 U8517 ( .A1(n4312), .A2(n9618), .ZN(n6614) );
  OAI211_X1 U8518 ( .C1(n5651), .C2(n6616), .A(n6615), .B(n6614), .ZN(n9355)
         );
  NAND2_X1 U8519 ( .A1(n9355), .A2(P1_U3973), .ZN(n6617) );
  OAI21_X1 U8520 ( .B1(P1_U3973), .B2(n6618), .A(n6617), .ZN(P1_U3585) );
  INV_X1 U8521 ( .A(n9311), .ZN(n6667) );
  OAI222_X1 U8522 ( .A1(n9766), .A2(n6619), .B1(n9769), .B2(n6621), .C1(
        P1_U3086), .C2(n6667), .ZN(P1_U3350) );
  OAI222_X1 U8523 ( .A1(n8800), .A2(n6622), .B1(n8803), .B2(n6621), .C1(
        P2_U3151), .C2(n6620), .ZN(P2_U3290) );
  INV_X1 U8524 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6631) );
  NAND2_X1 U8525 ( .A1(n6624), .A2(n6623), .ZN(n6650) );
  INV_X1 U8526 ( .A(n6650), .ZN(n6629) );
  NAND2_X1 U8527 ( .A1(n6646), .A2(n4992), .ZN(n6625) );
  NAND2_X1 U8528 ( .A1(n6649), .A2(n6625), .ZN(n9272) );
  AOI21_X1 U8529 ( .B1(n9763), .B2(n6626), .A(n9272), .ZN(n6627) );
  XNOR2_X1 U8530 ( .A(n6627), .B(n9271), .ZN(n6628) );
  AOI22_X1 U8531 ( .A1(n6629), .A2(n6628), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n6630) );
  OAI21_X1 U8532 ( .B1(n9904), .B2(n6631), .A(n6630), .ZN(P1_U3243) );
  INV_X1 U8533 ( .A(n9766), .ZN(n9759) );
  AOI22_X1 U8534 ( .A1(n6739), .A2(P1_STATE_REG_SCAN_IN), .B1(n9759), .B2(
        P2_DATAO_REG_6__SCAN_IN), .ZN(n6632) );
  OAI21_X1 U8535 ( .B1(n6634), .B2(n9769), .A(n6632), .ZN(P1_U3349) );
  OAI222_X1 U8536 ( .A1(n8800), .A2(n6635), .B1(n8788), .B2(n6634), .C1(
        P2_U3151), .C2(n6633), .ZN(P2_U3289) );
  AOI22_X1 U8537 ( .A1(n9792), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9759), .ZN(n6636) );
  OAI21_X1 U8538 ( .B1(n6656), .B2(n9769), .A(n6636), .ZN(P1_U3348) );
  XOR2_X1 U8539 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6671), .Z(n6643) );
  MUX2_X1 U8540 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6640), .S(n9278), .Z(n9281)
         );
  XNOR2_X1 U8541 ( .A(n9261), .B(n6637), .ZN(n9263) );
  NAND2_X1 U8542 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9270) );
  INV_X1 U8543 ( .A(n9270), .ZN(n9264) );
  NAND2_X1 U8544 ( .A1(n9263), .A2(n9264), .ZN(n9262) );
  OAI21_X1 U8545 ( .B1(n6638), .B2(n6637), .A(n9262), .ZN(n9280) );
  NAND2_X1 U8546 ( .A1(n9281), .A2(n9280), .ZN(n9279) );
  OAI21_X1 U8547 ( .B1(n6640), .B2(n6639), .A(n9279), .ZN(n6642) );
  NOR2_X1 U8548 ( .A1(n5716), .A2(n9763), .ZN(n9223) );
  INV_X1 U8549 ( .A(n9223), .ZN(n6641) );
  NAND2_X1 U8550 ( .A1(n6643), .A2(n6642), .ZN(n6663) );
  OAI211_X1 U8551 ( .C1(n6643), .C2(n6642), .A(n9883), .B(n6663), .ZN(n6644)
         );
  INV_X1 U8552 ( .A(n6644), .ZN(n6655) );
  XNOR2_X1 U8553 ( .A(n9261), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9258) );
  MUX2_X1 U8554 ( .A(n6645), .B(P1_REG1_REG_2__SCAN_IN), .S(n9278), .Z(n9283)
         );
  XNOR2_X1 U8555 ( .A(n6671), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n6647) );
  NOR2_X1 U8556 ( .A1(n6648), .A2(n6647), .ZN(n6670) );
  AOI211_X1 U8557 ( .C1(n6648), .C2(n6647), .A(n6670), .B(n9895), .ZN(n6654)
         );
  NAND2_X1 U8558 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n6652) );
  NAND2_X1 U8559 ( .A1(n9866), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n6651) );
  OAI211_X1 U8560 ( .C1(n9343), .C2(n6664), .A(n6652), .B(n6651), .ZN(n6653)
         );
  OR3_X1 U8561 ( .A1(n6655), .A2(n6654), .A3(n6653), .ZN(P1_U3246) );
  OAI222_X1 U8562 ( .A1(n8800), .A2(n6657), .B1(n8803), .B2(n6656), .C1(
        P2_U3151), .C2(n7072), .ZN(P2_U3288) );
  NOR2_X1 U8563 ( .A1(n6687), .A2(n8236), .ZN(P2_U3251) );
  NOR2_X1 U8564 ( .A1(n6687), .A2(n8138), .ZN(P2_U3245) );
  NOR2_X1 U8565 ( .A1(n6687), .A2(n8173), .ZN(P2_U3255) );
  NOR2_X1 U8566 ( .A1(n6687), .A2(n8219), .ZN(P2_U3257) );
  INV_X1 U8567 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n8152) );
  NOR2_X1 U8568 ( .A1(n6687), .A2(n8152), .ZN(P2_U3243) );
  AOI22_X1 U8569 ( .A1(n6798), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9759), .ZN(n6659) );
  OAI21_X1 U8570 ( .B1(n6661), .B2(n9769), .A(n6659), .ZN(P1_U3347) );
  OAI222_X1 U8571 ( .A1(n8800), .A2(n6662), .B1(n8788), .B2(n6661), .C1(
        P2_U3151), .C2(n6660), .ZN(P2_U3287) );
  OAI21_X1 U8572 ( .B1(n9921), .B2(n6664), .A(n6663), .ZN(n9298) );
  MUX2_X1 U8573 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6847), .S(n9292), .Z(n9299)
         );
  NAND2_X1 U8574 ( .A1(n9298), .A2(n9299), .ZN(n9297) );
  OAI21_X1 U8575 ( .B1(n6665), .B2(n6847), .A(n9297), .ZN(n9313) );
  MUX2_X1 U8576 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6666), .S(n9311), .Z(n9314)
         );
  NAND2_X1 U8577 ( .A1(n9313), .A2(n9314), .ZN(n9312) );
  OAI21_X1 U8578 ( .B1(n6667), .B2(n6666), .A(n9312), .ZN(n6668) );
  MUX2_X1 U8579 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7058), .S(n6739), .Z(n6669)
         );
  AND2_X1 U8580 ( .A1(n6668), .A2(n6669), .ZN(n6738) );
  OAI21_X1 U8581 ( .B1(n6669), .B2(n6668), .A(n9883), .ZN(n6681) );
  MUX2_X1 U8582 ( .A(n5054), .B(P1_REG1_REG_4__SCAN_IN), .S(n9292), .Z(n9294)
         );
  AOI21_X1 U8583 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9292), .A(n9293), .ZN(
        n9306) );
  XNOR2_X1 U8584 ( .A(n9311), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9305) );
  NOR2_X1 U8585 ( .A1(n9306), .A2(n9305), .ZN(n9304) );
  INV_X1 U8586 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6672) );
  MUX2_X1 U8587 ( .A(n6672), .B(P1_REG1_REG_6__SCAN_IN), .S(n6739), .Z(n6673)
         );
  NOR2_X1 U8588 ( .A1(n6674), .A2(n6673), .ZN(n6733) );
  AOI211_X1 U8589 ( .C1(n6674), .C2(n6673), .A(n9895), .B(n6733), .ZN(n6675)
         );
  INV_X1 U8590 ( .A(n6675), .ZN(n6680) );
  INV_X1 U8591 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6677) );
  NAND2_X1 U8592 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n6676) );
  OAI21_X1 U8593 ( .B1(n9904), .B2(n6677), .A(n6676), .ZN(n6678) );
  AOI21_X1 U8594 ( .B1(n6739), .B2(n9901), .A(n6678), .ZN(n6679) );
  OAI211_X1 U8595 ( .C1(n6738), .C2(n6681), .A(n6680), .B(n6679), .ZN(P1_U3249) );
  AND2_X1 U8596 ( .A1(n6682), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8597 ( .A1(n6682), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8598 ( .A1(n6682), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8599 ( .A1(n6682), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8600 ( .A1(n6682), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8601 ( .A1(n6682), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8602 ( .A1(n6682), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8603 ( .A1(n6682), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8604 ( .A1(n6682), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8605 ( .A1(n6682), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8606 ( .A1(n9256), .A2(n6684), .ZN(n9144) );
  OR2_X1 U8607 ( .A1(n9144), .A2(n6706), .ZN(n9092) );
  OAI21_X1 U8608 ( .B1(n9944), .B2(n9592), .A(n9092), .ZN(n6683) );
  NAND2_X1 U8609 ( .A1(n9255), .A2(n4309), .ZN(n6757) );
  OAI211_X1 U8610 ( .C1(n6685), .C2(n6684), .A(n6683), .B(n6757), .ZN(n6777)
         );
  NAND2_X1 U8611 ( .A1(n6777), .A2(n9959), .ZN(n6686) );
  OAI21_X1 U8612 ( .B1(n9959), .B2(n6626), .A(n6686), .ZN(P1_U3522) );
  AND2_X1 U8613 ( .A1(n6682), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8614 ( .A1(n6682), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8615 ( .A1(n6682), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8616 ( .A1(n6682), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8617 ( .A1(n6682), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8618 ( .A1(n6682), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8619 ( .A1(n6682), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8620 ( .A1(n6682), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8621 ( .A1(n6682), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8622 ( .A1(n6682), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8623 ( .A1(n6682), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8624 ( .A1(n6682), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8625 ( .A1(n6682), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8626 ( .A1(n6682), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8627 ( .A1(n6682), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  INV_X1 U8628 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6690) );
  INV_X1 U8629 ( .A(n6688), .ZN(n6689) );
  AOI22_X1 U8630 ( .A1(n6682), .A2(n6690), .B1(n6693), .B2(n6689), .ZN(
        P2_U3377) );
  INV_X1 U8631 ( .A(n6691), .ZN(n6692) );
  AOI22_X1 U8632 ( .A1(n6682), .A2(n5774), .B1(n6693), .B2(n6692), .ZN(
        P2_U3376) );
  INV_X1 U8633 ( .A(n6694), .ZN(n6697) );
  AOI22_X1 U8634 ( .A1(n7249), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9759), .ZN(n6695) );
  OAI21_X1 U8635 ( .B1(n6697), .B2(n9769), .A(n6695), .ZN(P1_U3346) );
  OAI222_X1 U8636 ( .A1(n8803), .A2(n6697), .B1(n7311), .B2(P2_U3151), .C1(
        n6696), .C2(n8800), .ZN(P2_U3286) );
  INV_X1 U8637 ( .A(n6698), .ZN(n6702) );
  AOI22_X1 U8638 ( .A1(n9780), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9759), .ZN(n6699) );
  OAI21_X1 U8639 ( .B1(n6702), .B2(n9769), .A(n6699), .ZN(P1_U3345) );
  OAI222_X1 U8640 ( .A1(n8803), .A2(n6702), .B1(n6701), .B2(P2_U3151), .C1(
        n6700), .C2(n8800), .ZN(P2_U3285) );
  OR2_X1 U8641 ( .A1(n6707), .A2(n6703), .ZN(n6704) );
  NAND2_X1 U8642 ( .A1(n6705), .A2(n6704), .ZN(n6858) );
  AOI211_X1 U8643 ( .C1(n6755), .C2(n4617), .A(n9548), .B(n7098), .ZN(n6854)
         );
  INV_X1 U8644 ( .A(n9589), .ZN(n7512) );
  NAND2_X1 U8645 ( .A1(n6858), .A2(n7512), .ZN(n6714) );
  INV_X1 U8646 ( .A(n6706), .ZN(n6708) );
  NAND2_X1 U8647 ( .A1(n6708), .A2(n6707), .ZN(n6710) );
  NAND2_X1 U8648 ( .A1(n6710), .A2(n6709), .ZN(n6711) );
  NAND2_X1 U8649 ( .A1(n6711), .A2(n9592), .ZN(n6713) );
  AOI22_X1 U8650 ( .A1(n9563), .A2(n9256), .B1(n9253), .B2(n4309), .ZN(n6712)
         );
  AND3_X1 U8651 ( .A1(n6714), .A2(n6713), .A3(n6712), .ZN(n6860) );
  INV_X1 U8652 ( .A(n6860), .ZN(n6715) );
  AOI211_X1 U8653 ( .C1(n7514), .C2(n6858), .A(n6854), .B(n6715), .ZN(n7030)
         );
  OAI22_X1 U8654 ( .A1(n9685), .A2(n9145), .B1(n9959), .B2(n4938), .ZN(n6716)
         );
  INV_X1 U8655 ( .A(n6716), .ZN(n6717) );
  OAI21_X1 U8656 ( .B1(n7030), .B2(n9957), .A(n6717), .ZN(P1_U3523) );
  XOR2_X1 U8657 ( .A(n6719), .B(n6718), .Z(n9269) );
  NAND2_X1 U8658 ( .A1(n9810), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6773) );
  AOI22_X1 U8659 ( .A1(n9269), .A2(n9806), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n6773), .ZN(n6721) );
  OR2_X1 U8661 ( .A1(n8955), .A2(n4308), .ZN(n8964) );
  INV_X1 U8662 ( .A(n8964), .ZN(n8904) );
  AOI22_X1 U8663 ( .A1(n8904), .A2(n9255), .B1(n6755), .B2(n8957), .ZN(n6720)
         );
  NAND2_X1 U8664 ( .A1(n6721), .A2(n6720), .ZN(P1_U3232) );
  INV_X1 U8665 ( .A(n6722), .ZN(n6731) );
  AOI22_X1 U8666 ( .A1(n9819), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9759), .ZN(n6723) );
  OAI21_X1 U8667 ( .B1(n6731), .B2(n9769), .A(n6723), .ZN(P1_U3344) );
  AOI21_X1 U8668 ( .B1(n6726), .B2(n6725), .A(n6724), .ZN(n6729) );
  AOI22_X1 U8669 ( .A1(n8904), .A2(n9253), .B1(n4617), .B2(n8957), .ZN(n6728)
         );
  NOR2_X1 U8670 ( .A1(n8955), .A2(n9583), .ZN(n8903) );
  AOI22_X1 U8671 ( .A1(n8903), .A2(n9256), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n6773), .ZN(n6727) );
  OAI211_X1 U8672 ( .C1(n6729), .C2(n8946), .A(n6728), .B(n6727), .ZN(P1_U3222) );
  OAI222_X1 U8673 ( .A1(n8800), .A2(n6732), .B1(n8788), .B2(n6731), .C1(
        P2_U3151), .C2(n6730), .ZN(P2_U3284) );
  AOI21_X1 U8674 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n6739), .A(n6733), .ZN(
        n9789) );
  MUX2_X1 U8675 ( .A(n6734), .B(P1_REG1_REG_7__SCAN_IN), .S(n9792), .Z(n9788)
         );
  NOR2_X1 U8676 ( .A1(n9789), .A2(n9788), .ZN(n9787) );
  MUX2_X1 U8677 ( .A(n6735), .B(P1_REG1_REG_8__SCAN_IN), .S(n6798), .Z(n6736)
         );
  NOR2_X1 U8678 ( .A1(n6737), .A2(n6736), .ZN(n6789) );
  AOI211_X1 U8679 ( .C1(n6737), .C2(n6736), .A(n9895), .B(n6789), .ZN(n6747)
         );
  NAND2_X1 U8680 ( .A1(n9792), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6740) );
  OAI21_X1 U8681 ( .B1(n9792), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6740), .ZN(
        n9785) );
  NOR2_X1 U8682 ( .A1(n9786), .A2(n9785), .ZN(n9784) );
  AOI21_X1 U8683 ( .B1(n9792), .B2(P1_REG2_REG_7__SCAN_IN), .A(n9784), .ZN(
        n6742) );
  XNOR2_X1 U8684 ( .A(n6798), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6741) );
  NOR2_X1 U8685 ( .A1(n6742), .A2(n6741), .ZN(n6797) );
  AOI211_X1 U8686 ( .C1(n6742), .C2(n6741), .A(n9889), .B(n6797), .ZN(n6746)
         );
  INV_X1 U8687 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6744) );
  NAND2_X1 U8688 ( .A1(n9901), .A2(n6798), .ZN(n6743) );
  NAND2_X1 U8689 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8854) );
  OAI211_X1 U8690 ( .C1(n6744), .C2(n9904), .A(n6743), .B(n8854), .ZN(n6745)
         );
  OR3_X1 U8691 ( .A1(n6747), .A2(n6746), .A3(n6745), .ZN(P1_U3251) );
  AND3_X1 U8692 ( .A1(n6749), .A2(P1_STATE_REG_SCAN_IN), .A3(n6748), .ZN(n6750) );
  NAND3_X1 U8693 ( .A1(n6752), .A2(n6751), .A3(n6750), .ZN(n6753) );
  INV_X2 U8694 ( .A(n9934), .ZN(n9922) );
  NOR2_X1 U8695 ( .A1(n9928), .A2(n9548), .ZN(n9603) );
  OAI21_X1 U8696 ( .B1(n9603), .B2(n9925), .A(n6755), .ZN(n6762) );
  INV_X1 U8697 ( .A(n9092), .ZN(n6759) );
  INV_X1 U8698 ( .A(n9920), .ZN(n9908) );
  NAND2_X1 U8699 ( .A1(n9908), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6756) );
  OAI211_X1 U8700 ( .C1(n6759), .C2(n6758), .A(n6757), .B(n6756), .ZN(n6760)
         );
  NAND2_X1 U8701 ( .A1(n9922), .A2(n6760), .ZN(n6761) );
  OAI211_X1 U8702 ( .C1(n4992), .C2(n9922), .A(n6762), .B(n6761), .ZN(P1_U3293) );
  OAI21_X1 U8703 ( .B1(n6765), .B2(n6764), .A(n6763), .ZN(n9930) );
  INV_X1 U8704 ( .A(n9930), .ZN(n6768) );
  OAI21_X1 U8705 ( .B1(n9094), .B2(n8983), .A(n6766), .ZN(n6767) );
  OAI22_X1 U8706 ( .A1(n6504), .A2(n4308), .B1(n6499), .B2(n9583), .ZN(n6782)
         );
  AOI21_X1 U8707 ( .B1(n6767), .B2(n9592), .A(n6782), .ZN(n9933) );
  OAI211_X1 U8708 ( .C1(n4522), .C2(n4523), .A(n9698), .B(n6807), .ZN(n9927)
         );
  OAI211_X1 U8709 ( .C1(n6768), .C2(n9953), .A(n9933), .B(n9927), .ZN(n7050)
         );
  OAI22_X1 U8710 ( .A1(n9685), .A2(n4523), .B1(n9959), .B2(n5031), .ZN(n6769)
         );
  AOI21_X1 U8711 ( .B1(n7050), .B2(n9959), .A(n6769), .ZN(n6770) );
  INV_X1 U8712 ( .A(n6770), .ZN(P1_U3525) );
  XOR2_X1 U8713 ( .A(n6772), .B(n6771), .Z(n6776) );
  AOI22_X1 U8714 ( .A1(n8904), .A2(n9252), .B1(n7101), .B2(n8957), .ZN(n6775)
         );
  AOI22_X1 U8715 ( .A1(n8903), .A2(n9255), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n6773), .ZN(n6774) );
  OAI211_X1 U8716 ( .C1(n6776), .C2(n8946), .A(n6775), .B(n6774), .ZN(P1_U3237) );
  INV_X1 U8717 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6779) );
  NAND2_X1 U8718 ( .A1(n6777), .A2(n9946), .ZN(n6778) );
  OAI21_X1 U8719 ( .B1(n9946), .B2(n6779), .A(n6778), .ZN(P1_U3453) );
  XOR2_X1 U8720 ( .A(n6781), .B(n6780), .Z(n6785) );
  INV_X1 U8721 ( .A(n8955), .ZN(n9801) );
  AOI22_X1 U8722 ( .A1(n9801), .A2(n6782), .B1(n8957), .B2(n9924), .ZN(n6784)
         );
  MUX2_X1 U8723 ( .A(n9810), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n6783) );
  OAI211_X1 U8724 ( .C1(n6785), .C2(n8946), .A(n6784), .B(n6783), .ZN(P1_U3218) );
  INV_X1 U8725 ( .A(n6786), .ZN(n6813) );
  OAI222_X1 U8726 ( .A1(n8788), .A2(n6813), .B1(n6788), .B2(P2_U3151), .C1(
        n6787), .C2(n8800), .ZN(P2_U3283) );
  MUX2_X1 U8727 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n6790), .S(n7249), .Z(n6791)
         );
  OAI21_X1 U8728 ( .B1(n6792), .B2(n6791), .A(n7248), .ZN(n6796) );
  INV_X1 U8729 ( .A(n7249), .ZN(n6794) );
  NAND2_X1 U8730 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7399) );
  NAND2_X1 U8731 ( .A1(n9866), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n6793) );
  OAI211_X1 U8732 ( .C1(n9343), .C2(n6794), .A(n7399), .B(n6793), .ZN(n6795)
         );
  AOI21_X1 U8733 ( .B1(n6796), .B2(n9880), .A(n6795), .ZN(n6804) );
  MUX2_X1 U8734 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n6799), .S(n7249), .Z(n6800)
         );
  NAND2_X1 U8735 ( .A1(n6801), .A2(n6800), .ZN(n7244) );
  OAI21_X1 U8736 ( .B1(n6801), .B2(n6800), .A(n7244), .ZN(n6802) );
  NAND2_X1 U8737 ( .A1(n6802), .A2(n9883), .ZN(n6803) );
  NAND2_X1 U8738 ( .A1(n6804), .A2(n6803), .ZN(P1_U3252) );
  OAI21_X1 U8739 ( .B1(n6806), .B2(n8988), .A(n6805), .ZN(n6842) );
  NAND2_X1 U8740 ( .A1(n6807), .A2(n8914), .ZN(n6808) );
  NAND2_X1 U8741 ( .A1(n6808), .A2(n9698), .ZN(n6809) );
  NOR2_X1 U8742 ( .A1(n6903), .A2(n6809), .ZN(n6849) );
  XNOR2_X1 U8743 ( .A(n6810), .B(n8988), .ZN(n6811) );
  AOI22_X1 U8744 ( .A1(n4309), .A2(n9250), .B1(n9252), .B2(n9563), .ZN(n8915)
         );
  OAI21_X1 U8745 ( .B1(n6811), .B2(n9544), .A(n8915), .ZN(n6845) );
  AOI211_X1 U8746 ( .C1(n9944), .C2(n6842), .A(n6849), .B(n6845), .ZN(n7023)
         );
  INV_X1 U8747 ( .A(n9685), .ZN(n7619) );
  AOI22_X1 U8748 ( .A1(n7619), .A2(n8914), .B1(n9957), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n6812) );
  OAI21_X1 U8749 ( .B1(n7023), .B2(n9957), .A(n6812), .ZN(P1_U3526) );
  INV_X1 U8750 ( .A(n9331), .ZN(n7258) );
  OAI222_X1 U8751 ( .A1(n9766), .A2(n6814), .B1(n9769), .B2(n6813), .C1(n7258), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8752 ( .A(n6815), .ZN(n6818) );
  AOI22_X1 U8753 ( .A1(n7671), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n8786), .ZN(n6816) );
  OAI21_X1 U8754 ( .B1(n6818), .B2(n8788), .A(n6816), .ZN(P2_U3282) );
  AOI22_X1 U8755 ( .A1(n9831), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9759), .ZN(n6817) );
  OAI21_X1 U8756 ( .B1(n6818), .B2(n9769), .A(n6817), .ZN(P1_U3342) );
  NAND2_X1 U8757 ( .A1(n6819), .A2(P1_U3973), .ZN(n6820) );
  OAI21_X1 U8758 ( .B1(n6462), .B2(P1_U3973), .A(n6820), .ZN(P1_U3583) );
  INV_X1 U8759 ( .A(n6821), .ZN(n6825) );
  OAI21_X1 U8760 ( .B1(n6872), .B2(n6823), .A(n6822), .ZN(n6824) );
  NAND3_X1 U8761 ( .A1(n6825), .A2(n10001), .A3(n6824), .ZN(n6840) );
  NOR2_X1 U8762 ( .A1(n4632), .A2(n6827), .ZN(n6830) );
  INV_X1 U8763 ( .A(n6828), .ZN(n6829) );
  AOI21_X1 U8764 ( .B1(n6830), .B2(n6862), .A(n6829), .ZN(n6831) );
  NAND2_X1 U8765 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7014) );
  OAI21_X1 U8766 ( .B1(n9967), .B2(n6831), .A(n7014), .ZN(n6838) );
  INV_X1 U8767 ( .A(n6832), .ZN(n6834) );
  NAND3_X1 U8768 ( .A1(n6865), .A2(n6834), .A3(n6833), .ZN(n6835) );
  AOI21_X1 U8769 ( .B1(n6836), .B2(n6835), .A(n10024), .ZN(n6837) );
  AOI211_X1 U8770 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n10013), .A(n6838), .B(
        n6837), .ZN(n6839) );
  OAI211_X1 U8771 ( .C1(n7312), .C2(n6841), .A(n6840), .B(n6839), .ZN(P2_U3186) );
  INV_X1 U8772 ( .A(n6842), .ZN(n6852) );
  NOR2_X2 U8773 ( .A1(n9934), .A2(n6844), .ZN(n9931) );
  INV_X1 U8774 ( .A(n6845), .ZN(n6846) );
  MUX2_X1 U8775 ( .A(n6847), .B(n6846), .S(n9922), .Z(n6851) );
  OAI22_X1 U8776 ( .A1(n9913), .A2(n6503), .B1(n9920), .B2(n8912), .ZN(n6848)
         );
  AOI21_X1 U8777 ( .B1(n9905), .B2(n6849), .A(n6848), .ZN(n6850) );
  OAI211_X1 U8778 ( .C1(n6852), .C2(n9556), .A(n6851), .B(n6850), .ZN(P1_U3289) );
  INV_X1 U8779 ( .A(n6843), .ZN(n6853) );
  NAND2_X1 U8780 ( .A1(n9922), .A2(n6853), .ZN(n9600) );
  INV_X1 U8781 ( .A(n9600), .ZN(n9916) );
  AOI22_X1 U8782 ( .A1(n9934), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9908), .ZN(n6856) );
  NAND2_X1 U8783 ( .A1(n9905), .A2(n6854), .ZN(n6855) );
  OAI211_X1 U8784 ( .C1(n9913), .C2(n9145), .A(n6856), .B(n6855), .ZN(n6857)
         );
  AOI21_X1 U8785 ( .B1(n9916), .B2(n6858), .A(n6857), .ZN(n6859) );
  OAI21_X1 U8786 ( .B1(n9910), .B2(n6860), .A(n6859), .ZN(P1_U3292) );
  OAI21_X1 U8787 ( .B1(n6863), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6862), .ZN(
        n6864) );
  INV_X1 U8788 ( .A(n6864), .ZN(n6871) );
  INV_X1 U8789 ( .A(n10024), .ZN(n6928) );
  OAI21_X1 U8790 ( .B1(n6866), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6865), .ZN(
        n6867) );
  AOI22_X1 U8791 ( .A1(n6928), .A2(n6867), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3151), .ZN(n6870) );
  INV_X1 U8792 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6868) );
  OR2_X1 U8793 ( .A1(n9982), .A2(n6868), .ZN(n6869) );
  OAI211_X1 U8794 ( .C1(n6871), .C2(n9967), .A(n6870), .B(n6869), .ZN(n6877)
         );
  AOI21_X1 U8795 ( .B1(n6874), .B2(n6873), .A(n6872), .ZN(n6875) );
  NOR2_X1 U8796 ( .A1(n6875), .A2(n10019), .ZN(n6876) );
  AOI211_X1 U8797 ( .C1(n10011), .C2(n4717), .A(n6877), .B(n6876), .ZN(n6878)
         );
  INV_X1 U8798 ( .A(n6878), .ZN(P2_U3185) );
  INV_X1 U8799 ( .A(n6879), .ZN(n6880) );
  AOI21_X1 U8800 ( .B1(n7753), .B2(n6882), .A(n6880), .ZN(n7328) );
  OAI21_X1 U8801 ( .B1(n6883), .B2(n6882), .A(n6881), .ZN(n6884) );
  AOI222_X1 U8802 ( .A1(n8627), .A2(n6884), .B1(n8346), .B2(n8622), .C1(n8349), 
        .C2(n8624), .ZN(n7324) );
  OAI21_X1 U8803 ( .B1(n7328), .B2(n10090), .A(n7324), .ZN(n6889) );
  INV_X1 U8804 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6885) );
  OAI22_X1 U8805 ( .A1(n7323), .A2(n8766), .B1(n10110), .B2(n6885), .ZN(n6886)
         );
  AOI21_X1 U8806 ( .B1(n6889), .B2(n10110), .A(n6886), .ZN(n6887) );
  INV_X1 U8807 ( .A(n6887), .ZN(P2_U3393) );
  OAI22_X1 U8808 ( .A1(n8656), .A2(n7323), .B1(n10124), .B2(n9962), .ZN(n6888)
         );
  AOI21_X1 U8809 ( .B1(n6889), .B2(n10124), .A(n6888), .ZN(n6890) );
  INV_X1 U8810 ( .A(n6890), .ZN(P2_U3460) );
  INV_X1 U8811 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6900) );
  INV_X1 U8812 ( .A(n6891), .ZN(n6896) );
  MUX2_X1 U8813 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n6892), .Z(n6894) );
  NAND2_X1 U8814 ( .A1(n6894), .A2(n6893), .ZN(n6895) );
  AOI22_X1 U8815 ( .A1(n10019), .A2(n6896), .B1(n9978), .B2(n6895), .ZN(n6897)
         );
  AOI21_X1 U8816 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n6897), .ZN(
        n6899) );
  NAND2_X1 U8817 ( .A1(n10011), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6898) );
  OAI211_X1 U8818 ( .C1(n9982), .C2(n6900), .A(n6899), .B(n6898), .ZN(P2_U3182) );
  OAI21_X1 U8819 ( .B1(n6902), .B2(n6909), .A(n6901), .ZN(n6918) );
  INV_X1 U8820 ( .A(n6918), .ZN(n6915) );
  INV_X1 U8821 ( .A(n6903), .ZN(n6904) );
  AOI211_X1 U8822 ( .C1(n6905), .C2(n6904), .A(n9548), .B(n7059), .ZN(n6917)
         );
  OAI22_X1 U8823 ( .A1(n9922), .A2(n6666), .B1(n6906), .B2(n9920), .ZN(n6908)
         );
  NOR2_X1 U8824 ( .A1(n9913), .A2(n6506), .ZN(n6907) );
  AOI211_X1 U8825 ( .C1(n6917), .C2(n9905), .A(n6908), .B(n6907), .ZN(n6914)
         );
  XNOR2_X1 U8826 ( .A(n6910), .B(n6909), .ZN(n6912) );
  OAI21_X1 U8827 ( .B1(n6912), .B2(n9544), .A(n6911), .ZN(n6916) );
  NAND2_X1 U8828 ( .A1(n6916), .A2(n9922), .ZN(n6913) );
  OAI211_X1 U8829 ( .C1(n6915), .C2(n9556), .A(n6914), .B(n6913), .ZN(P1_U3288) );
  AOI211_X1 U8830 ( .C1(n9944), .C2(n6918), .A(n6917), .B(n6916), .ZN(n7026)
         );
  INV_X1 U8831 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6919) );
  OAI22_X1 U8832 ( .A1(n9685), .A2(n6506), .B1(n9959), .B2(n6919), .ZN(n6920)
         );
  INV_X1 U8833 ( .A(n6920), .ZN(n6921) );
  OAI21_X1 U8834 ( .B1(n7026), .B2(n9957), .A(n6921), .ZN(P1_U3527) );
  OAI21_X1 U8835 ( .B1(n6922), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6949), .ZN(
        n6923) );
  INV_X1 U8836 ( .A(n6923), .ZN(n6932) );
  INV_X1 U8837 ( .A(n6944), .ZN(n6926) );
  NAND2_X1 U8838 ( .A1(n6924), .A2(n7408), .ZN(n6925) );
  NAND2_X1 U8839 ( .A1(n6926), .A2(n6925), .ZN(n6927) );
  AND2_X1 U8840 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7083) );
  AOI21_X1 U8841 ( .B1(n6928), .B2(n6927), .A(n7083), .ZN(n6931) );
  INV_X1 U8842 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6929) );
  OR2_X1 U8843 ( .A1(n9982), .A2(n6929), .ZN(n6930) );
  OAI211_X1 U8844 ( .C1(n6932), .C2(n9967), .A(n6931), .B(n6930), .ZN(n6937)
         );
  XNOR2_X1 U8845 ( .A(n6934), .B(n6933), .ZN(n6935) );
  NOR2_X1 U8846 ( .A1(n6935), .A2(n10019), .ZN(n6936) );
  AOI211_X1 U8847 ( .C1(n10011), .C2(n4727), .A(n6937), .B(n6936), .ZN(n6938)
         );
  INV_X1 U8848 ( .A(n6938), .ZN(P2_U3187) );
  AOI21_X1 U8849 ( .B1(n6941), .B2(n6940), .A(n6939), .ZN(n6958) );
  OR3_X1 U8850 ( .A1(n6944), .A2(n6943), .A3(n6942), .ZN(n6945) );
  AOI21_X1 U8851 ( .B1(n6946), .B2(n6945), .A(n10024), .ZN(n6954) );
  AND3_X1 U8852 ( .A1(n6949), .A2(n6948), .A3(n6947), .ZN(n6950) );
  INV_X1 U8853 ( .A(n9967), .ZN(n10014) );
  OAI21_X1 U8854 ( .B1(n6951), .B2(n6950), .A(n10014), .ZN(n6952) );
  NAND2_X1 U8855 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7154) );
  NAND2_X1 U8856 ( .A1(n6952), .A2(n7154), .ZN(n6953) );
  AOI211_X1 U8857 ( .C1(n10013), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n6954), .B(
        n6953), .ZN(n6957) );
  NAND2_X1 U8858 ( .A1(n10011), .A2(n6955), .ZN(n6956) );
  OAI211_X1 U8859 ( .C1(n6958), .C2(n10019), .A(n6957), .B(n6956), .ZN(
        P2_U3188) );
  NOR2_X1 U8860 ( .A1(n8317), .A2(P2_U3151), .ZN(n7007) );
  INV_X1 U8861 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6961) );
  NAND2_X1 U8862 ( .A1(n8349), .A2(n6975), .ZN(n7750) );
  NAND2_X1 U8863 ( .A1(n7753), .A2(n7750), .ZN(n10048) );
  OAI22_X1 U8864 ( .A1(n8332), .A2(n6975), .B1(n8324), .B2(n6981), .ZN(n6959)
         );
  AOI21_X1 U8865 ( .B1(n8320), .B2(n10048), .A(n6959), .ZN(n6960) );
  OAI21_X1 U8866 ( .B1(n7007), .B2(n6961), .A(n6960), .ZN(P2_U3172) );
  INV_X1 U8867 ( .A(n6962), .ZN(n6967) );
  INV_X1 U8868 ( .A(n7038), .ZN(n6968) );
  NOR2_X1 U8869 ( .A1(n6969), .A2(n10081), .ZN(n6970) );
  NOR2_X1 U8870 ( .A1(n6981), .A2(n10039), .ZN(n10052) );
  AOI21_X1 U8871 ( .B1(n6970), .B2(n10048), .A(n10052), .ZN(n6972) );
  MUX2_X1 U8872 ( .A(n6972), .B(n6971), .S(n8634), .Z(n6974) );
  NAND2_X1 U8873 ( .A1(n8604), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6973) );
  OAI211_X1 U8874 ( .C1(n10043), .C2(n6975), .A(n6974), .B(n6973), .ZN(
        P2_U3233) );
  OAI21_X1 U8875 ( .B1(n6979), .B2(n6976), .A(n6977), .ZN(n6980) );
  NAND2_X1 U8876 ( .A1(n6980), .A2(n8320), .ZN(n6984) );
  OAI22_X1 U8877 ( .A1(n8288), .A2(n6981), .B1(n10055), .B2(n8332), .ZN(n6982)
         );
  AOI21_X1 U8878 ( .B1(n8283), .B2(n6209), .A(n6982), .ZN(n6983) );
  OAI211_X1 U8879 ( .C1(n7007), .C2(n9986), .A(n6984), .B(n6983), .ZN(P2_U3177) );
  INV_X1 U8880 ( .A(n6986), .ZN(n6987) );
  AOI211_X1 U8881 ( .C1(n6988), .C2(n6985), .A(n8305), .B(n6987), .ZN(n6993)
         );
  MUX2_X1 U8882 ( .A(n8326), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n6990) );
  AOI22_X1 U8883 ( .A1(n8329), .A2(n8346), .B1(n7387), .B2(n8303), .ZN(n6989)
         );
  OAI211_X1 U8884 ( .C1(n6991), .C2(n8324), .A(n6990), .B(n6989), .ZN(n6992)
         );
  OR2_X1 U8885 ( .A1(n6993), .A2(n6992), .ZN(P2_U3158) );
  INV_X1 U8886 ( .A(n6994), .ZN(n6997) );
  INV_X1 U8887 ( .A(n9843), .ZN(n9332) );
  OAI222_X1 U8888 ( .A1(n9766), .A2(n6995), .B1(n9769), .B2(n6997), .C1(
        P1_U3086), .C2(n9332), .ZN(P1_U3341) );
  OAI222_X1 U8889 ( .A1(n8800), .A2(n6998), .B1(n8788), .B2(n6997), .C1(
        P2_U3151), .C2(n6996), .ZN(P2_U3281) );
  INV_X1 U8890 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7322) );
  INV_X1 U8891 ( .A(n8349), .ZN(n6999) );
  OAI22_X1 U8892 ( .A1(n8288), .A2(n6999), .B1(n7323), .B2(n8332), .ZN(n7000)
         );
  AOI21_X1 U8893 ( .B1(n8283), .B2(n8346), .A(n7000), .ZN(n7006) );
  OAI21_X1 U8894 ( .B1(n7001), .B2(n7003), .A(n7002), .ZN(n7004) );
  NAND2_X1 U8895 ( .A1(n7004), .A2(n8320), .ZN(n7005) );
  OAI211_X1 U8896 ( .C1(n7007), .C2(n7322), .A(n7006), .B(n7005), .ZN(P2_U3162) );
  INV_X1 U8897 ( .A(n7008), .ZN(n7033) );
  AOI22_X1 U8898 ( .A1(n9857), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n9759), .ZN(n7009) );
  OAI21_X1 U8899 ( .B1(n7033), .B2(n9769), .A(n7009), .ZN(P1_U3340) );
  INV_X1 U8900 ( .A(n7011), .ZN(n7012) );
  AOI21_X1 U8901 ( .B1(n7010), .B2(n7013), .A(n7012), .ZN(n7020) );
  AOI22_X1 U8902 ( .A1(n8283), .A2(n8344), .B1(n8329), .B2(n6209), .ZN(n7017)
         );
  INV_X1 U8903 ( .A(n7014), .ZN(n7015) );
  AOI21_X1 U8904 ( .B1(n8303), .B2(n7335), .A(n7015), .ZN(n7016) );
  OAI211_X1 U8905 ( .C1(n8326), .C2(n7333), .A(n7017), .B(n7016), .ZN(n7018)
         );
  INV_X1 U8906 ( .A(n7018), .ZN(n7019) );
  OAI21_X1 U8907 ( .B1(n7020), .B2(n8305), .A(n7019), .ZN(P2_U3170) );
  INV_X1 U8908 ( .A(n9946), .ZN(n9955) );
  OAI22_X1 U8909 ( .A1(n9747), .A2(n6503), .B1(n9946), .B2(n5055), .ZN(n7021)
         );
  INV_X1 U8910 ( .A(n7021), .ZN(n7022) );
  OAI21_X1 U8911 ( .B1(n7023), .B2(n9955), .A(n7022), .ZN(P1_U3465) );
  OAI22_X1 U8912 ( .A1(n9747), .A2(n6506), .B1(n9946), .B2(n5093), .ZN(n7024)
         );
  INV_X1 U8913 ( .A(n7024), .ZN(n7025) );
  OAI21_X1 U8914 ( .B1(n7026), .B2(n9955), .A(n7025), .ZN(P1_U3468) );
  INV_X1 U8915 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7027) );
  OAI22_X1 U8916 ( .A1(n9747), .A2(n9145), .B1(n9946), .B2(n7027), .ZN(n7028)
         );
  INV_X1 U8917 ( .A(n7028), .ZN(n7029) );
  OAI21_X1 U8918 ( .B1(n7030), .B2(n9955), .A(n7029), .ZN(P1_U3456) );
  OAI222_X1 U8919 ( .A1(n8788), .A2(n7033), .B1(n7032), .B2(P2_U3151), .C1(
        n7031), .C2(n8800), .ZN(P2_U3280) );
  OR2_X1 U8920 ( .A1(n7034), .A2(n7927), .ZN(n7036) );
  AND2_X1 U8921 ( .A1(n7036), .A2(n7377), .ZN(n10056) );
  OR2_X1 U8922 ( .A1(n7919), .A2(n7749), .ZN(n7037) );
  NOR2_X1 U8923 ( .A1(n7038), .A2(n7037), .ZN(n8449) );
  INV_X1 U8924 ( .A(n8449), .ZN(n7469) );
  AOI22_X1 U8925 ( .A1(n6209), .A2(n8622), .B1(n8624), .B2(n8348), .ZN(n7043)
         );
  INV_X1 U8926 ( .A(n7381), .ZN(n7041) );
  AND3_X1 U8927 ( .A1(n6881), .A2(n7927), .A3(n7039), .ZN(n7040) );
  OAI21_X1 U8928 ( .B1(n7041), .B2(n7040), .A(n8627), .ZN(n7042) );
  OAI211_X1 U8929 ( .C1(n10056), .C2(n6485), .A(n7043), .B(n7042), .ZN(n10058)
         );
  INV_X1 U8930 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9986) );
  OAI22_X1 U8931 ( .A1(n10040), .A2(n9986), .B1(n10055), .B2(n8615), .ZN(n7044) );
  NOR2_X1 U8932 ( .A1(n10058), .A2(n7044), .ZN(n7045) );
  MUX2_X1 U8933 ( .A(n7045), .B(n6372), .S(n8634), .Z(n7046) );
  OAI21_X1 U8934 ( .B1(n10056), .B2(n7469), .A(n7046), .ZN(P2_U3231) );
  NAND2_X1 U8935 ( .A1(n8347), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7047) );
  OAI21_X1 U8936 ( .B1(n8024), .B2(n8347), .A(n7047), .ZN(P2_U3520) );
  INV_X1 U8937 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7048) );
  OAI22_X1 U8938 ( .A1(n9747), .A2(n4523), .B1(n9946), .B2(n7048), .ZN(n7049)
         );
  AOI21_X1 U8939 ( .B1(n7050), .B2(n9946), .A(n7049), .ZN(n7051) );
  INV_X1 U8940 ( .A(n7051), .ZN(P1_U3462) );
  OAI21_X1 U8941 ( .B1(n7053), .B2(n7056), .A(n7052), .ZN(n7054) );
  INV_X1 U8942 ( .A(n7054), .ZN(n9952) );
  XOR2_X1 U8943 ( .A(n7055), .B(n7056), .Z(n7057) );
  AOI222_X1 U8944 ( .A1(n9592), .A2(n7057), .B1(n9248), .B2(n4309), .C1(n9250), 
        .C2(n9563), .ZN(n9951) );
  MUX2_X1 U8945 ( .A(n7058), .B(n9951), .S(n9922), .Z(n7064) );
  INV_X1 U8946 ( .A(n7059), .ZN(n7061) );
  INV_X1 U8947 ( .A(n7169), .ZN(n7060) );
  AOI211_X1 U8948 ( .C1(n9948), .C2(n7061), .A(n9548), .B(n7060), .ZN(n9947)
         );
  OAI22_X1 U8949 ( .A1(n9913), .A2(n6508), .B1(n9920), .B2(n7110), .ZN(n7062)
         );
  AOI21_X1 U8950 ( .B1(n9947), .B2(n9905), .A(n7062), .ZN(n7063) );
  OAI211_X1 U8951 ( .C1(n9952), .C2(n9556), .A(n7064), .B(n7063), .ZN(P1_U3287) );
  AOI21_X1 U8952 ( .B1(n7067), .B2(n7066), .A(n7065), .ZN(n7077) );
  OAI21_X1 U8953 ( .B1(n7068), .B2(P2_REG1_REG_7__SCAN_IN), .A(n10008), .ZN(
        n7075) );
  XNOR2_X1 U8954 ( .A(n7069), .B(n5926), .ZN(n7070) );
  NOR2_X1 U8955 ( .A1(n7070), .A2(n10024), .ZN(n7074) );
  NAND2_X1 U8956 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7215) );
  NAND2_X1 U8957 ( .A1(n10013), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7071) );
  OAI211_X1 U8958 ( .C1(n7312), .C2(n7072), .A(n7215), .B(n7071), .ZN(n7073)
         );
  AOI211_X1 U8959 ( .C1(n7075), .C2(n10014), .A(n7074), .B(n7073), .ZN(n7076)
         );
  OAI21_X1 U8960 ( .B1(n7077), .B2(n10019), .A(n7076), .ZN(P2_U3189) );
  INV_X1 U8961 ( .A(n7079), .ZN(n7081) );
  NAND3_X1 U8962 ( .A1(n7011), .A2(n7081), .A3(n7080), .ZN(n7082) );
  AOI21_X1 U8963 ( .B1(n7078), .B2(n7082), .A(n8305), .ZN(n7088) );
  AOI22_X1 U8964 ( .A1(n8283), .A2(n8343), .B1(n8329), .B2(n8345), .ZN(n7086)
         );
  AOI21_X1 U8965 ( .B1(n8303), .B2(n7084), .A(n7083), .ZN(n7085) );
  OAI211_X1 U8966 ( .C1(n8326), .C2(n7409), .A(n7086), .B(n7085), .ZN(n7087)
         );
  OR2_X1 U8967 ( .A1(n7088), .A2(n7087), .ZN(P2_U3167) );
  INV_X1 U8968 ( .A(n7089), .ZN(n7090) );
  XNOR2_X1 U8969 ( .A(n7091), .B(n7090), .ZN(n7092) );
  NAND2_X1 U8970 ( .A1(n7092), .A2(n9592), .ZN(n7094) );
  AOI22_X1 U8971 ( .A1(n9563), .A2(n9255), .B1(n9252), .B2(n4309), .ZN(n7093)
         );
  NAND2_X1 U8972 ( .A1(n7094), .A2(n7093), .ZN(n9941) );
  INV_X1 U8973 ( .A(n9941), .ZN(n7105) );
  OAI21_X1 U8974 ( .B1(n7096), .B2(n7089), .A(n7095), .ZN(n9943) );
  OAI211_X1 U8975 ( .C1(n7098), .C2(n9940), .A(n9698), .B(n7097), .ZN(n9938)
         );
  NAND2_X1 U8976 ( .A1(n9910), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7099) );
  OAI21_X1 U8977 ( .B1(n9920), .B2(n9275), .A(n7099), .ZN(n7100) );
  AOI21_X1 U8978 ( .B1(n9925), .B2(n7101), .A(n7100), .ZN(n7102) );
  OAI21_X1 U8979 ( .B1(n9928), .B2(n9938), .A(n7102), .ZN(n7103) );
  AOI21_X1 U8980 ( .B1(n9931), .B2(n9943), .A(n7103), .ZN(n7104) );
  OAI21_X1 U8981 ( .B1(n9910), .B2(n7105), .A(n7104), .ZN(P1_U3291) );
  AOI21_X1 U8982 ( .B1(n7108), .B2(n7107), .A(n7106), .ZN(n7116) );
  OAI22_X1 U8983 ( .A1(n9810), .A2(n7110), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7109), .ZN(n7114) );
  INV_X1 U8984 ( .A(n8903), .ZN(n8967) );
  OAI22_X1 U8985 ( .A1(n8967), .A2(n7112), .B1(n7111), .B2(n8964), .ZN(n7113)
         );
  AOI211_X1 U8986 ( .C1(n9948), .C2(n8957), .A(n7114), .B(n7113), .ZN(n7115)
         );
  OAI21_X1 U8987 ( .B1(n7116), .B2(n8946), .A(n7115), .ZN(P1_U3239) );
  AND2_X1 U8988 ( .A1(n7117), .A2(n8993), .ZN(n7164) );
  INV_X1 U8989 ( .A(n7161), .ZN(n8995) );
  NAND2_X1 U8990 ( .A1(n7164), .A2(n8995), .ZN(n7163) );
  NAND2_X1 U8991 ( .A1(n7163), .A2(n7118), .ZN(n7233) );
  XNOR2_X1 U8992 ( .A(n7233), .B(n7124), .ZN(n7122) );
  NAND2_X1 U8993 ( .A1(n9246), .A2(n4309), .ZN(n7120) );
  NAND2_X1 U8994 ( .A1(n9248), .A2(n9563), .ZN(n7119) );
  NAND2_X1 U8995 ( .A1(n7120), .A2(n7119), .ZN(n8856) );
  INV_X1 U8996 ( .A(n8856), .ZN(n7121) );
  OAI21_X1 U8997 ( .B1(n7122), .B2(n9544), .A(n7121), .ZN(n7180) );
  INV_X1 U8998 ( .A(n7180), .ZN(n7132) );
  OAI21_X1 U8999 ( .B1(n7125), .B2(n7124), .A(n7123), .ZN(n7182) );
  INV_X1 U9000 ( .A(n7226), .ZN(n7126) );
  AOI211_X1 U9001 ( .C1(n8857), .C2(n7168), .A(n9548), .B(n7126), .ZN(n7181)
         );
  NAND2_X1 U9002 ( .A1(n7181), .A2(n9905), .ZN(n7129) );
  INV_X1 U9003 ( .A(n8858), .ZN(n7127) );
  AOI22_X1 U9004 ( .A1(n9934), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7127), .B2(
        n9908), .ZN(n7128) );
  OAI211_X1 U9005 ( .C1(n4520), .C2(n9913), .A(n7129), .B(n7128), .ZN(n7130)
         );
  AOI21_X1 U9006 ( .B1(n7182), .B2(n9931), .A(n7130), .ZN(n7131) );
  OAI21_X1 U9007 ( .B1(n7132), .B2(n9910), .A(n7131), .ZN(P1_U3285) );
  INV_X1 U9008 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10131) );
  INV_X1 U9009 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9887) );
  INV_X1 U9010 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8410) );
  AOI22_X1 U9011 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n9887), .B2(n8410), .ZN(n10137) );
  NOR2_X1 U9012 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7133) );
  AOI21_X1 U9013 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7133), .ZN(n10140) );
  INV_X1 U9014 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8377) );
  INV_X1 U9015 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9860) );
  AOI22_X1 U9016 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .B1(n8377), .B2(n9860), .ZN(n10143) );
  NOR2_X1 U9017 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7134) );
  AOI21_X1 U9018 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7134), .ZN(n10146) );
  NOR2_X1 U9019 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7135) );
  AOI21_X1 U9020 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7135), .ZN(n10149) );
  NOR2_X1 U9021 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7136) );
  AOI21_X1 U9022 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7136), .ZN(n10152) );
  NOR2_X1 U9023 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7137) );
  AOI21_X1 U9024 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7137), .ZN(n10155) );
  NOR2_X1 U9025 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7138) );
  AOI21_X1 U9026 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7138), .ZN(n10158) );
  NOR2_X1 U9027 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7139) );
  AOI21_X1 U9028 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7139), .ZN(n10167) );
  NOR2_X1 U9029 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7140) );
  AOI21_X1 U9030 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7140), .ZN(n10173) );
  NOR2_X1 U9031 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(P2_ADDR_REG_7__SCAN_IN), 
        .ZN(n7141) );
  AOI21_X1 U9032 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n7141), .ZN(n10170) );
  NOR2_X1 U9033 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7142) );
  AOI21_X1 U9034 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7142), .ZN(n10161) );
  NOR2_X1 U9035 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7143) );
  AOI21_X1 U9036 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7143), .ZN(n10164) );
  AND2_X1 U9037 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7144) );
  NOR2_X1 U9038 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7144), .ZN(n10126) );
  INV_X1 U9039 ( .A(n10126), .ZN(n10127) );
  INV_X1 U9040 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10129) );
  NAND3_X1 U9041 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10128) );
  NAND2_X1 U9042 ( .A1(n10129), .A2(n10128), .ZN(n10125) );
  NAND2_X1 U9043 ( .A1(n10127), .A2(n10125), .ZN(n10176) );
  NAND2_X1 U9044 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7145) );
  OAI21_X1 U9045 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7145), .ZN(n10175) );
  NOR2_X1 U9046 ( .A1(n10176), .A2(n10175), .ZN(n10174) );
  AOI21_X1 U9047 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10174), .ZN(n10179) );
  NAND2_X1 U9048 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7146) );
  OAI21_X1 U9049 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7146), .ZN(n10178) );
  NOR2_X1 U9050 ( .A1(n10179), .A2(n10178), .ZN(n10177) );
  AOI21_X1 U9051 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10177), .ZN(n10182) );
  NOR2_X1 U9052 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n7147) );
  AOI21_X1 U9053 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n7147), .ZN(n10181) );
  NAND2_X1 U9054 ( .A1(n10182), .A2(n10181), .ZN(n10180) );
  OAI21_X1 U9055 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10180), .ZN(n10163) );
  NAND2_X1 U9056 ( .A1(n10164), .A2(n10163), .ZN(n10162) );
  OAI21_X1 U9057 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10162), .ZN(n10160) );
  NAND2_X1 U9058 ( .A1(n10161), .A2(n10160), .ZN(n10159) );
  OAI21_X1 U9059 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10159), .ZN(n10169) );
  NAND2_X1 U9060 ( .A1(n10170), .A2(n10169), .ZN(n10168) );
  OAI21_X1 U9061 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n10168), .ZN(n10172) );
  NAND2_X1 U9062 ( .A1(n10173), .A2(n10172), .ZN(n10171) );
  OAI21_X1 U9063 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10171), .ZN(n10166) );
  NAND2_X1 U9064 ( .A1(n10167), .A2(n10166), .ZN(n10165) );
  OAI21_X1 U9065 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10165), .ZN(n10157) );
  NAND2_X1 U9066 ( .A1(n10158), .A2(n10157), .ZN(n10156) );
  OAI21_X1 U9067 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10156), .ZN(n10154) );
  NAND2_X1 U9068 ( .A1(n10155), .A2(n10154), .ZN(n10153) );
  OAI21_X1 U9069 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10153), .ZN(n10151) );
  NAND2_X1 U9070 ( .A1(n10152), .A2(n10151), .ZN(n10150) );
  OAI21_X1 U9071 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10150), .ZN(n10148) );
  NAND2_X1 U9072 ( .A1(n10149), .A2(n10148), .ZN(n10147) );
  OAI21_X1 U9073 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10147), .ZN(n10145) );
  NAND2_X1 U9074 ( .A1(n10146), .A2(n10145), .ZN(n10144) );
  OAI21_X1 U9075 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10144), .ZN(n10142) );
  NAND2_X1 U9076 ( .A1(n10143), .A2(n10142), .ZN(n10141) );
  OAI21_X1 U9077 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10141), .ZN(n10139) );
  NAND2_X1 U9078 ( .A1(n10140), .A2(n10139), .ZN(n10138) );
  OAI21_X1 U9079 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10138), .ZN(n10136) );
  NAND2_X1 U9080 ( .A1(n10137), .A2(n10136), .ZN(n10135) );
  OAI21_X1 U9081 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10135), .ZN(n10132) );
  NOR2_X1 U9082 ( .A1(n10131), .A2(n10132), .ZN(n7148) );
  NAND2_X1 U9083 ( .A1(n10131), .A2(n10132), .ZN(n10130) );
  OAI21_X1 U9084 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7148), .A(n10130), .ZN(
        n7151) );
  XNOR2_X1 U9085 ( .A(n7149), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7150) );
  XNOR2_X1 U9086 ( .A(n7151), .B(n7150), .ZN(ADD_1068_U4) );
  OAI211_X1 U9087 ( .C1(n4413), .C2(n7153), .A(n7152), .B(n8320), .ZN(n7159)
         );
  INV_X1 U9088 ( .A(n7154), .ZN(n7157) );
  NAND2_X1 U9089 ( .A1(n8329), .A2(n8344), .ZN(n7155) );
  OAI21_X1 U9090 ( .B1(n10038), .B2(n8324), .A(n7155), .ZN(n7156) );
  AOI211_X1 U9091 ( .C1(n10080), .C2(n8303), .A(n7157), .B(n7156), .ZN(n7158)
         );
  OAI211_X1 U9092 ( .C1(n10041), .C2(n8326), .A(n7159), .B(n7158), .ZN(
        P2_U3179) );
  OAI21_X1 U9093 ( .B1(n7162), .B2(n7161), .A(n7160), .ZN(n7190) );
  INV_X1 U9094 ( .A(n7190), .ZN(n7175) );
  OAI21_X1 U9095 ( .B1(n8995), .B2(n7164), .A(n7163), .ZN(n7166) );
  OAI22_X1 U9096 ( .A1(n7205), .A2(n9583), .B1(n6509), .B2(n4308), .ZN(n7165)
         );
  AOI21_X1 U9097 ( .B1(n7166), .B2(n9592), .A(n7165), .ZN(n7167) );
  OAI21_X1 U9098 ( .B1(n7175), .B2(n9589), .A(n7167), .ZN(n7188) );
  NAND2_X1 U9099 ( .A1(n7188), .A2(n9922), .ZN(n7174) );
  AOI211_X1 U9100 ( .C1(n7208), .C2(n7169), .A(n9548), .B(n4521), .ZN(n7189)
         );
  NOR2_X1 U9101 ( .A1(n9913), .A2(n4462), .ZN(n7172) );
  OAI22_X1 U9102 ( .A1(n9922), .A2(n7170), .B1(n7204), .B2(n9920), .ZN(n7171)
         );
  AOI211_X1 U9103 ( .C1(n7189), .C2(n9905), .A(n7172), .B(n7171), .ZN(n7173)
         );
  OAI211_X1 U9104 ( .C1(n7175), .C2(n9600), .A(n7174), .B(n7173), .ZN(P1_U3286) );
  INV_X1 U9105 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7177) );
  INV_X1 U9106 ( .A(n7176), .ZN(n7179) );
  INV_X1 U9107 ( .A(n9870), .ZN(n9337) );
  OAI222_X1 U9108 ( .A1(n9766), .A2(n7177), .B1(n9769), .B2(n7179), .C1(
        P1_U3086), .C2(n9337), .ZN(P1_U3339) );
  INV_X1 U9109 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n8162) );
  OAI222_X1 U9110 ( .A1(n8800), .A2(n8162), .B1(n8788), .B2(n7179), .C1(
        P2_U3151), .C2(n7178), .ZN(P2_U3279) );
  AOI211_X1 U9111 ( .C1(n9944), .C2(n7182), .A(n7181), .B(n7180), .ZN(n7187)
         );
  INV_X1 U9112 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7183) );
  OAI22_X1 U9113 ( .A1(n4520), .A2(n9747), .B1(n9946), .B2(n7183), .ZN(n7184)
         );
  INV_X1 U9114 ( .A(n7184), .ZN(n7185) );
  OAI21_X1 U9115 ( .B1(n7187), .B2(n9955), .A(n7185), .ZN(P1_U3477) );
  AOI22_X1 U9116 ( .A1(n7619), .A2(n8857), .B1(n9957), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n7186) );
  OAI21_X1 U9117 ( .B1(n7187), .B2(n9957), .A(n7186), .ZN(P1_U3530) );
  AOI211_X1 U9118 ( .C1(n7514), .C2(n7190), .A(n7189), .B(n7188), .ZN(n7195)
         );
  INV_X1 U9119 ( .A(n9747), .ZN(n7617) );
  INV_X1 U9120 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7191) );
  NOR2_X1 U9121 ( .A1(n9946), .A2(n7191), .ZN(n7192) );
  AOI21_X1 U9122 ( .B1(n7617), .B2(n7208), .A(n7192), .ZN(n7193) );
  OAI21_X1 U9123 ( .B1(n7195), .B2(n9955), .A(n7193), .ZN(P1_U3474) );
  AOI22_X1 U9124 ( .A1(n7619), .A2(n7208), .B1(n9957), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7194) );
  OAI21_X1 U9125 ( .B1(n7195), .B2(n9957), .A(n7194), .ZN(P1_U3529) );
  INV_X1 U9126 ( .A(n7196), .ZN(n7199) );
  AOI22_X1 U9127 ( .A1(n8412), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n8786), .ZN(n7197) );
  OAI21_X1 U9128 ( .B1(n7199), .B2(n8788), .A(n7197), .ZN(P2_U3278) );
  AOI22_X1 U9129 ( .A1(n9882), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9759), .ZN(n7198) );
  OAI21_X1 U9130 ( .B1(n7199), .B2(n9769), .A(n7198), .ZN(P1_U3338) );
  XNOR2_X1 U9131 ( .A(n7201), .B(n7200), .ZN(n7202) );
  XNOR2_X1 U9132 ( .A(n4407), .B(n7202), .ZN(n7210) );
  INV_X1 U9133 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7203) );
  OAI22_X1 U9134 ( .A1(n9810), .A2(n7204), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7203), .ZN(n7207) );
  OAI22_X1 U9135 ( .A1(n8967), .A2(n7205), .B1(n6509), .B2(n8964), .ZN(n7206)
         );
  AOI211_X1 U9136 ( .C1(n7208), .C2(n8957), .A(n7207), .B(n7206), .ZN(n7209)
         );
  OAI21_X1 U9137 ( .B1(n7210), .B2(n8946), .A(n7209), .ZN(P1_U3213) );
  OAI21_X1 U9138 ( .B1(n7211), .B2(n7214), .A(n7212), .ZN(n7220) );
  AOI22_X1 U9139 ( .A1(n8283), .A2(n8341), .B1(n8329), .B2(n8343), .ZN(n7218)
         );
  INV_X1 U9140 ( .A(n7215), .ZN(n7216) );
  AOI21_X1 U9141 ( .B1(n8303), .B2(n7344), .A(n7216), .ZN(n7217) );
  OAI211_X1 U9142 ( .C1(n8326), .C2(n7342), .A(n7218), .B(n7217), .ZN(n7219)
         );
  AOI21_X1 U9143 ( .B1(n7220), .B2(n8320), .A(n7219), .ZN(n7221) );
  INV_X1 U9144 ( .A(n7221), .ZN(P2_U3153) );
  INV_X1 U9145 ( .A(n7222), .ZN(n7292) );
  AOI22_X1 U9146 ( .A1(n9900), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9759), .ZN(n7223) );
  OAI21_X1 U9147 ( .B1(n7292), .B2(n9769), .A(n7223), .ZN(P1_U3337) );
  OAI21_X1 U9148 ( .B1(n7225), .B2(n7235), .A(n7224), .ZN(n9606) );
  NAND2_X1 U9149 ( .A1(n7226), .A2(n9610), .ZN(n7227) );
  NAND2_X1 U9150 ( .A1(n7227), .A2(n9698), .ZN(n7231) );
  NAND2_X1 U9151 ( .A1(n9247), .A2(n9563), .ZN(n7229) );
  NAND2_X1 U9152 ( .A1(n9245), .A2(n4309), .ZN(n7228) );
  NAND2_X1 U9153 ( .A1(n7229), .A2(n7228), .ZN(n7398) );
  INV_X1 U9154 ( .A(n7398), .ZN(n7230) );
  OAI21_X1 U9155 ( .B1(n7270), .B2(n7231), .A(n7230), .ZN(n9611) );
  INV_X1 U9156 ( .A(n9000), .ZN(n7232) );
  OAI21_X1 U9157 ( .B1(n7233), .B2(n7232), .A(n8997), .ZN(n7234) );
  XOR2_X1 U9158 ( .A(n7235), .B(n7234), .Z(n7236) );
  NOR2_X1 U9159 ( .A1(n7236), .A2(n9544), .ZN(n9605) );
  AOI211_X1 U9160 ( .C1(n9944), .C2(n9606), .A(n9611), .B(n9605), .ZN(n7241)
         );
  AOI22_X1 U9161 ( .A1(n9610), .A2(n7619), .B1(n9957), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7237) );
  OAI21_X1 U9162 ( .B1(n7241), .B2(n9957), .A(n7237), .ZN(P1_U3531) );
  INV_X1 U9163 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7238) );
  NOR2_X1 U9164 ( .A1(n9946), .A2(n7238), .ZN(n7239) );
  AOI21_X1 U9165 ( .B1(n9610), .B2(n7617), .A(n7239), .ZN(n7240) );
  OAI21_X1 U9166 ( .B1(n7241), .B2(n9955), .A(n7240), .ZN(P1_U3480) );
  NOR2_X1 U9167 ( .A1(n9331), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7242) );
  AOI21_X1 U9168 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9331), .A(n7242), .ZN(
        n7247) );
  NAND2_X1 U9169 ( .A1(n9780), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7243) );
  OAI21_X1 U9170 ( .B1(n9780), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7243), .ZN(
        n9773) );
  OAI21_X1 U9171 ( .B1(n7249), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7244), .ZN(
        n9774) );
  NOR2_X1 U9172 ( .A1(n9773), .A2(n9774), .ZN(n9772) );
  NAND2_X1 U9173 ( .A1(n9819), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7245) );
  OAI21_X1 U9174 ( .B1(n9819), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7245), .ZN(
        n9812) );
  NOR2_X1 U9175 ( .A1(n9813), .A2(n9812), .ZN(n9811) );
  AOI21_X1 U9176 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9819), .A(n9811), .ZN(
        n7246) );
  NAND2_X1 U9177 ( .A1(n7247), .A2(n7246), .ZN(n9330) );
  OAI21_X1 U9178 ( .B1(n7247), .B2(n7246), .A(n9330), .ZN(n7260) );
  OAI21_X1 U9179 ( .B1(n7249), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7248), .ZN(
        n9776) );
  MUX2_X1 U9180 ( .A(n7250), .B(P1_REG1_REG_10__SCAN_IN), .S(n9780), .Z(n9777)
         );
  NOR2_X1 U9181 ( .A1(n9776), .A2(n9777), .ZN(n9775) );
  MUX2_X1 U9182 ( .A(n7251), .B(P1_REG1_REG_11__SCAN_IN), .S(n9819), .Z(n9815)
         );
  NOR2_X1 U9183 ( .A1(n9816), .A2(n9815), .ZN(n9814) );
  AOI22_X1 U9184 ( .A1(n9331), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n5270), .B2(
        n7258), .ZN(n7252) );
  NAND2_X1 U9185 ( .A1(n7253), .A2(n7252), .ZN(n9319) );
  OAI21_X1 U9186 ( .B1(n7253), .B2(n7252), .A(n9319), .ZN(n7254) );
  NAND2_X1 U9187 ( .A1(n7254), .A2(n9880), .ZN(n7257) );
  NOR2_X1 U9188 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7255), .ZN(n9799) );
  AOI21_X1 U9189 ( .B1(n9866), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9799), .ZN(
        n7256) );
  OAI211_X1 U9190 ( .C1(n9343), .C2(n7258), .A(n7257), .B(n7256), .ZN(n7259)
         );
  AOI21_X1 U9191 ( .B1(n9883), .B2(n7260), .A(n7259), .ZN(n7261) );
  INV_X1 U9192 ( .A(n7261), .ZN(P1_U3255) );
  OAI21_X1 U9193 ( .B1(n7263), .B2(n9091), .A(n7262), .ZN(n7297) );
  INV_X1 U9194 ( .A(n7297), .ZN(n7278) );
  INV_X1 U9195 ( .A(n7264), .ZN(n7265) );
  AOI21_X1 U9196 ( .B1(n9091), .B2(n7266), .A(n7265), .ZN(n7269) );
  NAND2_X1 U9197 ( .A1(n9246), .A2(n9563), .ZN(n7268) );
  NAND2_X1 U9198 ( .A1(n9244), .A2(n4309), .ZN(n7267) );
  AND2_X1 U9199 ( .A1(n7268), .A2(n7267), .ZN(n7562) );
  OAI21_X1 U9200 ( .B1(n7269), .B2(n9544), .A(n7562), .ZN(n7295) );
  INV_X1 U9201 ( .A(n7270), .ZN(n7272) );
  INV_X1 U9202 ( .A(n7505), .ZN(n7271) );
  AOI211_X1 U9203 ( .C1(n7301), .C2(n7272), .A(n9548), .B(n7271), .ZN(n7296)
         );
  NAND2_X1 U9204 ( .A1(n7296), .A2(n9905), .ZN(n7275) );
  INV_X1 U9205 ( .A(n7273), .ZN(n7564) );
  AOI22_X1 U9206 ( .A1(n9934), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7564), .B2(
        n9908), .ZN(n7274) );
  OAI211_X1 U9207 ( .C1(n6514), .C2(n9913), .A(n7275), .B(n7274), .ZN(n7276)
         );
  AOI21_X1 U9208 ( .B1(n7295), .B2(n9922), .A(n7276), .ZN(n7277) );
  OAI21_X1 U9209 ( .B1(n7278), .B2(n9556), .A(n7277), .ZN(P1_U3283) );
  INV_X1 U9210 ( .A(n7280), .ZN(n7282) );
  NAND3_X1 U9211 ( .A1(n7212), .A2(n7282), .A3(n7281), .ZN(n7283) );
  AOI21_X1 U9212 ( .B1(n7279), .B2(n7283), .A(n8305), .ZN(n7291) );
  INV_X1 U9213 ( .A(n7366), .ZN(n7284) );
  NAND2_X1 U9214 ( .A1(n8317), .A2(n7284), .ZN(n7289) );
  NAND2_X1 U9215 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10028) );
  INV_X1 U9216 ( .A(n10028), .ZN(n7285) );
  AOI21_X1 U9217 ( .B1(n8329), .B2(n8342), .A(n7285), .ZN(n7288) );
  NAND2_X1 U9218 ( .A1(n8303), .A2(n7368), .ZN(n7287) );
  OR2_X1 U9219 ( .A1(n7460), .A2(n8324), .ZN(n7286) );
  NAND4_X1 U9220 ( .A1(n7289), .A2(n7288), .A3(n7287), .A4(n7286), .ZN(n7290)
         );
  OR2_X1 U9221 ( .A1(n7291), .A2(n7290), .ZN(P2_U3161) );
  OAI222_X1 U9222 ( .A1(n8800), .A2(n7294), .B1(n7293), .B2(P2_U3151), .C1(
        n8803), .C2(n7292), .ZN(P2_U3277) );
  AOI211_X1 U9223 ( .C1(n7297), .C2(n9944), .A(n7296), .B(n7295), .ZN(n7303)
         );
  INV_X1 U9224 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7298) );
  OAI22_X1 U9225 ( .A1(n6514), .A2(n9747), .B1(n9946), .B2(n7298), .ZN(n7299)
         );
  INV_X1 U9226 ( .A(n7299), .ZN(n7300) );
  OAI21_X1 U9227 ( .B1(n7303), .B2(n9955), .A(n7300), .ZN(P1_U3483) );
  AOI22_X1 U9228 ( .A1(n7301), .A2(n7619), .B1(n9957), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7302) );
  OAI21_X1 U9229 ( .B1(n7303), .B2(n9957), .A(n7302), .ZN(P1_U3532) );
  AOI21_X1 U9230 ( .B1(n7306), .B2(n7305), .A(n7304), .ZN(n7320) );
  INV_X1 U9231 ( .A(n7307), .ZN(n7308) );
  OAI21_X1 U9232 ( .B1(n7309), .B2(P2_REG1_REG_9__SCAN_IN), .A(n7308), .ZN(
        n7318) );
  AND2_X1 U9233 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7444) );
  AOI21_X1 U9234 ( .B1(n10013), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7444), .ZN(
        n7310) );
  OAI21_X1 U9235 ( .B1(n7312), .B2(n7311), .A(n7310), .ZN(n7317) );
  AOI21_X1 U9236 ( .B1(n7314), .B2(n7355), .A(n7313), .ZN(n7315) );
  NOR2_X1 U9237 ( .A1(n7315), .A2(n10024), .ZN(n7316) );
  AOI211_X1 U9238 ( .C1(n10014), .C2(n7318), .A(n7317), .B(n7316), .ZN(n7319)
         );
  OAI21_X1 U9239 ( .B1(n7320), .B2(n10019), .A(n7319), .ZN(P2_U3191) );
  OR2_X1 U9240 ( .A1(n8449), .A2(n10100), .ZN(n7321) );
  OAI22_X1 U9241 ( .A1(n10043), .A2(n7323), .B1(n10040), .B2(n7322), .ZN(n7326) );
  NOR2_X1 U9242 ( .A1(n7324), .A2(n8634), .ZN(n7325) );
  AOI211_X1 U9243 ( .C1(n8634), .C2(P2_REG2_REG_1__SCAN_IN), .A(n7326), .B(
        n7325), .ZN(n7327) );
  OAI21_X1 U9244 ( .B1(n10047), .B2(n7328), .A(n7327), .ZN(P2_U3232) );
  AND2_X1 U9245 ( .A1(n7768), .A2(n7783), .ZN(n7928) );
  XNOR2_X1 U9246 ( .A(n7329), .B(n7928), .ZN(n10069) );
  INV_X1 U9247 ( .A(n10069), .ZN(n7338) );
  XOR2_X1 U9248 ( .A(n7928), .B(n7330), .Z(n7331) );
  AOI222_X1 U9249 ( .A1(n8627), .A2(n7331), .B1(n8344), .B2(n8622), .C1(n6209), 
        .C2(n8624), .ZN(n10066) );
  MUX2_X1 U9250 ( .A(n7332), .B(n10066), .S(n8616), .Z(n7337) );
  INV_X1 U9251 ( .A(n7333), .ZN(n7334) );
  AOI22_X1 U9252 ( .A1(n8605), .A2(n7335), .B1(n8604), .B2(n7334), .ZN(n7336)
         );
  OAI211_X1 U9253 ( .C1(n10047), .C2(n7338), .A(n7337), .B(n7336), .ZN(
        P2_U3229) );
  INV_X1 U9254 ( .A(n7364), .ZN(n7340) );
  AOI21_X1 U9255 ( .B1(n7346), .B2(n7341), .A(n7340), .ZN(n10087) );
  INV_X1 U9256 ( .A(n10087), .ZN(n10084) );
  OAI22_X1 U9257 ( .A1(n8616), .A2(n5926), .B1(n7342), .B2(n10040), .ZN(n7343)
         );
  AOI21_X1 U9258 ( .B1(n8605), .B2(n7344), .A(n7343), .ZN(n7351) );
  INV_X1 U9259 ( .A(n7346), .ZN(n7934) );
  XNOR2_X1 U9260 ( .A(n7345), .B(n7934), .ZN(n7347) );
  NAND2_X1 U9261 ( .A1(n7347), .A2(n8627), .ZN(n7349) );
  AOI22_X1 U9262 ( .A1(n8343), .A2(n8624), .B1(n8622), .B2(n8341), .ZN(n7348)
         );
  NAND2_X1 U9263 ( .A1(n7349), .A2(n7348), .ZN(n10086) );
  NAND2_X1 U9264 ( .A1(n10086), .A2(n8616), .ZN(n7350) );
  OAI211_X1 U9265 ( .C1(n10084), .C2(n10047), .A(n7351), .B(n7350), .ZN(
        P2_U3226) );
  INV_X1 U9266 ( .A(n7352), .ZN(n7353) );
  AOI21_X1 U9267 ( .B1(n7354), .B2(n7938), .A(n7353), .ZN(n10099) );
  INV_X1 U9268 ( .A(n10099), .ZN(n10096) );
  OAI22_X1 U9269 ( .A1(n8616), .A2(n7355), .B1(n7442), .B2(n10040), .ZN(n7356)
         );
  AOI21_X1 U9270 ( .B1(n8605), .B2(n7453), .A(n7356), .ZN(n7362) );
  XNOR2_X1 U9271 ( .A(n7357), .B(n7938), .ZN(n7358) );
  NAND2_X1 U9272 ( .A1(n7358), .A2(n8627), .ZN(n7360) );
  AOI22_X1 U9273 ( .A1(n8624), .A2(n8341), .B1(n8339), .B2(n8622), .ZN(n7359)
         );
  NAND2_X1 U9274 ( .A1(n7360), .A2(n7359), .ZN(n10098) );
  NAND2_X1 U9275 ( .A1(n10098), .A2(n8616), .ZN(n7361) );
  OAI211_X1 U9276 ( .C1(n10096), .C2(n10047), .A(n7362), .B(n7361), .ZN(
        P2_U3224) );
  NAND2_X1 U9277 ( .A1(n7791), .A2(n7775), .ZN(n7936) );
  NAND2_X1 U9278 ( .A1(n7364), .A2(n7363), .ZN(n7365) );
  XOR2_X1 U9279 ( .A(n7936), .B(n7365), .Z(n10091) );
  OAI22_X1 U9280 ( .A1(n8616), .A2(n6382), .B1(n7366), .B2(n10040), .ZN(n7367)
         );
  AOI21_X1 U9281 ( .B1(n8605), .B2(n7368), .A(n7367), .ZN(n7375) );
  INV_X1 U9282 ( .A(n7936), .ZN(n7370) );
  XNOR2_X1 U9283 ( .A(n7369), .B(n7370), .ZN(n7371) );
  NAND2_X1 U9284 ( .A1(n7371), .A2(n8627), .ZN(n7373) );
  AOI22_X1 U9285 ( .A1(n8342), .A2(n8624), .B1(n8622), .B2(n8340), .ZN(n7372)
         );
  NAND2_X1 U9286 ( .A1(n7373), .A2(n7372), .ZN(n10092) );
  NAND2_X1 U9287 ( .A1(n10092), .A2(n8616), .ZN(n7374) );
  OAI211_X1 U9288 ( .C1(n10091), .C2(n10047), .A(n7375), .B(n7374), .ZN(
        P2_U3225) );
  NAND3_X1 U9289 ( .A1(n7377), .A2(n7758), .A3(n7376), .ZN(n7378) );
  AND2_X1 U9290 ( .A1(n7379), .A2(n7378), .ZN(n10062) );
  NAND3_X1 U9291 ( .A1(n7381), .A2(n7929), .A3(n7380), .ZN(n7382) );
  NAND2_X1 U9292 ( .A1(n7383), .A2(n7382), .ZN(n7384) );
  AOI222_X1 U9293 ( .A1(n8627), .A2(n7384), .B1(n8345), .B2(n8622), .C1(n8346), 
        .C2(n8624), .ZN(n10060) );
  MUX2_X1 U9294 ( .A(n7385), .B(n10060), .S(n8616), .Z(n7389) );
  INV_X1 U9295 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7386) );
  AOI22_X1 U9296 ( .A1(n8605), .A2(n7387), .B1(n8604), .B2(n7386), .ZN(n7388)
         );
  OAI211_X1 U9297 ( .C1(n10062), .C2(n10047), .A(n7389), .B(n7388), .ZN(
        P2_U3230) );
  INV_X1 U9298 ( .A(n7390), .ZN(n7392) );
  OAI222_X1 U9299 ( .A1(n8800), .A2(n7391), .B1(n8803), .B2(n7392), .C1(
        P2_U3151), .C2(n4314), .ZN(P2_U3276) );
  OAI222_X1 U9300 ( .A1(n9766), .A2(n7393), .B1(n9769), .B2(n7392), .C1(
        P1_U3086), .C2(n4315), .ZN(P1_U3336) );
  INV_X1 U9301 ( .A(n7394), .ZN(n7395) );
  NOR2_X1 U9302 ( .A1(n7396), .A2(n7395), .ZN(n7397) );
  XNOR2_X1 U9303 ( .A(n4408), .B(n7397), .ZN(n7403) );
  NAND2_X1 U9304 ( .A1(n9801), .A2(n7398), .ZN(n7400) );
  OAI211_X1 U9305 ( .C1(n9810), .C2(n9608), .A(n7400), .B(n7399), .ZN(n7401)
         );
  AOI21_X1 U9306 ( .B1(n9610), .B2(n8957), .A(n7401), .ZN(n7402) );
  OAI21_X1 U9307 ( .B1(n7403), .B2(n8946), .A(n7402), .ZN(P1_U3231) );
  INV_X1 U9308 ( .A(n10030), .ZN(n7405) );
  OR2_X1 U9309 ( .A1(n7405), .A2(n7767), .ZN(n7930) );
  XNOR2_X1 U9310 ( .A(n7404), .B(n7930), .ZN(n7406) );
  AOI222_X1 U9311 ( .A1(n8627), .A2(n7406), .B1(n8343), .B2(n8622), .C1(n8345), 
        .C2(n8624), .ZN(n10071) );
  XOR2_X1 U9312 ( .A(n7407), .B(n7930), .Z(n10075) );
  INV_X1 U9313 ( .A(n10047), .ZN(n7412) );
  NOR2_X1 U9314 ( .A1(n8616), .A2(n7408), .ZN(n7411) );
  OAI22_X1 U9315 ( .A1(n10043), .A2(n10072), .B1(n7409), .B2(n10040), .ZN(
        n7410) );
  AOI211_X1 U9316 ( .C1(n10075), .C2(n7412), .A(n7411), .B(n7410), .ZN(n7413)
         );
  OAI21_X1 U9317 ( .B1(n10071), .B2(n8634), .A(n7413), .ZN(P2_U3228) );
  OAI211_X1 U9318 ( .C1(n7415), .C2(n9104), .A(n4441), .B(n9592), .ZN(n7419)
         );
  NAND2_X1 U9319 ( .A1(n9244), .A2(n9563), .ZN(n7417) );
  NAND2_X1 U9320 ( .A1(n9242), .A2(n4309), .ZN(n7416) );
  NAND2_X1 U9321 ( .A1(n7417), .A2(n7416), .ZN(n9800) );
  INV_X1 U9322 ( .A(n9800), .ZN(n7418) );
  NAND2_X1 U9323 ( .A1(n7419), .A2(n7418), .ZN(n7431) );
  INV_X1 U9324 ( .A(n7431), .ZN(n7430) );
  OAI21_X1 U9325 ( .B1(n7422), .B2(n7421), .A(n7420), .ZN(n7433) );
  NAND2_X1 U9326 ( .A1(n7433), .A2(n9931), .ZN(n7429) );
  INV_X1 U9327 ( .A(n7504), .ZN(n7424) );
  INV_X1 U9328 ( .A(n7491), .ZN(n7423) );
  AOI211_X1 U9329 ( .C1(n7434), .C2(n7424), .A(n9548), .B(n7423), .ZN(n7432)
         );
  NOR2_X1 U9330 ( .A1(n9804), .A2(n9913), .ZN(n7427) );
  OAI22_X1 U9331 ( .A1(n9922), .A2(n7425), .B1(n9809), .B2(n9920), .ZN(n7426)
         );
  AOI211_X1 U9332 ( .C1(n7432), .C2(n9905), .A(n7427), .B(n7426), .ZN(n7428)
         );
  OAI211_X1 U9333 ( .C1(n9910), .C2(n7430), .A(n7429), .B(n7428), .ZN(P1_U3281) );
  AOI211_X1 U9334 ( .C1(n7433), .C2(n9944), .A(n7432), .B(n7431), .ZN(n7439)
         );
  AOI22_X1 U9335 ( .A1(n7434), .A2(n7619), .B1(n9957), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7435) );
  OAI21_X1 U9336 ( .B1(n7439), .B2(n9957), .A(n7435), .ZN(P1_U3534) );
  INV_X1 U9337 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7436) );
  OAI22_X1 U9338 ( .A1(n9804), .A2(n9747), .B1(n9946), .B2(n7436), .ZN(n7437)
         );
  INV_X1 U9339 ( .A(n7437), .ZN(n7438) );
  OAI21_X1 U9340 ( .B1(n7439), .B2(n9955), .A(n7438), .ZN(P1_U3489) );
  INV_X1 U9341 ( .A(n7440), .ZN(n7456) );
  OAI222_X1 U9342 ( .A1(n8803), .A2(n7456), .B1(n7441), .B2(P2_U3151), .C1(
        n8164), .C2(n8800), .ZN(P2_U3275) );
  INV_X1 U9343 ( .A(n7442), .ZN(n7443) );
  NAND2_X1 U9344 ( .A1(n8317), .A2(n7443), .ZN(n7446) );
  AOI21_X1 U9345 ( .B1(n8329), .B2(n8341), .A(n7444), .ZN(n7445) );
  OAI211_X1 U9346 ( .C1(n8287), .C2(n8324), .A(n7446), .B(n7445), .ZN(n7452)
         );
  INV_X1 U9347 ( .A(n7448), .ZN(n7449) );
  AOI211_X1 U9348 ( .C1(n7450), .C2(n7447), .A(n8305), .B(n7449), .ZN(n7451)
         );
  AOI211_X1 U9349 ( .C1(n7453), .C2(n8303), .A(n7452), .B(n7451), .ZN(n7454)
         );
  INV_X1 U9350 ( .A(n7454), .ZN(P2_U3171) );
  INV_X1 U9351 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7455) );
  OAI222_X1 U9352 ( .A1(P1_U3086), .A2(n9126), .B1(n9769), .B2(n7456), .C1(
        n7455), .C2(n9766), .ZN(P1_U3335) );
  NAND2_X1 U9353 ( .A1(n7799), .A2(n7798), .ZN(n7937) );
  XOR2_X1 U9354 ( .A(n7937), .B(n7458), .Z(n10105) );
  XNOR2_X1 U9355 ( .A(n7459), .B(n7937), .ZN(n7462) );
  OAI22_X1 U9356 ( .A1(n7460), .A2(n10037), .B1(n7535), .B2(n10039), .ZN(n7461) );
  AOI21_X1 U9357 ( .B1(n7462), .B2(n8627), .A(n7461), .ZN(n7463) );
  OAI21_X1 U9358 ( .B1(n10105), .B2(n6485), .A(n7463), .ZN(n10107) );
  NAND2_X1 U9359 ( .A1(n10107), .A2(n8616), .ZN(n7468) );
  OAI22_X1 U9360 ( .A1(n8616), .A2(n7464), .B1(n7525), .B2(n10040), .ZN(n7465)
         );
  AOI21_X1 U9361 ( .B1(n8605), .B2(n7466), .A(n7465), .ZN(n7467) );
  OAI211_X1 U9362 ( .C1(n10105), .C2(n7469), .A(n7468), .B(n7467), .ZN(
        P2_U3223) );
  OAI21_X1 U9363 ( .B1(n7470), .B2(n7940), .A(n8627), .ZN(n7472) );
  OR2_X1 U9364 ( .A1(n7472), .A2(n4547), .ZN(n7474) );
  AOI22_X1 U9365 ( .A1(n8622), .A2(n8625), .B1(n8339), .B2(n8624), .ZN(n7473)
         );
  NAND2_X1 U9366 ( .A1(n7474), .A2(n7473), .ZN(n7481) );
  MUX2_X1 U9367 ( .A(n7481), .B(P2_REG0_REG_11__SCAN_IN), .S(n10108), .Z(n7477) );
  XNOR2_X1 U9368 ( .A(n7475), .B(n7940), .ZN(n7486) );
  INV_X1 U9369 ( .A(n8294), .ZN(n7478) );
  OAI22_X1 U9370 ( .A1(n7486), .A2(n8782), .B1(n7478), .B2(n8766), .ZN(n7476)
         );
  OR2_X1 U9371 ( .A1(n7477), .A2(n7476), .ZN(P2_U3423) );
  MUX2_X1 U9372 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7481), .S(n10124), .Z(n7480) );
  OAI22_X1 U9373 ( .A1(n7486), .A2(n8694), .B1(n7478), .B2(n8656), .ZN(n7479)
         );
  OR2_X1 U9374 ( .A1(n7480), .A2(n7479), .ZN(P2_U3470) );
  MUX2_X1 U9375 ( .A(n7481), .B(P2_REG2_REG_11__SCAN_IN), .S(n8634), .Z(n7482)
         );
  INV_X1 U9376 ( .A(n7482), .ZN(n7485) );
  INV_X1 U9377 ( .A(n7483), .ZN(n8284) );
  AOI22_X1 U9378 ( .A1(n8605), .A2(n8294), .B1(n8604), .B2(n8284), .ZN(n7484)
         );
  OAI211_X1 U9379 ( .C1(n7486), .C2(n10047), .A(n7485), .B(n7484), .ZN(
        P2_U3222) );
  OAI21_X1 U9380 ( .B1(n7488), .B2(n9106), .A(n7487), .ZN(n7489) );
  INV_X1 U9381 ( .A(n7489), .ZN(n9702) );
  INV_X1 U9382 ( .A(n9595), .ZN(n7490) );
  AOI21_X1 U9383 ( .B1(n9697), .B2(n7491), .A(n7490), .ZN(n9699) );
  INV_X1 U9384 ( .A(n7492), .ZN(n7589) );
  AOI22_X1 U9385 ( .A1(n9934), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7589), .B2(
        n9908), .ZN(n7493) );
  OAI21_X1 U9386 ( .B1(n4531), .B2(n9913), .A(n7493), .ZN(n7499) );
  OAI21_X1 U9387 ( .B1(n7496), .B2(n7495), .A(n7494), .ZN(n7497) );
  AOI222_X1 U9388 ( .A1(n9592), .A2(n7497), .B1(n9243), .B2(n9563), .C1(n9241), 
        .C2(n4309), .ZN(n9701) );
  NOR2_X1 U9389 ( .A1(n9701), .A2(n9910), .ZN(n7498) );
  AOI211_X1 U9390 ( .C1(n9699), .C2(n9603), .A(n7499), .B(n7498), .ZN(n7500)
         );
  OAI21_X1 U9391 ( .B1(n9702), .B2(n9556), .A(n7500), .ZN(P1_U3280) );
  INV_X1 U9392 ( .A(n7501), .ZN(n7520) );
  OAI222_X1 U9393 ( .A1(n8803), .A2(n7520), .B1(n7749), .B2(P2_U3151), .C1(
        n8239), .C2(n8800), .ZN(P2_U3274) );
  OAI21_X1 U9394 ( .B1(n7503), .B2(n7506), .A(n7502), .ZN(n9917) );
  AOI211_X1 U9395 ( .C1(n7632), .C2(n7505), .A(n9548), .B(n7504), .ZN(n9906)
         );
  XNOR2_X1 U9396 ( .A(n7507), .B(n7506), .ZN(n7508) );
  NOR2_X1 U9397 ( .A1(n7508), .A2(n9544), .ZN(n7511) );
  NAND2_X1 U9398 ( .A1(n9243), .A2(n4309), .ZN(n7510) );
  NAND2_X1 U9399 ( .A1(n9245), .A2(n9563), .ZN(n7509) );
  NAND2_X1 U9400 ( .A1(n7510), .A2(n7509), .ZN(n7629) );
  AOI211_X1 U9401 ( .C1(n9917), .C2(n7512), .A(n7511), .B(n7629), .ZN(n9919)
         );
  INV_X1 U9402 ( .A(n9919), .ZN(n7513) );
  AOI211_X1 U9403 ( .C1(n7514), .C2(n9917), .A(n9906), .B(n7513), .ZN(n7519)
         );
  INV_X1 U9404 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7515) );
  OAI22_X1 U9405 ( .A1(n9914), .A2(n9747), .B1(n9946), .B2(n7515), .ZN(n7516)
         );
  INV_X1 U9406 ( .A(n7516), .ZN(n7517) );
  OAI21_X1 U9407 ( .B1(n7519), .B2(n9955), .A(n7517), .ZN(P1_U3486) );
  AOI22_X1 U9408 ( .A1(n7632), .A2(n7619), .B1(n9957), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7518) );
  OAI21_X1 U9409 ( .B1(n7519), .B2(n9957), .A(n7518), .ZN(P1_U3533) );
  OAI222_X1 U9410 ( .A1(P1_U3086), .A2(n4316), .B1(n9769), .B2(n7520), .C1(
        n8221), .C2(n9766), .ZN(P1_U3334) );
  OAI21_X1 U9411 ( .B1(n7521), .B2(n7523), .A(n7522), .ZN(n7524) );
  NAND2_X1 U9412 ( .A1(n7524), .A2(n8320), .ZN(n7532) );
  INV_X1 U9413 ( .A(n7525), .ZN(n7526) );
  NAND2_X1 U9414 ( .A1(n8317), .A2(n7526), .ZN(n7529) );
  INV_X1 U9415 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7527) );
  NOR2_X1 U9416 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7527), .ZN(n7545) );
  AOI21_X1 U9417 ( .B1(n8329), .B2(n8340), .A(n7545), .ZN(n7528) );
  OAI211_X1 U9418 ( .C1(n7535), .C2(n8324), .A(n7529), .B(n7528), .ZN(n7530)
         );
  INV_X1 U9419 ( .A(n7530), .ZN(n7531) );
  OAI211_X1 U9420 ( .C1(n10103), .C2(n8332), .A(n7532), .B(n7531), .ZN(
        P2_U3157) );
  XNOR2_X1 U9421 ( .A(n7533), .B(n7942), .ZN(n8783) );
  XNOR2_X1 U9422 ( .A(n4917), .B(n7942), .ZN(n7534) );
  OAI222_X1 U9423 ( .A1(n10039), .A2(n8612), .B1(n10037), .B2(n7535), .C1(
        n7534), .C2(n10050), .ZN(n8690) );
  NAND2_X1 U9424 ( .A1(n8690), .A2(n8616), .ZN(n7539) );
  OAI22_X1 U9425 ( .A1(n8616), .A2(n7536), .B1(n8069), .B2(n10040), .ZN(n7537)
         );
  AOI21_X1 U9426 ( .B1(n8605), .B2(n8691), .A(n7537), .ZN(n7538) );
  OAI211_X1 U9427 ( .C1(n8783), .C2(n10047), .A(n7539), .B(n7538), .ZN(
        P2_U3221) );
  AOI21_X1 U9428 ( .B1(n4410), .B2(n7541), .A(n7540), .ZN(n7556) );
  AOI21_X1 U9429 ( .B1(n7544), .B2(n7543), .A(n7542), .ZN(n7547) );
  AOI21_X1 U9430 ( .B1(n10013), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7545), .ZN(
        n7546) );
  OAI21_X1 U9431 ( .B1(n7547), .B2(n10019), .A(n7546), .ZN(n7553) );
  AOI21_X1 U9432 ( .B1(n7550), .B2(n7549), .A(n7548), .ZN(n7551) );
  NOR2_X1 U9433 ( .A1(n7551), .A2(n9967), .ZN(n7552) );
  AOI211_X1 U9434 ( .C1(n10011), .C2(n7554), .A(n7553), .B(n7552), .ZN(n7555)
         );
  OAI21_X1 U9435 ( .B1(n7556), .B2(n10024), .A(n7555), .ZN(P2_U3192) );
  XOR2_X1 U9436 ( .A(n7557), .B(n7626), .Z(n7560) );
  INV_X1 U9437 ( .A(n7558), .ZN(n7559) );
  NAND2_X1 U9438 ( .A1(n7560), .A2(n7559), .ZN(n7625) );
  OAI211_X1 U9439 ( .C1(n7560), .C2(n7559), .A(n7625), .B(n9806), .ZN(n7566)
         );
  OAI22_X1 U9440 ( .A1(n8955), .A2(n7562), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7561), .ZN(n7563) );
  AOI21_X1 U9441 ( .B1(n7564), .B2(n8971), .A(n7563), .ZN(n7565) );
  OAI211_X1 U9442 ( .C1(n6514), .C2(n9803), .A(n7566), .B(n7565), .ZN(P1_U3217) );
  XNOR2_X1 U9443 ( .A(n7567), .B(n9108), .ZN(n7616) );
  INV_X1 U9444 ( .A(n7616), .ZN(n7578) );
  INV_X1 U9445 ( .A(n9027), .ZN(n9167) );
  NOR2_X1 U9446 ( .A1(n9108), .A2(n9167), .ZN(n7571) );
  INV_X1 U9447 ( .A(n7568), .ZN(n7569) );
  AOI21_X1 U9448 ( .B1(n7571), .B2(n7570), .A(n7569), .ZN(n7572) );
  OAI222_X1 U9449 ( .A1(n4308), .A2(n8965), .B1(n9583), .B2(n8966), .C1(n9544), 
        .C2(n7572), .ZN(n7614) );
  INV_X1 U9450 ( .A(n7677), .ZN(n7573) );
  AOI211_X1 U9451 ( .C1(n8981), .C2(n4532), .A(n9548), .B(n7573), .ZN(n7615)
         );
  NAND2_X1 U9452 ( .A1(n7615), .A2(n9905), .ZN(n7575) );
  AOI22_X1 U9453 ( .A1(n9934), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8970), .B2(
        n9908), .ZN(n7574) );
  OAI211_X1 U9454 ( .C1(n8974), .C2(n9913), .A(n7575), .B(n7574), .ZN(n7576)
         );
  AOI21_X1 U9455 ( .B1(n7614), .B2(n9922), .A(n7576), .ZN(n7577) );
  OAI21_X1 U9456 ( .B1(n7578), .B2(n9556), .A(n7577), .ZN(P1_U3278) );
  INV_X1 U9457 ( .A(n7579), .ZN(n7710) );
  OAI222_X1 U9458 ( .A1(n8800), .A2(n7581), .B1(n8788), .B2(n7710), .C1(
        P2_U3151), .C2(n7580), .ZN(P2_U3273) );
  OAI21_X1 U9459 ( .B1(n7584), .B2(n7583), .A(n7582), .ZN(n7585) );
  NAND2_X1 U9460 ( .A1(n7585), .A2(n9806), .ZN(n7591) );
  NAND2_X1 U9461 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9832) );
  INV_X1 U9462 ( .A(n9832), .ZN(n7588) );
  OAI22_X1 U9463 ( .A1(n8967), .A2(n7586), .B1(n8966), .B2(n8964), .ZN(n7587)
         );
  AOI211_X1 U9464 ( .C1(n7589), .C2(n8971), .A(n7588), .B(n7587), .ZN(n7590)
         );
  OAI211_X1 U9465 ( .C1(n4531), .C2(n9803), .A(n7591), .B(n7590), .ZN(P1_U3234) );
  AOI21_X1 U9466 ( .B1(n7594), .B2(n7593), .A(n7592), .ZN(n7613) );
  INV_X1 U9467 ( .A(n7595), .ZN(n7596) );
  NAND2_X1 U9468 ( .A1(n7597), .A2(n7596), .ZN(n7598) );
  XNOR2_X1 U9469 ( .A(n7599), .B(n7598), .ZN(n7600) );
  NAND2_X1 U9470 ( .A1(n7600), .A2(n10001), .ZN(n7612) );
  INV_X1 U9471 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7603) );
  INV_X1 U9472 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7601) );
  NOR2_X1 U9473 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7601), .ZN(n8071) );
  INV_X1 U9474 ( .A(n8071), .ZN(n7602) );
  OAI21_X1 U9475 ( .B1(n9982), .B2(n7603), .A(n7602), .ZN(n7609) );
  AOI21_X1 U9476 ( .B1(n7606), .B2(n7605), .A(n7604), .ZN(n7607) );
  NOR2_X1 U9477 ( .A1(n7607), .A2(n10024), .ZN(n7608) );
  AOI211_X1 U9478 ( .C1(n10011), .C2(n7610), .A(n7609), .B(n7608), .ZN(n7611)
         );
  OAI211_X1 U9479 ( .C1(n7613), .C2(n9967), .A(n7612), .B(n7611), .ZN(P2_U3194) );
  AOI211_X1 U9480 ( .C1(n7616), .C2(n9944), .A(n7615), .B(n7614), .ZN(n7621)
         );
  AOI22_X1 U9481 ( .A1(n8981), .A2(n7617), .B1(P1_REG0_REG_15__SCAN_IN), .B2(
        n9955), .ZN(n7618) );
  OAI21_X1 U9482 ( .B1(n7621), .B2(n9955), .A(n7618), .ZN(P1_U3498) );
  AOI22_X1 U9483 ( .A1(n8981), .A2(n7619), .B1(P1_REG1_REG_15__SCAN_IN), .B2(
        n9957), .ZN(n7620) );
  OAI21_X1 U9484 ( .B1(n7621), .B2(n9957), .A(n7620), .ZN(P1_U3537) );
  OAI21_X1 U9485 ( .B1(n7624), .B2(n7623), .A(n7622), .ZN(n7628) );
  OAI21_X1 U9486 ( .B1(n7626), .B2(n7557), .A(n7625), .ZN(n7627) );
  XOR2_X1 U9487 ( .A(n7628), .B(n7627), .Z(n7634) );
  AOI22_X1 U9488 ( .A1(n9801), .A2(n7629), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n7630) );
  OAI21_X1 U9489 ( .B1(n9907), .B2(n9810), .A(n7630), .ZN(n7631) );
  AOI21_X1 U9490 ( .B1(n7632), .B2(n8957), .A(n7631), .ZN(n7633) );
  OAI21_X1 U9491 ( .B1(n7634), .B2(n8946), .A(n7633), .ZN(P1_U3236) );
  INV_X1 U9492 ( .A(n7637), .ZN(n7636) );
  NAND2_X1 U9493 ( .A1(n9759), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7635) );
  OAI211_X1 U9494 ( .C1(n7636), .C2(n9769), .A(n9123), .B(n7635), .ZN(P1_U3332) );
  NAND2_X1 U9495 ( .A1(n7637), .A2(n8795), .ZN(n7639) );
  OR2_X1 U9496 ( .A1(n7638), .A2(P2_U3151), .ZN(n7983) );
  OAI211_X1 U9497 ( .C1(n7640), .C2(n8800), .A(n7639), .B(n7983), .ZN(P2_U3272) );
  AOI21_X1 U9498 ( .B1(n7643), .B2(n7642), .A(n7641), .ZN(n7657) );
  AOI21_X1 U9499 ( .B1(n7646), .B2(n7645), .A(n7644), .ZN(n7648) );
  INV_X1 U9500 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8238) );
  NOR2_X1 U9501 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8238), .ZN(n8282) );
  AOI21_X1 U9502 ( .B1(n10013), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8282), .ZN(
        n7647) );
  OAI21_X1 U9503 ( .B1(n7648), .B2(n10019), .A(n7647), .ZN(n7654) );
  AOI21_X1 U9504 ( .B1(n7651), .B2(n7650), .A(n7649), .ZN(n7652) );
  NOR2_X1 U9505 ( .A1(n7652), .A2(n9967), .ZN(n7653) );
  AOI211_X1 U9506 ( .C1(n10011), .C2(n7655), .A(n7654), .B(n7653), .ZN(n7656)
         );
  OAI21_X1 U9507 ( .B1(n7657), .B2(n10024), .A(n7656), .ZN(P2_U3193) );
  AOI21_X1 U9508 ( .B1(n8685), .B2(n7659), .A(n7658), .ZN(n7674) );
  OAI21_X1 U9509 ( .B1(n7662), .B2(n7661), .A(n7660), .ZN(n7663) );
  NAND2_X1 U9510 ( .A1(n7663), .A2(n10001), .ZN(n7673) );
  AOI21_X1 U9511 ( .B1(n7666), .B2(n7665), .A(n7664), .ZN(n7669) );
  NAND2_X1 U9512 ( .A1(n10013), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7668) );
  AND2_X1 U9513 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8268) );
  INV_X1 U9514 ( .A(n8268), .ZN(n7667) );
  OAI211_X1 U9515 ( .C1(n7669), .C2(n10024), .A(n7668), .B(n7667), .ZN(n7670)
         );
  AOI21_X1 U9516 ( .B1(n10011), .B2(n7671), .A(n7670), .ZN(n7672) );
  OAI211_X1 U9517 ( .C1(n7674), .C2(n9967), .A(n7673), .B(n7672), .ZN(P2_U3195) );
  XNOR2_X1 U9518 ( .A(n7676), .B(n7675), .ZN(n9690) );
  AOI211_X1 U9519 ( .C1(n9687), .C2(n7677), .A(n9548), .B(n9570), .ZN(n9686)
         );
  INV_X1 U9520 ( .A(n9687), .ZN(n8889) );
  INV_X1 U9521 ( .A(n7678), .ZN(n8886) );
  AOI22_X1 U9522 ( .A1(n9934), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n8886), .B2(
        n9908), .ZN(n7679) );
  OAI21_X1 U9523 ( .B1(n8889), .B2(n9913), .A(n7679), .ZN(n7683) );
  OAI21_X1 U9524 ( .B1(n9109), .B2(n7680), .A(n9558), .ZN(n7681) );
  AOI222_X1 U9525 ( .A1(n9592), .A2(n7681), .B1(n9239), .B2(n4309), .C1(n9240), 
        .C2(n9563), .ZN(n9689) );
  NOR2_X1 U9526 ( .A1(n9689), .A2(n9910), .ZN(n7682) );
  AOI211_X1 U9527 ( .C1(n9686), .C2(n9905), .A(n7683), .B(n7682), .ZN(n7684)
         );
  OAI21_X1 U9528 ( .B1(n9690), .B2(n9556), .A(n7684), .ZN(P1_U3277) );
  INV_X1 U9529 ( .A(n7685), .ZN(n7689) );
  OAI222_X1 U9530 ( .A1(n7687), .A2(P1_U3086), .B1(n9769), .B2(n7689), .C1(
        n7686), .C2(n9766), .ZN(P1_U3331) );
  OAI222_X1 U9531 ( .A1(n8803), .A2(n7689), .B1(P2_U3151), .B2(n5775), .C1(
        n7688), .C2(n8800), .ZN(P2_U3271) );
  INV_X1 U9532 ( .A(n7690), .ZN(n7693) );
  OAI222_X1 U9533 ( .A1(n8803), .A2(n7693), .B1(P2_U3151), .B2(n6144), .C1(
        n7691), .C2(n8800), .ZN(P2_U3270) );
  OAI222_X1 U9534 ( .A1(n7694), .A2(P1_U3086), .B1(n9769), .B2(n7693), .C1(
        n7692), .C2(n9766), .ZN(P1_U3330) );
  INV_X1 U9535 ( .A(n6533), .ZN(n8790) );
  OAI222_X1 U9536 ( .A1(n9766), .A2(n7696), .B1(n9769), .B2(n8790), .C1(n7695), 
        .C2(P1_U3086), .ZN(P1_U3326) );
  INV_X1 U9537 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7706) );
  INV_X1 U9538 ( .A(SI_29_), .ZN(n7700) );
  INV_X1 U9539 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7714) );
  MUX2_X1 U9540 ( .A(n7706), .B(n7714), .S(n4701), .Z(n7702) );
  NAND2_X1 U9541 ( .A1(n7702), .A2(n8151), .ZN(n7724) );
  INV_X1 U9542 ( .A(n7702), .ZN(n7703) );
  NAND2_X1 U9543 ( .A1(n7703), .A2(SI_30_), .ZN(n7704) );
  NAND2_X1 U9544 ( .A1(n7724), .A2(n7704), .ZN(n7725) );
  INV_X1 U9545 ( .A(n7713), .ZN(n7708) );
  OAI222_X1 U9546 ( .A1(n9766), .A2(n7706), .B1(n9769), .B2(n7708), .C1(
        P1_U3086), .C2(n7705), .ZN(P1_U3325) );
  OAI222_X1 U9547 ( .A1(n8800), .A2(n7714), .B1(n8788), .B2(n7708), .C1(
        P2_U3151), .C2(n7707), .ZN(P2_U3265) );
  OAI222_X1 U9548 ( .A1(n9766), .A2(n7711), .B1(n9769), .B2(n7710), .C1(
        P1_U3086), .C2(n7709), .ZN(P1_U3333) );
  OR2_X1 U9549 ( .A1(n6083), .A2(n7714), .ZN(n7715) );
  INV_X1 U9550 ( .A(n8334), .ZN(n7735) );
  NAND2_X1 U9551 ( .A1(n8699), .A2(n7735), .ZN(n7960) );
  AND2_X1 U9552 ( .A1(n7960), .A2(n7901), .ZN(n7716) );
  NAND2_X1 U9553 ( .A1(n5839), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7721) );
  NAND2_X1 U9554 ( .A1(n6475), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7720) );
  NAND2_X1 U9555 ( .A1(n7718), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7719) );
  AND3_X1 U9556 ( .A1(n7721), .A2(n7720), .A3(n7719), .ZN(n7722) );
  NAND2_X1 U9557 ( .A1(n7723), .A2(n7722), .ZN(n8439) );
  INV_X1 U9558 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7728) );
  MUX2_X1 U9559 ( .A(n7728), .B(n6618), .S(n4701), .Z(n7729) );
  XNOR2_X1 U9560 ( .A(n7729), .B(SI_31_), .ZN(n7730) );
  NAND2_X1 U9561 ( .A1(n8975), .A2(n7732), .ZN(n7734) );
  OR2_X1 U9562 ( .A1(n6083), .A2(n6618), .ZN(n7733) );
  INV_X1 U9563 ( .A(n8439), .ZN(n7914) );
  NOR2_X1 U9564 ( .A1(n7973), .A2(n7971), .ZN(n7738) );
  MUX2_X1 U9565 ( .A(n7901), .B(n7903), .S(n7894), .Z(n7897) );
  AND2_X1 U9566 ( .A1(n8503), .A2(n7740), .ZN(n7744) );
  INV_X1 U9567 ( .A(n7741), .ZN(n7742) );
  NOR2_X1 U9568 ( .A1(n7925), .A2(n7742), .ZN(n7743) );
  MUX2_X1 U9569 ( .A(n7744), .B(n7743), .S(n7910), .Z(n7870) );
  AND2_X1 U9570 ( .A1(n7869), .A2(n7847), .ZN(n7840) );
  INV_X1 U9571 ( .A(n7840), .ZN(n7745) );
  AND2_X1 U9572 ( .A1(n7745), .A2(n7894), .ZN(n7862) );
  AND2_X1 U9573 ( .A1(n7847), .A2(n7854), .ZN(n7843) );
  INV_X1 U9574 ( .A(n7746), .ZN(n7747) );
  NOR2_X1 U9575 ( .A1(n8551), .A2(n7747), .ZN(n7748) );
  MUX2_X1 U9576 ( .A(n7843), .B(n7748), .S(n7894), .Z(n7861) );
  AOI21_X1 U9577 ( .B1(n7754), .B2(n7980), .A(n7749), .ZN(n7751) );
  MUX2_X1 U9578 ( .A(n7910), .B(n7751), .S(n7750), .Z(n7757) );
  OAI21_X1 U9579 ( .B1(n7753), .B2(n7752), .A(n6208), .ZN(n7756) );
  MUX2_X1 U9580 ( .A(n6208), .B(n7754), .S(n7894), .Z(n7755) );
  OAI211_X1 U9581 ( .C1(n7757), .C2(n7756), .A(n7755), .B(n7927), .ZN(n7765)
         );
  NAND2_X1 U9582 ( .A1(n7782), .A2(n7758), .ZN(n7762) );
  NAND2_X1 U9583 ( .A1(n7759), .A2(n7760), .ZN(n7761) );
  MUX2_X1 U9584 ( .A(n7762), .B(n7761), .S(n7910), .Z(n7763) );
  INV_X1 U9585 ( .A(n7763), .ZN(n7764) );
  NAND2_X1 U9586 ( .A1(n7765), .A2(n7764), .ZN(n7766) );
  NAND2_X1 U9587 ( .A1(n7766), .A2(n7928), .ZN(n7785) );
  INV_X1 U9588 ( .A(n7759), .ZN(n7769) );
  OAI211_X1 U9589 ( .C1(n7785), .C2(n7769), .A(n6211), .B(n7768), .ZN(n7771)
         );
  NAND2_X1 U9590 ( .A1(n7771), .A2(n7770), .ZN(n7772) );
  NAND3_X1 U9591 ( .A1(n7772), .A2(n7786), .A3(n7934), .ZN(n7774) );
  NAND2_X1 U9592 ( .A1(n7774), .A2(n7773), .ZN(n7781) );
  NAND2_X1 U9593 ( .A1(n7779), .A2(n7775), .ZN(n7777) );
  NAND2_X1 U9594 ( .A1(n7791), .A2(n7792), .ZN(n7776) );
  MUX2_X1 U9595 ( .A(n7777), .B(n7776), .S(n7894), .Z(n7778) );
  INV_X1 U9596 ( .A(n7778), .ZN(n7794) );
  NAND2_X1 U9597 ( .A1(n7799), .A2(n7779), .ZN(n7780) );
  AOI21_X1 U9598 ( .B1(n7781), .B2(n7794), .A(n7780), .ZN(n7797) );
  INV_X1 U9599 ( .A(n7782), .ZN(n7784) );
  OAI211_X1 U9600 ( .C1(n7785), .C2(n7784), .A(n10030), .B(n7783), .ZN(n7787)
         );
  NAND3_X1 U9601 ( .A1(n7787), .A2(n6211), .A3(n7786), .ZN(n7789) );
  NAND2_X1 U9602 ( .A1(n7798), .A2(n7792), .ZN(n7793) );
  AOI21_X1 U9603 ( .B1(n7795), .B2(n7794), .A(n7793), .ZN(n7796) );
  NAND2_X1 U9604 ( .A1(n7802), .A2(n7798), .ZN(n7801) );
  NAND2_X1 U9605 ( .A1(n7803), .A2(n7799), .ZN(n7800) );
  MUX2_X1 U9606 ( .A(n7801), .B(n7800), .S(n7910), .Z(n7805) );
  MUX2_X1 U9607 ( .A(n7803), .B(n7802), .S(n7910), .Z(n7804) );
  OAI211_X1 U9608 ( .C1(n7806), .C2(n7805), .A(n7942), .B(n7804), .ZN(n7810)
         );
  MUX2_X1 U9609 ( .A(n7808), .B(n7807), .S(n7910), .Z(n7809) );
  NAND2_X1 U9610 ( .A1(n7810), .A2(n7809), .ZN(n7816) );
  INV_X1 U9611 ( .A(n7811), .ZN(n7820) );
  OR2_X1 U9612 ( .A1(n7819), .A2(n7820), .ZN(n7945) );
  OAI21_X1 U9613 ( .B1(n7816), .B2(n7812), .A(n8610), .ZN(n7818) );
  INV_X1 U9614 ( .A(n7813), .ZN(n7815) );
  MUX2_X1 U9615 ( .A(n8337), .B(n8773), .S(n7894), .Z(n7814) );
  AOI21_X1 U9616 ( .B1(n7816), .B2(n7815), .A(n7814), .ZN(n7817) );
  MUX2_X1 U9617 ( .A(n7820), .B(n7819), .S(n7910), .Z(n7821) );
  INV_X1 U9618 ( .A(n7821), .ZN(n7822) );
  NAND2_X1 U9619 ( .A1(n7823), .A2(n7822), .ZN(n7825) );
  INV_X1 U9620 ( .A(n7824), .ZN(n7833) );
  NAND2_X1 U9621 ( .A1(n7825), .A2(n7988), .ZN(n7834) );
  NAND3_X1 U9622 ( .A1(n7834), .A2(n8597), .A3(n7826), .ZN(n7829) );
  XNOR2_X1 U9623 ( .A(n7827), .B(n7910), .ZN(n7828) );
  AOI21_X1 U9624 ( .B1(n7829), .B2(n7828), .A(n8586), .ZN(n7842) );
  AND2_X1 U9625 ( .A1(n7831), .A2(n7830), .ZN(n7950) );
  INV_X1 U9626 ( .A(n7950), .ZN(n7832) );
  AND2_X1 U9627 ( .A1(n7832), .A2(n7910), .ZN(n7841) );
  NAND2_X1 U9628 ( .A1(n7834), .A2(n7833), .ZN(n7836) );
  OAI21_X1 U9629 ( .B1(n7910), .B2(n8560), .A(n8751), .ZN(n7837) );
  OAI21_X1 U9630 ( .B1(n8560), .B2(n8751), .A(n7837), .ZN(n7838) );
  OAI211_X1 U9631 ( .C1(n7842), .C2(n7841), .A(n7840), .B(n7839), .ZN(n7860)
         );
  INV_X1 U9632 ( .A(n7843), .ZN(n7846) );
  OAI21_X1 U9633 ( .B1(n8590), .B2(n7947), .A(n8751), .ZN(n7844) );
  NAND2_X1 U9634 ( .A1(n7947), .A2(n8590), .ZN(n7848) );
  NAND4_X1 U9635 ( .A1(n7844), .A2(n7894), .A3(n8553), .A4(n7848), .ZN(n7845)
         );
  OAI21_X1 U9636 ( .B1(n7846), .B2(n7845), .A(n8738), .ZN(n7858) );
  INV_X1 U9637 ( .A(n7847), .ZN(n7856) );
  NAND3_X1 U9638 ( .A1(n7849), .A2(n7894), .A3(n7848), .ZN(n7852) );
  INV_X1 U9639 ( .A(n7947), .ZN(n7850) );
  NAND3_X1 U9640 ( .A1(n7850), .A2(n7894), .A3(n8560), .ZN(n7851) );
  NAND3_X1 U9641 ( .A1(n7852), .A2(n8528), .A3(n7851), .ZN(n7853) );
  OAI21_X1 U9642 ( .B1(n7854), .B2(n8553), .A(n7853), .ZN(n7855) );
  AOI21_X1 U9643 ( .B1(n7856), .B2(n8528), .A(n7855), .ZN(n7857) );
  NAND2_X1 U9644 ( .A1(n7858), .A2(n7857), .ZN(n7859) );
  OAI211_X1 U9645 ( .C1(n7862), .C2(n7861), .A(n7860), .B(n7859), .ZN(n7867)
         );
  NAND2_X1 U9646 ( .A1(n7864), .A2(n7863), .ZN(n7865) );
  NAND2_X1 U9647 ( .A1(n7865), .A2(n7910), .ZN(n7866) );
  NAND2_X1 U9648 ( .A1(n7867), .A2(n7866), .ZN(n7868) );
  AND2_X1 U9649 ( .A1(n6227), .A2(n7923), .ZN(n7872) );
  INV_X1 U9650 ( .A(n7922), .ZN(n7871) );
  AOI21_X1 U9651 ( .B1(n7875), .B2(n7872), .A(n7871), .ZN(n7877) );
  INV_X1 U9652 ( .A(n7923), .ZN(n7873) );
  AOI21_X1 U9653 ( .B1(n7875), .B2(n7874), .A(n7873), .ZN(n7876) );
  MUX2_X1 U9654 ( .A(n7879), .B(n7878), .S(n7910), .Z(n7880) );
  INV_X1 U9655 ( .A(n7882), .ZN(n7886) );
  INV_X1 U9656 ( .A(n8476), .ZN(n7883) );
  NAND2_X1 U9657 ( .A1(n7884), .A2(n7883), .ZN(n7893) );
  MUX2_X1 U9658 ( .A(n7886), .B(n7885), .S(n7910), .Z(n7887) );
  INV_X1 U9659 ( .A(n7887), .ZN(n7888) );
  AND2_X1 U9660 ( .A1(n7888), .A2(n8469), .ZN(n7892) );
  AND2_X1 U9661 ( .A1(n8478), .A2(n7894), .ZN(n7890) );
  NOR2_X1 U9662 ( .A1(n8478), .A2(n7894), .ZN(n7889) );
  MUX2_X1 U9663 ( .A(n7890), .B(n7889), .S(n8028), .Z(n7891) );
  MUX2_X1 U9664 ( .A(n8335), .B(n8458), .S(n7894), .Z(n7895) );
  OR2_X1 U9665 ( .A1(n7902), .A2(n7895), .ZN(n7896) );
  NAND2_X1 U9666 ( .A1(n7897), .A2(n7896), .ZN(n7904) );
  NAND3_X1 U9667 ( .A1(n7903), .A2(n7902), .A3(n8458), .ZN(n7898) );
  AND3_X1 U9668 ( .A1(n7960), .A2(n7901), .A3(n7898), .ZN(n7899) );
  OAI21_X1 U9669 ( .B1(n7904), .B2(n8335), .A(n7899), .ZN(n7900) );
  NAND2_X1 U9670 ( .A1(n7900), .A2(n7894), .ZN(n7907) );
  AND2_X1 U9671 ( .A1(n7909), .A2(n7960), .ZN(n7908) );
  NAND2_X1 U9672 ( .A1(n7908), .A2(n7910), .ZN(n7913) );
  NAND2_X1 U9673 ( .A1(n7913), .A2(n7912), .ZN(n7916) );
  NOR2_X1 U9674 ( .A1(n8695), .A2(n7914), .ZN(n7964) );
  INV_X1 U9675 ( .A(n7964), .ZN(n7915) );
  NOR2_X1 U9676 ( .A1(n7966), .A2(n7917), .ZN(n7918) );
  INV_X1 U9677 ( .A(n8503), .ZN(n7924) );
  INV_X1 U9678 ( .A(n8551), .ZN(n8549) );
  AND4_X1 U9679 ( .A1(n7929), .A2(n7928), .A3(n7927), .A4(n7926), .ZN(n7935)
         );
  NOR2_X1 U9680 ( .A1(n7930), .A2(n10048), .ZN(n7933) );
  NAND2_X1 U9681 ( .A1(n7932), .A2(n7931), .ZN(n10034) );
  NAND4_X1 U9682 ( .A1(n7935), .A2(n7934), .A3(n7933), .A4(n10034), .ZN(n7939)
         );
  NOR4_X1 U9683 ( .A1(n7939), .A2(n7938), .A3(n7937), .A4(n7936), .ZN(n7943)
         );
  INV_X1 U9684 ( .A(n7940), .ZN(n7941) );
  NAND4_X1 U9685 ( .A1(n7943), .A2(n7942), .A3(n7941), .A4(n8632), .ZN(n7944)
         );
  NOR2_X1 U9686 ( .A1(n7945), .A2(n7944), .ZN(n7946) );
  AND4_X1 U9687 ( .A1(n8597), .A2(n7947), .A3(n7988), .A4(n7946), .ZN(n7949)
         );
  NAND3_X1 U9688 ( .A1(n7950), .A2(n7949), .A3(n7948), .ZN(n7951) );
  NOR2_X1 U9689 ( .A1(n7952), .A2(n7951), .ZN(n7953) );
  NAND3_X1 U9690 ( .A1(n8539), .A2(n8549), .A3(n7953), .ZN(n7954) );
  NOR2_X1 U9691 ( .A1(n8523), .A2(n7954), .ZN(n7955) );
  NAND4_X1 U9692 ( .A1(n8488), .A2(n8505), .A3(n8511), .A4(n7955), .ZN(n7956)
         );
  NOR2_X1 U9693 ( .A1(n8476), .A2(n7956), .ZN(n7957) );
  NAND4_X1 U9694 ( .A1(n7958), .A2(n7957), .A3(n8469), .A4(n8019), .ZN(n7963)
         );
  INV_X1 U9695 ( .A(n7959), .ZN(n7962) );
  INV_X1 U9696 ( .A(n7960), .ZN(n7961) );
  NOR4_X1 U9697 ( .A1(n7964), .A2(n7963), .A3(n7962), .A4(n7961), .ZN(n7969)
         );
  INV_X1 U9698 ( .A(n7968), .ZN(n7965) );
  NAND4_X1 U9699 ( .A1(n7969), .A2(n7967), .A3(n4314), .A4(n7965), .ZN(n7970)
         );
  INV_X1 U9700 ( .A(n7966), .ZN(n7967) );
  INV_X1 U9701 ( .A(n7971), .ZN(n7972) );
  NAND3_X1 U9702 ( .A1(n7974), .A2(n7973), .A3(n7972), .ZN(n7975) );
  NOR3_X1 U9703 ( .A1(n7979), .A2(n7978), .A3(n7977), .ZN(n7982) );
  OAI21_X1 U9704 ( .B1(n7983), .B2(n7980), .A(P2_B_REG_SCAN_IN), .ZN(n7981) );
  OAI22_X1 U9705 ( .A1(n7984), .A2(n7983), .B1(n7982), .B2(n7981), .ZN(
        P2_U3296) );
  INV_X1 U9706 ( .A(n8791), .ZN(n7985) );
  OAI222_X1 U9707 ( .A1(n9766), .A2(n7986), .B1(n9769), .B2(n7985), .C1(n5716), 
        .C2(P1_U3086), .ZN(P1_U3327) );
  XOR2_X1 U9708 ( .A(n7988), .B(n7987), .Z(n8001) );
  INV_X1 U9709 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7991) );
  XNOR2_X1 U9710 ( .A(n7989), .B(n7988), .ZN(n7990) );
  AOI222_X1 U9711 ( .A1(n8627), .A2(n7990), .B1(n6044), .B2(n8622), .C1(n8623), 
        .C2(n8624), .ZN(n7996) );
  MUX2_X1 U9712 ( .A(n7991), .B(n7996), .S(n10110), .Z(n7993) );
  NAND2_X1 U9713 ( .A1(n7998), .A2(n8774), .ZN(n7992) );
  OAI211_X1 U9714 ( .C1(n8001), .C2(n8782), .A(n7993), .B(n7992), .ZN(P2_U3435) );
  MUX2_X1 U9715 ( .A(n8380), .B(n7996), .S(n10124), .Z(n7995) );
  NAND2_X1 U9716 ( .A1(n7998), .A2(n8686), .ZN(n7994) );
  OAI211_X1 U9717 ( .C1(n8694), .C2(n8001), .A(n7995), .B(n7994), .ZN(P2_U3474) );
  MUX2_X1 U9718 ( .A(n8369), .B(n7996), .S(n8616), .Z(n8000) );
  INV_X1 U9719 ( .A(n8325), .ZN(n7997) );
  AOI22_X1 U9720 ( .A1(n7998), .A2(n8605), .B1(n8604), .B2(n7997), .ZN(n7999)
         );
  OAI211_X1 U9721 ( .C1(n8001), .C2(n10047), .A(n8000), .B(n7999), .ZN(
        P2_U3218) );
  NAND2_X1 U9722 ( .A1(n8002), .A2(n4914), .ZN(n8006) );
  NAND2_X1 U9723 ( .A1(n8004), .A2(n8003), .ZN(n8005) );
  NAND3_X1 U9724 ( .A1(n8006), .A2(n8005), .A3(n8080), .ZN(n8010) );
  XNOR2_X1 U9725 ( .A(n8717), .B(n8018), .ZN(n8007) );
  NAND2_X1 U9726 ( .A1(n8007), .A2(n8500), .ZN(n8307) );
  INV_X1 U9727 ( .A(n8007), .ZN(n8008) );
  NAND2_X1 U9728 ( .A1(n8008), .A2(n8479), .ZN(n8009) );
  NAND2_X1 U9729 ( .A1(n8010), .A2(n8082), .ZN(n8083) );
  NAND2_X1 U9730 ( .A1(n8083), .A2(n8307), .ZN(n8011) );
  XNOR2_X1 U9731 ( .A(n8483), .B(n8018), .ZN(n8012) );
  XNOR2_X1 U9732 ( .A(n8012), .B(n8491), .ZN(n8308) );
  NAND2_X1 U9733 ( .A1(n8012), .A2(n8462), .ZN(n8013) );
  XNOR2_X1 U9734 ( .A(n8028), .B(n8018), .ZN(n8015) );
  XNOR2_X1 U9735 ( .A(n8015), .B(n8315), .ZN(n8029) );
  INV_X1 U9736 ( .A(n8029), .ZN(n8014) );
  INV_X1 U9737 ( .A(n8015), .ZN(n8016) );
  NAND2_X1 U9738 ( .A1(n8016), .A2(n8478), .ZN(n8017) );
  NAND2_X1 U9739 ( .A1(n8031), .A2(n8017), .ZN(n8021) );
  XNOR2_X1 U9740 ( .A(n8019), .B(n8018), .ZN(n8020) );
  XNOR2_X1 U9741 ( .A(n8021), .B(n8020), .ZN(n8027) );
  AOI22_X1 U9742 ( .A1(n8478), .A2(n8329), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8023) );
  NAND2_X1 U9743 ( .A1(n8452), .A2(n8317), .ZN(n8022) );
  OAI211_X1 U9744 ( .C1(n8024), .C2(n8324), .A(n8023), .B(n8022), .ZN(n8025)
         );
  AOI21_X1 U9745 ( .B1(n8458), .B2(n8303), .A(n8025), .ZN(n8026) );
  OAI21_X1 U9746 ( .B1(n8027), .B2(n8305), .A(n8026), .ZN(P2_U3160) );
  AOI21_X1 U9747 ( .B1(n8030), .B2(n8029), .A(n8305), .ZN(n8033) );
  NAND2_X1 U9748 ( .A1(n8033), .A2(n8031), .ZN(n8037) );
  NOR2_X1 U9749 ( .A1(n8462), .A2(n8288), .ZN(n8035) );
  INV_X1 U9750 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8213) );
  OAI22_X1 U9751 ( .A1(n8463), .A2(n8324), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8213), .ZN(n8034) );
  AOI211_X1 U9752 ( .C1(n8468), .C2(n8317), .A(n8035), .B(n8034), .ZN(n8036)
         );
  OAI211_X1 U9753 ( .C1(n8708), .C2(n8332), .A(n8037), .B(n8036), .ZN(P2_U3154) );
  XOR2_X1 U9754 ( .A(n4404), .B(n8038), .Z(n8043) );
  NAND2_X1 U9755 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8357) );
  OAI21_X1 U9756 ( .B1(n8324), .B2(n8613), .A(n8357), .ZN(n8039) );
  AOI21_X1 U9757 ( .B1(n8329), .B2(n8337), .A(n8039), .ZN(n8040) );
  OAI21_X1 U9758 ( .B1(n8614), .B2(n8326), .A(n8040), .ZN(n8041) );
  AOI21_X1 U9759 ( .B1(n8682), .B2(n8303), .A(n8041), .ZN(n8042) );
  OAI21_X1 U9760 ( .B1(n8043), .B2(n8305), .A(n8042), .ZN(P2_U3155) );
  AOI21_X1 U9761 ( .B1(n8336), .B2(n8045), .A(n8044), .ZN(n8050) );
  AOI22_X1 U9762 ( .A1(n8329), .A2(n8542), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8047) );
  NAND2_X1 U9763 ( .A1(n8317), .A2(n8517), .ZN(n8046) );
  OAI211_X1 U9764 ( .C1(n8088), .C2(n8324), .A(n8047), .B(n8046), .ZN(n8048)
         );
  AOI21_X1 U9765 ( .B1(n6296), .B2(n8303), .A(n8048), .ZN(n8049) );
  OAI21_X1 U9766 ( .B1(n8050), .B2(n8305), .A(n8049), .ZN(P2_U3156) );
  INV_X1 U9767 ( .A(n8566), .ZN(n8669) );
  OAI211_X1 U9768 ( .C1(n8052), .C2(n8051), .A(n8253), .B(n8320), .ZN(n8057)
         );
  OAI21_X1 U9769 ( .B1(n8324), .B2(n8063), .A(n8053), .ZN(n8055) );
  NOR2_X1 U9770 ( .A1(n8326), .A2(n8563), .ZN(n8054) );
  AOI211_X1 U9771 ( .C1(n8329), .C2(n8560), .A(n8055), .B(n8054), .ZN(n8056)
         );
  OAI211_X1 U9772 ( .C1(n8669), .C2(n8332), .A(n8057), .B(n8056), .ZN(P2_U3159) );
  INV_X1 U9773 ( .A(n8738), .ZN(n8068) );
  AND3_X1 U9774 ( .A1(n8250), .A2(n8059), .A3(n8058), .ZN(n8060) );
  OAI21_X1 U9775 ( .B1(n4361), .B2(n8060), .A(n8320), .ZN(n8067) );
  OAI22_X1 U9776 ( .A1(n8324), .A2(n8062), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8061), .ZN(n8065) );
  NOR2_X1 U9777 ( .A1(n8288), .A2(n8063), .ZN(n8064) );
  AOI211_X1 U9778 ( .C1(n8545), .C2(n8317), .A(n8065), .B(n8064), .ZN(n8066)
         );
  OAI211_X1 U9779 ( .C1(n8068), .C2(n8332), .A(n8067), .B(n8066), .ZN(P2_U3163) );
  INV_X1 U9780 ( .A(n8069), .ZN(n8070) );
  NAND2_X1 U9781 ( .A1(n8317), .A2(n8070), .ZN(n8073) );
  AOI21_X1 U9782 ( .B1(n8329), .B2(n8338), .A(n8071), .ZN(n8072) );
  OAI211_X1 U9783 ( .C1(n8612), .C2(n8324), .A(n8073), .B(n8072), .ZN(n8078)
         );
  XNOR2_X1 U9784 ( .A(n8075), .B(n8074), .ZN(n8076) );
  NOR2_X1 U9785 ( .A1(n8076), .A2(n8305), .ZN(n8077) );
  AOI211_X1 U9786 ( .C1(n8691), .C2(n8303), .A(n8078), .B(n8077), .ZN(n8079)
         );
  INV_X1 U9787 ( .A(n8079), .ZN(P2_U3164) );
  INV_X1 U9788 ( .A(n8080), .ZN(n8081) );
  NOR2_X1 U9789 ( .A1(n8082), .A2(n8081), .ZN(n8084) );
  INV_X1 U9790 ( .A(n8083), .ZN(n8310) );
  AOI21_X1 U9791 ( .B1(n8085), .B2(n8084), .A(n8310), .ZN(n8091) );
  AOI22_X1 U9792 ( .A1(n8491), .A2(n8283), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8087) );
  NAND2_X1 U9793 ( .A1(n8317), .A2(n8495), .ZN(n8086) );
  OAI211_X1 U9794 ( .C1(n8088), .C2(n8288), .A(n8087), .B(n8086), .ZN(n8089)
         );
  AOI21_X1 U9795 ( .B1(n8717), .B2(n8303), .A(n8089), .ZN(n8090) );
  OAI21_X1 U9796 ( .B1(n8091), .B2(n8305), .A(n8090), .ZN(P2_U3165) );
  OAI211_X1 U9797 ( .C1(n8094), .C2(n8093), .A(n8092), .B(n8320), .ZN(n8098)
         );
  NAND2_X1 U9798 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8394) );
  OAI21_X1 U9799 ( .B1(n8324), .B2(n8101), .A(n8394), .ZN(n8096) );
  NOR2_X1 U9800 ( .A1(n8326), .A2(n8602), .ZN(n8095) );
  AOI211_X1 U9801 ( .C1(n8329), .C2(n6029), .A(n8096), .B(n8095), .ZN(n8097)
         );
  OAI211_X1 U9802 ( .C1(n8099), .C2(n8332), .A(n8098), .B(n8097), .ZN(P2_U3166) );
  XNOR2_X1 U9803 ( .A(n8102), .B(n8101), .ZN(n8103) );
  XNOR2_X1 U9804 ( .A(n8100), .B(n8103), .ZN(n8108) );
  NOR2_X1 U9805 ( .A1(n8326), .A2(n8591), .ZN(n8106) );
  NAND2_X1 U9806 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8409) );
  NAND2_X1 U9807 ( .A1(n8283), .A2(n8560), .ZN(n8104) );
  OAI211_X1 U9808 ( .C1(n8288), .C2(n8589), .A(n8409), .B(n8104), .ZN(n8105)
         );
  AOI211_X1 U9809 ( .C1(n8674), .C2(n8303), .A(n8106), .B(n8105), .ZN(n8107)
         );
  OAI21_X1 U9810 ( .B1(n8108), .B2(n8305), .A(n8107), .ZN(n8249) );
  NOR2_X1 U9811 ( .A1(keyinput24), .A2(keyinput10), .ZN(n8115) );
  NAND2_X1 U9812 ( .A1(keyinput5), .A2(keyinput22), .ZN(n8113) );
  NOR3_X1 U9813 ( .A1(keyinput15), .A2(keyinput7), .A3(keyinput48), .ZN(n8111)
         );
  INV_X1 U9814 ( .A(keyinput6), .ZN(n8109) );
  NOR3_X1 U9815 ( .A1(keyinput50), .A2(keyinput39), .A3(n8109), .ZN(n8110) );
  NAND4_X1 U9816 ( .A1(keyinput14), .A2(n8111), .A3(keyinput33), .A4(n8110), 
        .ZN(n8112) );
  NOR4_X1 U9817 ( .A1(keyinput44), .A2(keyinput3), .A3(n8113), .A4(n8112), 
        .ZN(n8114) );
  NAND4_X1 U9818 ( .A1(keyinput38), .A2(keyinput17), .A3(n8115), .A4(n8114), 
        .ZN(n8247) );
  NOR3_X1 U9819 ( .A1(keyinput52), .A2(keyinput28), .A3(keyinput20), .ZN(n8117) );
  NOR3_X1 U9820 ( .A1(keyinput47), .A2(keyinput1), .A3(keyinput12), .ZN(n8116)
         );
  NAND4_X1 U9821 ( .A1(keyinput26), .A2(n8117), .A3(keyinput56), .A4(n8116), 
        .ZN(n8119) );
  NAND2_X1 U9822 ( .A1(keyinput36), .A2(keyinput13), .ZN(n8118) );
  OR4_X1 U9823 ( .A1(n8119), .A2(keyinput23), .A3(n8118), .A4(keyinput32), 
        .ZN(n8135) );
  NOR2_X1 U9824 ( .A1(keyinput42), .A2(keyinput54), .ZN(n8122) );
  INV_X1 U9825 ( .A(keyinput31), .ZN(n8120) );
  NOR4_X1 U9826 ( .A1(keyinput62), .A2(keyinput11), .A3(keyinput19), .A4(n8120), .ZN(n8121) );
  NAND4_X1 U9827 ( .A1(keyinput51), .A2(keyinput63), .A3(n8122), .A4(n8121), 
        .ZN(n8134) );
  NOR2_X1 U9828 ( .A1(keyinput8), .A2(keyinput30), .ZN(n8126) );
  NAND3_X1 U9829 ( .A1(keyinput46), .A2(keyinput40), .A3(keyinput61), .ZN(
        n8124) );
  NAND3_X1 U9830 ( .A1(keyinput60), .A2(keyinput55), .A3(keyinput43), .ZN(
        n8123) );
  NOR4_X1 U9831 ( .A1(keyinput49), .A2(keyinput37), .A3(n8124), .A4(n8123), 
        .ZN(n8125) );
  NAND4_X1 U9832 ( .A1(keyinput25), .A2(keyinput0), .A3(n8126), .A4(n8125), 
        .ZN(n8133) );
  NOR3_X1 U9833 ( .A1(keyinput59), .A2(keyinput4), .A3(keyinput57), .ZN(n8131)
         );
  NOR4_X1 U9834 ( .A1(keyinput34), .A2(keyinput45), .A3(keyinput53), .A4(
        keyinput58), .ZN(n8130) );
  NAND2_X1 U9835 ( .A1(keyinput18), .A2(keyinput41), .ZN(n8128) );
  NAND4_X1 U9836 ( .A1(keyinput29), .A2(keyinput27), .A3(keyinput35), .A4(
        keyinput9), .ZN(n8127) );
  NOR4_X1 U9837 ( .A1(keyinput16), .A2(keyinput21), .A3(n8128), .A4(n8127), 
        .ZN(n8129) );
  NAND4_X1 U9838 ( .A1(keyinput2), .A2(n8131), .A3(n8130), .A4(n8129), .ZN(
        n8132) );
  OR4_X1 U9839 ( .A1(n8135), .A2(n8134), .A3(n8133), .A4(n8132), .ZN(n8246) );
  INV_X1 U9840 ( .A(keyinput23), .ZN(n8137) );
  AOI22_X1 U9841 ( .A1(n8138), .A2(keyinput32), .B1(P2_WR_REG_SCAN_IN), .B2(
        n8137), .ZN(n8136) );
  OAI221_X1 U9842 ( .B1(n8138), .B2(keyinput32), .C1(n8137), .C2(
        P2_WR_REG_SCAN_IN), .A(n8136), .ZN(n8149) );
  INV_X1 U9843 ( .A(keyinput17), .ZN(n8140) );
  AOI22_X1 U9844 ( .A1(n8141), .A2(keyinput10), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n8140), .ZN(n8139) );
  OAI221_X1 U9845 ( .B1(n8141), .B2(keyinput10), .C1(n8140), .C2(
        P1_ADDR_REG_15__SCAN_IN), .A(n8139), .ZN(n8148) );
  INV_X1 U9846 ( .A(keyinput45), .ZN(n8143) );
  AOI22_X1 U9847 ( .A1(n8868), .A2(keyinput34), .B1(P1_ADDR_REG_7__SCAN_IN), 
        .B2(n8143), .ZN(n8142) );
  OAI221_X1 U9848 ( .B1(n8868), .B2(keyinput34), .C1(n8143), .C2(
        P1_ADDR_REG_7__SCAN_IN), .A(n8142), .ZN(n8147) );
  INV_X1 U9849 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8145) );
  AOI22_X1 U9850 ( .A1(n6734), .A2(keyinput19), .B1(keyinput31), .B2(n8145), 
        .ZN(n8144) );
  OAI221_X1 U9851 ( .B1(n6734), .B2(keyinput19), .C1(n8145), .C2(keyinput31), 
        .A(n8144), .ZN(n8146) );
  NOR4_X1 U9852 ( .A1(n8149), .A2(n8148), .A3(n8147), .A4(n8146), .ZN(n8170)
         );
  INV_X1 U9853 ( .A(SI_30_), .ZN(n8151) );
  AOI22_X1 U9854 ( .A1(n8152), .A2(keyinput46), .B1(keyinput49), .B2(n8151), 
        .ZN(n8150) );
  OAI221_X1 U9855 ( .B1(n8152), .B2(keyinput46), .C1(n8151), .C2(keyinput49), 
        .A(n8150), .ZN(n8157) );
  INV_X1 U9856 ( .A(keyinput18), .ZN(n8155) );
  INV_X1 U9857 ( .A(keyinput41), .ZN(n8154) );
  AOI22_X1 U9858 ( .A1(n8155), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P2_ADDR_REG_4__SCAN_IN), .B2(n8154), .ZN(n8153) );
  OAI221_X1 U9859 ( .B1(n8155), .B2(P1_ADDR_REG_1__SCAN_IN), .C1(n8154), .C2(
        P2_ADDR_REG_4__SCAN_IN), .A(n8153), .ZN(n8156) );
  NOR2_X1 U9860 ( .A1(n8157), .A2(n8156), .ZN(n8169) );
  INV_X1 U9861 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8159) );
  INV_X1 U9862 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10094) );
  AOI22_X1 U9863 ( .A1(n8159), .A2(keyinput39), .B1(keyinput6), .B2(n10094), 
        .ZN(n8158) );
  OAI221_X1 U9864 ( .B1(n8159), .B2(keyinput39), .C1(n10094), .C2(keyinput6), 
        .A(n8158), .ZN(n8167) );
  INV_X1 U9865 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8161) );
  AOI22_X1 U9866 ( .A1(n8162), .A2(keyinput24), .B1(keyinput38), .B2(n8161), 
        .ZN(n8160) );
  OAI221_X1 U9867 ( .B1(n8162), .B2(keyinput24), .C1(n8161), .C2(keyinput38), 
        .A(n8160), .ZN(n8166) );
  AOI22_X1 U9868 ( .A1(n9683), .A2(keyinput40), .B1(n8164), .B2(keyinput61), 
        .ZN(n8163) );
  OAI221_X1 U9869 ( .B1(n9683), .B2(keyinput40), .C1(n8164), .C2(keyinput61), 
        .A(n8163), .ZN(n8165) );
  NOR3_X1 U9870 ( .A1(n8167), .A2(n8166), .A3(n8165), .ZN(n8168) );
  NAND3_X1 U9871 ( .A1(n8170), .A2(n8169), .A3(n8168), .ZN(n8231) );
  INV_X1 U9872 ( .A(SI_15_), .ZN(n8172) );
  AOI22_X1 U9873 ( .A1(n8173), .A2(keyinput26), .B1(n8172), .B2(keyinput20), 
        .ZN(n8171) );
  OAI221_X1 U9874 ( .B1(n8173), .B2(keyinput26), .C1(n8172), .C2(keyinput20), 
        .A(n8171), .ZN(n8179) );
  XNOR2_X1 U9875 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput56), .ZN(n8177) );
  XNOR2_X1 U9876 ( .A(P2_REG2_REG_0__SCAN_IN), .B(keyinput1), .ZN(n8176) );
  XNOR2_X1 U9877 ( .A(keyinput53), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n8175) );
  XNOR2_X1 U9878 ( .A(keyinput11), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n8174) );
  NAND4_X1 U9879 ( .A1(n8177), .A2(n8176), .A3(n8175), .A4(n8174), .ZN(n8178)
         );
  NOR2_X1 U9880 ( .A1(n8179), .A2(n8178), .ZN(n8210) );
  INV_X1 U9881 ( .A(keyinput33), .ZN(n8180) );
  XNOR2_X1 U9882 ( .A(n8180), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n8186) );
  XNOR2_X1 U9883 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput58), .ZN(n8184) );
  XNOR2_X1 U9884 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput9), .ZN(n8183) );
  XNOR2_X1 U9885 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput50), .ZN(n8182) );
  XNOR2_X1 U9886 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput22), .ZN(n8181) );
  NAND4_X1 U9887 ( .A1(n8184), .A2(n8183), .A3(n8182), .A4(n8181), .ZN(n8185)
         );
  NOR2_X1 U9888 ( .A1(n8186), .A2(n8185), .ZN(n8209) );
  XNOR2_X1 U9889 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput5), .ZN(n8190) );
  XNOR2_X1 U9890 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput7), .ZN(n8189) );
  XNOR2_X1 U9891 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput21), .ZN(n8188) );
  XNOR2_X1 U9892 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput35), .ZN(n8187) );
  NAND4_X1 U9893 ( .A1(n8190), .A2(n8189), .A3(n8188), .A4(n8187), .ZN(n8196)
         );
  XNOR2_X1 U9894 ( .A(P2_REG1_REG_29__SCAN_IN), .B(keyinput44), .ZN(n8194) );
  XNOR2_X1 U9895 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput3), .ZN(n8193) );
  XNOR2_X1 U9896 ( .A(P2_REG1_REG_31__SCAN_IN), .B(keyinput15), .ZN(n8192) );
  XNOR2_X1 U9897 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput12), .ZN(n8191) );
  NAND4_X1 U9898 ( .A1(n8194), .A2(n8193), .A3(n8192), .A4(n8191), .ZN(n8195)
         );
  NOR2_X1 U9899 ( .A1(n8196), .A2(n8195), .ZN(n8208) );
  XNOR2_X1 U9900 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput52), .ZN(n8200) );
  XNOR2_X1 U9901 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput42), .ZN(n8199) );
  XNOR2_X1 U9902 ( .A(P1_REG0_REG_16__SCAN_IN), .B(keyinput51), .ZN(n8198) );
  XNOR2_X1 U9903 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput13), .ZN(n8197) );
  NAND4_X1 U9904 ( .A1(n8200), .A2(n8199), .A3(n8198), .A4(n8197), .ZN(n8206)
         );
  XNOR2_X1 U9905 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput62), .ZN(n8204) );
  XNOR2_X1 U9906 ( .A(P2_REG1_REG_18__SCAN_IN), .B(keyinput36), .ZN(n8203) );
  XNOR2_X1 U9907 ( .A(P2_IR_REG_2__SCAN_IN), .B(keyinput28), .ZN(n8202) );
  XNOR2_X1 U9908 ( .A(P2_REG1_REG_23__SCAN_IN), .B(keyinput47), .ZN(n8201) );
  NAND4_X1 U9909 ( .A1(n8204), .A2(n8203), .A3(n8202), .A4(n8201), .ZN(n8205)
         );
  NOR2_X1 U9910 ( .A1(n8206), .A2(n8205), .ZN(n8207) );
  NAND4_X1 U9911 ( .A1(n8210), .A2(n8209), .A3(n8208), .A4(n8207), .ZN(n8230)
         );
  AOI22_X1 U9912 ( .A1(n5223), .A2(keyinput4), .B1(keyinput57), .B2(n6666), 
        .ZN(n8211) );
  OAI221_X1 U9913 ( .B1(n5223), .B2(keyinput4), .C1(n6666), .C2(keyinput57), 
        .A(n8211), .ZN(n8217) );
  AOI22_X1 U9914 ( .A1(n8213), .A2(keyinput2), .B1(keyinput59), .B2(n8675), 
        .ZN(n8212) );
  OAI221_X1 U9915 ( .B1(n8213), .B2(keyinput2), .C1(n8675), .C2(keyinput59), 
        .A(n8212), .ZN(n8216) );
  INV_X1 U9916 ( .A(keyinput16), .ZN(n8214) );
  XNOR2_X1 U9917 ( .A(n8214), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(n8215) );
  OR3_X1 U9918 ( .A1(n8217), .A2(n8216), .A3(n8215), .ZN(n8228) );
  AOI22_X1 U9919 ( .A1(n8219), .A2(keyinput54), .B1(keyinput63), .B2(n6405), 
        .ZN(n8218) );
  OAI221_X1 U9920 ( .B1(n8219), .B2(keyinput54), .C1(n6405), .C2(keyinput63), 
        .A(n8218), .ZN(n8227) );
  AOI22_X1 U9921 ( .A1(n8222), .A2(keyinput48), .B1(keyinput14), .B2(n8221), 
        .ZN(n8220) );
  OAI221_X1 U9922 ( .B1(n8222), .B2(keyinput48), .C1(n8221), .C2(keyinput14), 
        .A(n8220), .ZN(n8226) );
  AOI22_X1 U9923 ( .A1(n8224), .A2(keyinput29), .B1(keyinput27), .B2(n8685), 
        .ZN(n8223) );
  OAI221_X1 U9924 ( .B1(n8224), .B2(keyinput29), .C1(n8685), .C2(keyinput27), 
        .A(n8223), .ZN(n8225) );
  OR4_X1 U9925 ( .A1(n8228), .A2(n8227), .A3(n8226), .A4(n8225), .ZN(n8229) );
  NOR3_X1 U9926 ( .A1(n8231), .A2(n8230), .A3(n8229), .ZN(n8245) );
  INV_X1 U9927 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9745) );
  AOI22_X1 U9928 ( .A1(n9745), .A2(keyinput37), .B1(keyinput43), .B2(n8233), 
        .ZN(n8232) );
  OAI221_X1 U9929 ( .B1(n9745), .B2(keyinput37), .C1(n8233), .C2(keyinput43), 
        .A(n8232), .ZN(n8243) );
  INV_X1 U9930 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9935) );
  AOI22_X1 U9931 ( .A1(n9935), .A2(keyinput60), .B1(keyinput55), .B2(n5926), 
        .ZN(n8234) );
  OAI221_X1 U9932 ( .B1(n9935), .B2(keyinput60), .C1(n5926), .C2(keyinput55), 
        .A(n8234), .ZN(n8242) );
  AOI22_X1 U9933 ( .A1(n8236), .A2(keyinput30), .B1(keyinput0), .B2(n8481), 
        .ZN(n8235) );
  OAI221_X1 U9934 ( .B1(n8236), .B2(keyinput30), .C1(n8481), .C2(keyinput0), 
        .A(n8235), .ZN(n8241) );
  AOI22_X1 U9935 ( .A1(n8239), .A2(keyinput25), .B1(keyinput8), .B2(n8238), 
        .ZN(n8237) );
  OAI221_X1 U9936 ( .B1(n8239), .B2(keyinput25), .C1(n8238), .C2(keyinput8), 
        .A(n8237), .ZN(n8240) );
  NOR4_X1 U9937 ( .A1(n8243), .A2(n8242), .A3(n8241), .A4(n8240), .ZN(n8244)
         );
  OAI211_X1 U9938 ( .C1(n8247), .C2(n8246), .A(n8245), .B(n8244), .ZN(n8248)
         );
  XNOR2_X1 U9939 ( .A(n8249), .B(n8248), .ZN(P2_U3168) );
  INV_X1 U9940 ( .A(n8250), .ZN(n8255) );
  AOI21_X1 U9941 ( .B1(n8253), .B2(n8252), .A(n8251), .ZN(n8254) );
  OAI21_X1 U9942 ( .B1(n8255), .B2(n8254), .A(n8320), .ZN(n8259) );
  AOI22_X1 U9943 ( .A1(n8283), .A2(n8553), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8256) );
  OAI21_X1 U9944 ( .B1(n8300), .B2(n8288), .A(n8256), .ZN(n8257) );
  AOI21_X1 U9945 ( .B1(n8556), .B2(n8317), .A(n8257), .ZN(n8258) );
  OAI211_X1 U9946 ( .C1(n8260), .C2(n8332), .A(n8259), .B(n8258), .ZN(P2_U3173) );
  INV_X1 U9947 ( .A(n8261), .ZN(n8262) );
  NOR2_X1 U9948 ( .A1(n8263), .A2(n8262), .ZN(n8264) );
  XNOR2_X1 U9949 ( .A(n8265), .B(n8264), .ZN(n8272) );
  NOR2_X1 U9950 ( .A1(n8324), .A2(n8266), .ZN(n8267) );
  AOI211_X1 U9951 ( .C1(n8329), .C2(n8625), .A(n8268), .B(n8267), .ZN(n8269)
         );
  OAI21_X1 U9952 ( .B1(n8620), .B2(n8326), .A(n8269), .ZN(n8270) );
  AOI21_X1 U9953 ( .B1(n8773), .B2(n8303), .A(n8270), .ZN(n8271) );
  OAI21_X1 U9954 ( .B1(n8272), .B2(n8305), .A(n8271), .ZN(P2_U3174) );
  INV_X1 U9955 ( .A(n8533), .ZN(n8732) );
  INV_X1 U9956 ( .A(n8273), .ZN(n8277) );
  NOR3_X1 U9957 ( .A1(n4361), .A2(n8275), .A3(n8274), .ZN(n8276) );
  OAI21_X1 U9958 ( .B1(n8277), .B2(n8276), .A(n8320), .ZN(n8281) );
  AOI22_X1 U9959 ( .A1(n8329), .A2(n8553), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8278) );
  OAI21_X1 U9960 ( .B1(n8529), .B2(n8324), .A(n8278), .ZN(n8279) );
  AOI21_X1 U9961 ( .B1(n8532), .B2(n8317), .A(n8279), .ZN(n8280) );
  OAI211_X1 U9962 ( .C1(n8732), .C2(n8332), .A(n8281), .B(n8280), .ZN(P2_U3175) );
  AOI21_X1 U9963 ( .B1(n8283), .B2(n8625), .A(n8282), .ZN(n8286) );
  NAND2_X1 U9964 ( .A1(n8317), .A2(n8284), .ZN(n8285) );
  OAI211_X1 U9965 ( .C1(n8288), .C2(n8287), .A(n8286), .B(n8285), .ZN(n8293)
         );
  AOI211_X1 U9966 ( .C1(n8291), .C2(n8289), .A(n8305), .B(n8290), .ZN(n8292)
         );
  AOI211_X1 U9967 ( .C1(n8294), .C2(n8303), .A(n8293), .B(n8292), .ZN(n8295)
         );
  INV_X1 U9968 ( .A(n8295), .ZN(P2_U3176) );
  AOI21_X1 U9969 ( .B1(n8298), .B2(n8296), .A(n8297), .ZN(n8306) );
  NOR2_X1 U9970 ( .A1(n8326), .A2(n8580), .ZN(n8302) );
  NAND2_X1 U9971 ( .A1(n8329), .A2(n8599), .ZN(n8299) );
  NAND2_X1 U9972 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8433) );
  OAI211_X1 U9973 ( .C1(n8300), .C2(n8324), .A(n8299), .B(n8433), .ZN(n8301)
         );
  AOI211_X1 U9974 ( .C1(n8751), .C2(n8303), .A(n8302), .B(n8301), .ZN(n8304)
         );
  OAI21_X1 U9975 ( .B1(n8306), .B2(n8305), .A(n8304), .ZN(P2_U3178) );
  INV_X1 U9976 ( .A(n8307), .ZN(n8309) );
  NOR3_X1 U9977 ( .A1(n8310), .A2(n8309), .A3(n8308), .ZN(n8313) );
  INV_X1 U9978 ( .A(n8311), .ZN(n8312) );
  OAI21_X1 U9979 ( .B1(n8313), .B2(n8312), .A(n8320), .ZN(n8319) );
  AOI22_X1 U9980 ( .A1(n8479), .A2(n8329), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8314) );
  OAI21_X1 U9981 ( .B1(n8315), .B2(n8324), .A(n8314), .ZN(n8316) );
  AOI21_X1 U9982 ( .B1(n8482), .B2(n8317), .A(n8316), .ZN(n8318) );
  OAI211_X1 U9983 ( .C1(n8714), .C2(n8332), .A(n8319), .B(n8318), .ZN(P2_U3180) );
  OAI211_X1 U9984 ( .C1(n8323), .C2(n8322), .A(n8321), .B(n8320), .ZN(n8331)
         );
  NAND2_X1 U9985 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8375) );
  OAI21_X1 U9986 ( .B1(n8324), .B2(n8589), .A(n8375), .ZN(n8328) );
  NOR2_X1 U9987 ( .A1(n8326), .A2(n8325), .ZN(n8327) );
  AOI211_X1 U9988 ( .C1(n8329), .C2(n8623), .A(n8328), .B(n8327), .ZN(n8330)
         );
  OAI211_X1 U9989 ( .C1(n8333), .C2(n8332), .A(n8331), .B(n8330), .ZN(P2_U3181) );
  MUX2_X1 U9990 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8439), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9991 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8334), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9992 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8335), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9993 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8478), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9994 ( .A(n8491), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8347), .Z(
        P2_U3517) );
  MUX2_X1 U9995 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8479), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9996 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8514), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9997 ( .A(n8336), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8347), .Z(
        P2_U3514) );
  MUX2_X1 U9998 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8542), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9999 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8553), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10000 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8561), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10001 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8577), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10002 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8560), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10003 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8599), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10004 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n6044), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10005 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n6029), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10006 ( .A(n8623), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8347), .Z(
        P2_U3505) );
  MUX2_X1 U10007 ( .A(n8337), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8347), .Z(
        P2_U3504) );
  MUX2_X1 U10008 ( .A(n8625), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8347), .Z(
        P2_U3503) );
  MUX2_X1 U10009 ( .A(n8338), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8347), .Z(
        P2_U3502) );
  MUX2_X1 U10010 ( .A(n8339), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8347), .Z(
        P2_U3501) );
  MUX2_X1 U10011 ( .A(n8340), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8347), .Z(
        P2_U3500) );
  MUX2_X1 U10012 ( .A(n8341), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8347), .Z(
        P2_U3499) );
  MUX2_X1 U10013 ( .A(n8342), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8347), .Z(
        P2_U3498) );
  MUX2_X1 U10014 ( .A(n8343), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8347), .Z(
        P2_U3497) );
  MUX2_X1 U10015 ( .A(n8344), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8347), .Z(
        P2_U3496) );
  MUX2_X1 U10016 ( .A(n8345), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8347), .Z(
        P2_U3495) );
  MUX2_X1 U10017 ( .A(n6209), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8347), .Z(
        P2_U3494) );
  MUX2_X1 U10018 ( .A(n8346), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8347), .Z(
        P2_U3493) );
  MUX2_X1 U10019 ( .A(n8348), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8347), .Z(
        P2_U3492) );
  MUX2_X1 U10020 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8349), .S(P2_U3893), .Z(
        P2_U3491) );
  AOI21_X1 U10021 ( .B1(n8352), .B2(n8351), .A(n8350), .ZN(n8367) );
  OAI21_X1 U10022 ( .B1(n8355), .B2(n8354), .A(n8353), .ZN(n8365) );
  INV_X1 U10023 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8359) );
  NAND2_X1 U10024 ( .A1(n10011), .A2(n8356), .ZN(n8358) );
  OAI211_X1 U10025 ( .C1(n9982), .C2(n8359), .A(n8358), .B(n8357), .ZN(n8364)
         );
  AOI21_X1 U10026 ( .B1(n4364), .B2(n8361), .A(n8360), .ZN(n8362) );
  NOR2_X1 U10027 ( .A1(n8362), .A2(n9967), .ZN(n8363) );
  AOI211_X1 U10028 ( .C1(n10001), .C2(n8365), .A(n8364), .B(n8363), .ZN(n8366)
         );
  OAI21_X1 U10029 ( .B1(n8367), .B2(n10024), .A(n8366), .ZN(P2_U3196) );
  AOI21_X1 U10030 ( .B1(n8370), .B2(n8369), .A(n8368), .ZN(n8386) );
  OAI21_X1 U10031 ( .B1(n8373), .B2(n8372), .A(n8371), .ZN(n8384) );
  NAND2_X1 U10032 ( .A1(n10011), .A2(n8374), .ZN(n8376) );
  OAI211_X1 U10033 ( .C1(n9982), .C2(n8377), .A(n8376), .B(n8375), .ZN(n8383)
         );
  AOI21_X1 U10034 ( .B1(n8380), .B2(n8379), .A(n8378), .ZN(n8381) );
  NOR2_X1 U10035 ( .A1(n8381), .A2(n9967), .ZN(n8382) );
  AOI211_X1 U10036 ( .C1(n10001), .C2(n8384), .A(n8383), .B(n8382), .ZN(n8385)
         );
  OAI21_X1 U10037 ( .B1(n8386), .B2(n10024), .A(n8385), .ZN(P2_U3197) );
  AOI21_X1 U10038 ( .B1(n8389), .B2(n8388), .A(n8387), .ZN(n8405) );
  OAI21_X1 U10039 ( .B1(n8392), .B2(n8391), .A(n8390), .ZN(n8403) );
  INV_X1 U10040 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8396) );
  NAND2_X1 U10041 ( .A1(n10011), .A2(n8393), .ZN(n8395) );
  OAI211_X1 U10042 ( .C1(n9982), .C2(n8396), .A(n8395), .B(n8394), .ZN(n8402)
         );
  AOI21_X1 U10043 ( .B1(n8399), .B2(n8398), .A(n8397), .ZN(n8400) );
  NOR2_X1 U10044 ( .A1(n8400), .A2(n9967), .ZN(n8401) );
  AOI211_X1 U10045 ( .C1(n10001), .C2(n8403), .A(n8402), .B(n8401), .ZN(n8404)
         );
  OAI21_X1 U10046 ( .B1(n8405), .B2(n10024), .A(n8404), .ZN(P2_U3198) );
  AOI21_X1 U10047 ( .B1(n8675), .B2(n8407), .A(n8406), .ZN(n8419) );
  NOR2_X1 U10048 ( .A1(n9982), .A2(n8410), .ZN(n8411) );
  OAI21_X1 U10049 ( .B1(n8415), .B2(n8414), .A(n8413), .ZN(n8416) );
  NAND2_X1 U10050 ( .A1(n8416), .A2(n10001), .ZN(n8417) );
  OAI211_X1 U10051 ( .C1(n8419), .C2(n9967), .A(n8418), .B(n8417), .ZN(
        P2_U3199) );
  AOI21_X1 U10052 ( .B1(n4397), .B2(n8421), .A(n8420), .ZN(n8437) );
  NOR2_X1 U10053 ( .A1(n8424), .A2(n9967), .ZN(n8436) );
  INV_X1 U10054 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10133) );
  INV_X1 U10055 ( .A(n8429), .ZN(n8428) );
  NAND2_X1 U10056 ( .A1(n8428), .A2(n10001), .ZN(n8432) );
  OAI211_X1 U10057 ( .C1(n10133), .C2(n9982), .A(n8434), .B(n8433), .ZN(n8435)
         );
  NAND2_X1 U10058 ( .A1(n8445), .A2(n8604), .ZN(n8440) );
  NAND2_X1 U10059 ( .A1(n8439), .A2(n8438), .ZN(n8696) );
  AOI21_X1 U10060 ( .B1(n8440), .B2(n8696), .A(n8634), .ZN(n8442) );
  AOI21_X1 U10061 ( .B1(n8634), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8442), .ZN(
        n8441) );
  OAI21_X1 U10062 ( .B1(n8637), .B2(n10043), .A(n8441), .ZN(P2_U3202) );
  INV_X1 U10063 ( .A(n8699), .ZN(n8640) );
  AOI21_X1 U10064 ( .B1(n8634), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8442), .ZN(
        n8443) );
  OAI21_X1 U10065 ( .B1(n8640), .B2(n10043), .A(n8443), .ZN(P2_U3203) );
  AOI22_X1 U10066 ( .A1(n8445), .A2(n8604), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n8634), .ZN(n8446) );
  OAI21_X1 U10067 ( .B1(n8447), .B2(n10043), .A(n8446), .ZN(n8448) );
  AOI21_X1 U10068 ( .B1(n8450), .B2(n8449), .A(n8448), .ZN(n8451) );
  OAI21_X1 U10069 ( .B1(n8444), .B2(n8634), .A(n8451), .ZN(P2_U3204) );
  INV_X1 U10070 ( .A(n8452), .ZN(n8454) );
  OAI22_X1 U10071 ( .A1(n8454), .A2(n10040), .B1(n8616), .B2(n8453), .ZN(n8457) );
  NOR2_X1 U10072 ( .A1(n8455), .A2(n10047), .ZN(n8456) );
  AOI211_X1 U10073 ( .C1(n8605), .C2(n8458), .A(n8457), .B(n8456), .ZN(n8459)
         );
  OAI21_X1 U10074 ( .B1(n8460), .B2(n8634), .A(n8459), .ZN(P2_U3205) );
  AOI21_X1 U10075 ( .B1(n8461), .B2(n8469), .A(n10050), .ZN(n8466) );
  OAI22_X1 U10076 ( .A1(n8463), .A2(n10039), .B1(n8462), .B2(n10037), .ZN(
        n8464) );
  AOI21_X1 U10077 ( .B1(n8466), .B2(n8465), .A(n8464), .ZN(n8703) );
  INV_X1 U10078 ( .A(n8703), .ZN(n8467) );
  AOI21_X1 U10079 ( .B1(n8604), .B2(n8468), .A(n8467), .ZN(n8474) );
  XNOR2_X1 U10080 ( .A(n8470), .B(n8469), .ZN(n8705) );
  OAI22_X1 U10081 ( .A1(n8708), .A2(n10043), .B1(n8471), .B2(n8616), .ZN(n8472) );
  AOI21_X1 U10082 ( .B1(n8705), .B2(n7412), .A(n8472), .ZN(n8473) );
  OAI21_X1 U10083 ( .B1(n8474), .B2(n8634), .A(n8473), .ZN(P2_U3206) );
  XNOR2_X1 U10084 ( .A(n8475), .B(n8476), .ZN(n8711) );
  INV_X1 U10085 ( .A(n8711), .ZN(n8486) );
  XNOR2_X1 U10086 ( .A(n8477), .B(n8476), .ZN(n8480) );
  AOI222_X1 U10087 ( .A1(n8627), .A2(n8480), .B1(n8479), .B2(n8624), .C1(n8478), .C2(n8622), .ZN(n8709) );
  MUX2_X1 U10088 ( .A(n8481), .B(n8709), .S(n8616), .Z(n8485) );
  AOI22_X1 U10089 ( .A1(n8483), .A2(n8605), .B1(n8604), .B2(n8482), .ZN(n8484)
         );
  OAI211_X1 U10090 ( .C1(n8486), .C2(n10047), .A(n8485), .B(n8484), .ZN(
        P2_U3207) );
  XNOR2_X1 U10091 ( .A(n8487), .B(n8488), .ZN(n8720) );
  OAI21_X1 U10092 ( .B1(n8490), .B2(n6300), .A(n8489), .ZN(n8492) );
  AOI222_X1 U10093 ( .A1(n8627), .A2(n8492), .B1(n8491), .B2(n8622), .C1(n8514), .C2(n8624), .ZN(n8715) );
  OAI21_X1 U10094 ( .B1(n8493), .B2(n8615), .A(n8715), .ZN(n8494) );
  NAND2_X1 U10095 ( .A1(n8494), .A2(n8616), .ZN(n8497) );
  AOI22_X1 U10096 ( .A1(n8604), .A2(n8495), .B1(n8634), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8496) );
  OAI211_X1 U10097 ( .C1(n8720), .C2(n10047), .A(n8497), .B(n8496), .ZN(
        P2_U3208) );
  NOR2_X1 U10098 ( .A1(n8722), .A2(n8615), .ZN(n8501) );
  XOR2_X1 U10099 ( .A(n8498), .B(n8505), .Z(n8499) );
  OAI222_X1 U10100 ( .A1(n10039), .A2(n8500), .B1(n10037), .B2(n8529), .C1(
        n10050), .C2(n8499), .ZN(n8721) );
  AOI211_X1 U10101 ( .C1(n8604), .C2(n8502), .A(n8501), .B(n8721), .ZN(n8508)
         );
  NAND2_X1 U10102 ( .A1(n8504), .A2(n8503), .ZN(n8506) );
  XNOR2_X1 U10103 ( .A(n8506), .B(n8505), .ZN(n8650) );
  AOI22_X1 U10104 ( .A1(n8650), .A2(n7412), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n8634), .ZN(n8507) );
  OAI21_X1 U10105 ( .B1(n8508), .B2(n8634), .A(n8507), .ZN(P2_U3209) );
  XNOR2_X1 U10106 ( .A(n8510), .B(n8511), .ZN(n8730) );
  XNOR2_X1 U10107 ( .A(n8512), .B(n8513), .ZN(n8515) );
  AOI222_X1 U10108 ( .A1(n8627), .A2(n8515), .B1(n8514), .B2(n8622), .C1(n8542), .C2(n8624), .ZN(n8726) );
  MUX2_X1 U10109 ( .A(n8516), .B(n8726), .S(n8616), .Z(n8519) );
  AOI22_X1 U10110 ( .A1(n6296), .A2(n8605), .B1(n8604), .B2(n8517), .ZN(n8518)
         );
  OAI211_X1 U10111 ( .C1(n8730), .C2(n10047), .A(n8519), .B(n8518), .ZN(
        P2_U3210) );
  XNOR2_X1 U10112 ( .A(n8520), .B(n4561), .ZN(n8733) );
  INV_X1 U10113 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8531) );
  INV_X1 U10114 ( .A(n8521), .ZN(n8526) );
  NOR3_X1 U10115 ( .A1(n8522), .A2(n8524), .A3(n8523), .ZN(n8525) );
  NOR2_X1 U10116 ( .A1(n8526), .A2(n8525), .ZN(n8527) );
  OAI222_X1 U10117 ( .A1(n10039), .A2(n8529), .B1(n10037), .B2(n8528), .C1(
        n10050), .C2(n8527), .ZN(n8731) );
  INV_X1 U10118 ( .A(n8731), .ZN(n8530) );
  MUX2_X1 U10119 ( .A(n8531), .B(n8530), .S(n8616), .Z(n8535) );
  AOI22_X1 U10120 ( .A1(n8533), .A2(n8605), .B1(n8604), .B2(n8532), .ZN(n8534)
         );
  OAI211_X1 U10121 ( .C1(n8733), .C2(n10047), .A(n8535), .B(n8534), .ZN(
        P2_U3211) );
  XOR2_X1 U10122 ( .A(n8539), .B(n8536), .Z(n8741) );
  INV_X1 U10123 ( .A(n8522), .ZN(n8541) );
  NAND3_X1 U10124 ( .A1(n8537), .A2(n8539), .A3(n8538), .ZN(n8540) );
  NAND2_X1 U10125 ( .A1(n8541), .A2(n8540), .ZN(n8543) );
  AOI222_X1 U10126 ( .A1(n8627), .A2(n8543), .B1(n8542), .B2(n8622), .C1(n8561), .C2(n8624), .ZN(n8736) );
  MUX2_X1 U10127 ( .A(n8544), .B(n8736), .S(n8616), .Z(n8547) );
  AOI22_X1 U10128 ( .A1(n8738), .A2(n8605), .B1(n8604), .B2(n8545), .ZN(n8546)
         );
  OAI211_X1 U10129 ( .C1(n8741), .C2(n10047), .A(n8547), .B(n8546), .ZN(
        P2_U3212) );
  XNOR2_X1 U10130 ( .A(n8550), .B(n8549), .ZN(n8747) );
  OAI21_X1 U10131 ( .B1(n8552), .B2(n8551), .A(n8537), .ZN(n8554) );
  AOI222_X1 U10132 ( .A1(n8627), .A2(n8554), .B1(n8553), .B2(n8622), .C1(n8577), .C2(n8624), .ZN(n8742) );
  MUX2_X1 U10133 ( .A(n8555), .B(n8742), .S(n8616), .Z(n8558) );
  AOI22_X1 U10134 ( .A1(n8744), .A2(n8605), .B1(n8604), .B2(n8556), .ZN(n8557)
         );
  OAI211_X1 U10135 ( .C1(n8747), .C2(n10047), .A(n8558), .B(n8557), .ZN(
        P2_U3213) );
  XNOR2_X1 U10136 ( .A(n8559), .B(n8567), .ZN(n8562) );
  AOI222_X1 U10137 ( .A1(n8627), .A2(n8562), .B1(n8561), .B2(n8622), .C1(n8560), .C2(n8624), .ZN(n8668) );
  OAI22_X1 U10138 ( .A1(n8616), .A2(n8564), .B1(n8563), .B2(n10040), .ZN(n8565) );
  AOI21_X1 U10139 ( .B1(n8566), .B2(n8605), .A(n8565), .ZN(n8570) );
  OR2_X1 U10140 ( .A1(n8568), .A2(n8567), .ZN(n8666) );
  NAND3_X1 U10141 ( .A1(n8666), .A2(n8665), .A3(n7412), .ZN(n8569) );
  OAI211_X1 U10142 ( .C1(n8668), .C2(n8634), .A(n8570), .B(n8569), .ZN(
        P2_U3214) );
  INV_X1 U10143 ( .A(n8571), .ZN(n8584) );
  OAI21_X1 U10144 ( .B1(n8584), .B2(n8572), .A(n8575), .ZN(n8574) );
  NAND2_X1 U10145 ( .A1(n8574), .A2(n8573), .ZN(n8754) );
  XNOR2_X1 U10146 ( .A(n8576), .B(n8575), .ZN(n8578) );
  AOI222_X1 U10147 ( .A1(n8627), .A2(n8578), .B1(n8577), .B2(n8622), .C1(n8599), .C2(n8624), .ZN(n8749) );
  MUX2_X1 U10148 ( .A(n8579), .B(n8749), .S(n8616), .Z(n8583) );
  INV_X1 U10149 ( .A(n8580), .ZN(n8581) );
  AOI22_X1 U10150 ( .A1(n8751), .A2(n8605), .B1(n8604), .B2(n8581), .ZN(n8582)
         );
  OAI211_X1 U10151 ( .C1(n8754), .C2(n10047), .A(n8583), .B(n8582), .ZN(
        P2_U3215) );
  AOI21_X1 U10152 ( .B1(n8586), .B2(n8585), .A(n8584), .ZN(n8758) );
  XNOR2_X1 U10153 ( .A(n8587), .B(n8586), .ZN(n8588) );
  OAI222_X1 U10154 ( .A1(n10039), .A2(n8590), .B1(n10037), .B2(n8589), .C1(
        n8588), .C2(n10050), .ZN(n8673) );
  NAND2_X1 U10155 ( .A1(n8673), .A2(n8616), .ZN(n8595) );
  OAI22_X1 U10156 ( .A1(n8616), .A2(n8592), .B1(n8591), .B2(n10040), .ZN(n8593) );
  AOI21_X1 U10157 ( .B1(n8674), .B2(n8605), .A(n8593), .ZN(n8594) );
  OAI211_X1 U10158 ( .C1(n8758), .C2(n10047), .A(n8595), .B(n8594), .ZN(
        P2_U3216) );
  XNOR2_X1 U10159 ( .A(n8596), .B(n8597), .ZN(n8764) );
  XOR2_X1 U10160 ( .A(n8598), .B(n8597), .Z(n8600) );
  AOI222_X1 U10161 ( .A1(n8627), .A2(n8600), .B1(n8599), .B2(n8622), .C1(n6029), .C2(n8624), .ZN(n8759) );
  MUX2_X1 U10162 ( .A(n8601), .B(n8759), .S(n8616), .Z(n8607) );
  INV_X1 U10163 ( .A(n8602), .ZN(n8603) );
  AOI22_X1 U10164 ( .A1(n8761), .A2(n8605), .B1(n8604), .B2(n8603), .ZN(n8606)
         );
  OAI211_X1 U10165 ( .C1(n8764), .C2(n10047), .A(n8607), .B(n8606), .ZN(
        P2_U3217) );
  XNOR2_X1 U10166 ( .A(n8608), .B(n8610), .ZN(n8768) );
  XNOR2_X1 U10167 ( .A(n8609), .B(n8610), .ZN(n8611) );
  OAI222_X1 U10168 ( .A1(n10039), .A2(n8613), .B1(n10037), .B2(n8612), .C1(
        n10050), .C2(n8611), .ZN(n8765) );
  OAI22_X1 U10169 ( .A1(n8767), .A2(n8615), .B1(n8614), .B2(n10040), .ZN(n8617) );
  OAI21_X1 U10170 ( .B1(n8765), .B2(n8617), .A(n8616), .ZN(n8619) );
  NAND2_X1 U10171 ( .A1(n8634), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8618) );
  OAI211_X1 U10172 ( .C1(n8768), .C2(n10047), .A(n8619), .B(n8618), .ZN(
        P2_U3219) );
  NOR2_X1 U10173 ( .A1(n10040), .A2(n8620), .ZN(n8629) );
  XNOR2_X1 U10174 ( .A(n8621), .B(n8632), .ZN(n8626) );
  AOI222_X1 U10175 ( .A1(n8627), .A2(n8626), .B1(n8625), .B2(n8624), .C1(n8623), .C2(n8622), .ZN(n8771) );
  INV_X1 U10176 ( .A(n8771), .ZN(n8628) );
  AOI211_X1 U10177 ( .C1(n8630), .C2(n8773), .A(n8629), .B(n8628), .ZN(n8635)
         );
  XOR2_X1 U10178 ( .A(n8631), .B(n8632), .Z(n8776) );
  AOI22_X1 U10179 ( .A1(n8776), .A2(n7412), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n8634), .ZN(n8633) );
  OAI21_X1 U10180 ( .B1(n8635), .B2(n8634), .A(n8633), .ZN(P2_U3220) );
  NOR2_X1 U10181 ( .A1(n8696), .A2(n10122), .ZN(n8638) );
  AOI21_X1 U10182 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10122), .A(n8638), .ZN(
        n8636) );
  OAI21_X1 U10183 ( .B1(n8637), .B2(n8656), .A(n8636), .ZN(P2_U3490) );
  AOI21_X1 U10184 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n10122), .A(n8638), .ZN(
        n8639) );
  OAI21_X1 U10185 ( .B1(n8640), .B2(n8656), .A(n8639), .ZN(P2_U3489) );
  INV_X1 U10186 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8641) );
  MUX2_X1 U10187 ( .A(n8641), .B(n8703), .S(n10124), .Z(n8643) );
  NAND2_X1 U10188 ( .A1(n8705), .A2(n8687), .ZN(n8642) );
  OAI211_X1 U10189 ( .C1(n8708), .C2(n8656), .A(n8643), .B(n8642), .ZN(
        P2_U3486) );
  INV_X1 U10190 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8644) );
  MUX2_X1 U10191 ( .A(n8644), .B(n8709), .S(n10124), .Z(n8646) );
  NAND2_X1 U10192 ( .A1(n8711), .A2(n8687), .ZN(n8645) );
  OAI211_X1 U10193 ( .C1(n8714), .C2(n8656), .A(n8646), .B(n8645), .ZN(
        P2_U3485) );
  INV_X1 U10194 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8647) );
  MUX2_X1 U10195 ( .A(n8647), .B(n8715), .S(n10124), .Z(n8649) );
  NAND2_X1 U10196 ( .A1(n8717), .A2(n8686), .ZN(n8648) );
  OAI211_X1 U10197 ( .C1(n8720), .C2(n8694), .A(n8649), .B(n8648), .ZN(
        P2_U3484) );
  MUX2_X1 U10198 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8721), .S(n10124), .Z(
        n8652) );
  INV_X1 U10199 ( .A(n8650), .ZN(n8723) );
  OAI22_X1 U10200 ( .A1(n8723), .A2(n8694), .B1(n8722), .B2(n8656), .ZN(n8651)
         );
  OR2_X1 U10201 ( .A1(n8652), .A2(n8651), .ZN(P2_U3483) );
  INV_X1 U10202 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8653) );
  MUX2_X1 U10203 ( .A(n8653), .B(n8726), .S(n10124), .Z(n8655) );
  NAND2_X1 U10204 ( .A1(n6296), .A2(n8686), .ZN(n8654) );
  OAI211_X1 U10205 ( .C1(n8730), .C2(n8694), .A(n8655), .B(n8654), .ZN(
        P2_U3482) );
  MUX2_X1 U10206 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8731), .S(n10124), .Z(
        n8658) );
  OAI22_X1 U10207 ( .A1(n8733), .A2(n8694), .B1(n8732), .B2(n8656), .ZN(n8657)
         );
  OR2_X1 U10208 ( .A1(n8658), .A2(n8657), .ZN(P2_U3481) );
  MUX2_X1 U10209 ( .A(n8659), .B(n8736), .S(n10124), .Z(n8661) );
  NAND2_X1 U10210 ( .A1(n8738), .A2(n8686), .ZN(n8660) );
  OAI211_X1 U10211 ( .C1(n8694), .C2(n8741), .A(n8661), .B(n8660), .ZN(
        P2_U3480) );
  MUX2_X1 U10212 ( .A(n8662), .B(n8742), .S(n10124), .Z(n8664) );
  NAND2_X1 U10213 ( .A1(n8744), .A2(n8686), .ZN(n8663) );
  OAI211_X1 U10214 ( .C1(n8747), .C2(n8694), .A(n8664), .B(n8663), .ZN(
        P2_U3479) );
  NAND3_X1 U10215 ( .A1(n8666), .A2(n8665), .A3(n10074), .ZN(n8667) );
  OAI211_X1 U10216 ( .C1(n8669), .C2(n10102), .A(n8668), .B(n8667), .ZN(n8748)
         );
  MUX2_X1 U10217 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8748), .S(n10124), .Z(
        P2_U3478) );
  MUX2_X1 U10218 ( .A(n8670), .B(n8749), .S(n10124), .Z(n8672) );
  NAND2_X1 U10219 ( .A1(n8751), .A2(n8686), .ZN(n8671) );
  OAI211_X1 U10220 ( .C1(n8694), .C2(n8754), .A(n8672), .B(n8671), .ZN(
        P2_U3477) );
  AOI21_X1 U10221 ( .B1(n10081), .B2(n8674), .A(n8673), .ZN(n8755) );
  MUX2_X1 U10222 ( .A(n8675), .B(n8755), .S(n10124), .Z(n8676) );
  OAI21_X1 U10223 ( .B1(n8758), .B2(n8694), .A(n8676), .ZN(P2_U3476) );
  MUX2_X1 U10224 ( .A(n8677), .B(n8759), .S(n10124), .Z(n8679) );
  NAND2_X1 U10225 ( .A1(n8761), .A2(n8686), .ZN(n8678) );
  OAI211_X1 U10226 ( .C1(n8764), .C2(n8694), .A(n8679), .B(n8678), .ZN(
        P2_U3475) );
  INV_X1 U10227 ( .A(n8765), .ZN(n8680) );
  MUX2_X1 U10228 ( .A(n8681), .B(n8680), .S(n10124), .Z(n8684) );
  NAND2_X1 U10229 ( .A1(n8682), .A2(n8686), .ZN(n8683) );
  OAI211_X1 U10230 ( .C1(n8768), .C2(n8694), .A(n8684), .B(n8683), .ZN(
        P2_U3473) );
  MUX2_X1 U10231 ( .A(n8685), .B(n8771), .S(n10124), .Z(n8689) );
  AOI22_X1 U10232 ( .A1(n8776), .A2(n8687), .B1(n8686), .B2(n8773), .ZN(n8688)
         );
  NAND2_X1 U10233 ( .A1(n8689), .A2(n8688), .ZN(P2_U3472) );
  AOI21_X1 U10234 ( .B1(n10081), .B2(n8691), .A(n8690), .ZN(n8779) );
  MUX2_X1 U10235 ( .A(n8692), .B(n8779), .S(n10124), .Z(n8693) );
  OAI21_X1 U10236 ( .B1(n8783), .B2(n8694), .A(n8693), .ZN(P2_U3471) );
  INV_X1 U10237 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8698) );
  NAND2_X1 U10238 ( .A1(n8695), .A2(n8774), .ZN(n8697) );
  OR2_X1 U10239 ( .A1(n8696), .A2(n10108), .ZN(n8700) );
  OAI211_X1 U10240 ( .C1(n8698), .C2(n10110), .A(n8697), .B(n8700), .ZN(
        P2_U3458) );
  INV_X1 U10241 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8702) );
  NAND2_X1 U10242 ( .A1(n8699), .A2(n8774), .ZN(n8701) );
  OAI211_X1 U10243 ( .C1(n8702), .C2(n10110), .A(n8701), .B(n8700), .ZN(
        P2_U3457) );
  INV_X1 U10244 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8704) );
  MUX2_X1 U10245 ( .A(n8704), .B(n8703), .S(n10110), .Z(n8707) );
  INV_X1 U10246 ( .A(n8782), .ZN(n8775) );
  NAND2_X1 U10247 ( .A1(n8705), .A2(n8775), .ZN(n8706) );
  OAI211_X1 U10248 ( .C1(n8708), .C2(n8766), .A(n8707), .B(n8706), .ZN(
        P2_U3454) );
  INV_X1 U10249 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8710) );
  MUX2_X1 U10250 ( .A(n8710), .B(n8709), .S(n10110), .Z(n8713) );
  NAND2_X1 U10251 ( .A1(n8711), .A2(n8775), .ZN(n8712) );
  OAI211_X1 U10252 ( .C1(n8714), .C2(n8766), .A(n8713), .B(n8712), .ZN(
        P2_U3453) );
  INV_X1 U10253 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8716) );
  MUX2_X1 U10254 ( .A(n8716), .B(n8715), .S(n10110), .Z(n8719) );
  NAND2_X1 U10255 ( .A1(n8717), .A2(n8774), .ZN(n8718) );
  OAI211_X1 U10256 ( .C1(n8720), .C2(n8782), .A(n8719), .B(n8718), .ZN(
        P2_U3452) );
  MUX2_X1 U10257 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8721), .S(n10110), .Z(
        n8725) );
  OAI22_X1 U10258 ( .A1(n8723), .A2(n8782), .B1(n8722), .B2(n8766), .ZN(n8724)
         );
  OR2_X1 U10259 ( .A1(n8725), .A2(n8724), .ZN(P2_U3451) );
  INV_X1 U10260 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8727) );
  MUX2_X1 U10261 ( .A(n8727), .B(n8726), .S(n10110), .Z(n8729) );
  NAND2_X1 U10262 ( .A1(n6296), .A2(n8774), .ZN(n8728) );
  OAI211_X1 U10263 ( .C1(n8730), .C2(n8782), .A(n8729), .B(n8728), .ZN(
        P2_U3450) );
  MUX2_X1 U10264 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8731), .S(n10110), .Z(
        n8735) );
  OAI22_X1 U10265 ( .A1(n8733), .A2(n8782), .B1(n8732), .B2(n8766), .ZN(n8734)
         );
  OR2_X1 U10266 ( .A1(n8735), .A2(n8734), .ZN(P2_U3449) );
  MUX2_X1 U10267 ( .A(n8737), .B(n8736), .S(n10110), .Z(n8740) );
  NAND2_X1 U10268 ( .A1(n8738), .A2(n8774), .ZN(n8739) );
  OAI211_X1 U10269 ( .C1(n8741), .C2(n8782), .A(n8740), .B(n8739), .ZN(
        P2_U3448) );
  MUX2_X1 U10270 ( .A(n8743), .B(n8742), .S(n10110), .Z(n8746) );
  NAND2_X1 U10271 ( .A1(n8744), .A2(n8774), .ZN(n8745) );
  OAI211_X1 U10272 ( .C1(n8747), .C2(n8782), .A(n8746), .B(n8745), .ZN(
        P2_U3447) );
  MUX2_X1 U10273 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8748), .S(n10110), .Z(
        P2_U3446) );
  INV_X1 U10274 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8750) );
  MUX2_X1 U10275 ( .A(n8750), .B(n8749), .S(n10110), .Z(n8753) );
  NAND2_X1 U10276 ( .A1(n8751), .A2(n8774), .ZN(n8752) );
  OAI211_X1 U10277 ( .C1(n8754), .C2(n8782), .A(n8753), .B(n8752), .ZN(
        P2_U3444) );
  INV_X1 U10278 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8756) );
  MUX2_X1 U10279 ( .A(n8756), .B(n8755), .S(n10110), .Z(n8757) );
  OAI21_X1 U10280 ( .B1(n8758), .B2(n8782), .A(n8757), .ZN(P2_U3441) );
  INV_X1 U10281 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8760) );
  MUX2_X1 U10282 ( .A(n8760), .B(n8759), .S(n10110), .Z(n8763) );
  NAND2_X1 U10283 ( .A1(n8761), .A2(n8774), .ZN(n8762) );
  OAI211_X1 U10284 ( .C1(n8764), .C2(n8782), .A(n8763), .B(n8762), .ZN(
        P2_U3438) );
  MUX2_X1 U10285 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8765), .S(n10110), .Z(
        n8770) );
  OAI22_X1 U10286 ( .A1(n8768), .A2(n8782), .B1(n8767), .B2(n8766), .ZN(n8769)
         );
  OR2_X1 U10287 ( .A1(n8770), .A2(n8769), .ZN(P2_U3432) );
  INV_X1 U10288 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8772) );
  MUX2_X1 U10289 ( .A(n8772), .B(n8771), .S(n10110), .Z(n8778) );
  AOI22_X1 U10290 ( .A1(n8776), .A2(n8775), .B1(n8774), .B2(n8773), .ZN(n8777)
         );
  NAND2_X1 U10291 ( .A1(n8778), .A2(n8777), .ZN(P2_U3429) );
  INV_X1 U10292 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8780) );
  MUX2_X1 U10293 ( .A(n8780), .B(n8779), .S(n10110), .Z(n8781) );
  OAI21_X1 U10294 ( .B1(n8783), .B2(n8782), .A(n8781), .ZN(P2_U3426) );
  INV_X1 U10295 ( .A(n8975), .ZN(n9761) );
  NOR4_X1 U10296 ( .A1(n4581), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n8784), .ZN(n8785) );
  AOI21_X1 U10297 ( .B1(n8786), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8785), .ZN(
        n8787) );
  OAI21_X1 U10298 ( .B1(n9761), .B2(n8788), .A(n8787), .ZN(P2_U3264) );
  OAI222_X1 U10299 ( .A1(n8803), .A2(n8790), .B1(n8800), .B2(n6462), .C1(
        P2_U3151), .C2(n8789), .ZN(P2_U3266) );
  NAND2_X1 U10300 ( .A1(n8791), .A2(n8795), .ZN(n8793) );
  OAI211_X1 U10301 ( .C1(n8800), .C2(n8794), .A(n8793), .B(n8792), .ZN(
        P2_U3267) );
  NAND2_X1 U10302 ( .A1(n9762), .A2(n8795), .ZN(n8797) );
  OAI211_X1 U10303 ( .C1(n8800), .C2(n8798), .A(n8797), .B(n8796), .ZN(
        P2_U3268) );
  INV_X1 U10304 ( .A(n8799), .ZN(n9768) );
  OAI222_X1 U10305 ( .A1(n8803), .A2(n9768), .B1(P2_U3151), .B2(n8802), .C1(
        n8801), .C2(n8800), .ZN(P2_U3269) );
  MUX2_X1 U10306 ( .A(n8804), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI21_X1 U10307 ( .B1(n8951), .B2(n8806), .A(n8805), .ZN(n8808) );
  OAI21_X1 U10308 ( .B1(n8808), .B2(n8807), .A(n9806), .ZN(n8814) );
  AND2_X1 U10309 ( .A1(n9234), .A2(n9563), .ZN(n8809) );
  AOI21_X1 U10310 ( .B1(n9232), .B2(n4309), .A(n8809), .ZN(n9397) );
  INV_X1 U10311 ( .A(n8810), .ZN(n9403) );
  AOI22_X1 U10312 ( .A1(n9403), .A2(n8971), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n8811) );
  OAI21_X1 U10313 ( .B1(n9397), .B2(n8955), .A(n8811), .ZN(n8812) );
  AOI21_X1 U10314 ( .B1(n9402), .B2(n8957), .A(n8812), .ZN(n8813) );
  NAND2_X1 U10315 ( .A1(n8814), .A2(n8813), .ZN(P1_U3214) );
  NAND2_X1 U10316 ( .A1(n8816), .A2(n8815), .ZN(n8818) );
  XNOR2_X1 U10317 ( .A(n8818), .B(n8817), .ZN(n8823) );
  OAI22_X1 U10318 ( .A1(n9810), .A2(n9596), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8819), .ZN(n8821) );
  OAI22_X1 U10319 ( .A1(n8967), .A2(n9584), .B1(n9586), .B2(n8964), .ZN(n8820)
         );
  AOI211_X1 U10320 ( .C1(n9691), .C2(n8957), .A(n8821), .B(n8820), .ZN(n8822)
         );
  OAI21_X1 U10321 ( .B1(n8823), .B2(n8946), .A(n8822), .ZN(P1_U3215) );
  INV_X1 U10322 ( .A(n8824), .ZN(n8931) );
  INV_X1 U10323 ( .A(n8825), .ZN(n8827) );
  NOR3_X1 U10324 ( .A1(n8931), .A2(n8827), .A3(n8826), .ZN(n8830) );
  INV_X1 U10325 ( .A(n8828), .ZN(n8829) );
  OAI21_X1 U10326 ( .B1(n8830), .B2(n8829), .A(n9806), .ZN(n8836) );
  NAND2_X1 U10327 ( .A1(n9235), .A2(n4309), .ZN(n8832) );
  NAND2_X1 U10328 ( .A1(n9236), .A2(n9563), .ZN(n8831) );
  NAND2_X1 U10329 ( .A1(n8832), .A2(n8831), .ZN(n9649) );
  OAI22_X1 U10330 ( .A1(n9464), .A2(n9810), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8833), .ZN(n8834) );
  AOI21_X1 U10331 ( .B1(n9649), .B2(n9801), .A(n8834), .ZN(n8835) );
  OAI211_X1 U10332 ( .C1(n4480), .C2(n9803), .A(n8836), .B(n8835), .ZN(
        P1_U3216) );
  XOR2_X1 U10333 ( .A(n8837), .B(n8838), .Z(n8940) );
  AOI22_X1 U10334 ( .A1(n8940), .A2(n8941), .B1(n8838), .B2(n8837), .ZN(n8841)
         );
  NOR2_X1 U10335 ( .A1(n8924), .A2(n8839), .ZN(n8840) );
  XNOR2_X1 U10336 ( .A(n8841), .B(n8840), .ZN(n8849) );
  INV_X1 U10337 ( .A(n9532), .ZN(n8843) );
  OAI22_X1 U10338 ( .A1(n9810), .A2(n8843), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8842), .ZN(n8847) );
  OAI22_X1 U10339 ( .A1(n8967), .A2(n8845), .B1(n8844), .B2(n8964), .ZN(n8846)
         );
  AOI211_X1 U10340 ( .C1(n9531), .C2(n8957), .A(n8847), .B(n8846), .ZN(n8848)
         );
  OAI21_X1 U10341 ( .B1(n8849), .B2(n8946), .A(n8848), .ZN(P1_U3219) );
  AOI21_X1 U10342 ( .B1(n8852), .B2(n8851), .A(n8850), .ZN(n8853) );
  OR2_X1 U10343 ( .A1(n8853), .A2(n8946), .ZN(n8862) );
  INV_X1 U10344 ( .A(n8854), .ZN(n8855) );
  AOI21_X1 U10345 ( .B1(n9801), .B2(n8856), .A(n8855), .ZN(n8861) );
  NAND2_X1 U10346 ( .A1(n8957), .A2(n8857), .ZN(n8860) );
  OR2_X1 U10347 ( .A1(n9810), .A2(n8858), .ZN(n8859) );
  NAND4_X1 U10348 ( .A1(n8862), .A2(n8861), .A3(n8860), .A4(n8859), .ZN(
        P1_U3221) );
  OAI21_X1 U10349 ( .B1(n8865), .B2(n8863), .A(n8864), .ZN(n8866) );
  NAND2_X1 U10350 ( .A1(n8866), .A2(n9806), .ZN(n8871) );
  AND2_X1 U10351 ( .A1(n9525), .A2(n9563), .ZN(n8867) );
  AOI21_X1 U10352 ( .B1(n9236), .B2(n4309), .A(n8867), .ZN(n9493) );
  OAI22_X1 U10353 ( .A1(n9493), .A2(n8955), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8868), .ZN(n8869) );
  AOI21_X1 U10354 ( .B1(n9496), .B2(n8971), .A(n8869), .ZN(n8870) );
  OAI211_X1 U10355 ( .C1(n4536), .C2(n9803), .A(n8871), .B(n8870), .ZN(
        P1_U3223) );
  OAI21_X1 U10356 ( .B1(n8874), .B2(n8873), .A(n8872), .ZN(n8879) );
  AND2_X1 U10357 ( .A1(n9235), .A2(n9563), .ZN(n8875) );
  AOI21_X1 U10358 ( .B1(n9234), .B2(n4309), .A(n8875), .ZN(n9429) );
  NAND2_X1 U10359 ( .A1(n9436), .A2(n8957), .ZN(n8877) );
  AOI22_X1 U10360 ( .A1(n9437), .A2(n8971), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n8876) );
  OAI211_X1 U10361 ( .C1(n9429), .C2(n8955), .A(n8877), .B(n8876), .ZN(n8878)
         );
  AOI21_X1 U10362 ( .B1(n8879), .B2(n9806), .A(n8878), .ZN(n8880) );
  INV_X1 U10363 ( .A(n8880), .ZN(P1_U3225) );
  OAI21_X1 U10364 ( .B1(n8883), .B2(n8882), .A(n8881), .ZN(n8884) );
  NAND2_X1 U10365 ( .A1(n8884), .A2(n9806), .ZN(n8888) );
  AND2_X1 U10366 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9865) );
  OAI22_X1 U10367 ( .A1(n8967), .A2(n9586), .B1(n9545), .B2(n8964), .ZN(n8885)
         );
  AOI211_X1 U10368 ( .C1(n8971), .C2(n8886), .A(n9865), .B(n8885), .ZN(n8887)
         );
  OAI211_X1 U10369 ( .C1(n8889), .C2(n9803), .A(n8888), .B(n8887), .ZN(
        P1_U3226) );
  NAND2_X1 U10370 ( .A1(n8890), .A2(n9806), .ZN(n8897) );
  AOI21_X1 U10371 ( .B1(n8881), .B2(n8892), .A(n8891), .ZN(n8896) );
  AOI22_X1 U10372 ( .A1(n8903), .A2(n9562), .B1(n8904), .B2(n9565), .ZN(n8893)
         );
  NAND2_X1 U10373 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9885) );
  OAI211_X1 U10374 ( .C1(n9810), .C2(n9575), .A(n8893), .B(n9885), .ZN(n8894)
         );
  AOI21_X1 U10375 ( .B1(n9574), .B2(n8957), .A(n8894), .ZN(n8895) );
  OAI21_X1 U10376 ( .B1(n8897), .B2(n8896), .A(n8895), .ZN(P1_U3228) );
  INV_X1 U10377 ( .A(n8899), .ZN(n8900) );
  NAND3_X1 U10378 ( .A1(n8828), .A2(n8901), .A3(n8900), .ZN(n8902) );
  AOI21_X1 U10379 ( .B1(n8898), .B2(n8902), .A(n8946), .ZN(n8908) );
  AOI22_X1 U10380 ( .A1(n9453), .A2(n8971), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8906) );
  AOI22_X1 U10381 ( .A1(n9449), .A2(n8904), .B1(n8903), .B2(n9448), .ZN(n8905)
         );
  OAI211_X1 U10382 ( .C1(n9456), .C2(n9803), .A(n8906), .B(n8905), .ZN(n8907)
         );
  OR2_X1 U10383 ( .A1(n8908), .A2(n8907), .ZN(P1_U3229) );
  OAI211_X1 U10384 ( .C1(n8911), .C2(n8910), .A(n8909), .B(n9806), .ZN(n8918)
         );
  INV_X1 U10385 ( .A(n8912), .ZN(n8913) );
  AOI22_X1 U10386 ( .A1(n8914), .A2(n8957), .B1(n8971), .B2(n8913), .ZN(n8917)
         );
  NAND2_X1 U10387 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9289) );
  OR2_X1 U10388 ( .A1(n8955), .A2(n8915), .ZN(n8916) );
  NAND4_X1 U10389 ( .A1(n8918), .A2(n8917), .A3(n9289), .A4(n8916), .ZN(
        P1_U3230) );
  NAND2_X1 U10390 ( .A1(n9237), .A2(n4309), .ZN(n8920) );
  NAND2_X1 U10391 ( .A1(n9238), .A2(n9563), .ZN(n8919) );
  NAND2_X1 U10392 ( .A1(n8920), .A2(n8919), .ZN(n9505) );
  AOI22_X1 U10393 ( .A1(n9505), .A2(n9801), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n8921) );
  OAI21_X1 U10394 ( .B1(n9513), .B2(n9810), .A(n8921), .ZN(n8929) );
  INV_X1 U10395 ( .A(n8922), .ZN(n8925) );
  OAI21_X1 U10396 ( .B1(n8925), .B2(n8924), .A(n8923), .ZN(n8927) );
  AOI21_X1 U10397 ( .B1(n8927), .B2(n8926), .A(n8946), .ZN(n8928) );
  AOI211_X1 U10398 ( .C1(n9512), .C2(n8957), .A(n8929), .B(n8928), .ZN(n8930)
         );
  INV_X1 U10399 ( .A(n8930), .ZN(P1_U3233) );
  AOI21_X1 U10400 ( .B1(n8933), .B2(n8932), .A(n8931), .ZN(n8939) );
  NAND2_X1 U10401 ( .A1(n9448), .A2(n4309), .ZN(n8935) );
  NAND2_X1 U10402 ( .A1(n9237), .A2(n9563), .ZN(n8934) );
  NAND2_X1 U10403 ( .A1(n8935), .A2(n8934), .ZN(n9474) );
  AOI22_X1 U10404 ( .A1(n9474), .A2(n9801), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n8936) );
  OAI21_X1 U10405 ( .B1(n9479), .B2(n9810), .A(n8936), .ZN(n8937) );
  AOI21_X1 U10406 ( .B1(n9484), .B2(n8957), .A(n8937), .ZN(n8938) );
  OAI21_X1 U10407 ( .B1(n8939), .B2(n8946), .A(n8938), .ZN(P1_U3235) );
  XOR2_X1 U10408 ( .A(n8941), .B(n8940), .Z(n8947) );
  OAI22_X1 U10409 ( .A1(n9810), .A2(n9549), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8942), .ZN(n8944) );
  OAI22_X1 U10410 ( .A1(n8967), .A2(n9545), .B1(n9546), .B2(n8964), .ZN(n8943)
         );
  AOI211_X1 U10411 ( .C1(n9677), .C2(n8957), .A(n8944), .B(n8943), .ZN(n8945)
         );
  OAI21_X1 U10412 ( .B1(n8947), .B2(n8946), .A(n8945), .ZN(P1_U3238) );
  INV_X1 U10413 ( .A(n8872), .ZN(n8950) );
  OAI21_X1 U10414 ( .B1(n8950), .B2(n8949), .A(n8948), .ZN(n8952) );
  NAND3_X1 U10415 ( .A1(n8952), .A2(n9806), .A3(n8951), .ZN(n8959) );
  AND2_X1 U10416 ( .A1(n9449), .A2(n9563), .ZN(n8953) );
  AOI21_X1 U10417 ( .B1(n9233), .B2(n4309), .A(n8953), .ZN(n9411) );
  AOI22_X1 U10418 ( .A1(n9418), .A2(n8971), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n8954) );
  OAI21_X1 U10419 ( .B1(n9411), .B2(n8955), .A(n8954), .ZN(n8956) );
  AOI21_X1 U10420 ( .B1(n9417), .B2(n8957), .A(n8956), .ZN(n8958) );
  NAND2_X1 U10421 ( .A1(n8959), .A2(n8958), .ZN(P1_U3240) );
  OAI21_X1 U10422 ( .B1(n8962), .B2(n8961), .A(n8960), .ZN(n8963) );
  NAND2_X1 U10423 ( .A1(n8963), .A2(n9806), .ZN(n8973) );
  NAND2_X1 U10424 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9858) );
  INV_X1 U10425 ( .A(n9858), .ZN(n8969) );
  OAI22_X1 U10426 ( .A1(n8967), .A2(n8966), .B1(n8965), .B2(n8964), .ZN(n8968)
         );
  AOI211_X1 U10427 ( .C1(n8971), .C2(n8970), .A(n8969), .B(n8968), .ZN(n8972)
         );
  OAI211_X1 U10428 ( .C1(n8974), .C2(n9803), .A(n8973), .B(n8972), .ZN(
        P1_U3241) );
  NAND2_X1 U10429 ( .A1(n8975), .A2(n9080), .ZN(n8977) );
  NAND2_X1 U10430 ( .A1(n5037), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8976) );
  INV_X1 U10431 ( .A(n9706), .ZN(n8978) );
  INV_X1 U10432 ( .A(n9355), .ZN(n9203) );
  AOI21_X1 U10433 ( .B1(n9355), .B2(n4627), .A(n9213), .ZN(n9086) );
  NOR2_X1 U10434 ( .A1(n9738), .A2(n9525), .ZN(n9048) );
  NOR2_X1 U10435 ( .A1(n9048), .A2(n4710), .ZN(n9040) );
  INV_X1 U10436 ( .A(n9031), .ZN(n8979) );
  NOR2_X1 U10437 ( .A1(n8979), .A2(n9166), .ZN(n9029) );
  INV_X1 U10438 ( .A(n9029), .ZN(n8980) );
  OAI211_X1 U10439 ( .C1(n8981), .C2(n4628), .A(n8980), .B(n9557), .ZN(n9036)
         );
  OAI21_X1 U10440 ( .B1(n9030), .B2(n9586), .A(n9125), .ZN(n9035) );
  INV_X1 U10441 ( .A(n9149), .ZN(n8984) );
  NOR3_X1 U10442 ( .A1(n8989), .A2(n8988), .A3(n8984), .ZN(n8986) );
  NAND2_X1 U10443 ( .A1(n8990), .A2(n8985), .ZN(n9152) );
  OAI211_X1 U10444 ( .C1(n8986), .C2(n9152), .A(n9155), .B(n8993), .ZN(n8987)
         );
  NAND2_X1 U10445 ( .A1(n6503), .A2(n9251), .ZN(n9150) );
  NAND2_X1 U10446 ( .A1(n9155), .A2(n9150), .ZN(n8991) );
  OAI211_X1 U10447 ( .C1(n8992), .C2(n8991), .A(n9097), .B(n8990), .ZN(n8994)
         );
  AND2_X1 U10448 ( .A1(n8997), .A2(n8996), .ZN(n8998) );
  MUX2_X1 U10449 ( .A(n8999), .B(n8998), .S(n9125), .Z(n9004) );
  NAND2_X1 U10450 ( .A1(n9005), .A2(n9000), .ZN(n9001) );
  MUX2_X1 U10451 ( .A(n9002), .B(n9001), .S(n9125), .Z(n9003) );
  INV_X1 U10452 ( .A(n9005), .ZN(n9006) );
  NAND2_X1 U10453 ( .A1(n9015), .A2(n9009), .ZN(n9161) );
  NOR3_X1 U10454 ( .A1(n9011), .A2(n9006), .A3(n9161), .ZN(n9007) );
  OAI211_X1 U10455 ( .C1(n9161), .C2(n9013), .A(n9017), .B(n9012), .ZN(n9165)
         );
  OAI21_X1 U10456 ( .B1(n9007), .B2(n9165), .A(n9162), .ZN(n9020) );
  INV_X1 U10457 ( .A(n9008), .ZN(n9010) );
  OAI21_X1 U10458 ( .B1(n9011), .B2(n9010), .A(n9009), .ZN(n9014) );
  NAND3_X1 U10459 ( .A1(n9014), .A2(n9013), .A3(n9012), .ZN(n9016) );
  NAND3_X1 U10460 ( .A1(n9016), .A2(n9162), .A3(n9015), .ZN(n9018) );
  NAND2_X1 U10461 ( .A1(n9018), .A2(n9017), .ZN(n9019) );
  MUX2_X1 U10462 ( .A(n9020), .B(n9019), .S(n9125), .Z(n9024) );
  NAND2_X1 U10463 ( .A1(n9026), .A2(n9027), .ZN(n9090) );
  AOI211_X1 U10464 ( .C1(n9024), .C2(n9025), .A(n4697), .B(n9090), .ZN(n9023)
         );
  INV_X1 U10465 ( .A(n9026), .ZN(n9022) );
  NAND2_X1 U10466 ( .A1(n9031), .A2(n9021), .ZN(n9170) );
  NOR3_X1 U10467 ( .A1(n9023), .A2(n9022), .A3(n9170), .ZN(n9034) );
  AND2_X1 U10468 ( .A1(n9024), .A2(n9163), .ZN(n9028) );
  NAND2_X1 U10469 ( .A1(n9026), .A2(n9025), .ZN(n9143) );
  OAI21_X1 U10470 ( .B1(n9028), .B2(n9143), .A(n9027), .ZN(n9032) );
  AOI211_X1 U10471 ( .C1(n9032), .C2(n9031), .A(n9030), .B(n9029), .ZN(n9033)
         );
  NAND2_X1 U10472 ( .A1(n9175), .A2(n9037), .ZN(n9172) );
  AND3_X1 U10473 ( .A1(n9038), .A2(n9047), .A3(n9174), .ZN(n9039) );
  MUX2_X1 U10474 ( .A(n9040), .B(n9039), .S(n9125), .Z(n9052) );
  NAND2_X1 U10475 ( .A1(n9042), .A2(n9041), .ZN(n9176) );
  INV_X1 U10476 ( .A(n9175), .ZN(n9043) );
  NOR2_X1 U10477 ( .A1(n9043), .A2(n9125), .ZN(n9044) );
  OAI211_X1 U10478 ( .C1(n9045), .C2(n9176), .A(n9044), .B(n9174), .ZN(n9051)
         );
  OR2_X1 U10479 ( .A1(n9495), .A2(n9046), .ZN(n9132) );
  NAND2_X1 U10480 ( .A1(n9132), .A2(n9047), .ZN(n9178) );
  INV_X1 U10481 ( .A(n9048), .ZN(n9049) );
  NAND2_X1 U10482 ( .A1(n9053), .A2(n9049), .ZN(n9131) );
  MUX2_X1 U10483 ( .A(n9178), .B(n9131), .S(n9125), .Z(n9050) );
  INV_X1 U10484 ( .A(n9053), .ZN(n9055) );
  INV_X1 U10485 ( .A(n9132), .ZN(n9054) );
  MUX2_X1 U10486 ( .A(n9055), .B(n9054), .S(n9125), .Z(n9056) );
  NAND2_X1 U10487 ( .A1(n9060), .A2(n9057), .ZN(n9130) );
  NAND2_X1 U10488 ( .A1(n9130), .A2(n9059), .ZN(n9062) );
  NAND2_X1 U10489 ( .A1(n9059), .A2(n9058), .ZN(n9061) );
  NAND2_X1 U10490 ( .A1(n9061), .A2(n9060), .ZN(n9133) );
  MUX2_X1 U10491 ( .A(n9062), .B(n9133), .S(n9125), .Z(n9063) );
  MUX2_X1 U10492 ( .A(n9134), .B(n9424), .S(n9125), .Z(n9064) );
  INV_X1 U10493 ( .A(n9139), .ZN(n9065) );
  NOR2_X1 U10494 ( .A1(n9069), .A2(n9065), .ZN(n9067) );
  NAND2_X1 U10495 ( .A1(n9127), .A2(n9137), .ZN(n9068) );
  OAI21_X1 U10496 ( .B1(n9067), .B2(n9068), .A(n9066), .ZN(n9072) );
  AOI21_X1 U10497 ( .B1(n9069), .B2(n9139), .A(n9068), .ZN(n9070) );
  NOR2_X1 U10498 ( .A1(n9070), .A2(n9197), .ZN(n9071) );
  NAND2_X1 U10499 ( .A1(n9074), .A2(n9073), .ZN(n9141) );
  OAI21_X1 U10500 ( .B1(n9141), .B2(n9075), .A(n9183), .ZN(n9076) );
  MUX2_X1 U10501 ( .A(n9184), .B(n9186), .S(n9125), .Z(n9077) );
  OAI21_X1 U10502 ( .B1(n9079), .B2(n9078), .A(n9077), .ZN(n9083) );
  NAND2_X1 U10503 ( .A1(n7713), .A2(n9080), .ZN(n9082) );
  NAND2_X1 U10504 ( .A1(n5037), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9081) );
  MUX2_X1 U10505 ( .A(n9083), .B(n9125), .S(n9620), .Z(n9085) );
  INV_X1 U10506 ( .A(n9083), .ZN(n9084) );
  AOI21_X1 U10507 ( .B1(n9189), .B2(n9125), .A(n9089), .ZN(n9231) );
  INV_X1 U10508 ( .A(n9087), .ZN(n9124) );
  NOR2_X1 U10509 ( .A1(n9123), .A2(n9088), .ZN(n9224) );
  OAI211_X1 U10510 ( .C1(n9190), .C2(n4315), .A(n9124), .B(n9224), .ZN(n9230)
         );
  OR2_X1 U10511 ( .A1(n9620), .A2(n9119), .ZN(n9207) );
  INV_X1 U10512 ( .A(n9431), .ZN(n9117) );
  INV_X1 U10513 ( .A(n9542), .ZN(n9112) );
  INV_X1 U10514 ( .A(n9090), .ZN(n9587) );
  NOR3_X1 U10515 ( .A1(n9092), .A2(n5692), .A3(n7089), .ZN(n9096) );
  NAND4_X1 U10516 ( .A1(n9096), .A2(n9095), .A3(n9094), .A4(n9093), .ZN(n9100)
         );
  NAND2_X1 U10517 ( .A1(n9098), .A2(n9097), .ZN(n9099) );
  OR3_X1 U10518 ( .A1(n9101), .A2(n9100), .A3(n9099), .ZN(n9102) );
  NOR2_X1 U10519 ( .A1(n9159), .A2(n9102), .ZN(n9103) );
  NAND4_X1 U10520 ( .A1(n9104), .A2(n4781), .A3(n4778), .A4(n9103), .ZN(n9105)
         );
  NOR2_X1 U10521 ( .A1(n9106), .A2(n9105), .ZN(n9107) );
  NAND4_X1 U10522 ( .A1(n9109), .A2(n9587), .A3(n9108), .A4(n9107), .ZN(n9110)
         );
  NOR2_X1 U10523 ( .A1(n9110), .A2(n9568), .ZN(n9111) );
  NAND3_X1 U10524 ( .A1(n9523), .A2(n9112), .A3(n9111), .ZN(n9113) );
  NOR2_X1 U10525 ( .A1(n9508), .A2(n9113), .ZN(n9114) );
  NAND4_X1 U10526 ( .A1(n9466), .A2(n9478), .A3(n9114), .A4(n4711), .ZN(n9115)
         );
  NOR2_X1 U10527 ( .A1(n9445), .A2(n9115), .ZN(n9116) );
  NAND3_X1 U10528 ( .A1(n9413), .A2(n9117), .A3(n9116), .ZN(n9118) );
  NAND2_X1 U10529 ( .A1(n9620), .A2(n9119), .ZN(n9187) );
  AND4_X1 U10530 ( .A1(n9120), .A2(n9207), .A3(n4389), .A4(n9187), .ZN(n9121)
         );
  INV_X1 U10531 ( .A(n9189), .ZN(n9211) );
  NAND3_X1 U10532 ( .A1(n9190), .A2(n9121), .A3(n9211), .ZN(n9215) );
  NOR2_X1 U10533 ( .A1(n9215), .A2(n4340), .ZN(n9122) );
  AOI211_X1 U10534 ( .C1(n9125), .C2(n9124), .A(n9123), .B(n9122), .ZN(n9221)
         );
  NAND2_X1 U10535 ( .A1(n9126), .A2(n9347), .ZN(n9193) );
  INV_X1 U10536 ( .A(n9127), .ZN(n9128) );
  NOR2_X1 U10537 ( .A1(n9377), .A2(n9128), .ZN(n9199) );
  INV_X1 U10538 ( .A(n9134), .ZN(n9129) );
  AOI211_X1 U10539 ( .C1(n9132), .C2(n9131), .A(n9130), .B(n9129), .ZN(n9140)
         );
  INV_X1 U10540 ( .A(n9133), .ZN(n9135) );
  OAI21_X1 U10541 ( .B1(n9136), .B2(n9135), .A(n9134), .ZN(n9138) );
  NAND2_X1 U10542 ( .A1(n9138), .A2(n9137), .ZN(n9179) );
  OAI21_X1 U10543 ( .B1(n9140), .B2(n9179), .A(n9139), .ZN(n9142) );
  AOI21_X1 U10544 ( .B1(n9199), .B2(n9142), .A(n9141), .ZN(n9200) );
  INV_X1 U10545 ( .A(n9143), .ZN(n9169) );
  INV_X1 U10546 ( .A(n9144), .ZN(n9147) );
  NAND2_X1 U10547 ( .A1(n9255), .A2(n9145), .ZN(n9146) );
  AND4_X1 U10548 ( .A1(n9148), .A2(n9147), .A3(n5692), .A4(n9146), .ZN(n9151)
         );
  OAI211_X1 U10549 ( .C1(n4609), .C2(n9151), .A(n9150), .B(n9149), .ZN(n9154)
         );
  INV_X1 U10550 ( .A(n9152), .ZN(n9153) );
  NAND2_X1 U10551 ( .A1(n9154), .A2(n9153), .ZN(n9156) );
  AOI21_X1 U10552 ( .B1(n9156), .B2(n9155), .A(n4621), .ZN(n9158) );
  OAI21_X1 U10553 ( .B1(n9159), .B2(n9158), .A(n9157), .ZN(n9160) );
  NOR2_X1 U10554 ( .A1(n9161), .A2(n9160), .ZN(n9164) );
  OAI211_X1 U10555 ( .C1(n9165), .C2(n9164), .A(n9163), .B(n9162), .ZN(n9168)
         );
  AOI211_X1 U10556 ( .C1(n9169), .C2(n9168), .A(n9167), .B(n4694), .ZN(n9171)
         );
  OR2_X1 U10557 ( .A1(n9171), .A2(n9170), .ZN(n9173) );
  AOI21_X1 U10558 ( .B1(n9557), .B2(n9173), .A(n9172), .ZN(n9177) );
  OAI211_X1 U10559 ( .C1(n9177), .C2(n9176), .A(n9175), .B(n9174), .ZN(n9180)
         );
  OR2_X1 U10560 ( .A1(n9179), .A2(n9178), .ZN(n9196) );
  AOI21_X1 U10561 ( .B1(n9181), .B2(n9180), .A(n9196), .ZN(n9182) );
  OAI21_X1 U10562 ( .B1(n9197), .B2(n9182), .A(n9199), .ZN(n9185) );
  NAND2_X1 U10563 ( .A1(n9184), .A2(n9183), .ZN(n9195) );
  AOI21_X1 U10564 ( .B1(n9200), .B2(n9185), .A(n9195), .ZN(n9188) );
  NAND2_X1 U10565 ( .A1(n9187), .A2(n9186), .ZN(n9206) );
  OAI21_X1 U10566 ( .B1(n9188), .B2(n9206), .A(n9207), .ZN(n9191) );
  AOI21_X1 U10567 ( .B1(n9191), .B2(n9190), .A(n9189), .ZN(n9192) );
  MUX2_X1 U10568 ( .A(n9194), .B(n9193), .S(n9192), .Z(n9220) );
  INV_X1 U10569 ( .A(n9195), .ZN(n9205) );
  INV_X1 U10570 ( .A(n9196), .ZN(n9198) );
  AOI21_X1 U10571 ( .B1(n9198), .B2(n9503), .A(n9197), .ZN(n9202) );
  INV_X1 U10572 ( .A(n9199), .ZN(n9201) );
  OAI21_X1 U10573 ( .B1(n9202), .B2(n9201), .A(n9200), .ZN(n9204) );
  AOI22_X1 U10574 ( .A1(n9205), .A2(n9204), .B1(n9203), .B2(n9620), .ZN(n9210)
         );
  INV_X1 U10575 ( .A(n9206), .ZN(n9209) );
  INV_X1 U10576 ( .A(n9207), .ZN(n9208) );
  AOI22_X1 U10577 ( .A1(n9210), .A2(n9209), .B1(n9208), .B2(n9355), .ZN(n9214)
         );
  OAI211_X1 U10578 ( .C1(n9214), .C2(n9213), .A(n9212), .B(n9211), .ZN(n9218)
         );
  NAND4_X1 U10579 ( .A1(n9218), .A2(n9217), .A3(n4315), .A4(n9215), .ZN(n9219)
         );
  NAND4_X1 U10580 ( .A1(n9222), .A2(n9221), .A3(n9220), .A4(n9219), .ZN(n9229)
         );
  NAND2_X1 U10581 ( .A1(n9752), .A2(n9223), .ZN(n9227) );
  INV_X1 U10582 ( .A(n9224), .ZN(n9225) );
  OAI211_X1 U10583 ( .C1(n9227), .C2(n9226), .A(P1_B_REG_SCAN_IN), .B(n9225), 
        .ZN(n9228) );
  OAI211_X1 U10584 ( .C1(n9231), .C2(n9230), .A(n9229), .B(n9228), .ZN(
        P1_U3242) );
  MUX2_X1 U10585 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n4627), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10586 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9232), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10587 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9233), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10588 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9234), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10589 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9449), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10590 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9235), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10591 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9448), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10592 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9236), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10593 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9237), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10594 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9525), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10595 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9238), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10596 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9565), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10597 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9239), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10598 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9562), .S(P1_U3973), .Z(
        P1_U3570) );
  INV_X1 U10599 ( .A(P1_U3973), .ZN(n9254) );
  MUX2_X1 U10600 ( .A(n9240), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9254), .Z(
        P1_U3569) );
  MUX2_X1 U10601 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9241), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10602 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9242), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10603 ( .A(n9243), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9254), .Z(
        P1_U3566) );
  MUX2_X1 U10604 ( .A(n9244), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9254), .Z(
        P1_U3565) );
  MUX2_X1 U10605 ( .A(n9245), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9254), .Z(
        P1_U3564) );
  MUX2_X1 U10606 ( .A(n9246), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9254), .Z(
        P1_U3563) );
  MUX2_X1 U10607 ( .A(n9247), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9254), .Z(
        P1_U3562) );
  MUX2_X1 U10608 ( .A(n9248), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9254), .Z(
        P1_U3561) );
  MUX2_X1 U10609 ( .A(n9249), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9254), .Z(
        P1_U3560) );
  MUX2_X1 U10610 ( .A(n9250), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9254), .Z(
        P1_U3559) );
  MUX2_X1 U10611 ( .A(n9251), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9254), .Z(
        P1_U3558) );
  MUX2_X1 U10612 ( .A(n9252), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9254), .Z(
        P1_U3557) );
  MUX2_X1 U10613 ( .A(n9253), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9254), .Z(
        P1_U3556) );
  MUX2_X1 U10614 ( .A(n9255), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9254), .Z(
        P1_U3555) );
  MUX2_X1 U10615 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9256), .S(P1_U3973), .Z(
        P1_U3554) );
  NAND2_X1 U10616 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9259) );
  AOI211_X1 U10617 ( .C1(n9259), .C2(n9258), .A(n9257), .B(n9895), .ZN(n9260)
         );
  INV_X1 U10618 ( .A(n9260), .ZN(n9268) );
  AOI22_X1 U10619 ( .A1(n9866), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9267) );
  NAND2_X1 U10620 ( .A1(n9901), .A2(n9261), .ZN(n9266) );
  OAI211_X1 U10621 ( .C1(n9264), .C2(n9263), .A(n9883), .B(n9262), .ZN(n9265)
         );
  NAND4_X1 U10622 ( .A1(n9268), .A2(n9267), .A3(n9266), .A4(n9265), .ZN(
        P1_U3244) );
  MUX2_X1 U10623 ( .A(n9270), .B(n9269), .S(n9763), .Z(n9274) );
  NAND2_X1 U10624 ( .A1(n9272), .A2(n9271), .ZN(n9273) );
  OAI211_X1 U10625 ( .C1(n9274), .C2(n5716), .A(P1_U3973), .B(n9273), .ZN(
        n9303) );
  INV_X1 U10626 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9276) );
  OAI22_X1 U10627 ( .A1(n9904), .A2(n9276), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9275), .ZN(n9277) );
  AOI21_X1 U10628 ( .B1(n9278), .B2(n9901), .A(n9277), .ZN(n9288) );
  OAI211_X1 U10629 ( .C1(n9281), .C2(n9280), .A(n9883), .B(n9279), .ZN(n9287)
         );
  AOI211_X1 U10630 ( .C1(n9284), .C2(n9283), .A(n9282), .B(n9895), .ZN(n9285)
         );
  INV_X1 U10631 ( .A(n9285), .ZN(n9286) );
  NAND4_X1 U10632 ( .A1(n9303), .A2(n9288), .A3(n9287), .A4(n9286), .ZN(
        P1_U3245) );
  INV_X1 U10633 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9290) );
  OAI21_X1 U10634 ( .B1(n9904), .B2(n9290), .A(n9289), .ZN(n9291) );
  AOI21_X1 U10635 ( .B1(n9901), .B2(n9292), .A(n9291), .ZN(n9302) );
  AOI211_X1 U10636 ( .C1(n9295), .C2(n9294), .A(n9895), .B(n9293), .ZN(n9296)
         );
  INV_X1 U10637 ( .A(n9296), .ZN(n9301) );
  OAI211_X1 U10638 ( .C1(n9299), .C2(n9298), .A(n9883), .B(n9297), .ZN(n9300)
         );
  NAND4_X1 U10639 ( .A1(n9303), .A2(n9302), .A3(n9301), .A4(n9300), .ZN(
        P1_U3247) );
  AOI211_X1 U10640 ( .C1(n9306), .C2(n9305), .A(n9895), .B(n9304), .ZN(n9307)
         );
  INV_X1 U10641 ( .A(n9307), .ZN(n9317) );
  INV_X1 U10642 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9309) );
  NAND2_X1 U10643 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9308) );
  OAI21_X1 U10644 ( .B1(n9904), .B2(n9309), .A(n9308), .ZN(n9310) );
  AOI21_X1 U10645 ( .B1(n9311), .B2(n9901), .A(n9310), .ZN(n9316) );
  OAI211_X1 U10646 ( .C1(n9314), .C2(n9313), .A(n9883), .B(n9312), .ZN(n9315)
         );
  NAND3_X1 U10647 ( .A1(n9317), .A2(n9316), .A3(n9315), .ZN(P1_U3248) );
  INV_X1 U10648 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9351) );
  OR2_X1 U10649 ( .A1(n9882), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9323) );
  XNOR2_X1 U10650 ( .A(n9882), .B(n9683), .ZN(n9878) );
  AOI22_X1 U10651 ( .A1(n9870), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9318), .B2(
        n9337), .ZN(n9869) );
  NAND2_X1 U10652 ( .A1(n9843), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9320) );
  XNOR2_X1 U10653 ( .A(n9831), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9824) );
  OAI21_X1 U10654 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n9331), .A(n9319), .ZN(
        n9825) );
  NOR2_X1 U10655 ( .A1(n9824), .A2(n9825), .ZN(n9823) );
  XNOR2_X1 U10656 ( .A(n9843), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9839) );
  NAND2_X1 U10657 ( .A1(n9320), .A2(n9842), .ZN(n9321) );
  NAND2_X1 U10658 ( .A1(n9869), .A2(n9868), .ZN(n9867) );
  NAND2_X1 U10659 ( .A1(n9878), .A2(n9879), .ZN(n9877) );
  NAND2_X1 U10660 ( .A1(n9323), .A2(n9877), .ZN(n9897) );
  INV_X1 U10661 ( .A(n9897), .ZN(n9325) );
  NAND2_X1 U10662 ( .A1(n9900), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9326) );
  OAI21_X1 U10663 ( .B1(n9900), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9326), .ZN(
        n9896) );
  INV_X1 U10664 ( .A(n9896), .ZN(n9324) );
  NAND2_X1 U10665 ( .A1(n9325), .A2(n9324), .ZN(n9893) );
  NAND2_X1 U10666 ( .A1(n9893), .A2(n9326), .ZN(n9327) );
  INV_X1 U10667 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9673) );
  XNOR2_X1 U10668 ( .A(n9327), .B(n9673), .ZN(n9342) );
  NAND2_X1 U10669 ( .A1(n9900), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9339) );
  OAI21_X1 U10670 ( .B1(n9900), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9339), .ZN(
        n9891) );
  NOR2_X1 U10671 ( .A1(n9882), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9328) );
  AOI21_X1 U10672 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n9882), .A(n9328), .ZN(
        n9875) );
  NAND2_X1 U10673 ( .A1(n9831), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9329) );
  OAI21_X1 U10674 ( .B1(n9831), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9329), .ZN(
        n9827) );
  OAI21_X1 U10675 ( .B1(n9331), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9330), .ZN(
        n9828) );
  NOR2_X1 U10676 ( .A1(n9827), .A2(n9828), .ZN(n9826) );
  AOI22_X1 U10677 ( .A1(n9843), .A2(n5323), .B1(P1_REG2_REG_14__SCAN_IN), .B2(
        n9332), .ZN(n9836) );
  NOR2_X1 U10678 ( .A1(n9837), .A2(n9836), .ZN(n9835) );
  INV_X1 U10679 ( .A(n9857), .ZN(n9333) );
  NOR2_X1 U10680 ( .A1(n9334), .A2(n9333), .ZN(n9336) );
  AOI21_X1 U10681 ( .B1(n9334), .B2(n9333), .A(n9336), .ZN(n9335) );
  INV_X1 U10682 ( .A(n9335), .ZN(n9854) );
  NOR2_X1 U10683 ( .A1(n9336), .A2(n9853), .ZN(n9863) );
  AOI22_X1 U10684 ( .A1(n9870), .A2(n9338), .B1(P1_REG2_REG_16__SCAN_IN), .B2(
        n9337), .ZN(n9862) );
  AOI21_X1 U10685 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9870), .A(n9861), .ZN(
        n9876) );
  XNOR2_X1 U10686 ( .A(n9341), .B(n9340), .ZN(n9344) );
  AOI22_X1 U10687 ( .A1(n9342), .A2(n9880), .B1(n9883), .B2(n9344), .ZN(n9348)
         );
  INV_X1 U10688 ( .A(n9342), .ZN(n9346) );
  OAI21_X1 U10689 ( .B1(n9889), .B2(n9344), .A(n9343), .ZN(n9345) );
  NAND2_X1 U10690 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9349) );
  OAI211_X1 U10691 ( .C1(n9904), .C2(n9351), .A(n9350), .B(n9349), .ZN(
        P1_U3262) );
  NAND2_X1 U10692 ( .A1(n9617), .A2(n9905), .ZN(n9357) );
  INV_X1 U10693 ( .A(n9353), .ZN(n9354) );
  AND2_X1 U10694 ( .A1(n9355), .A2(n9354), .ZN(n9616) );
  INV_X1 U10695 ( .A(n9616), .ZN(n9621) );
  NOR2_X1 U10696 ( .A1(n9934), .A2(n9621), .ZN(n9362) );
  AOI21_X1 U10697 ( .B1(n9910), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9362), .ZN(
        n9356) );
  OAI211_X1 U10698 ( .C1(n9706), .C2(n9913), .A(n9357), .B(n9356), .ZN(
        P1_U3263) );
  NAND2_X1 U10699 ( .A1(n9620), .A2(n9358), .ZN(n9359) );
  NAND2_X1 U10700 ( .A1(n9359), .A2(n9698), .ZN(n9360) );
  NOR2_X1 U10701 ( .A1(n9922), .A2(n9361), .ZN(n9363) );
  AOI211_X1 U10702 ( .C1(n9620), .C2(n9925), .A(n9363), .B(n9362), .ZN(n9364)
         );
  OAI21_X1 U10703 ( .B1(n9622), .B2(n9928), .A(n9364), .ZN(P1_U3264) );
  OR2_X1 U10704 ( .A1(n9920), .A2(n9365), .ZN(n9367) );
  OAI22_X1 U10705 ( .A1(n9368), .A2(n9367), .B1(n9366), .B2(n9922), .ZN(n9369)
         );
  AOI21_X1 U10706 ( .B1(n9370), .B2(n9925), .A(n9369), .ZN(n9371) );
  OAI21_X1 U10707 ( .B1(n9372), .B2(n9928), .A(n9371), .ZN(n9373) );
  AOI21_X1 U10708 ( .B1(n9374), .B2(n9931), .A(n9373), .ZN(n9375) );
  OAI21_X1 U10709 ( .B1(n9376), .B2(n9910), .A(n9375), .ZN(P1_U3356) );
  INV_X1 U10710 ( .A(n9378), .ZN(n9379) );
  INV_X1 U10711 ( .A(n9627), .ZN(n9391) );
  AOI21_X1 U10712 ( .B1(n9387), .B2(n9401), .A(n9548), .ZN(n9385) );
  NAND2_X1 U10713 ( .A1(n9385), .A2(n9384), .ZN(n9625) );
  AOI22_X1 U10714 ( .A1(n9386), .A2(n9908), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9934), .ZN(n9389) );
  NAND2_X1 U10715 ( .A1(n9387), .A2(n9925), .ZN(n9388) );
  OAI211_X1 U10716 ( .C1(n9625), .C2(n9928), .A(n9389), .B(n9388), .ZN(n9390)
         );
  AOI21_X1 U10717 ( .B1(n9391), .B2(n9931), .A(n9390), .ZN(n9392) );
  OAI21_X1 U10718 ( .B1(n9626), .B2(n9910), .A(n9392), .ZN(P1_U3265) );
  OAI21_X1 U10719 ( .B1(n9394), .B2(n9393), .A(n9592), .ZN(n9396) );
  NAND2_X1 U10720 ( .A1(n9398), .A2(n9397), .ZN(n9628) );
  INV_X1 U10721 ( .A(n9628), .ZN(n9408) );
  XNOR2_X1 U10722 ( .A(n9400), .B(n9399), .ZN(n9630) );
  NAND2_X1 U10723 ( .A1(n9630), .A2(n9931), .ZN(n9407) );
  AOI211_X1 U10724 ( .C1(n9402), .C2(n9415), .A(n9548), .B(n9383), .ZN(n9629)
         );
  AOI22_X1 U10725 ( .A1(n9403), .A2(n9908), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9910), .ZN(n9404) );
  OAI21_X1 U10726 ( .B1(n9715), .B2(n9913), .A(n9404), .ZN(n9405) );
  AOI21_X1 U10727 ( .B1(n9629), .B2(n9905), .A(n9405), .ZN(n9406) );
  OAI211_X1 U10728 ( .C1(n9408), .C2(n9934), .A(n9407), .B(n9406), .ZN(
        P1_U3266) );
  XNOR2_X1 U10729 ( .A(n9409), .B(n9413), .ZN(n9410) );
  NAND2_X1 U10730 ( .A1(n9410), .A2(n9592), .ZN(n9412) );
  NAND2_X1 U10731 ( .A1(n9412), .A2(n9411), .ZN(n9633) );
  INV_X1 U10732 ( .A(n9633), .ZN(n9423) );
  XNOR2_X1 U10733 ( .A(n9414), .B(n9413), .ZN(n9635) );
  NAND2_X1 U10734 ( .A1(n9635), .A2(n9931), .ZN(n9422) );
  INV_X1 U10735 ( .A(n9415), .ZN(n9416) );
  AOI211_X1 U10736 ( .C1(n9417), .C2(n9433), .A(n9548), .B(n9416), .ZN(n9634)
         );
  AOI22_X1 U10737 ( .A1(n9418), .A2(n9908), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9910), .ZN(n9419) );
  OAI21_X1 U10738 ( .B1(n9719), .B2(n9913), .A(n9419), .ZN(n9420) );
  AOI21_X1 U10739 ( .B1(n9634), .B2(n9905), .A(n9420), .ZN(n9421) );
  OAI211_X1 U10740 ( .C1(n9910), .C2(n9423), .A(n9422), .B(n9421), .ZN(
        P1_U3267) );
  NAND2_X1 U10741 ( .A1(n9446), .A2(n9424), .ZN(n9425) );
  NAND2_X1 U10742 ( .A1(n9425), .A2(n9431), .ZN(n9427) );
  NAND2_X1 U10743 ( .A1(n9427), .A2(n9426), .ZN(n9428) );
  NAND2_X1 U10744 ( .A1(n9428), .A2(n9592), .ZN(n9430) );
  NAND2_X1 U10745 ( .A1(n9430), .A2(n9429), .ZN(n9638) );
  INV_X1 U10746 ( .A(n9638), .ZN(n9442) );
  XNOR2_X1 U10747 ( .A(n9432), .B(n9431), .ZN(n9640) );
  NAND2_X1 U10748 ( .A1(n9640), .A2(n9931), .ZN(n9441) );
  INV_X1 U10749 ( .A(n9452), .ZN(n9435) );
  INV_X1 U10750 ( .A(n9433), .ZN(n9434) );
  AOI211_X1 U10751 ( .C1(n9436), .C2(n9435), .A(n9548), .B(n9434), .ZN(n9639)
         );
  AOI22_X1 U10752 ( .A1(n9437), .A2(n9908), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9910), .ZN(n9438) );
  OAI21_X1 U10753 ( .B1(n9723), .B2(n9913), .A(n9438), .ZN(n9439) );
  AOI21_X1 U10754 ( .B1(n9639), .B2(n9905), .A(n9439), .ZN(n9440) );
  OAI211_X1 U10755 ( .C1(n9910), .C2(n9442), .A(n9441), .B(n9440), .ZN(
        P1_U3268) );
  XNOR2_X1 U10756 ( .A(n9443), .B(n9445), .ZN(n9647) );
  INV_X1 U10757 ( .A(n9444), .ZN(n9447) );
  OAI211_X1 U10758 ( .C1(n9447), .C2(n4602), .A(n9446), .B(n9592), .ZN(n9451)
         );
  AOI22_X1 U10759 ( .A1(n9449), .A2(n4309), .B1(n9563), .B2(n9448), .ZN(n9450)
         );
  NAND2_X1 U10760 ( .A1(n9451), .A2(n9450), .ZN(n9643) );
  AOI211_X1 U10761 ( .C1(n9645), .C2(n9460), .A(n9548), .B(n9452), .ZN(n9644)
         );
  NAND2_X1 U10762 ( .A1(n9644), .A2(n9905), .ZN(n9455) );
  AOI22_X1 U10763 ( .A1(n9453), .A2(n9908), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9934), .ZN(n9454) );
  OAI211_X1 U10764 ( .C1(n9456), .C2(n9913), .A(n9455), .B(n9454), .ZN(n9457)
         );
  AOI21_X1 U10765 ( .B1(n9922), .B2(n9643), .A(n9457), .ZN(n9458) );
  OAI21_X1 U10766 ( .B1(n9647), .B2(n9556), .A(n9458), .ZN(P1_U3269) );
  XOR2_X1 U10767 ( .A(n9466), .B(n9459), .Z(n9648) );
  INV_X1 U10768 ( .A(n9460), .ZN(n9461) );
  AOI211_X1 U10769 ( .C1(n9462), .C2(n9481), .A(n9548), .B(n9461), .ZN(n9650)
         );
  OAI22_X1 U10770 ( .A1(n4480), .A2(n9913), .B1(n9463), .B2(n9922), .ZN(n9471)
         );
  INV_X1 U10771 ( .A(n9464), .ZN(n9468) );
  XOR2_X1 U10772 ( .A(n9465), .B(n9466), .Z(n9467) );
  NOR2_X1 U10773 ( .A1(n9467), .A2(n9544), .ZN(n9651) );
  AOI211_X1 U10774 ( .C1(n9908), .C2(n9468), .A(n9649), .B(n9651), .ZN(n9469)
         );
  NOR2_X1 U10775 ( .A1(n9469), .A2(n9910), .ZN(n9470) );
  AOI211_X1 U10776 ( .C1(n9650), .C2(n9905), .A(n9471), .B(n9470), .ZN(n9472)
         );
  OAI21_X1 U10777 ( .B1(n9648), .B2(n9556), .A(n9472), .ZN(P1_U3270) );
  XNOR2_X1 U10778 ( .A(n9473), .B(n9478), .ZN(n9475) );
  AOI21_X1 U10779 ( .B1(n9475), .B2(n9592), .A(n9474), .ZN(n9656) );
  INV_X1 U10780 ( .A(n9476), .ZN(n9477) );
  XOR2_X1 U10781 ( .A(n9478), .B(n9477), .Z(n9657) );
  OR2_X1 U10782 ( .A1(n9657), .A2(n9556), .ZN(n9486) );
  OAI22_X1 U10783 ( .A1(n9480), .A2(n9922), .B1(n9479), .B2(n9920), .ZN(n9483)
         );
  OAI211_X1 U10784 ( .C1(n9731), .C2(n4401), .A(n9698), .B(n9481), .ZN(n9655)
         );
  NOR2_X1 U10785 ( .A1(n9655), .A2(n9928), .ZN(n9482) );
  AOI211_X1 U10786 ( .C1(n9925), .C2(n9484), .A(n9483), .B(n9482), .ZN(n9485)
         );
  OAI211_X1 U10787 ( .C1(n9910), .C2(n9656), .A(n9486), .B(n9485), .ZN(
        P1_U3271) );
  XNOR2_X1 U10788 ( .A(n9487), .B(n4711), .ZN(n9662) );
  INV_X1 U10789 ( .A(n9662), .ZN(n9501) );
  NAND2_X1 U10790 ( .A1(n9489), .A2(n9488), .ZN(n9490) );
  NAND2_X1 U10791 ( .A1(n9491), .A2(n9490), .ZN(n9492) );
  NAND2_X1 U10792 ( .A1(n9492), .A2(n9592), .ZN(n9494) );
  NAND2_X1 U10793 ( .A1(n9494), .A2(n9493), .ZN(n9660) );
  NAND2_X1 U10794 ( .A1(n9661), .A2(n9905), .ZN(n9498) );
  AOI22_X1 U10795 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(n9934), .B1(n9496), .B2(
        n9908), .ZN(n9497) );
  OAI211_X1 U10796 ( .C1(n4536), .C2(n9913), .A(n9498), .B(n9497), .ZN(n9499)
         );
  AOI21_X1 U10797 ( .B1(n9922), .B2(n9660), .A(n9499), .ZN(n9500) );
  OAI21_X1 U10798 ( .B1(n9501), .B2(n9556), .A(n9500), .ZN(P1_U3272) );
  INV_X1 U10799 ( .A(n9508), .ZN(n9502) );
  XNOR2_X1 U10800 ( .A(n9503), .B(n9502), .ZN(n9504) );
  NAND2_X1 U10801 ( .A1(n9504), .A2(n9592), .ZN(n9507) );
  INV_X1 U10802 ( .A(n9505), .ZN(n9506) );
  NAND2_X1 U10803 ( .A1(n9507), .A2(n9506), .ZN(n9665) );
  INV_X1 U10804 ( .A(n9665), .ZN(n9519) );
  XOR2_X1 U10805 ( .A(n9509), .B(n9508), .Z(n9667) );
  NAND2_X1 U10806 ( .A1(n9667), .A2(n9931), .ZN(n9518) );
  INV_X1 U10807 ( .A(n9510), .ZN(n9511) );
  AOI211_X1 U10808 ( .C1(n9512), .C2(n9529), .A(n9548), .B(n9511), .ZN(n9666)
         );
  NOR2_X1 U10809 ( .A1(n9738), .A2(n9913), .ZN(n9516) );
  OAI22_X1 U10810 ( .A1(n9922), .A2(n9514), .B1(n9513), .B2(n9920), .ZN(n9515)
         );
  AOI211_X1 U10811 ( .C1(n9666), .C2(n9905), .A(n9516), .B(n9515), .ZN(n9517)
         );
  OAI211_X1 U10812 ( .C1(n9910), .C2(n9519), .A(n9518), .B(n9517), .ZN(
        P1_U3273) );
  XOR2_X1 U10813 ( .A(n9520), .B(n9523), .Z(n9672) );
  INV_X1 U10814 ( .A(n9672), .ZN(n9537) );
  OAI21_X1 U10815 ( .B1(n9523), .B2(n9522), .A(n9521), .ZN(n9524) );
  NAND2_X1 U10816 ( .A1(n9524), .A2(n9592), .ZN(n9527) );
  AOI22_X1 U10817 ( .A1(n9525), .A2(n4309), .B1(n9563), .B2(n9565), .ZN(n9526)
         );
  NAND2_X1 U10818 ( .A1(n9527), .A2(n9526), .ZN(n9670) );
  INV_X1 U10819 ( .A(n9528), .ZN(n9547) );
  INV_X1 U10820 ( .A(n9529), .ZN(n9530) );
  AOI211_X1 U10821 ( .C1(n9531), .C2(n9547), .A(n9548), .B(n9530), .ZN(n9671)
         );
  NAND2_X1 U10822 ( .A1(n9671), .A2(n9905), .ZN(n9534) );
  AOI22_X1 U10823 ( .A1(n9934), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9532), .B2(
        n9908), .ZN(n9533) );
  OAI211_X1 U10824 ( .C1(n9742), .C2(n9913), .A(n9534), .B(n9533), .ZN(n9535)
         );
  AOI21_X1 U10825 ( .B1(n9922), .B2(n9670), .A(n9535), .ZN(n9536) );
  OAI21_X1 U10826 ( .B1(n9537), .B2(n9556), .A(n9536), .ZN(P1_U3274) );
  XNOR2_X1 U10827 ( .A(n9538), .B(n9542), .ZN(n9679) );
  INV_X1 U10828 ( .A(n9539), .ZN(n9540) );
  AOI21_X1 U10829 ( .B1(n9542), .B2(n9541), .A(n9540), .ZN(n9543) );
  OAI222_X1 U10830 ( .A1(n4308), .A2(n9546), .B1(n9583), .B2(n9545), .C1(n9544), .C2(n9543), .ZN(n9675) );
  INV_X1 U10831 ( .A(n9677), .ZN(n9553) );
  AOI211_X1 U10832 ( .C1(n9677), .C2(n9571), .A(n9548), .B(n9528), .ZN(n9676)
         );
  NAND2_X1 U10833 ( .A1(n9676), .A2(n9905), .ZN(n9552) );
  INV_X1 U10834 ( .A(n9549), .ZN(n9550) );
  AOI22_X1 U10835 ( .A1(n9910), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9550), .B2(
        n9908), .ZN(n9551) );
  OAI211_X1 U10836 ( .C1(n9553), .C2(n9913), .A(n9552), .B(n9551), .ZN(n9554)
         );
  AOI21_X1 U10837 ( .B1(n9675), .B2(n9922), .A(n9554), .ZN(n9555) );
  OAI21_X1 U10838 ( .B1(n9679), .B2(n9556), .A(n9555), .ZN(P1_U3275) );
  NAND2_X1 U10839 ( .A1(n9558), .A2(n9557), .ZN(n9560) );
  INV_X1 U10840 ( .A(n9568), .ZN(n9559) );
  XNOR2_X1 U10841 ( .A(n9560), .B(n9559), .ZN(n9561) );
  NAND2_X1 U10842 ( .A1(n9561), .A2(n9592), .ZN(n9567) );
  AOI22_X1 U10843 ( .A1(n9565), .A2(n4309), .B1(n9563), .B2(n9562), .ZN(n9566)
         );
  NAND2_X1 U10844 ( .A1(n9567), .A2(n9566), .ZN(n9680) );
  INV_X1 U10845 ( .A(n9680), .ZN(n9581) );
  XNOR2_X1 U10846 ( .A(n9569), .B(n9568), .ZN(n9682) );
  NAND2_X1 U10847 ( .A1(n9682), .A2(n9931), .ZN(n9580) );
  INV_X1 U10848 ( .A(n9570), .ZN(n9573) );
  INV_X1 U10849 ( .A(n9571), .ZN(n9572) );
  AOI211_X1 U10850 ( .C1(n9574), .C2(n9573), .A(n9548), .B(n9572), .ZN(n9681)
         );
  NOR2_X1 U10851 ( .A1(n9748), .A2(n9913), .ZN(n9578) );
  INV_X1 U10852 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9576) );
  OAI22_X1 U10853 ( .A1(n9922), .A2(n9576), .B1(n9575), .B2(n9920), .ZN(n9577)
         );
  AOI211_X1 U10854 ( .C1(n9681), .C2(n9905), .A(n9578), .B(n9577), .ZN(n9579)
         );
  OAI211_X1 U10855 ( .C1(n9910), .C2(n9581), .A(n9580), .B(n9579), .ZN(
        P1_U3276) );
  XNOR2_X1 U10856 ( .A(n9582), .B(n9587), .ZN(n9593) );
  OAI22_X1 U10857 ( .A1(n9586), .A2(n4308), .B1(n9584), .B2(n9583), .ZN(n9591)
         );
  XNOR2_X1 U10858 ( .A(n9588), .B(n9587), .ZN(n9696) );
  NOR2_X1 U10859 ( .A1(n9696), .A2(n9589), .ZN(n9590) );
  AOI211_X1 U10860 ( .C1(n9593), .C2(n9592), .A(n9591), .B(n9590), .ZN(n9694)
         );
  AOI21_X1 U10861 ( .B1(n9691), .B2(n9595), .A(n9594), .ZN(n9692) );
  INV_X1 U10862 ( .A(n9596), .ZN(n9597) );
  AOI22_X1 U10863 ( .A1(n9934), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9597), .B2(
        n9908), .ZN(n9598) );
  OAI21_X1 U10864 ( .B1(n9599), .B2(n9913), .A(n9598), .ZN(n9602) );
  NOR2_X1 U10865 ( .A1(n9696), .A2(n9600), .ZN(n9601) );
  AOI211_X1 U10866 ( .C1(n9692), .C2(n9603), .A(n9602), .B(n9601), .ZN(n9604)
         );
  OAI21_X1 U10867 ( .B1(n9694), .B2(n9910), .A(n9604), .ZN(P1_U3279) );
  NAND2_X1 U10868 ( .A1(n9605), .A2(n9922), .ZN(n9615) );
  NAND2_X1 U10869 ( .A1(n9606), .A2(n9931), .ZN(n9614) );
  NAND2_X1 U10870 ( .A1(n9910), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9607) );
  OAI21_X1 U10871 ( .B1(n9920), .B2(n9608), .A(n9607), .ZN(n9609) );
  AOI21_X1 U10872 ( .B1(n9610), .B2(n9925), .A(n9609), .ZN(n9613) );
  NAND2_X1 U10873 ( .A1(n9611), .A2(n9905), .ZN(n9612) );
  NAND4_X1 U10874 ( .A1(n9615), .A2(n9614), .A3(n9613), .A4(n9612), .ZN(
        P1_U3284) );
  NOR2_X1 U10875 ( .A1(n9617), .A2(n9616), .ZN(n9703) );
  MUX2_X1 U10876 ( .A(n9618), .B(n9703), .S(n9959), .Z(n9619) );
  OAI21_X1 U10877 ( .B1(n9706), .B2(n9685), .A(n9619), .ZN(P1_U3553) );
  MUX2_X1 U10878 ( .A(n9623), .B(n9708), .S(n9959), .Z(n9624) );
  OAI21_X1 U10879 ( .B1(n4529), .B2(n9685), .A(n9624), .ZN(P1_U3552) );
  INV_X1 U10880 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9631) );
  AOI211_X1 U10881 ( .C1(n9630), .C2(n9944), .A(n9629), .B(n9628), .ZN(n9712)
         );
  MUX2_X1 U10882 ( .A(n9631), .B(n9712), .S(n9959), .Z(n9632) );
  OAI21_X1 U10883 ( .B1(n9715), .B2(n9685), .A(n9632), .ZN(P1_U3549) );
  INV_X1 U10884 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9636) );
  AOI211_X1 U10885 ( .C1(n9635), .C2(n9944), .A(n9634), .B(n9633), .ZN(n9716)
         );
  MUX2_X1 U10886 ( .A(n9636), .B(n9716), .S(n9959), .Z(n9637) );
  OAI21_X1 U10887 ( .B1(n9719), .B2(n9685), .A(n9637), .ZN(P1_U3548) );
  INV_X1 U10888 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9641) );
  AOI211_X1 U10889 ( .C1(n9640), .C2(n9944), .A(n9639), .B(n9638), .ZN(n9720)
         );
  MUX2_X1 U10890 ( .A(n9641), .B(n9720), .S(n9959), .Z(n9642) );
  OAI21_X1 U10891 ( .B1(n9723), .B2(n9685), .A(n9642), .ZN(P1_U3547) );
  AOI211_X1 U10892 ( .C1(n9949), .C2(n9645), .A(n9644), .B(n9643), .ZN(n9646)
         );
  OAI21_X1 U10893 ( .B1(n9647), .B2(n9953), .A(n9646), .ZN(n9724) );
  MUX2_X1 U10894 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9724), .S(n9959), .Z(
        P1_U3546) );
  INV_X1 U10895 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9653) );
  NOR2_X1 U10896 ( .A1(n9648), .A2(n9953), .ZN(n9652) );
  NOR4_X1 U10897 ( .A1(n9652), .A2(n9651), .A3(n9650), .A4(n9649), .ZN(n9725)
         );
  MUX2_X1 U10898 ( .A(n9653), .B(n9725), .S(n9959), .Z(n9654) );
  OAI21_X1 U10899 ( .B1(n4480), .B2(n9685), .A(n9654), .ZN(P1_U3545) );
  OAI211_X1 U10900 ( .C1(n9657), .C2(n9953), .A(n9656), .B(n9655), .ZN(n9728)
         );
  MUX2_X1 U10901 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9728), .S(n9959), .Z(n9658) );
  INV_X1 U10902 ( .A(n9658), .ZN(n9659) );
  OAI21_X1 U10903 ( .B1(n9731), .B2(n9685), .A(n9659), .ZN(P1_U3544) );
  INV_X1 U10904 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9663) );
  AOI211_X1 U10905 ( .C1(n9662), .C2(n9944), .A(n9661), .B(n9660), .ZN(n9732)
         );
  MUX2_X1 U10906 ( .A(n9663), .B(n9732), .S(n9959), .Z(n9664) );
  OAI21_X1 U10907 ( .B1(n4536), .B2(n9685), .A(n9664), .ZN(P1_U3543) );
  INV_X1 U10908 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9668) );
  AOI211_X1 U10909 ( .C1(n9667), .C2(n9944), .A(n9666), .B(n9665), .ZN(n9735)
         );
  MUX2_X1 U10910 ( .A(n9668), .B(n9735), .S(n9959), .Z(n9669) );
  OAI21_X1 U10911 ( .B1(n9738), .B2(n9685), .A(n9669), .ZN(P1_U3542) );
  AOI211_X1 U10912 ( .C1(n9672), .C2(n9944), .A(n9671), .B(n9670), .ZN(n9739)
         );
  MUX2_X1 U10913 ( .A(n9673), .B(n9739), .S(n9959), .Z(n9674) );
  OAI21_X1 U10914 ( .B1(n9742), .B2(n9685), .A(n9674), .ZN(P1_U3541) );
  AOI211_X1 U10915 ( .C1(n9949), .C2(n9677), .A(n9676), .B(n9675), .ZN(n9678)
         );
  OAI21_X1 U10916 ( .B1(n9679), .B2(n9953), .A(n9678), .ZN(n9743) );
  MUX2_X1 U10917 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9743), .S(n9959), .Z(
        P1_U3540) );
  AOI211_X1 U10918 ( .C1(n9682), .C2(n9944), .A(n9681), .B(n9680), .ZN(n9744)
         );
  MUX2_X1 U10919 ( .A(n9683), .B(n9744), .S(n9959), .Z(n9684) );
  OAI21_X1 U10920 ( .B1(n9748), .B2(n9685), .A(n9684), .ZN(P1_U3539) );
  AOI21_X1 U10921 ( .B1(n9949), .B2(n9687), .A(n9686), .ZN(n9688) );
  OAI211_X1 U10922 ( .C1(n9690), .C2(n9953), .A(n9689), .B(n9688), .ZN(n9749)
         );
  MUX2_X1 U10923 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9749), .S(n9959), .Z(
        P1_U3538) );
  AOI22_X1 U10924 ( .A1(n9692), .A2(n9698), .B1(n9949), .B2(n9691), .ZN(n9693)
         );
  OAI211_X1 U10925 ( .C1(n9696), .C2(n9695), .A(n9694), .B(n9693), .ZN(n9750)
         );
  MUX2_X1 U10926 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9750), .S(n9959), .Z(
        P1_U3536) );
  AOI22_X1 U10927 ( .A1(n9699), .A2(n9698), .B1(n9949), .B2(n9697), .ZN(n9700)
         );
  OAI211_X1 U10928 ( .C1(n9702), .C2(n9953), .A(n9701), .B(n9700), .ZN(n9751)
         );
  MUX2_X1 U10929 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9751), .S(n9959), .Z(
        P1_U3535) );
  INV_X1 U10930 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9704) );
  MUX2_X1 U10931 ( .A(n9704), .B(n9703), .S(n9946), .Z(n9705) );
  OAI21_X1 U10932 ( .B1(n9706), .B2(n9747), .A(n9705), .ZN(P1_U3521) );
  INV_X1 U10933 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9707) );
  MUX2_X1 U10934 ( .A(n9708), .B(n9707), .S(n9955), .Z(n9709) );
  OAI21_X1 U10935 ( .B1(n4529), .B2(n9747), .A(n9709), .ZN(P1_U3520) );
  OAI21_X1 U10936 ( .B1(n9711), .B2(n9747), .A(n4311), .ZN(P1_U3518) );
  INV_X1 U10937 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9713) );
  MUX2_X1 U10938 ( .A(n9713), .B(n9712), .S(n9946), .Z(n9714) );
  OAI21_X1 U10939 ( .B1(n9715), .B2(n9747), .A(n9714), .ZN(P1_U3517) );
  INV_X1 U10940 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9717) );
  MUX2_X1 U10941 ( .A(n9717), .B(n9716), .S(n9946), .Z(n9718) );
  OAI21_X1 U10942 ( .B1(n9719), .B2(n9747), .A(n9718), .ZN(P1_U3516) );
  INV_X1 U10943 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9721) );
  MUX2_X1 U10944 ( .A(n9721), .B(n9720), .S(n9946), .Z(n9722) );
  OAI21_X1 U10945 ( .B1(n9723), .B2(n9747), .A(n9722), .ZN(P1_U3515) );
  MUX2_X1 U10946 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9724), .S(n9946), .Z(
        P1_U3514) );
  INV_X1 U10947 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9726) );
  MUX2_X1 U10948 ( .A(n9726), .B(n9725), .S(n9946), .Z(n9727) );
  OAI21_X1 U10949 ( .B1(n4480), .B2(n9747), .A(n9727), .ZN(P1_U3513) );
  MUX2_X1 U10950 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9728), .S(n9946), .Z(n9729) );
  INV_X1 U10951 ( .A(n9729), .ZN(n9730) );
  OAI21_X1 U10952 ( .B1(n9731), .B2(n9747), .A(n9730), .ZN(P1_U3512) );
  INV_X1 U10953 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9733) );
  MUX2_X1 U10954 ( .A(n9733), .B(n9732), .S(n9946), .Z(n9734) );
  OAI21_X1 U10955 ( .B1(n4536), .B2(n9747), .A(n9734), .ZN(P1_U3511) );
  INV_X1 U10956 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9736) );
  MUX2_X1 U10957 ( .A(n9736), .B(n9735), .S(n9946), .Z(n9737) );
  OAI21_X1 U10958 ( .B1(n9738), .B2(n9747), .A(n9737), .ZN(P1_U3510) );
  INV_X1 U10959 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9740) );
  MUX2_X1 U10960 ( .A(n9740), .B(n9739), .S(n9946), .Z(n9741) );
  OAI21_X1 U10961 ( .B1(n9742), .B2(n9747), .A(n9741), .ZN(P1_U3509) );
  MUX2_X1 U10962 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9743), .S(n9946), .Z(
        P1_U3507) );
  MUX2_X1 U10963 ( .A(n9745), .B(n9744), .S(n9946), .Z(n9746) );
  OAI21_X1 U10964 ( .B1(n9748), .B2(n9747), .A(n9746), .ZN(P1_U3504) );
  MUX2_X1 U10965 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9749), .S(n9946), .Z(
        P1_U3501) );
  MUX2_X1 U10966 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9750), .S(n9946), .Z(
        P1_U3495) );
  MUX2_X1 U10967 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9751), .S(n9946), .Z(
        P1_U3492) );
  AND2_X1 U10968 ( .A1(n9753), .A2(n9752), .ZN(n9936) );
  MUX2_X1 U10969 ( .A(P1_D_REG_1__SCAN_IN), .B(n9754), .S(n9936), .Z(P1_U3440)
         );
  MUX2_X1 U10970 ( .A(P1_D_REG_0__SCAN_IN), .B(n9755), .S(n9936), .Z(P1_U3439)
         );
  NOR4_X1 U10971 ( .A1(n9757), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9756), .A4(
        P1_U3086), .ZN(n9758) );
  AOI21_X1 U10972 ( .B1(n9759), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9758), .ZN(
        n9760) );
  OAI21_X1 U10973 ( .B1(n9761), .B2(n9769), .A(n9760), .ZN(P1_U3324) );
  INV_X1 U10974 ( .A(n9762), .ZN(n9764) );
  OAI222_X1 U10975 ( .A1(n9766), .A2(n9765), .B1(n9769), .B2(n9764), .C1(n9763), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U10976 ( .A1(n9770), .A2(P1_U3086), .B1(n9769), .B2(n9768), .C1(
        n9767), .C2(n9766), .ZN(P1_U3329) );
  MUX2_X1 U10977 ( .A(n9771), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10978 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9783) );
  AOI211_X1 U10979 ( .C1(n9774), .C2(n9773), .A(n9772), .B(n9889), .ZN(n9779)
         );
  AOI211_X1 U10980 ( .C1(n9777), .C2(n9776), .A(n9895), .B(n9775), .ZN(n9778)
         );
  AOI211_X1 U10981 ( .C1(n9901), .C2(n9780), .A(n9779), .B(n9778), .ZN(n9782)
         );
  NAND2_X1 U10982 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9781) );
  OAI211_X1 U10983 ( .C1(n9904), .C2(n9783), .A(n9782), .B(n9781), .ZN(
        P1_U3253) );
  INV_X1 U10984 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9795) );
  AOI211_X1 U10985 ( .C1(n9786), .C2(n9785), .A(n9889), .B(n9784), .ZN(n9791)
         );
  AOI211_X1 U10986 ( .C1(n9789), .C2(n9788), .A(n9895), .B(n9787), .ZN(n9790)
         );
  AOI211_X1 U10987 ( .C1(n9901), .C2(n9792), .A(n9791), .B(n9790), .ZN(n9794)
         );
  NAND2_X1 U10988 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9793) );
  OAI211_X1 U10989 ( .C1(n9904), .C2(n9795), .A(n9794), .B(n9793), .ZN(
        P1_U3250) );
  OAI21_X1 U10990 ( .B1(n9798), .B2(n9797), .A(n9796), .ZN(n9807) );
  AOI21_X1 U10991 ( .B1(n9801), .B2(n9800), .A(n9799), .ZN(n9802) );
  OAI21_X1 U10992 ( .B1(n9804), .B2(n9803), .A(n9802), .ZN(n9805) );
  AOI21_X1 U10993 ( .B1(n9807), .B2(n9806), .A(n9805), .ZN(n9808) );
  OAI21_X1 U10994 ( .B1(n9810), .B2(n9809), .A(n9808), .ZN(P1_U3224) );
  XNOR2_X1 U10995 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10996 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10997 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9822) );
  AOI211_X1 U10998 ( .C1(n9813), .C2(n9812), .A(n9811), .B(n9889), .ZN(n9818)
         );
  AOI211_X1 U10999 ( .C1(n9816), .C2(n9815), .A(n9814), .B(n9895), .ZN(n9817)
         );
  AOI211_X1 U11000 ( .C1(n9901), .C2(n9819), .A(n9818), .B(n9817), .ZN(n9821)
         );
  NAND2_X1 U11001 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9820) );
  OAI211_X1 U11002 ( .C1(n9904), .C2(n9822), .A(n9821), .B(n9820), .ZN(
        P1_U3254) );
  INV_X1 U11003 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9834) );
  AOI211_X1 U11004 ( .C1(n9825), .C2(n9824), .A(n9823), .B(n9895), .ZN(n9830)
         );
  AOI211_X1 U11005 ( .C1(n9828), .C2(n9827), .A(n9826), .B(n9889), .ZN(n9829)
         );
  AOI211_X1 U11006 ( .C1(n9901), .C2(n9831), .A(n9830), .B(n9829), .ZN(n9833)
         );
  OAI211_X1 U11007 ( .C1(n9904), .C2(n9834), .A(n9833), .B(n9832), .ZN(
        P1_U3256) );
  INV_X1 U11008 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9849) );
  AOI21_X1 U11009 ( .B1(n9837), .B2(n9836), .A(n9835), .ZN(n9838) );
  NAND2_X1 U11010 ( .A1(n9883), .A2(n9838), .ZN(n9846) );
  NAND2_X1 U11011 ( .A1(n9840), .A2(n9839), .ZN(n9841) );
  NAND3_X1 U11012 ( .A1(n9880), .A2(n9842), .A3(n9841), .ZN(n9845) );
  NAND2_X1 U11013 ( .A1(n9901), .A2(n9843), .ZN(n9844) );
  AND3_X1 U11014 ( .A1(n9846), .A2(n9845), .A3(n9844), .ZN(n9848) );
  NAND2_X1 U11015 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9847) );
  OAI211_X1 U11016 ( .C1(n9904), .C2(n9849), .A(n9848), .B(n9847), .ZN(
        P1_U3257) );
  AOI211_X1 U11017 ( .C1(n9852), .C2(n9851), .A(n9895), .B(n9850), .ZN(n9856)
         );
  AOI211_X1 U11018 ( .C1(n9854), .C2(n5344), .A(n9853), .B(n9889), .ZN(n9855)
         );
  AOI211_X1 U11019 ( .C1(n9901), .C2(n9857), .A(n9856), .B(n9855), .ZN(n9859)
         );
  OAI211_X1 U11020 ( .C1(n9860), .C2(n9904), .A(n9859), .B(n9858), .ZN(
        P1_U3258) );
  AOI211_X1 U11021 ( .C1(n9863), .C2(n9862), .A(n9861), .B(n9889), .ZN(n9864)
         );
  AOI211_X1 U11022 ( .C1(n9866), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9865), .B(
        n9864), .ZN(n9873) );
  OAI21_X1 U11023 ( .B1(n9869), .B2(n9868), .A(n9867), .ZN(n9871) );
  AOI22_X1 U11024 ( .A1(n9871), .A2(n9880), .B1(n9870), .B2(n9901), .ZN(n9872)
         );
  NAND2_X1 U11025 ( .A1(n9873), .A2(n9872), .ZN(P1_U3259) );
  OAI21_X1 U11026 ( .B1(n9876), .B2(n9875), .A(n9874), .ZN(n9884) );
  OAI21_X1 U11027 ( .B1(n9879), .B2(n9878), .A(n9877), .ZN(n9881) );
  AOI222_X1 U11028 ( .A1(n9884), .A2(n9883), .B1(n9882), .B2(n9901), .C1(n9881), .C2(n9880), .ZN(n9886) );
  OAI211_X1 U11029 ( .C1(n9904), .C2(n9887), .A(n9886), .B(n9885), .ZN(
        P1_U3260) );
  INV_X1 U11030 ( .A(n9888), .ZN(n9890) );
  AOI211_X1 U11031 ( .C1(n9892), .C2(n9891), .A(n9890), .B(n9889), .ZN(n9899)
         );
  INV_X1 U11032 ( .A(n9893), .ZN(n9894) );
  AOI211_X1 U11033 ( .C1(n9897), .C2(n9896), .A(n9895), .B(n9894), .ZN(n9898)
         );
  AOI211_X1 U11034 ( .C1(n9901), .C2(n9900), .A(n9899), .B(n9898), .ZN(n9903)
         );
  NAND2_X1 U11035 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9902) );
  OAI211_X1 U11036 ( .C1(n9904), .C2(n10131), .A(n9903), .B(n9902), .ZN(
        P1_U3261) );
  NAND2_X1 U11037 ( .A1(n9906), .A2(n9905), .ZN(n9912) );
  INV_X1 U11038 ( .A(n9907), .ZN(n9909) );
  AOI22_X1 U11039 ( .A1(n9910), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9909), .B2(
        n9908), .ZN(n9911) );
  OAI211_X1 U11040 ( .C1(n9914), .C2(n9913), .A(n9912), .B(n9911), .ZN(n9915)
         );
  AOI21_X1 U11041 ( .B1(n9917), .B2(n9916), .A(n9915), .ZN(n9918) );
  OAI21_X1 U11042 ( .B1(n9934), .B2(n9919), .A(n9918), .ZN(P1_U3282) );
  OAI22_X1 U11043 ( .A1(n9922), .A2(n9921), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9920), .ZN(n9923) );
  AOI21_X1 U11044 ( .B1(n9925), .B2(n9924), .A(n9923), .ZN(n9926) );
  OAI21_X1 U11045 ( .B1(n9928), .B2(n9927), .A(n9926), .ZN(n9929) );
  AOI21_X1 U11046 ( .B1(n9931), .B2(n9930), .A(n9929), .ZN(n9932) );
  OAI21_X1 U11047 ( .B1(n9934), .B2(n9933), .A(n9932), .ZN(P1_U3290) );
  AND2_X1 U11048 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9937), .ZN(P1_U3294) );
  AND2_X1 U11049 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9937), .ZN(P1_U3295) );
  AND2_X1 U11050 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9937), .ZN(P1_U3296) );
  AND2_X1 U11051 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9937), .ZN(P1_U3297) );
  AND2_X1 U11052 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9937), .ZN(P1_U3298) );
  AND2_X1 U11053 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9937), .ZN(P1_U3299) );
  AND2_X1 U11054 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9937), .ZN(P1_U3300) );
  AND2_X1 U11055 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9937), .ZN(P1_U3301) );
  AND2_X1 U11056 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9937), .ZN(P1_U3302) );
  AND2_X1 U11057 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9937), .ZN(P1_U3303) );
  AND2_X1 U11058 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9937), .ZN(P1_U3304) );
  AND2_X1 U11059 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9937), .ZN(P1_U3305) );
  AND2_X1 U11060 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9937), .ZN(P1_U3306) );
  AND2_X1 U11061 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9937), .ZN(P1_U3307) );
  AND2_X1 U11062 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9937), .ZN(P1_U3308) );
  AND2_X1 U11063 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9937), .ZN(P1_U3309) );
  AND2_X1 U11064 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9937), .ZN(P1_U3310) );
  AND2_X1 U11065 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9937), .ZN(P1_U3311) );
  AND2_X1 U11066 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9937), .ZN(P1_U3312) );
  AND2_X1 U11067 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9937), .ZN(P1_U3313) );
  AND2_X1 U11068 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9937), .ZN(P1_U3314) );
  AND2_X1 U11069 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9937), .ZN(P1_U3315) );
  NOR2_X1 U11070 ( .A1(n9936), .A2(n9935), .ZN(P1_U3316) );
  AND2_X1 U11071 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9937), .ZN(P1_U3317) );
  AND2_X1 U11072 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9937), .ZN(P1_U3318) );
  AND2_X1 U11073 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9937), .ZN(P1_U3319) );
  AND2_X1 U11074 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9937), .ZN(P1_U3320) );
  AND2_X1 U11075 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9937), .ZN(P1_U3321) );
  AND2_X1 U11076 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9937), .ZN(P1_U3322) );
  AND2_X1 U11077 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9937), .ZN(P1_U3323) );
  OAI21_X1 U11078 ( .B1(n9940), .B2(n9939), .A(n9938), .ZN(n9942) );
  AOI211_X1 U11079 ( .C1(n9944), .C2(n9943), .A(n9942), .B(n9941), .ZN(n9956)
         );
  INV_X1 U11080 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9945) );
  AOI22_X1 U11081 ( .A1(n9946), .A2(n9956), .B1(n9945), .B2(n9955), .ZN(
        P1_U3459) );
  AOI21_X1 U11082 ( .B1(n9949), .B2(n9948), .A(n9947), .ZN(n9950) );
  OAI211_X1 U11083 ( .C1(n9953), .C2(n9952), .A(n9951), .B(n9950), .ZN(n9954)
         );
  INV_X1 U11084 ( .A(n9954), .ZN(n9958) );
  AOI22_X1 U11085 ( .A1(n9946), .A2(n9958), .B1(n5111), .B2(n9955), .ZN(
        P1_U3471) );
  AOI22_X1 U11086 ( .A1(n9959), .A2(n9956), .B1(n6645), .B2(n9957), .ZN(
        P1_U3524) );
  AOI22_X1 U11087 ( .A1(n9959), .A2(n9958), .B1(n6672), .B2(n9957), .ZN(
        P1_U3528) );
  INV_X1 U11088 ( .A(n4426), .ZN(n9961) );
  NAND2_X1 U11089 ( .A1(n10011), .A2(n9961), .ZN(n9976) );
  NAND2_X1 U11090 ( .A1(n9963), .A2(n9962), .ZN(n9964) );
  AND2_X1 U11091 ( .A1(n9965), .A2(n9964), .ZN(n9966) );
  OR2_X1 U11092 ( .A1(n9967), .A2(n9966), .ZN(n9975) );
  NAND2_X1 U11093 ( .A1(n9969), .A2(n9968), .ZN(n9970) );
  AND2_X1 U11094 ( .A1(n9971), .A2(n9970), .ZN(n9972) );
  OR2_X1 U11095 ( .A1(n10024), .A2(n9972), .ZN(n9974) );
  NAND2_X1 U11096 ( .A1(P2_U3151), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9973) );
  AND4_X1 U11097 ( .A1(n9976), .A2(n9975), .A3(n9974), .A4(n9973), .ZN(n9981)
         );
  XOR2_X1 U11098 ( .A(n9978), .B(n9977), .Z(n9979) );
  NAND2_X1 U11099 ( .A1(n9979), .A2(n10001), .ZN(n9980) );
  OAI211_X1 U11100 ( .C1(n10129), .C2(n9982), .A(n9981), .B(n9980), .ZN(
        P2_U3183) );
  OAI21_X1 U11101 ( .B1(n9985), .B2(n9984), .A(n9983), .ZN(n9988) );
  NOR2_X1 U11102 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9986), .ZN(n9987) );
  AOI21_X1 U11103 ( .B1(n10014), .B2(n9988), .A(n9987), .ZN(n9998) );
  NAND2_X1 U11104 ( .A1(n10011), .A2(n9989), .ZN(n9997) );
  NAND2_X1 U11105 ( .A1(n10013), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n9996) );
  OAI21_X1 U11106 ( .B1(n9992), .B2(n9991), .A(n9990), .ZN(n9993) );
  INV_X1 U11107 ( .A(n9993), .ZN(n9994) );
  OR2_X1 U11108 ( .A1(n10024), .A2(n9994), .ZN(n9995) );
  AND4_X1 U11109 ( .A1(n9998), .A2(n9997), .A3(n9996), .A4(n9995), .ZN(n10004)
         );
  XOR2_X1 U11110 ( .A(n10000), .B(n9999), .Z(n10002) );
  NAND2_X1 U11111 ( .A1(n10002), .A2(n10001), .ZN(n10003) );
  NAND2_X1 U11112 ( .A1(n10004), .A2(n10003), .ZN(P2_U3184) );
  INV_X1 U11113 ( .A(n10005), .ZN(n10010) );
  NAND3_X1 U11114 ( .A1(n10008), .A2(n10007), .A3(n10006), .ZN(n10009) );
  NAND2_X1 U11115 ( .A1(n10010), .A2(n10009), .ZN(n10015) );
  AOI222_X1 U11116 ( .A1(n10015), .A2(n10014), .B1(n10013), .B2(
        P2_ADDR_REG_8__SCAN_IN), .C1(n10012), .C2(n10011), .ZN(n10029) );
  AOI21_X1 U11117 ( .B1(n10018), .B2(n10017), .A(n10016), .ZN(n10020) );
  OR2_X1 U11118 ( .A1(n10020), .A2(n10019), .ZN(n10027) );
  AOI21_X1 U11119 ( .B1(n10023), .B2(n10022), .A(n10021), .ZN(n10025) );
  OR2_X1 U11120 ( .A1(n10025), .A2(n10024), .ZN(n10026) );
  NAND4_X1 U11121 ( .A1(n10029), .A2(n10028), .A3(n10027), .A4(n10026), .ZN(
        P2_U3190) );
  NAND2_X1 U11122 ( .A1(n10031), .A2(n10030), .ZN(n10032) );
  XNOR2_X1 U11123 ( .A(n10032), .B(n10034), .ZN(n10077) );
  XOR2_X1 U11124 ( .A(n10033), .B(n10034), .Z(n10035) );
  OAI222_X1 U11125 ( .A1(n10039), .A2(n10038), .B1(n10037), .B2(n10036), .C1(
        n10050), .C2(n10035), .ZN(n10078) );
  MUX2_X1 U11126 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10078), .S(n8616), .Z(
        n10045) );
  OAI22_X1 U11127 ( .A1(n10043), .A2(n10042), .B1(n10041), .B2(n10040), .ZN(
        n10044) );
  NOR2_X1 U11128 ( .A1(n10045), .A2(n10044), .ZN(n10046) );
  OAI21_X1 U11129 ( .B1(n10047), .B2(n10077), .A(n10046), .ZN(P2_U3227) );
  INV_X1 U11130 ( .A(n10048), .ZN(n10049) );
  AOI21_X1 U11131 ( .B1(n10090), .B2(n10050), .A(n10049), .ZN(n10051) );
  AOI211_X1 U11132 ( .C1(n10081), .C2(n10053), .A(n10052), .B(n10051), .ZN(
        n10111) );
  INV_X1 U11133 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10054) );
  AOI22_X1 U11134 ( .A1(n10110), .A2(n10111), .B1(n10054), .B2(n10108), .ZN(
        P2_U3390) );
  OAI22_X1 U11135 ( .A1(n10056), .A2(n10104), .B1(n10055), .B2(n10102), .ZN(
        n10057) );
  NOR2_X1 U11136 ( .A1(n10058), .A2(n10057), .ZN(n10113) );
  INV_X1 U11137 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10059) );
  AOI22_X1 U11138 ( .A1(n10110), .A2(n10113), .B1(n10059), .B2(n10108), .ZN(
        P2_U3396) );
  INV_X1 U11139 ( .A(n10060), .ZN(n10064) );
  OAI22_X1 U11140 ( .A1(n10062), .A2(n10090), .B1(n10061), .B2(n10102), .ZN(
        n10063) );
  NOR2_X1 U11141 ( .A1(n10064), .A2(n10063), .ZN(n10114) );
  INV_X1 U11142 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10065) );
  AOI22_X1 U11143 ( .A1(n10110), .A2(n10114), .B1(n10065), .B2(n10108), .ZN(
        P2_U3399) );
  OAI21_X1 U11144 ( .B1(n10067), .B2(n10102), .A(n10066), .ZN(n10068) );
  AOI21_X1 U11145 ( .B1(n10069), .B2(n10074), .A(n10068), .ZN(n10115) );
  INV_X1 U11146 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10070) );
  AOI22_X1 U11147 ( .A1(n10110), .A2(n10115), .B1(n10070), .B2(n10108), .ZN(
        P2_U3402) );
  OAI21_X1 U11148 ( .B1(n10072), .B2(n10102), .A(n10071), .ZN(n10073) );
  AOI21_X1 U11149 ( .B1(n10075), .B2(n10074), .A(n10073), .ZN(n10116) );
  INV_X1 U11150 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10076) );
  AOI22_X1 U11151 ( .A1(n10110), .A2(n10116), .B1(n10076), .B2(n10108), .ZN(
        P2_U3405) );
  NOR2_X1 U11152 ( .A1(n10077), .A2(n10090), .ZN(n10079) );
  AOI211_X1 U11153 ( .C1(n10081), .C2(n10080), .A(n10079), .B(n10078), .ZN(
        n10117) );
  INV_X1 U11154 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10082) );
  AOI22_X1 U11155 ( .A1(n10110), .A2(n10117), .B1(n10082), .B2(n10108), .ZN(
        P2_U3408) );
  OAI22_X1 U11156 ( .A1(n10084), .A2(n10104), .B1(n10083), .B2(n10102), .ZN(
        n10085) );
  AOI211_X1 U11157 ( .C1(n10100), .C2(n10087), .A(n10086), .B(n10085), .ZN(
        n10118) );
  INV_X1 U11158 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10088) );
  AOI22_X1 U11159 ( .A1(n10110), .A2(n10118), .B1(n10088), .B2(n10108), .ZN(
        P2_U3411) );
  OAI22_X1 U11160 ( .A1(n10091), .A2(n10090), .B1(n10089), .B2(n10102), .ZN(
        n10093) );
  NOR2_X1 U11161 ( .A1(n10093), .A2(n10092), .ZN(n10119) );
  AOI22_X1 U11162 ( .A1(n10110), .A2(n10119), .B1(n10094), .B2(n10108), .ZN(
        P2_U3414) );
  OAI22_X1 U11163 ( .A1(n10096), .A2(n10104), .B1(n10095), .B2(n10102), .ZN(
        n10097) );
  AOI211_X1 U11164 ( .C1(n10100), .C2(n10099), .A(n10098), .B(n10097), .ZN(
        n10121) );
  INV_X1 U11165 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10101) );
  AOI22_X1 U11166 ( .A1(n10110), .A2(n10121), .B1(n10101), .B2(n10108), .ZN(
        P2_U3417) );
  OAI22_X1 U11167 ( .A1(n10105), .A2(n10104), .B1(n10103), .B2(n10102), .ZN(
        n10106) );
  NOR2_X1 U11168 ( .A1(n10107), .A2(n10106), .ZN(n10123) );
  INV_X1 U11169 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10109) );
  AOI22_X1 U11170 ( .A1(n10110), .A2(n10123), .B1(n10109), .B2(n10108), .ZN(
        P2_U3420) );
  AOI22_X1 U11171 ( .A1(n10124), .A2(n10111), .B1(n6405), .B2(n10122), .ZN(
        P2_U3459) );
  AOI22_X1 U11172 ( .A1(n10124), .A2(n10113), .B1(n10112), .B2(n10122), .ZN(
        P2_U3461) );
  AOI22_X1 U11173 ( .A1(n10124), .A2(n10114), .B1(n5853), .B2(n10122), .ZN(
        P2_U3462) );
  AOI22_X1 U11174 ( .A1(n10124), .A2(n10115), .B1(n6348), .B2(n10122), .ZN(
        P2_U3463) );
  AOI22_X1 U11175 ( .A1(n10124), .A2(n10116), .B1(n4643), .B2(n10122), .ZN(
        P2_U3464) );
  AOI22_X1 U11176 ( .A1(n10124), .A2(n10117), .B1(n6415), .B2(n10122), .ZN(
        P2_U3465) );
  AOI22_X1 U11177 ( .A1(n10124), .A2(n10118), .B1(n5922), .B2(n10122), .ZN(
        P2_U3466) );
  AOI22_X1 U11178 ( .A1(n10124), .A2(n10119), .B1(n6353), .B2(n10122), .ZN(
        P2_U3467) );
  AOI22_X1 U11179 ( .A1(n10124), .A2(n10121), .B1(n10120), .B2(n10122), .ZN(
        P2_U3468) );
  AOI22_X1 U11180 ( .A1(n10124), .A2(n10123), .B1(n6404), .B2(n10122), .ZN(
        P2_U3469) );
  OAI222_X1 U11181 ( .A1(n10129), .A2(n10128), .B1(n10129), .B2(n10127), .C1(
        n10126), .C2(n10125), .ZN(ADD_1068_U5) );
  XOR2_X1 U11182 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U11183 ( .B1(n10132), .B2(n10131), .A(n10130), .ZN(n10134) );
  XOR2_X1 U11184 ( .A(n10134), .B(n10133), .Z(ADD_1068_U55) );
  OAI21_X1 U11185 ( .B1(n10137), .B2(n10136), .A(n10135), .ZN(ADD_1068_U56) );
  OAI21_X1 U11186 ( .B1(n10140), .B2(n10139), .A(n10138), .ZN(ADD_1068_U57) );
  OAI21_X1 U11187 ( .B1(n10143), .B2(n10142), .A(n10141), .ZN(ADD_1068_U58) );
  OAI21_X1 U11188 ( .B1(n10146), .B2(n10145), .A(n10144), .ZN(ADD_1068_U59) );
  OAI21_X1 U11189 ( .B1(n10149), .B2(n10148), .A(n10147), .ZN(ADD_1068_U60) );
  OAI21_X1 U11190 ( .B1(n10152), .B2(n10151), .A(n10150), .ZN(ADD_1068_U61) );
  OAI21_X1 U11191 ( .B1(n10155), .B2(n10154), .A(n10153), .ZN(ADD_1068_U62) );
  OAI21_X1 U11192 ( .B1(n10158), .B2(n10157), .A(n10156), .ZN(ADD_1068_U63) );
  OAI21_X1 U11193 ( .B1(n10161), .B2(n10160), .A(n10159), .ZN(ADD_1068_U50) );
  OAI21_X1 U11194 ( .B1(n10164), .B2(n10163), .A(n10162), .ZN(ADD_1068_U51) );
  OAI21_X1 U11195 ( .B1(n10167), .B2(n10166), .A(n10165), .ZN(ADD_1068_U47) );
  OAI21_X1 U11196 ( .B1(n10170), .B2(n10169), .A(n10168), .ZN(ADD_1068_U49) );
  OAI21_X1 U11197 ( .B1(n10173), .B2(n10172), .A(n10171), .ZN(ADD_1068_U48) );
  AOI21_X1 U11198 ( .B1(n10176), .B2(n10175), .A(n10174), .ZN(ADD_1068_U54) );
  AOI21_X1 U11199 ( .B1(n10179), .B2(n10178), .A(n10177), .ZN(ADD_1068_U53) );
  OAI21_X1 U11200 ( .B1(n10182), .B2(n10181), .A(n10180), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4817 ( .A(n8004), .Z(n6141) );
  INV_X2 U4837 ( .A(n7894), .ZN(n7910) );
  CLKBUF_X1 U4848 ( .A(n5879), .Z(n6083) );
  CLKBUF_X1 U4877 ( .A(n5804), .Z(n7707) );
  CLKBUF_X1 U4986 ( .A(n6072), .Z(n4314) );
  CLKBUF_X1 U5186 ( .A(n4980), .Z(n4316) );
endmodule

