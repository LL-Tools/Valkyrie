

module b15_C_gen_AntiSAT_k_256_4 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66,
         keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71,
         keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76,
         keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81,
         keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86,
         keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91,
         keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96,
         keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145;

  CLKBUF_X2 U3599 ( .A(n3569), .Z(n4694) );
  AND2_X1 U3600 ( .A1(n3398), .A2(n4783), .ZN(n3694) );
  NAND4_X2 U3601 ( .A1(n3287), .A2(n3286), .A3(n3285), .A4(n3284), .ZN(n3385)
         );
  AND2_X1 U3602 ( .A1(n4695), .A2(n3243), .ZN(n3289) );
  AND2_X2 U3603 ( .A1(n4545), .A2(n3251), .ZN(n3546) );
  INV_X1 U3605 ( .A(n7145), .ZN(n3152) );
  NAND2_X1 U3606 ( .A1(n3366), .A2(n3398), .ZN(n3741) );
  AND2_X1 U3608 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4692) );
  AND4_X1 U3609 ( .A1(n3261), .A2(n3260), .A3(n3259), .A4(n3258), .ZN(n3267)
         );
  OR2_X1 U3610 ( .A1(n3936), .A2(n4659), .ZN(n4754) );
  INV_X2 U3611 ( .A(n4874), .ZN(n3859) );
  NAND2_X1 U3612 ( .A1(n3938), .A2(n3937), .ZN(n4752) );
  NAND2_X1 U3613 ( .A1(n5630), .A2(n5653), .ZN(n5647) );
  AOI221_X1 U3614 ( .B1(REIP_REG_26__SCAN_IN), .B2(n6005), .C1(n6004), .C2(
        n6005), .A(n6003), .ZN(n6006) );
  INV_X1 U3615 ( .A(n6267), .ZN(n6280) );
  OAI21_X1 U3616 ( .B1(n5630), .B2(n5653), .A(n5647), .ZN(n6002) );
  INV_X1 U3617 ( .A(n4217), .ZN(n3425) );
  INV_X2 U3618 ( .A(n4973), .ZN(n3998) );
  AOI21_X2 U3619 ( .B1(n5729), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5728), 
        .ZN(n5730) );
  XNOR2_X2 U3620 ( .A(n3560), .B(n4895), .ZN(n4798) );
  INV_X2 U3622 ( .A(n4727), .ZN(n5415) );
  AND2_X4 U3623 ( .A1(n3249), .A2(n4692), .ZN(n3459) );
  INV_X1 U3624 ( .A(n6100), .ZN(n6101) );
  NAND2_X2 U3625 ( .A1(n3511), .A2(n3510), .ZN(n4727) );
  NAND2_X1 U3626 ( .A1(n3494), .A2(n3507), .ZN(n3511) );
  AND2_X1 U3628 ( .A1(n3408), .A2(n3379), .ZN(n3389) );
  AND4_X1 U3629 ( .A1(n3407), .A2(n6653), .A3(n4698), .A4(n3406), .ZN(n3409)
         );
  AND2_X1 U3630 ( .A1(n3374), .A2(n3324), .ZN(n4540) );
  AND2_X2 U3631 ( .A1(n3685), .A2(n3153), .ZN(n3512) );
  OAI22_X1 U3632 ( .A1(n3425), .A2(n3296), .B1(n3295), .B2(n3294), .ZN(n3297)
         );
  CLKBUF_X2 U3633 ( .A(n3430), .Z(n4372) );
  BUF_X2 U3634 ( .A(n4384), .Z(n4351) );
  CLKBUF_X2 U3635 ( .A(n4380), .Z(n4229) );
  CLKBUF_X2 U3636 ( .A(n3351), .Z(n4356) );
  CLKBUF_X2 U3637 ( .A(n3288), .Z(n4234) );
  BUF_X2 U3638 ( .A(n3289), .Z(n4373) );
  CLKBUF_X2 U3639 ( .A(n3350), .Z(n4382) );
  BUF_X2 U3640 ( .A(n3348), .Z(n4374) );
  CLKBUF_X2 U3641 ( .A(n3349), .Z(n4381) );
  AOI22_X1 U3642 ( .A1(n5566), .A2(n5747), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5885), .ZN(n5567) );
  OAI21_X1 U3643 ( .B1(n5738), .B2(n5835), .A(n3903), .ZN(n3904) );
  NAND2_X1 U3644 ( .A1(n3901), .A2(n3900), .ZN(n5727) );
  NAND2_X1 U3645 ( .A1(n5777), .A2(n5778), .ZN(n5776) );
  NOR3_X1 U3646 ( .A1(n5989), .A2(n5988), .A3(n5987), .ZN(n5990) );
  AOI21_X1 U3647 ( .B1(n5783), .B2(n5784), .A(n3673), .ZN(n5777) );
  XNOR2_X1 U3648 ( .A(n4405), .B(n4404), .ZN(n5584) );
  OR3_X1 U3649 ( .A1(n5565), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n5755), 
        .ZN(n5747) );
  AND2_X1 U3650 ( .A1(n6092), .A2(n3672), .ZN(n5783) );
  OAI21_X1 U3651 ( .B1(n5570), .B2(n5571), .A(n5618), .ZN(n5576) );
  NOR2_X1 U3652 ( .A1(n5647), .A2(n3229), .ZN(n5619) );
  CLKBUF_X1 U3653 ( .A(n5628), .Z(n5629) );
  NAND2_X1 U3654 ( .A1(n3217), .A2(n3156), .ZN(n3216) );
  AND2_X1 U3655 ( .A1(n4096), .A2(n3173), .ZN(n5695) );
  OR2_X1 U3656 ( .A1(n5257), .A2(n4060), .ZN(n5543) );
  NAND2_X2 U3657 ( .A1(n3998), .A2(n3171), .ZN(n5257) );
  AND3_X1 U3658 ( .A1(n3206), .A2(n3207), .A3(n3662), .ZN(n3205) );
  AOI21_X1 U3659 ( .B1(n3965), .B2(n4087), .A(n3964), .ZN(n4956) );
  AND2_X1 U3660 ( .A1(n3537), .A2(n3536), .ZN(n6367) );
  XNOR2_X1 U3661 ( .A(n3640), .B(n3639), .ZN(n3965) );
  NAND2_X1 U3662 ( .A1(n3625), .A2(n3626), .ZN(n3640) );
  NAND2_X1 U3663 ( .A1(n4754), .A2(n4753), .ZN(n3938) );
  NOR2_X2 U3664 ( .A1(n6132), .A2(n6131), .ZN(n6133) );
  XNOR2_X1 U3665 ( .A(n3609), .B(n3611), .ZN(n3946) );
  NAND2_X1 U3666 ( .A1(n3945), .A2(n3944), .ZN(n4766) );
  NOR3_X1 U3667 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6262), .A3(n6543), .ZN(
        n6265) );
  BUF_X1 U3668 ( .A(n6346), .Z(n6337) );
  AND2_X1 U3669 ( .A1(n4895), .A2(n3611), .ZN(n3221) );
  NAND2_X1 U3670 ( .A1(n6111), .A2(n4410), .ZN(n6384) );
  NAND2_X2 U3671 ( .A1(n3559), .A2(n3558), .ZN(n4895) );
  NAND2_X1 U3672 ( .A1(n4690), .A2(n6656), .ZN(n3559) );
  NAND2_X1 U3673 ( .A1(n3511), .A2(n3496), .ZN(n3522) );
  NAND2_X1 U3674 ( .A1(n3181), .A2(n3180), .ZN(n5082) );
  INV_X1 U3675 ( .A(n4841), .ZN(n3181) );
  AND2_X1 U3676 ( .A1(n4664), .A2(n3783), .ZN(n4764) );
  OR2_X1 U3677 ( .A1(n3453), .A2(n3452), .ZN(n3525) );
  OR2_X1 U3678 ( .A1(n3467), .A2(n3466), .ZN(n3652) );
  OR2_X1 U3679 ( .A1(n3487), .A2(n3486), .ZN(n3524) );
  INV_X2 U3680 ( .A(n3380), .ZN(n3685) );
  NAND2_X2 U3681 ( .A1(n3312), .A2(n3162), .ZN(n4819) );
  NAND2_X2 U3682 ( .A1(n3161), .A2(n3322), .ZN(n3383) );
  AND4_X1 U3683 ( .A1(n3255), .A2(n3254), .A3(n3253), .A4(n3252), .ZN(n3256)
         );
  AND4_X1 U3684 ( .A1(n3307), .A2(n3306), .A3(n3305), .A4(n3304), .ZN(n3312)
         );
  AND4_X1 U3685 ( .A1(n3345), .A2(n3344), .A3(n3343), .A4(n3342), .ZN(n3346)
         );
  AND4_X1 U3686 ( .A1(n3321), .A2(n3320), .A3(n3319), .A4(n3318), .ZN(n3322)
         );
  AND4_X1 U3687 ( .A1(n3279), .A2(n3278), .A3(n3277), .A4(n3276), .ZN(n3285)
         );
  AND4_X1 U3688 ( .A1(n3328), .A2(n3327), .A3(n3326), .A4(n3325), .ZN(n3341)
         );
  AND4_X1 U3689 ( .A1(n3283), .A2(n3282), .A3(n3281), .A4(n3280), .ZN(n3284)
         );
  AND4_X1 U3690 ( .A1(n3271), .A2(n3270), .A3(n3269), .A4(n3268), .ZN(n3287)
         );
  AND4_X1 U3691 ( .A1(n3275), .A2(n3274), .A3(n3273), .A4(n3272), .ZN(n3286)
         );
  AND4_X1 U3692 ( .A1(n3265), .A2(n3264), .A3(n3263), .A4(n3262), .ZN(n3266)
         );
  NAND2_X2 U3693 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6713), .ZN(n6708) );
  AND2_X2 U3694 ( .A1(n3250), .A2(n4691), .ZN(n3545) );
  AND2_X2 U3695 ( .A1(n3250), .A2(n3251), .ZN(n4217) );
  AND2_X2 U3696 ( .A1(n4545), .A2(n3248), .ZN(n3569) );
  AND2_X2 U3697 ( .A1(n3248), .A2(n3250), .ZN(n4380) );
  AND2_X2 U3698 ( .A1(n3249), .A2(n3251), .ZN(n4384) );
  AND2_X2 U3699 ( .A1(n3251), .A2(n4544), .ZN(n3288) );
  AND2_X1 U3700 ( .A1(n3939), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3248)
         );
  AND2_X1 U3701 ( .A1(n3682), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3249)
         );
  AND2_X2 U3702 ( .A1(n3370), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3250)
         );
  NAND2_X1 U3703 ( .A1(n6722), .A2(n6655), .ZN(n6543) );
  AND2_X2 U3704 ( .A1(n4545), .A2(n4692), .ZN(n3356) );
  AND2_X2 U3705 ( .A1(n4544), .A2(n4692), .ZN(n3348) );
  NOR2_X2 U3706 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4691) );
  NOR2_X1 U3707 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3243) );
  INV_X1 U3708 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6722) );
  XNOR2_X1 U3709 ( .A(n3567), .B(n6444), .ZN(n6368) );
  NAND2_X1 U3710 ( .A1(n3566), .A2(n3565), .ZN(n3567) );
  NAND2_X2 U3711 ( .A1(n3899), .A2(n3239), .ZN(n3901) );
  AND2_X2 U3712 ( .A1(n5628), .A2(n5627), .ZN(n5630) );
  AND2_X2 U3713 ( .A1(n3390), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3415) );
  NAND2_X1 U3714 ( .A1(n3347), .A2(n3346), .ZN(n3153) );
  NAND2_X1 U3715 ( .A1(n3347), .A2(n3346), .ZN(n3154) );
  NOR2_X2 U3716 ( .A1(n4839), .A2(n4956), .ZN(n4972) );
  OR2_X1 U3717 ( .A1(n3741), .A2(n3385), .ZN(n3386) );
  AND3_X1 U3718 ( .A1(n3385), .A2(n4874), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3695) );
  AND2_X2 U3719 ( .A1(n3257), .A2(n3256), .ZN(n3365) );
  AND4_X1 U3720 ( .A1(n3247), .A2(n3246), .A3(n3245), .A4(n3244), .ZN(n3257)
         );
  NAND2_X1 U3721 ( .A1(n3640), .A2(n3651), .ZN(n3155) );
  OAI22_X2 U3722 ( .A1(n5812), .A2(n3666), .B1(n6101), .B2(n5813), .ZN(n5804)
         );
  OR2_X2 U3723 ( .A1(n3303), .A2(n3302), .ZN(n4832) );
  OAI21_X2 U3724 ( .B1(n4776), .B2(n4027), .A(n3919), .ZN(n3936) );
  NAND2_X2 U3725 ( .A1(n3501), .A2(n3560), .ZN(n4776) );
  NAND2_X4 U3726 ( .A1(n3772), .A2(n4874), .ZN(n4455) );
  NAND2_X4 U3727 ( .A1(n3347), .A2(n3346), .ZN(n4874) );
  OR2_X1 U3728 ( .A1(n3403), .A2(n3685), .ZN(n3407) );
  OR2_X1 U3729 ( .A1(n6101), .A2(n3896), .ZN(n3897) );
  INV_X1 U3730 ( .A(n5804), .ZN(n3217) );
  INV_X1 U3731 ( .A(n5521), .ZN(n3207) );
  INV_X1 U3732 ( .A(n5297), .ZN(n3213) );
  OR2_X1 U3733 ( .A1(n6741), .A2(n4433), .ZN(n5248) );
  AND2_X1 U3734 ( .A1(n5248), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4965) );
  NAND2_X1 U3735 ( .A1(n3233), .A2(n3230), .ZN(n3229) );
  INV_X1 U3736 ( .A(n5620), .ZN(n3233) );
  INV_X1 U3737 ( .A(n3231), .ZN(n3230) );
  NOR2_X1 U3738 ( .A1(n4496), .A2(n3833), .ZN(n4505) );
  AND2_X2 U3739 ( .A1(n4601), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3251)
         );
  CLKBUF_X2 U3740 ( .A(n3545), .Z(n4379) );
  INV_X1 U3741 ( .A(n3560), .ZN(n3222) );
  NAND2_X1 U3742 ( .A1(n3222), .A2(n4895), .ZN(n3609) );
  NAND2_X1 U3743 ( .A1(n3581), .A2(n3580), .ZN(n3611) );
  NOR2_X1 U3744 ( .A1(n3745), .A2(n3388), .ZN(n3403) );
  NAND2_X1 U3745 ( .A1(n5571), .A2(n3232), .ZN(n3231) );
  INV_X1 U3746 ( .A(n5648), .ZN(n3232) );
  INV_X1 U3747 ( .A(n4367), .ZN(n4393) );
  NAND2_X1 U3748 ( .A1(n4267), .A2(n3224), .ZN(n3223) );
  INV_X1 U3749 ( .A(n3226), .ZN(n3224) );
  NAND2_X1 U3750 ( .A1(n3227), .A2(n4216), .ZN(n3226) );
  INV_X1 U3751 ( .A(n4420), .ZN(n3227) );
  INV_X1 U3752 ( .A(n5670), .ZN(n4216) );
  INV_X1 U3753 ( .A(n6057), .ZN(n4164) );
  NAND2_X1 U3754 ( .A1(n4546), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4367) );
  NOR2_X1 U3755 ( .A1(n3999), .A2(n3981), .ZN(n4024) );
  AND2_X1 U3756 ( .A1(n3859), .A2(n4819), .ZN(n3503) );
  INV_X1 U3757 ( .A(n4397), .ZN(n4395) );
  NOR2_X2 U3758 ( .A1(n4805), .A2(n6655), .ZN(n4087) );
  AND2_X1 U3759 ( .A1(n5797), .A2(n3669), .ZN(n3670) );
  INV_X1 U3760 ( .A(n3628), .ZN(n3625) );
  NAND2_X1 U3761 ( .A1(n3778), .A2(EBX_REG_2__SCAN_IN), .ZN(n3184) );
  OR2_X1 U3762 ( .A1(n3436), .A2(n3435), .ZN(n3437) );
  AOI21_X1 U3763 ( .B1(n3415), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3419), 
        .ZN(n3422) );
  INV_X1 U3764 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6625) );
  NOR2_X1 U3765 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4782), .ZN(n5264) );
  NOR2_X1 U3766 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4397) );
  AND2_X1 U3767 ( .A1(n3828), .A2(n3827), .ZN(n5554) );
  NOR2_X2 U3768 ( .A1(n5082), .A2(n5081), .ZN(n5226) );
  NAND2_X1 U3769 ( .A1(n3737), .A2(n3736), .ZN(n5597) );
  NAND3_X1 U3770 ( .A1(n3734), .A2(n3733), .A3(n3732), .ZN(n3737) );
  OR2_X1 U3771 ( .A1(n4563), .A2(n5599), .ZN(n4515) );
  NOR2_X1 U3772 ( .A1(n4346), .A2(n5568), .ZN(n4347) );
  NAND2_X1 U3773 ( .A1(n4347), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4411)
         );
  NAND2_X1 U3774 ( .A1(n4246), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4285)
         );
  INV_X1 U3775 ( .A(n4196), .ZN(n4197) );
  NAND2_X1 U3776 ( .A1(n4198), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4245)
         );
  NOR2_X1 U3777 ( .A1(n3952), .A2(n6263), .ZN(n3951) );
  NAND2_X1 U3778 ( .A1(n5597), .A2(n6652), .ZN(n4563) );
  NOR2_X1 U3779 ( .A1(n5678), .A2(n5677), .ZN(n3186) );
  NAND2_X1 U3780 ( .A1(n3186), .A2(n3185), .ZN(n5668) );
  INV_X1 U3781 ( .A(n5665), .ZN(n3185) );
  OR3_X1 U3782 ( .A1(n5215), .A2(n3213), .A3(n3663), .ZN(n3206) );
  OR2_X1 U3783 ( .A1(n3658), .A2(n5357), .ZN(n3661) );
  NAND2_X1 U3784 ( .A1(n3210), .A2(n3209), .ZN(n3208) );
  INV_X1 U3785 ( .A(n3659), .ZN(n3210) );
  AND2_X1 U3786 ( .A1(n3807), .A2(n3806), .ZN(n4976) );
  AND2_X1 U3787 ( .A1(n4429), .A2(n4783), .ZN(n6617) );
  AND2_X1 U3788 ( .A1(n4712), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3761) );
  NAND2_X1 U3789 ( .A1(n4488), .A2(n4478), .ZN(n3179) );
  AND2_X1 U3790 ( .A1(n5248), .A2(n4871), .ZN(n6267) );
  AND2_X1 U3791 ( .A1(n4476), .A2(n4474), .ZN(n6260) );
  XNOR2_X1 U3792 ( .A(n4473), .B(n4472), .ZN(n5839) );
  AOI21_X1 U3793 ( .B1(n4501), .B2(n5617), .A(n4505), .ZN(n4473) );
  AND2_X1 U3794 ( .A1(n6314), .A2(n4677), .ZN(n6310) );
  AND2_X1 U3795 ( .A1(n6314), .A2(n4678), .ZN(n6307) );
  NAND2_X1 U3796 ( .A1(n5619), .A2(n4490), .ZN(n4405) );
  INV_X1 U3797 ( .A(n6111), .ZN(n6374) );
  OR2_X1 U3798 ( .A1(n4563), .A2(n6607), .ZN(n6164) );
  XNOR2_X1 U3799 ( .A(n3677), .B(n3676), .ZN(n4418) );
  NAND2_X1 U3800 ( .A1(n5762), .A2(n3675), .ZN(n3677) );
  AND2_X1 U3801 ( .A1(n3872), .A2(n3771), .ZN(n6454) );
  CLKBUF_X1 U3802 ( .A(n3920), .Z(n5964) );
  OR2_X1 U3803 ( .A1(n3680), .A2(n3683), .ZN(n3701) );
  AND2_X1 U3804 ( .A1(n3701), .A2(n3700), .ZN(n3703) );
  NAND2_X1 U3805 ( .A1(n3695), .A2(n3694), .ZN(n3731) );
  CLKBUF_X1 U3806 ( .A(n3546), .Z(n3476) );
  NAND2_X1 U3807 ( .A1(n3612), .A2(n3242), .ZN(n3628) );
  OR2_X1 U3808 ( .A1(n3598), .A2(n3597), .ZN(n3630) );
  OR2_X1 U3809 ( .A1(n3557), .A2(n3556), .ZN(n3582) );
  OAI21_X1 U3810 ( .B1(n3381), .B2(n4783), .A(n3859), .ZN(n3397) );
  AOI22_X1 U3811 ( .A1(n4217), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U3812 ( .A1(n3288), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3348), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U3813 ( .A1(n3459), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3255) );
  AOI22_X1 U3814 ( .A1(n4384), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3546), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3246) );
  AND2_X1 U3815 ( .A1(n4540), .A2(n4874), .ZN(n4428) );
  OR2_X1 U3816 ( .A1(n3725), .A2(n3724), .ZN(n3753) );
  NAND3_X1 U3817 ( .A1(n3410), .A2(n3409), .A3(n3408), .ZN(n3474) );
  INV_X1 U3818 ( .A(n3731), .ZN(n3735) );
  NAND2_X1 U3819 ( .A1(n3544), .A2(n3543), .ZN(n3730) );
  OR2_X1 U3820 ( .A1(n4261), .A2(n4260), .ZN(n4268) );
  NOR2_X1 U3821 ( .A1(n4245), .A2(n5772), .ZN(n4246) );
  INV_X1 U3822 ( .A(n6106), .ZN(n3219) );
  AND2_X1 U3823 ( .A1(n4112), .A2(n4095), .ZN(n3220) );
  INV_X1 U3824 ( .A(n5704), .ZN(n4112) );
  INV_X1 U3825 ( .A(n5223), .ZN(n3228) );
  INV_X1 U3826 ( .A(n5079), .ZN(n3997) );
  AND2_X1 U3827 ( .A1(n4767), .A2(n4838), .ZN(n3958) );
  AND2_X1 U3828 ( .A1(n4678), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3932) );
  NAND2_X1 U3829 ( .A1(n3694), .A2(n4492), .ZN(n3650) );
  INV_X1 U3830 ( .A(n4449), .ZN(n4462) );
  INV_X1 U3831 ( .A(n4438), .ZN(n4453) );
  NAND2_X1 U3832 ( .A1(n5685), .A2(n4465), .ZN(n4449) );
  INV_X1 U3833 ( .A(n3385), .ZN(n3399) );
  AOI21_X1 U3834 ( .B1(n3415), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3411), 
        .ZN(n3413) );
  AND2_X1 U3835 ( .A1(n3739), .A2(n3859), .ZN(n4429) );
  OR2_X1 U3836 ( .A1(n3741), .A2(n3738), .ZN(n6613) );
  NOR2_X1 U3837 ( .A1(n4819), .A2(n4832), .ZN(n4493) );
  NAND2_X1 U3838 ( .A1(n3332), .A2(n3331), .ZN(n3333) );
  AOI22_X1 U3839 ( .A1(n4380), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3265) );
  AOI22_X1 U3840 ( .A1(n3569), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U3841 ( .A1(n3481), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3348), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3259) );
  AOI22_X1 U3842 ( .A1(n4384), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3260) );
  AOI22_X1 U3843 ( .A1(n4217), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3258) );
  AOI22_X1 U3844 ( .A1(n3288), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3348), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3319) );
  AND2_X1 U3845 ( .A1(n6533), .A2(n3418), .ZN(n4996) );
  INV_X1 U3846 ( .A(n4428), .ZN(n5599) );
  NOR2_X1 U3847 ( .A1(n6271), .A2(n4480), .ZN(n6207) );
  INV_X1 U3848 ( .A(n5248), .ZN(n6262) );
  NAND2_X1 U3849 ( .A1(n4455), .A2(EBX_REG_1__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U3850 ( .A1(n4345), .A2(n4344), .B1(n4430), .B2(n5983), .ZN(n5571)
         );
  INV_X1 U3851 ( .A(n6348), .ZN(n4564) );
  AND2_X1 U3852 ( .A1(n6655), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4401) );
  AOI21_X1 U3853 ( .B1(n4400), .B2(n4399), .A(n4398), .ZN(n4490) );
  NAND2_X1 U3854 ( .A1(n4327), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4346)
         );
  AOI21_X1 U3855 ( .B1(n4308), .B2(n4307), .A(n4306), .ZN(n5653) );
  AND2_X1 U3856 ( .A1(n6000), .A2(n4430), .ZN(n4306) );
  AND2_X1 U3857 ( .A1(n4289), .A2(n4288), .ZN(n5627) );
  OR2_X1 U3858 ( .A1(n6017), .A2(n4395), .ZN(n4248) );
  INV_X1 U3859 ( .A(n5669), .ZN(n3225) );
  AND2_X1 U3860 ( .A1(n4200), .A2(n4199), .ZN(n5673) );
  CLKBUF_X1 U3861 ( .A(n5669), .Z(n5676) );
  NOR2_X1 U3862 ( .A1(n4146), .A2(n5794), .ZN(n4147) );
  NAND2_X1 U3863 ( .A1(n4147), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4196)
         );
  CLKBUF_X1 U3864 ( .A(n5680), .Z(n5681) );
  AND2_X1 U3865 ( .A1(n4145), .A2(n4144), .ZN(n5698) );
  AND2_X1 U3866 ( .A1(n4127), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4128)
         );
  CLKBUF_X1 U3867 ( .A(n5695), .Z(n5696) );
  NOR2_X1 U3868 ( .A1(n4061), .A2(n4045), .ZN(n4078) );
  CLKBUF_X1 U3869 ( .A(n5540), .Z(n5541) );
  NAND2_X1 U3870 ( .A1(n4044), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4061)
         );
  NOR2_X1 U3871 ( .A1(n4030), .A2(n4029), .ZN(n4044) );
  NAND2_X1 U3872 ( .A1(n4024), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4030)
         );
  NAND2_X1 U3873 ( .A1(n3980), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3999)
         );
  CLKBUF_X1 U3874 ( .A(n4973), .Z(n4974) );
  NOR2_X1 U3875 ( .A1(n3960), .A2(n3959), .ZN(n3961) );
  NAND2_X1 U3876 ( .A1(n3951), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3960)
         );
  NAND2_X1 U3877 ( .A1(n3956), .A2(n3955), .ZN(n4758) );
  CLKBUF_X1 U3878 ( .A(n4756), .Z(n4757) );
  INV_X1 U3879 ( .A(n3933), .ZN(n3940) );
  NAND2_X1 U3880 ( .A1(n3940), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3952)
         );
  NAND2_X1 U3881 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3933) );
  AOI21_X1 U3882 ( .B1(n3404), .B2(n4727), .A(n6655), .ZN(n4584) );
  NAND2_X1 U3883 ( .A1(n3155), .A2(n6115), .ZN(n3900) );
  NOR2_X1 U3884 ( .A1(n5651), .A2(n3176), .ZN(n3175) );
  INV_X1 U3885 ( .A(n5577), .ZN(n3176) );
  AND2_X1 U3886 ( .A1(n5655), .A2(n4452), .ZN(n5649) );
  OR2_X1 U3887 ( .A1(n3658), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5755)
         );
  NOR2_X1 U3888 ( .A1(n5668), .A2(n3853), .ZN(n5661) );
  NAND2_X1 U3889 ( .A1(n5661), .A2(n5660), .ZN(n5663) );
  NOR2_X1 U3890 ( .A1(n5761), .A2(n3194), .ZN(n3191) );
  NAND2_X1 U3891 ( .A1(n3216), .A2(n3214), .ZN(n3674) );
  NOR2_X1 U3892 ( .A1(n3166), .A2(n3215), .ZN(n3214) );
  INV_X1 U3893 ( .A(n3667), .ZN(n3215) );
  NOR2_X1 U3894 ( .A1(n3658), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5769)
         );
  NAND2_X1 U3895 ( .A1(n5505), .A2(n3169), .ZN(n5700) );
  AND2_X1 U3896 ( .A1(n3831), .A2(n3830), .ZN(n5699) );
  AND2_X1 U3897 ( .A1(n6101), .A2(n6099), .ZN(n5798) );
  AND2_X1 U3898 ( .A1(n5505), .A2(n5548), .ZN(n5555) );
  INV_X1 U3899 ( .A(n3168), .ZN(n3202) );
  NAND2_X1 U3900 ( .A1(n3205), .A2(n3212), .ZN(n3203) );
  NOR2_X1 U3901 ( .A1(n4959), .A2(n4976), .ZN(n3180) );
  OR2_X1 U3902 ( .A1(n6732), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4406) );
  INV_X1 U3903 ( .A(n5847), .ZN(n5939) );
  INV_X1 U3904 ( .A(n3608), .ZN(n3201) );
  NAND2_X1 U3905 ( .A1(n3181), .A2(n3803), .ZN(n4977) );
  NOR2_X2 U3906 ( .A1(n3174), .A2(n3796), .ZN(n4843) );
  NAND2_X1 U3907 ( .A1(n3785), .A2(n3182), .ZN(n4768) );
  OAI21_X1 U3908 ( .B1(n4438), .B2(EBX_REG_2__SCAN_IN), .A(n3184), .ZN(n3183)
         );
  INV_X1 U3909 ( .A(n6375), .ZN(n3535) );
  NAND2_X1 U3910 ( .A1(n3872), .A2(n5593), .ZN(n6453) );
  AND2_X1 U3911 ( .A1(n5685), .A2(n4455), .ZN(n4581) );
  NAND2_X1 U3912 ( .A1(n3516), .A2(n3515), .ZN(n4587) );
  XNOR2_X1 U3913 ( .A(n3187), .B(n3438), .ZN(n3500) );
  NAND2_X1 U3914 ( .A1(n3218), .A2(n3188), .ZN(n3187) );
  NAND2_X1 U3915 ( .A1(n3437), .A2(n3495), .ZN(n3188) );
  NAND2_X1 U3916 ( .A1(n3189), .A2(n3498), .ZN(n3499) );
  NAND2_X1 U3917 ( .A1(n3497), .A2(n3522), .ZN(n3189) );
  NAND2_X1 U3918 ( .A1(n3499), .A2(n3500), .ZN(n3560) );
  INV_X1 U3919 ( .A(n6613), .ZN(n4546) );
  NAND2_X1 U3920 ( .A1(n3739), .A2(n5596), .ZN(n4542) );
  AND3_X1 U3921 ( .A1(n4530), .A2(n4529), .A3(n4528), .ZN(n4708) );
  OR2_X1 U3922 ( .A1(n4776), .A2(n4895), .ZN(n5365) );
  OR2_X1 U3923 ( .A1(n6539), .A2(n5964), .ZN(n4804) );
  NAND2_X1 U3924 ( .A1(n4798), .A2(n4776), .ZN(n6539) );
  INV_X1 U3925 ( .A(n5964), .ZN(n5175) );
  NOR2_X1 U3926 ( .A1(n6719), .A2(n4782), .ZN(n4833) );
  NOR2_X1 U3927 ( .A1(n5176), .A2(n5964), .ZN(n4904) );
  INV_X1 U3928 ( .A(n6542), .ZN(n5180) );
  INV_X1 U3929 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4712) );
  OR2_X1 U3930 ( .A1(n3769), .A2(n3768), .ZN(n6607) );
  INV_X1 U3932 ( .A(n6180), .ZN(n6043) );
  INV_X1 U3933 ( .A(n6230), .ZN(n6279) );
  INV_X1 U3934 ( .A(n6265), .ZN(n6249) );
  AND2_X1 U3935 ( .A1(n4965), .A2(n4877), .ZN(n6282) );
  OR2_X1 U3936 ( .A1(n5844), .A2(n6293), .ZN(n4508) );
  INV_X1 U3937 ( .A(n6293), .ZN(n6065) );
  NAND2_X1 U3938 ( .A1(n4674), .A2(n4673), .ZN(n6314) );
  OAI21_X1 U3939 ( .B1(n4672), .B2(n4671), .A(n6652), .ZN(n4673) );
  INV_X1 U3941 ( .A(n4610), .ZN(n4650) );
  XNOR2_X1 U3942 ( .A(n4413), .B(n4412), .ZN(n4870) );
  OR2_X1 U3943 ( .A1(n4411), .A2(n5733), .ZN(n4413) );
  INV_X1 U3944 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5772) );
  OR2_X1 U3945 ( .A1(n5877), .A2(n5866), .ZN(n5856) );
  INV_X1 U3946 ( .A(n3186), .ZN(n5666) );
  AND2_X1 U3947 ( .A1(n3662), .A2(n3206), .ZN(n3211) );
  NAND2_X1 U3948 ( .A1(n5298), .A2(n5297), .ZN(n5356) );
  NAND2_X1 U3949 ( .A1(n6358), .A2(n3608), .ZN(n4940) );
  INV_X1 U3950 ( .A(n6454), .ZN(n6138) );
  INV_X1 U3951 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5407) );
  CLKBUF_X1 U3952 ( .A(n4536), .Z(n4537) );
  NAND2_X1 U3953 ( .A1(n3538), .A2(n3424), .ZN(n4591) );
  NAND2_X1 U3954 ( .A1(n6722), .A2(n4712), .ZN(n6732) );
  OAI21_X1 U3955 ( .B1(n5414), .B2(n5413), .A(n5412), .ZN(n5445) );
  OR3_X1 U3956 ( .A1(n6476), .A2(n6475), .A3(n6474), .ZN(n6510) );
  OR2_X1 U3957 ( .A1(n4804), .A2(n4727), .ZN(n5039) );
  INV_X1 U3958 ( .A(n6563), .ZN(n5424) );
  INV_X1 U3959 ( .A(n6577), .ZN(n5428) );
  INV_X1 U3960 ( .A(n6584), .ZN(n5440) );
  OAI211_X1 U3961 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6655), .A(n5320), .B(n5038), .ZN(n5061) );
  AOI21_X1 U3962 ( .B1(n5037), .B2(n6541), .A(n5035), .ZN(n5067) );
  INV_X1 U3963 ( .A(n6601), .ZN(n5420) );
  OR3_X1 U3964 ( .A1(n6539), .A2(n5175), .A3(n4727), .ZN(n6605) );
  NOR2_X1 U3965 ( .A1(n6847), .A2(n4993), .ZN(n6549) );
  NOR2_X1 U3966 ( .A1(n7029), .A2(n4993), .ZN(n6556) );
  NOR2_X1 U3967 ( .A1(n6862), .A2(n4993), .ZN(n6570) );
  NOR2_X1 U3968 ( .A1(n7095), .A2(n4993), .ZN(n6577) );
  NOR2_X1 U3969 ( .A1(n4869), .A2(n4993), .ZN(n6591) );
  NOR2_X2 U3970 ( .A1(n5185), .A2(n5415), .ZN(n5493) );
  AND2_X1 U3971 ( .A1(n6644), .A2(n6643), .ZN(n6661) );
  INV_X1 U3972 ( .A(n6661), .ZN(n6720) );
  OAI21_X1 U3973 ( .B1(n5839), .B2(n6286), .A(n3177), .ZN(U2796) );
  AOI21_X1 U3974 ( .B1(n5584), .B2(n6244), .A(n3178), .ZN(n3177) );
  OAI211_X1 U3975 ( .C1(n6384), .C2(n5573), .A(n5572), .B(n3160), .ZN(n5574)
         );
  OAI21_X1 U3976 ( .B1(n6019), .B2(n6108), .A(n4424), .ZN(n4425) );
  OAI21_X1 U3977 ( .B1(n3890), .B2(n6405), .A(n3889), .ZN(n3891) );
  AND2_X2 U3978 ( .A1(n4545), .A2(n4691), .ZN(n3350) );
  OR2_X1 U3979 ( .A1(n6101), .A2(n5942), .ZN(n3156) );
  NAND2_X1 U3980 ( .A1(n4096), .A2(n4095), .ZN(n5552) );
  NAND2_X1 U3981 ( .A1(n3225), .A2(n4216), .ZN(n4419) );
  INV_X2 U3982 ( .A(n3365), .ZN(n3398) );
  INV_X1 U3983 ( .A(n3437), .ZN(n3561) );
  AND2_X1 U3984 ( .A1(n3167), .A2(n5242), .ZN(n3157) );
  AND2_X1 U3985 ( .A1(n3998), .A2(n3167), .ZN(n5222) );
  INV_X1 U3986 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3939) );
  AND2_X2 U3987 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4545) );
  OR2_X1 U3988 ( .A1(n5663), .A2(n5636), .ZN(n3158) );
  INV_X1 U3989 ( .A(n3658), .ZN(n6100) );
  NAND2_X1 U3990 ( .A1(n3216), .A2(n3667), .ZN(n5789) );
  AND2_X1 U3991 ( .A1(n3636), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3159)
         );
  AND2_X1 U3992 ( .A1(n3366), .A2(n3383), .ZN(n3404) );
  OR2_X1 U3993 ( .A1(n5576), .A2(n6108), .ZN(n3160) );
  AND2_X1 U3994 ( .A1(n3377), .A2(n3376), .ZN(n3408) );
  AND4_X1 U3995 ( .A1(n3317), .A2(n3316), .A3(n3315), .A4(n3314), .ZN(n3161)
         );
  INV_X1 U3996 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4601) );
  NAND2_X1 U3997 ( .A1(n4096), .A2(n3220), .ZN(n5702) );
  AND2_X1 U3998 ( .A1(n3311), .A2(n3240), .ZN(n3162) );
  NAND2_X1 U3999 ( .A1(n3365), .A2(n4805), .ZN(n3382) );
  AND2_X1 U4000 ( .A1(n6101), .A2(n3869), .ZN(n3163) );
  XNOR2_X1 U4001 ( .A(n3601), .B(n3610), .ZN(n3905) );
  OR2_X1 U4002 ( .A1(n5669), .A2(n3226), .ZN(n3164) );
  OR2_X1 U4003 ( .A1(n5789), .A2(n5798), .ZN(n3165) );
  INV_X1 U4004 ( .A(n4959), .ZN(n3803) );
  NAND2_X1 U4005 ( .A1(n3382), .A2(n3399), .ZN(n3740) );
  OR2_X1 U4006 ( .A1(n5798), .A2(n3163), .ZN(n3166) );
  INV_X1 U4007 ( .A(n3212), .ZN(n3209) );
  OR2_X1 U4008 ( .A1(n3663), .A2(n3213), .ZN(n3212) );
  INV_X1 U4009 ( .A(n4832), .ZN(n3313) );
  OR2_X1 U4010 ( .A1(n5647), .A2(n3231), .ZN(n5618) );
  INV_X1 U4011 ( .A(n3926), .ZN(n4161) );
  BUF_X1 U4012 ( .A(n3459), .Z(n3460) );
  AND2_X1 U4013 ( .A1(n3998), .A2(n3157), .ZN(n5240) );
  NAND2_X1 U4014 ( .A1(n5248), .A2(n4434), .ZN(n6192) );
  NAND2_X1 U4015 ( .A1(n3998), .A2(n3997), .ZN(n5078) );
  NAND2_X1 U4016 ( .A1(n3659), .A2(n5215), .ZN(n5298) );
  NAND2_X1 U4017 ( .A1(n3208), .A2(n3211), .ZN(n5520) );
  AND2_X1 U4018 ( .A1(n3997), .A2(n3228), .ZN(n3167) );
  AND2_X1 U4019 ( .A1(n6101), .A2(n5534), .ZN(n3168) );
  OR2_X1 U4020 ( .A1(n3385), .A2(n6656), .ZN(n3543) );
  INV_X1 U4021 ( .A(n3543), .ZN(n3495) );
  AND2_X1 U4022 ( .A1(n5548), .A2(n5554), .ZN(n3169) );
  INV_X1 U4023 ( .A(n3194), .ZN(n3193) );
  NOR2_X1 U4024 ( .A1(n6100), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3194)
         );
  AND2_X1 U4025 ( .A1(n5778), .A2(n5769), .ZN(n3170) );
  AND2_X1 U4026 ( .A1(n3157), .A2(n5258), .ZN(n3171) );
  INV_X1 U4027 ( .A(n3833), .ZN(n5685) );
  NOR2_X1 U4028 ( .A1(n5244), .A2(n5245), .ZN(n5243) );
  NAND2_X1 U4029 ( .A1(n4843), .A2(n4842), .ZN(n4841) );
  NOR3_X1 U4030 ( .A1(n3863), .A2(n3862), .A3(n3861), .ZN(n3172) );
  AND2_X1 U4031 ( .A1(n5243), .A2(n3235), .ZN(n5505) );
  AND2_X1 U4032 ( .A1(n3219), .A2(n3220), .ZN(n3173) );
  INV_X1 U4033 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6656) );
  INV_X2 U4034 ( .A(n6108), .ZN(n6378) );
  AND2_X1 U4035 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4695) );
  INV_X1 U4036 ( .A(n3174), .ZN(n4793) );
  NAND2_X1 U4037 ( .A1(n4771), .A2(n3174), .ZN(n6438) );
  XNOR2_X1 U4038 ( .A(n3174), .B(n4792), .ZN(n6430) );
  NAND2_X1 U4039 ( .A1(n4764), .A2(n3789), .ZN(n3174) );
  NOR2_X4 U4040 ( .A1(n3158), .A2(n5654), .ZN(n5655) );
  NAND2_X2 U4041 ( .A1(n5655), .A2(n3175), .ZN(n4469) );
  NOR2_X2 U4042 ( .A1(n4469), .A2(n4468), .ZN(n4496) );
  NAND3_X1 U4043 ( .A1(n4489), .A2(n4477), .A3(n3179), .ZN(n3178) );
  OR2_X2 U4044 ( .A1(n5700), .A2(n5699), .ZN(n6132) );
  INV_X1 U4045 ( .A(n3183), .ZN(n3182) );
  NAND2_X2 U4046 ( .A1(n4465), .A2(n3833), .ZN(n4438) );
  INV_X4 U4047 ( .A(n4666), .ZN(n4465) );
  NAND2_X1 U4048 ( .A1(n5777), .A2(n3170), .ZN(n5762) );
  NAND2_X1 U4049 ( .A1(n5776), .A2(n3193), .ZN(n5771) );
  OAI21_X1 U4050 ( .B1(n5776), .B2(n3192), .A(n3190), .ZN(n5763) );
  NAND2_X1 U4051 ( .A1(n5776), .A2(n3191), .ZN(n3190) );
  NAND2_X1 U4052 ( .A1(n5769), .A2(n3676), .ZN(n3192) );
  OAI21_X1 U4053 ( .B1(n6358), .B2(n3196), .A(n3195), .ZN(n6352) );
  AOI21_X1 U4054 ( .B1(n4939), .B2(n3201), .A(n3159), .ZN(n3195) );
  INV_X1 U4055 ( .A(n4939), .ZN(n3196) );
  NAND2_X1 U4056 ( .A1(n3199), .A2(n3197), .ZN(n6350) );
  INV_X1 U4057 ( .A(n3198), .ZN(n3197) );
  OAI21_X1 U4058 ( .B1(n4939), .B2(n3159), .A(n6351), .ZN(n3198) );
  NAND2_X1 U4059 ( .A1(n6358), .A2(n3200), .ZN(n3199) );
  NOR2_X1 U4060 ( .A1(n3159), .A2(n3201), .ZN(n3200) );
  NAND2_X1 U4061 ( .A1(n4940), .A2(n4939), .ZN(n4938) );
  NAND2_X1 U4062 ( .A1(n3659), .A2(n3205), .ZN(n3204) );
  NAND3_X1 U4063 ( .A1(n3204), .A2(n3203), .A3(n3202), .ZN(n5818) );
  NAND3_X1 U4064 ( .A1(n3538), .A2(n6656), .A3(n3424), .ZN(n3218) );
  NAND2_X1 U4065 ( .A1(n3222), .A2(n3221), .ZN(n3601) );
  NOR2_X2 U4066 ( .A1(n5669), .A2(n3223), .ZN(n5628) );
  NOR2_X1 U4067 ( .A1(n5647), .A2(n5648), .ZN(n5570) );
  NAND2_X1 U4068 ( .A1(n3413), .A2(n3412), .ZN(n3440) );
  AND2_X1 U4069 ( .A1(n4508), .A2(n4507), .ZN(n3234) );
  NAND2_X1 U4070 ( .A1(n6297), .A2(n5582), .ZN(n6293) );
  AND2_X1 U4071 ( .A1(n6297), .A2(n3383), .ZN(n6066) );
  INV_X1 U4072 ( .A(n6297), .ZN(n4506) );
  NAND2_X1 U4073 ( .A1(n3395), .A2(n3394), .ZN(n3473) );
  AND2_X1 U4074 ( .A1(n5503), .A2(n5504), .ZN(n3235) );
  INV_X1 U4075 ( .A(n5243), .ZN(n5259) );
  NAND2_X1 U4076 ( .A1(n3781), .A2(n3780), .ZN(n3783) );
  NOR3_X1 U4077 ( .A1(n4798), .A2(n3502), .A3(n5964), .ZN(n3236) );
  AND4_X1 U4078 ( .A1(n3355), .A2(n3354), .A3(n3353), .A4(n3352), .ZN(n3237)
         );
  AND2_X1 U4079 ( .A1(n4380), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3238) );
  INV_X1 U4080 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6263) );
  INV_X1 U4081 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4097) );
  INV_X1 U4082 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3959) );
  INV_X1 U4083 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3534) );
  OR2_X1 U4084 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6157), .ZN(n7142) );
  XOR2_X1 U4085 ( .A(n3155), .B(n6115), .Z(n3239) );
  AND3_X1 U4086 ( .A1(n3310), .A2(n3309), .A3(n3308), .ZN(n3240) );
  AND4_X1 U4087 ( .A1(n3360), .A2(n3359), .A3(n3358), .A4(n3357), .ZN(n3241)
         );
  AND2_X1 U4088 ( .A1(n3611), .A2(n3610), .ZN(n3242) );
  INV_X1 U4089 ( .A(n3425), .ZN(n4228) );
  OR2_X1 U4090 ( .A1(n3699), .A2(n3698), .ZN(n3711) );
  AOI22_X1 U4091 ( .A1(n3695), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3468), 
        .B2(n3437), .ZN(n3438) );
  INV_X1 U4092 ( .A(n3703), .ZN(n3706) );
  OR2_X1 U4093 ( .A1(n3411), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3371)
         );
  AND2_X1 U4094 ( .A1(n3721), .A2(n3720), .ZN(n3723) );
  NAND2_X1 U4095 ( .A1(n3706), .A2(n3705), .ZN(n3718) );
  NOR2_X1 U4096 ( .A1(n3334), .A2(n3333), .ZN(n3340) );
  INV_X1 U4097 ( .A(n5659), .ZN(n4267) );
  OR2_X1 U4098 ( .A1(n3579), .A2(n3578), .ZN(n3629) );
  OR2_X1 U4099 ( .A1(n3622), .A2(n3621), .ZN(n3642) );
  INV_X1 U4100 ( .A(n3422), .ZN(n3420) );
  INV_X1 U4101 ( .A(n3695), .ZN(n3726) );
  AOI21_X1 U4102 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6630), .A(n3723), 
        .ZN(n3729) );
  NOR2_X1 U4103 ( .A1(n3383), .A2(n6655), .ZN(n3926) );
  OR2_X1 U4104 ( .A1(n6090), .A2(n4395), .ZN(n4288) );
  INV_X1 U4105 ( .A(n5551), .ZN(n4095) );
  INV_X1 U4106 ( .A(n3979), .ZN(n3980) );
  INV_X1 U4107 ( .A(n3932), .ZN(n3950) );
  AND2_X1 U4108 ( .A1(n4448), .A2(n4447), .ZN(n5654) );
  AND2_X1 U4109 ( .A1(n3819), .A2(n3818), .ZN(n5503) );
  NAND2_X1 U4110 ( .A1(n3473), .A2(n3474), .ZN(n3442) );
  NOR2_X1 U4111 ( .A1(n6197), .A2(n6200), .ZN(n6188) );
  INV_X1 U4112 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4029) );
  AND2_X1 U4113 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n4326), .ZN(n4327)
         );
  AND2_X1 U4114 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n4197), .ZN(n4198)
         );
  AND2_X1 U4115 ( .A1(n3155), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5564)
         );
  AND2_X1 U4116 ( .A1(n3852), .A2(n3851), .ZN(n5665) );
  NAND2_X1 U4117 ( .A1(n3640), .A2(n3651), .ZN(n3658) );
  AND2_X1 U4118 ( .A1(n5355), .A2(n3661), .ZN(n3662) );
  AOI21_X1 U4119 ( .B1(n6647), .B2(n4725), .A(n4722), .ZN(n4782) );
  AND2_X1 U4120 ( .A1(n5973), .A2(n5094), .ZN(n5324) );
  AND2_X1 U4121 ( .A1(n4799), .A2(n6537), .ZN(n4801) );
  INV_X1 U4122 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U4123 ( .A1(n3509), .A2(n3508), .ZN(n3510) );
  INV_X1 U4124 ( .A(n5596), .ZN(n4669) );
  NOR2_X1 U4125 ( .A1(n4098), .A2(n4097), .ZN(n4127) );
  OR3_X1 U4126 ( .A1(n6697), .A2(n4480), .A3(n6262), .ZN(n5557) );
  OR2_X1 U4127 ( .A1(n4432), .A2(n6645), .ZN(n4433) );
  AND2_X1 U4128 ( .A1(n4870), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4871) );
  AND2_X1 U4129 ( .A1(n4965), .A2(EBX_REG_31__SCAN_IN), .ZN(n4476) );
  INV_X1 U4130 ( .A(n4490), .ZN(n4491) );
  NOR2_X1 U4131 ( .A1(n4285), .A2(n4284), .ZN(n4286) );
  NAND2_X1 U4132 ( .A1(n4078), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4098)
         );
  OR2_X1 U4133 ( .A1(n5755), .A2(n5865), .ZN(n5739) );
  INV_X1 U4134 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3676) );
  NAND2_X1 U4135 ( .A1(n5947), .A2(n5952), .ZN(n5925) );
  AND2_X1 U4136 ( .A1(n3519), .A2(n3531), .ZN(n4680) );
  NAND2_X1 U4137 ( .A1(n3767), .A2(n3766), .ZN(n3872) );
  NOR2_X1 U4138 ( .A1(n5365), .A2(n5964), .ZN(n5416) );
  OR3_X1 U4139 ( .A1(n5365), .A2(n5175), .A3(n4727), .ZN(n6526) );
  INV_X1 U4140 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6630) );
  NAND2_X1 U4141 ( .A1(n3542), .A2(n3541), .ZN(n4990) );
  AND3_X1 U4142 ( .A1(n4901), .A2(n5180), .A3(n4900), .ZN(n4932) );
  OR2_X1 U4143 ( .A1(n5176), .A2(n5175), .ZN(n5185) );
  AND2_X1 U4144 ( .A1(n5597), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4722) );
  INV_X2 U4145 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6655) );
  AND2_X1 U4146 ( .A1(n4429), .A2(n5590), .ZN(n5598) );
  NAND2_X1 U4147 ( .A1(n4515), .A2(n5981), .ZN(n6741) );
  AND2_X1 U4148 ( .A1(n4481), .A2(n6043), .ZN(n6036) );
  NAND2_X1 U4149 ( .A1(n4128), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4146)
         );
  AND2_X1 U4150 ( .A1(n5248), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6230) );
  INV_X1 U4151 ( .A(n6192), .ZN(n6244) );
  NAND2_X1 U4152 ( .A1(n4965), .A2(n4436), .ZN(n6271) );
  INV_X1 U4153 ( .A(n3383), .ZN(n5582) );
  INV_X1 U4154 ( .A(n6314), .ZN(n6311) );
  NOR2_X1 U4155 ( .A1(n6638), .A2(n4564), .ZN(n6346) );
  INV_X1 U4156 ( .A(n4674), .ZN(n4637) );
  OAI21_X1 U4157 ( .B1(n3685), .B2(n5605), .A(n4513), .ZN(n4559) );
  NAND2_X1 U4158 ( .A1(n4286), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4325)
         );
  NAND2_X1 U4159 ( .A1(n3961), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3979)
         );
  INV_X1 U4160 ( .A(n6384), .ZN(n5808) );
  INV_X1 U4161 ( .A(n6164), .ZN(n6380) );
  NAND2_X1 U4162 ( .A1(n5684), .A2(n3847), .ZN(n5678) );
  NOR2_X1 U4163 ( .A1(n6156), .A2(n5924), .ZN(n6130) );
  OR2_X1 U4164 ( .A1(n5925), .A2(n6450), .ZN(n5847) );
  INV_X1 U4165 ( .A(n6453), .ZN(n6450) );
  INV_X1 U4166 ( .A(n5264), .ZN(n4993) );
  OAI21_X1 U4167 ( .B1(n5266), .B2(n5267), .A(n5265), .ZN(n5289) );
  INV_X1 U4168 ( .A(n5354), .ZN(n5317) );
  OAI221_X1 U4169 ( .B1(n5325), .B2(n6722), .C1(n5325), .C2(n5321), .A(n5320), 
        .ZN(n5347) );
  OAI211_X1 U4170 ( .C1(n6537), .C2(n5102), .A(n5101), .B(n5180), .ZN(n5125)
         );
  INV_X1 U4171 ( .A(n6477), .ZN(n6508) );
  OR2_X1 U4172 ( .A1(n5136), .A2(n5135), .ZN(n5162) );
  NOR2_X1 U4173 ( .A1(n4804), .A2(n5415), .ZN(n5129) );
  INV_X1 U4174 ( .A(n5039), .ZN(n5064) );
  INV_X1 U4175 ( .A(n6605), .ZN(n5029) );
  AND2_X1 U4176 ( .A1(n4904), .A2(n5415), .ZN(n5494) );
  NOR2_X1 U4177 ( .A1(n7036), .A2(n4993), .ZN(n6563) );
  NOR2_X1 U4178 ( .A1(n7085), .A2(n4993), .ZN(n6584) );
  NOR2_X1 U4179 ( .A1(n7042), .A2(n4993), .ZN(n6601) );
  AND2_X1 U4180 ( .A1(n3761), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6652) );
  NAND2_X1 U4181 ( .A1(n5598), .A2(n6652), .ZN(n5981) );
  OR2_X1 U4182 ( .A1(n5617), .A2(n5616), .ZN(n5861) );
  INV_X1 U4183 ( .A(n6282), .ZN(n6054) );
  INV_X1 U4184 ( .A(n6260), .ZN(n6286) );
  AND2_X2 U4185 ( .A1(n4495), .A2(n6652), .ZN(n6297) );
  OR2_X1 U4186 ( .A1(n4563), .A2(n4562), .ZN(n6348) );
  OR2_X1 U4187 ( .A1(n4515), .A2(n4514), .ZN(n4674) );
  INV_X1 U4188 ( .A(n4425), .ZN(n4426) );
  NAND2_X1 U4189 ( .A1(n6164), .A2(n4407), .ZN(n6111) );
  OR2_X1 U4190 ( .A1(n6663), .A2(n6543), .ZN(n6108) );
  OR2_X1 U4191 ( .A1(n4406), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6403) );
  NOR2_X1 U4192 ( .A1(n5955), .A2(n5533), .ZN(n6156) );
  INV_X1 U4193 ( .A(n6448), .ZN(n6405) );
  AND2_X1 U4194 ( .A1(n4723), .A2(n4993), .ZN(n6463) );
  NAND2_X1 U4195 ( .A1(n3236), .A2(n4727), .ZN(n5296) );
  NAND2_X1 U4196 ( .A1(n3236), .A2(n5415), .ZN(n5354) );
  OR2_X1 U4197 ( .A1(n5096), .A2(n4727), .ZN(n5404) );
  NAND3_X1 U4198 ( .A1(n4781), .A2(n4727), .A3(n5964), .ZN(n6532) );
  INV_X1 U4199 ( .A(n5129), .ZN(n5168) );
  INV_X1 U4200 ( .A(n6549), .ZN(n5451) );
  INV_X1 U4201 ( .A(n6556), .ZN(n5432) );
  INV_X1 U4202 ( .A(n6591), .ZN(n5444) );
  OR3_X1 U4203 ( .A1(n6539), .A2(n5415), .A3(n5175), .ZN(n6598) );
  NOR2_X1 U4204 ( .A1(n4995), .A2(n4994), .ZN(n5032) );
  NAND2_X1 U4205 ( .A1(n4904), .A2(n4727), .ZN(n5027) );
  INV_X1 U4206 ( .A(n5459), .ZN(n5498) );
  AOI21_X1 U4207 ( .B1(n5183), .B2(n5184), .A(n5182), .ZN(n5212) );
  AND2_X1 U4208 ( .A1(n6637), .A2(n6636), .ZN(n6651) );
  CLKBUF_X1 U4209 ( .A(n6698), .Z(n6709) );
  INV_X2 U4210 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4211 ( .A1(n4380), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3247) );
  INV_X1 U4212 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4213 ( .A1(n4217), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3245) );
  AOI22_X1 U4214 ( .A1(n3569), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3244) );
  NOR2_X4 U4215 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4544) );
  AND2_X2 U4216 ( .A1(n3248), .A2(n4544), .ZN(n3430) );
  AND2_X2 U4217 ( .A1(n3249), .A2(n4691), .ZN(n3351) );
  AOI22_X1 U4218 ( .A1(n3351), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3254) );
  AND2_X4 U4219 ( .A1(n4692), .A2(n3250), .ZN(n3481) );
  AND2_X2 U4220 ( .A1(n4691), .A2(n4544), .ZN(n3349) );
  AOI22_X1 U4221 ( .A1(n3481), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4222 ( .A1(n3430), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3261) );
  AOI22_X1 U4223 ( .A1(n3545), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3264) );
  AOI22_X1 U4224 ( .A1(n3546), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3262) );
  NAND2_X2 U4225 ( .A1(n3267), .A2(n3266), .ZN(n4805) );
  NAND2_X1 U4226 ( .A1(n4217), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3271) );
  NAND2_X1 U4227 ( .A1(n4380), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3270) );
  NAND2_X1 U4228 ( .A1(n3545), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3269) );
  NAND2_X1 U4229 ( .A1(n3289), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3268) );
  NAND2_X1 U4230 ( .A1(n4384), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3275)
         );
  NAND2_X1 U4231 ( .A1(n3569), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3274) );
  NAND2_X1 U4232 ( .A1(n3546), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3273)
         );
  NAND2_X1 U4233 ( .A1(n3356), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3272)
         );
  NAND2_X1 U4234 ( .A1(n3288), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3279) );
  NAND2_X1 U4235 ( .A1(n3351), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3278) );
  NAND2_X1 U4236 ( .A1(n3348), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3277)
         );
  NAND2_X1 U4237 ( .A1(n3350), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3276) );
  NAND2_X1 U4238 ( .A1(n3459), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3283)
         );
  NAND2_X1 U4239 ( .A1(n3430), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3282) );
  NAND2_X1 U4240 ( .A1(n3481), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3281)
         );
  NAND2_X1 U4241 ( .A1(n3349), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U4242 ( .A1(n4380), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3293) );
  AOI22_X1 U4243 ( .A1(n4384), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U4244 ( .A1(n3288), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4245 ( .A1(n3546), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3290) );
  NAND4_X1 U4246 ( .A1(n3293), .A2(n3292), .A3(n3291), .A4(n3290), .ZN(n3303)
         );
  INV_X1 U4247 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3296) );
  INV_X1 U4248 ( .A(n3348), .ZN(n3295) );
  INV_X1 U4249 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3294) );
  INV_X1 U4250 ( .A(n3297), .ZN(n3301) );
  AOI22_X1 U4251 ( .A1(n3459), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4252 ( .A1(n3430), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4253 ( .A1(n3481), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3298) );
  NAND4_X1 U4254 ( .A1(n3301), .A2(n3300), .A3(n3299), .A4(n3298), .ZN(n3302)
         );
  AOI22_X1 U4255 ( .A1(n3459), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U4256 ( .A1(n3481), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4257 ( .A1(n3288), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3348), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3305) );
  AOI22_X1 U4258 ( .A1(n3351), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3304) );
  AOI22_X1 U4259 ( .A1(n4217), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4260 ( .A1(n4380), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4261 ( .A1(n4384), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3546), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4262 ( .A1(n3569), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3308) );
  NAND2_X1 U4263 ( .A1(n3313), .A2(n4819), .ZN(n3323) );
  AOI22_X1 U4264 ( .A1(n4217), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4265 ( .A1(n4384), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3546), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4266 ( .A1(n4380), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4267 ( .A1(n3569), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4268 ( .A1(n3459), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3321) );
  AOI22_X1 U4269 ( .A1(n3481), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4270 ( .A1(n3351), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3318) );
  NAND2_X1 U4271 ( .A1(n3365), .A2(n3383), .ZN(n4676) );
  NOR2_X1 U4272 ( .A1(n3323), .A2(n4676), .ZN(n3324) );
  NAND2_X1 U4273 ( .A1(n3351), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3328) );
  NAND2_X1 U4274 ( .A1(n4217), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3327) );
  NAND2_X1 U4275 ( .A1(n3569), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3326) );
  NAND2_X1 U4276 ( .A1(n3545), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3325) );
  NAND2_X1 U4277 ( .A1(n3289), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3330) );
  NAND2_X1 U4278 ( .A1(n3349), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3329) );
  NAND2_X1 U4279 ( .A1(n3330), .A2(n3329), .ZN(n3334) );
  NAND2_X1 U4280 ( .A1(n3546), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3332)
         );
  NAND2_X1 U4281 ( .A1(n3356), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3331)
         );
  NAND2_X1 U4282 ( .A1(n3481), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3337)
         );
  NAND2_X1 U4283 ( .A1(n3459), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3336)
         );
  NAND2_X1 U4284 ( .A1(n3350), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3335) );
  NAND3_X1 U4285 ( .A1(n3337), .A2(n3336), .A3(n3335), .ZN(n3338) );
  NOR2_X1 U4286 ( .A1(n3238), .A2(n3338), .ZN(n3339) );
  AND3_X2 U4287 ( .A1(n3341), .A2(n3340), .A3(n3339), .ZN(n3347) );
  NAND2_X1 U4288 ( .A1(n4384), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3345)
         );
  NAND2_X1 U4289 ( .A1(n3430), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3344) );
  NAND2_X1 U4290 ( .A1(n3288), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3343) );
  NAND2_X1 U4291 ( .A1(n3348), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3342)
         );
  AOI22_X1 U4292 ( .A1(n3288), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3348), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4293 ( .A1(n3481), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4294 ( .A1(n3459), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4295 ( .A1(n3351), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3352) );
  AOI22_X1 U4296 ( .A1(n4384), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3546), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4297 ( .A1(n4380), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4298 ( .A1(n3569), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3357) );
  NAND2_X2 U4299 ( .A1(n3237), .A2(n3241), .ZN(n3380) );
  XNOR2_X1 U4300 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n3750) );
  NAND2_X1 U4301 ( .A1(n3685), .A2(n3750), .ZN(n3378) );
  AND2_X2 U4302 ( .A1(n3859), .A2(n3685), .ZN(n5596) );
  NAND3_X1 U4303 ( .A1(n5596), .A2(n4493), .A3(n3365), .ZN(n4538) );
  NAND2_X1 U4304 ( .A1(n4805), .A2(n3383), .ZN(n3858) );
  NOR2_X1 U4305 ( .A1(n4538), .A2(n3858), .ZN(n3854) );
  AOI21_X1 U4306 ( .B1(n4428), .B2(n3378), .A(n3854), .ZN(n3368) );
  INV_X1 U4307 ( .A(n4805), .ZN(n3366) );
  NOR2_X1 U4308 ( .A1(n3740), .A2(n3404), .ZN(n3364) );
  OAI21_X1 U4309 ( .B1(n3399), .B2(n4805), .A(n3382), .ZN(n3361) );
  OAI21_X1 U4310 ( .B1(n3361), .B2(n4832), .A(n3383), .ZN(n3362) );
  INV_X1 U4311 ( .A(n3362), .ZN(n3363) );
  OAI21_X1 U4312 ( .B1(n3364), .B2(n3313), .A(n3363), .ZN(n3381) );
  NAND2_X1 U4313 ( .A1(n3741), .A2(n4819), .ZN(n3405) );
  NAND2_X1 U4314 ( .A1(n3399), .A2(n3398), .ZN(n3768) );
  INV_X1 U4315 ( .A(n3768), .ZN(n3373) );
  NAND2_X1 U4316 ( .A1(n3405), .A2(n3373), .ZN(n3367) );
  NOR2_X1 U4317 ( .A1(n3381), .A2(n3367), .ZN(n3739) );
  NAND2_X1 U4318 ( .A1(n3368), .A2(n4542), .ZN(n3369) );
  NAND2_X1 U4319 ( .A1(n3369), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3412) );
  INV_X1 U4320 ( .A(n3412), .ZN(n3372) );
  XNOR2_X1 U4321 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5322) );
  OAI22_X1 U4322 ( .A1(n4406), .A2(n5322), .B1(n3761), .B2(n5370), .ZN(n3411)
         );
  NAND2_X1 U4323 ( .A1(n3372), .A2(n3371), .ZN(n3439) );
  AND2_X4 U4324 ( .A1(n4819), .A2(n3380), .ZN(n3833) );
  NAND2_X1 U4325 ( .A1(n3373), .A2(n3833), .ZN(n3377) );
  INV_X1 U4326 ( .A(n3740), .ZN(n3374) );
  NAND2_X1 U4327 ( .A1(n3374), .A2(n3383), .ZN(n3375) );
  NAND2_X1 U4328 ( .A1(n3375), .A2(n3512), .ZN(n3376) );
  AOI21_X1 U4329 ( .B1(n3378), .B2(n3365), .A(n4832), .ZN(n3379) );
  BUF_X4 U4330 ( .A(n3380), .Z(n4783) );
  AND2_X1 U4331 ( .A1(n4819), .A2(n3383), .ZN(n3384) );
  AND2_X1 U4332 ( .A1(n3382), .A2(n3384), .ZN(n3387) );
  NAND2_X1 U4333 ( .A1(n3387), .A2(n3386), .ZN(n3745) );
  AND2_X1 U4334 ( .A1(n3741), .A2(n3385), .ZN(n3388) );
  NAND3_X1 U4335 ( .A1(n3389), .A2(n3397), .A3(n3403), .ZN(n3390) );
  NAND2_X1 U4336 ( .A1(n3415), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3395) );
  INV_X1 U4337 ( .A(n3761), .ZN(n3392) );
  INV_X1 U4338 ( .A(n4406), .ZN(n3391) );
  MUX2_X1 U4339 ( .A(n3392), .B(n3391), .S(n5407), .Z(n3393) );
  INV_X1 U4340 ( .A(n3393), .ZN(n3394) );
  NAND2_X1 U4341 ( .A1(n3503), .A2(n3741), .ZN(n3396) );
  NAND2_X1 U4342 ( .A1(n3397), .A2(n3396), .ZN(n3400) );
  NAND2_X1 U4343 ( .A1(n3400), .A2(n3650), .ZN(n3402) );
  NAND2_X1 U4344 ( .A1(n4832), .A2(n4874), .ZN(n3401) );
  NAND2_X1 U4345 ( .A1(n3402), .A2(n3401), .ZN(n3863) );
  INV_X1 U4346 ( .A(n3863), .ZN(n3410) );
  NOR2_X1 U4347 ( .A1(n6732), .A2(n6656), .ZN(n6653) );
  NAND3_X1 U4348 ( .A1(n3404), .A2(n4493), .A3(n3385), .ZN(n4698) );
  NAND2_X1 U4349 ( .A1(n3405), .A2(n3512), .ZN(n3406) );
  NAND2_X1 U4350 ( .A1(n3439), .A2(n3442), .ZN(n3414) );
  NAND2_X1 U4351 ( .A1(n3414), .A2(n3440), .ZN(n3423) );
  INV_X1 U4352 ( .A(n3423), .ZN(n3421) );
  AND2_X1 U4353 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3416) );
  NAND2_X1 U4354 ( .A1(n3416), .A2(n6625), .ZN(n6533) );
  INV_X1 U4355 ( .A(n3416), .ZN(n3417) );
  NAND2_X1 U4356 ( .A1(n3417), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3418) );
  OAI22_X1 U4357 ( .A1(n4996), .A2(n4406), .B1(n3761), .B2(n6625), .ZN(n3419)
         );
  NAND2_X2 U4358 ( .A1(n3421), .A2(n3420), .ZN(n3538) );
  NAND2_X1 U4359 ( .A1(n3423), .A2(n3422), .ZN(n3424) );
  AOI22_X1 U4360 ( .A1(n4229), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4361 ( .A1(n4384), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4362 ( .A1(n4228), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3427) );
  INV_X1 U4363 ( .A(n3356), .ZN(n3447) );
  INV_X2 U4364 ( .A(n3447), .ZN(n4383) );
  AOI22_X1 U4365 ( .A1(n4694), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3426) );
  NAND4_X1 U4366 ( .A1(n3429), .A2(n3428), .A3(n3427), .A4(n3426), .ZN(n3436)
         );
  AOI22_X1 U4367 ( .A1(n3460), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3434) );
  AOI22_X1 U4368 ( .A1(n3461), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3433) );
  AOI22_X1 U4369 ( .A1(n4234), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3432) );
  AOI22_X1 U4370 ( .A1(n4356), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3431) );
  NAND4_X1 U4371 ( .A1(n3434), .A2(n3433), .A3(n3432), .A4(n3431), .ZN(n3435)
         );
  NAND2_X1 U4372 ( .A1(n3859), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3544) );
  INV_X1 U4373 ( .A(n3544), .ZN(n3468) );
  NAND2_X1 U4374 ( .A1(n3440), .A2(n3439), .ZN(n3441) );
  XNOR2_X1 U4375 ( .A(n3442), .B(n3441), .ZN(n4536) );
  AOI22_X1 U4376 ( .A1(n4380), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3446) );
  AOI22_X1 U4377 ( .A1(n3460), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3445) );
  AOI22_X1 U4378 ( .A1(n3545), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4379 ( .A1(n4374), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3443) );
  NAND4_X1 U4380 ( .A1(n3446), .A2(n3445), .A3(n3444), .A4(n3443), .ZN(n3453)
         );
  AOI22_X1 U4381 ( .A1(n4351), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4228), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4382 ( .A1(n4234), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4383 ( .A1(n3546), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4384 ( .A1(n4694), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3448) );
  NAND4_X1 U4385 ( .A1(n3451), .A2(n3450), .A3(n3449), .A4(n3448), .ZN(n3452)
         );
  NAND2_X1 U4386 ( .A1(n3495), .A2(n3525), .ZN(n3454) );
  OAI21_X2 U4387 ( .B1(n4536), .B2(STATE2_REG_0__SCAN_IN), .A(n3454), .ZN(
        n3521) );
  INV_X1 U4388 ( .A(n3521), .ZN(n3472) );
  AOI22_X1 U4389 ( .A1(n4372), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4228), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3458) );
  AOI22_X1 U4390 ( .A1(n4351), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3457) );
  AOI22_X1 U4391 ( .A1(n4229), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4234), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3456) );
  AOI22_X1 U4392 ( .A1(n4694), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3455) );
  NAND4_X1 U4393 ( .A1(n3458), .A2(n3457), .A3(n3456), .A4(n3455), .ZN(n3467)
         );
  AOI22_X1 U4394 ( .A1(n3460), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3546), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3465) );
  BUF_X1 U4395 ( .A(n3481), .Z(n3461) );
  AOI22_X1 U4396 ( .A1(n4356), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4397 ( .A1(n4383), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3463) );
  AOI22_X1 U4398 ( .A1(n3349), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3348), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3462) );
  NAND4_X1 U4399 ( .A1(n3465), .A2(n3464), .A3(n3463), .A4(n3462), .ZN(n3466)
         );
  NAND2_X1 U4400 ( .A1(n3695), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3470) );
  NAND2_X1 U4401 ( .A1(n3468), .A2(n3525), .ZN(n3469) );
  OAI211_X1 U4402 ( .C1(n3652), .C2(n3543), .A(n3470), .B(n3469), .ZN(n3520)
         );
  INV_X1 U4403 ( .A(n3520), .ZN(n3471) );
  NAND2_X1 U4404 ( .A1(n3472), .A2(n3471), .ZN(n3497) );
  INV_X1 U4405 ( .A(n3474), .ZN(n3475) );
  XNOR2_X1 U4406 ( .A(n3473), .B(n3475), .ZN(n3925) );
  NAND2_X1 U4407 ( .A1(n3925), .A2(n6656), .ZN(n3490) );
  AOI22_X1 U4408 ( .A1(n3460), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3480) );
  AOI22_X1 U4409 ( .A1(n4356), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4410 ( .A1(n4228), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4411 ( .A1(n4374), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3477) );
  NAND4_X1 U4412 ( .A1(n3480), .A2(n3479), .A3(n3478), .A4(n3477), .ZN(n3487)
         );
  AOI22_X1 U4413 ( .A1(n4694), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3485) );
  AOI22_X1 U4414 ( .A1(n4372), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4234), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3484) );
  AOI22_X1 U4415 ( .A1(n4351), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4416 ( .A1(n4229), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3482) );
  NAND4_X1 U4417 ( .A1(n3485), .A2(n3484), .A3(n3483), .A4(n3482), .ZN(n3486)
         );
  INV_X1 U4418 ( .A(n3524), .ZN(n3488) );
  XNOR2_X1 U4419 ( .A(n3488), .B(n3652), .ZN(n3489) );
  NAND2_X1 U4420 ( .A1(n3489), .A2(n3495), .ZN(n3508) );
  NAND2_X1 U4421 ( .A1(n3490), .A2(n3508), .ZN(n3494) );
  INV_X1 U4422 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3493) );
  AOI21_X1 U4423 ( .B1(n4492), .B2(n3652), .A(n6656), .ZN(n3492) );
  NAND2_X1 U4424 ( .A1(n3859), .A2(n3524), .ZN(n3491) );
  OAI211_X1 U4425 ( .C1(n3726), .C2(n3493), .A(n3492), .B(n3491), .ZN(n3507)
         );
  NAND2_X1 U4426 ( .A1(n3495), .A2(n3652), .ZN(n3496) );
  NAND2_X1 U4427 ( .A1(n3521), .A2(n3520), .ZN(n3498) );
  OR2_X1 U4428 ( .A1(n3500), .A2(n3499), .ZN(n3501) );
  INV_X1 U4429 ( .A(n4776), .ZN(n3502) );
  NAND2_X1 U4430 ( .A1(n3502), .A2(n3694), .ZN(n3506) );
  NAND2_X1 U4431 ( .A1(n3525), .A2(n3524), .ZN(n3562) );
  XNOR2_X1 U4432 ( .A(n3562), .B(n3561), .ZN(n3504) );
  AOI21_X1 U4433 ( .B1(n3504), .B2(n3512), .A(n3503), .ZN(n3505) );
  NAND2_X1 U4434 ( .A1(n3506), .A2(n3505), .ZN(n6375) );
  NAND2_X1 U4435 ( .A1(n6375), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3533)
         );
  INV_X1 U4436 ( .A(n3507), .ZN(n3509) );
  NAND2_X1 U4437 ( .A1(n5415), .A2(n3694), .ZN(n3516) );
  INV_X1 U4438 ( .A(n3512), .ZN(n6745) );
  INV_X1 U4439 ( .A(n3503), .ZN(n3513) );
  OAI21_X1 U4440 ( .B1(n6745), .B2(n3524), .A(n3513), .ZN(n3514) );
  INV_X1 U4441 ( .A(n3514), .ZN(n3515) );
  NAND2_X1 U4442 ( .A1(n4587), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3517)
         );
  INV_X1 U4443 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4684) );
  NAND2_X1 U4444 ( .A1(n3517), .A2(n4684), .ZN(n3519) );
  AND2_X1 U4445 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3518) );
  NAND2_X1 U4446 ( .A1(n4587), .A2(n3518), .ZN(n3531) );
  XNOR2_X1 U4447 ( .A(n3521), .B(n3520), .ZN(n3523) );
  XNOR2_X1 U4448 ( .A(n3523), .B(n3522), .ZN(n3920) );
  NAND2_X1 U4449 ( .A1(n3920), .A2(n3694), .ZN(n3530) );
  OAI21_X1 U4450 ( .B1(n3525), .B2(n3524), .A(n3562), .ZN(n3526) );
  INV_X1 U4451 ( .A(n3526), .ZN(n3528) );
  NAND3_X1 U4452 ( .A1(n3313), .A2(n3398), .A3(n4819), .ZN(n3527) );
  AOI21_X1 U4453 ( .B1(n3528), .B2(n3512), .A(n3527), .ZN(n3529) );
  NAND2_X1 U4454 ( .A1(n3530), .A2(n3529), .ZN(n4679) );
  INV_X1 U4455 ( .A(n3531), .ZN(n3532) );
  AOI21_X2 U4456 ( .B1(n4680), .B2(n4679), .A(n3532), .ZN(n6376) );
  NAND2_X1 U4457 ( .A1(n3533), .A2(n6376), .ZN(n3537) );
  NAND2_X1 U4458 ( .A1(n3535), .A2(n3534), .ZN(n3536) );
  NAND2_X1 U4459 ( .A1(n3415), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3542) );
  NAND3_X1 U4460 ( .A1(n6630), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6468) );
  INV_X1 U4461 ( .A(n6468), .ZN(n4780) );
  NAND2_X1 U4462 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4780), .ZN(n6525) );
  NAND2_X1 U4463 ( .A1(n6630), .A2(n6525), .ZN(n3539) );
  NAND3_X1 U4464 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5453) );
  INV_X1 U4465 ( .A(n5453), .ZN(n5181) );
  NAND2_X1 U4466 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5181), .ZN(n5178) );
  NAND2_X1 U4467 ( .A1(n3539), .A2(n5178), .ZN(n4992) );
  OAI22_X1 U4468 ( .A1(n4406), .A2(n4992), .B1(n3761), .B2(n6630), .ZN(n3540)
         );
  INV_X1 U4469 ( .A(n3540), .ZN(n3541) );
  XNOR2_X2 U4470 ( .A(n3538), .B(n4990), .ZN(n4690) );
  AOI22_X1 U4471 ( .A1(n4379), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4234), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3551) );
  AOI22_X1 U4472 ( .A1(n3982), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4473 ( .A1(n3460), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4475 ( .A1(n3547), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3548) );
  NAND4_X1 U4476 ( .A1(n3551), .A2(n3550), .A3(n3549), .A4(n3548), .ZN(n3557)
         );
  AOI22_X1 U4477 ( .A1(n4694), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3555) );
  AOI22_X1 U4478 ( .A1(n4229), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4479 ( .A1(n4356), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4480 ( .A1(n4351), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3552) );
  NAND4_X1 U4481 ( .A1(n3555), .A2(n3554), .A3(n3553), .A4(n3552), .ZN(n3556)
         );
  AOI22_X1 U4482 ( .A1(n3730), .A2(n3582), .B1(n3695), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3558) );
  NAND2_X1 U4483 ( .A1(n4798), .A2(n3694), .ZN(n3566) );
  NAND2_X1 U4484 ( .A1(n3562), .A2(n3561), .ZN(n3583) );
  INV_X1 U4485 ( .A(n3582), .ZN(n3563) );
  XNOR2_X1 U4486 ( .A(n3583), .B(n3563), .ZN(n3564) );
  NAND2_X1 U4487 ( .A1(n3564), .A2(n3512), .ZN(n3565) );
  INV_X1 U4488 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U4489 ( .A1(n6367), .A2(n6368), .ZN(n6366) );
  NAND2_X1 U4490 ( .A1(n3567), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3568)
         );
  NAND2_X1 U4491 ( .A1(n6366), .A2(n3568), .ZN(n4887) );
  AOI22_X1 U4492 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4351), .B1(n3982), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3573) );
  AOI22_X1 U4493 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4229), .B1(n3461), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3572) );
  AOI22_X1 U4494 ( .A1(n3547), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3571) );
  AOI22_X1 U4495 ( .A1(n4694), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3570) );
  NAND4_X1 U4496 ( .A1(n3573), .A2(n3572), .A3(n3571), .A4(n3570), .ZN(n3579)
         );
  AOI22_X1 U4497 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4372), .B1(n4356), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3577) );
  AOI22_X1 U4498 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3459), .B1(n4381), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4499 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4234), .B1(n4382), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4500 ( .A1(n4379), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3574) );
  NAND4_X1 U4501 ( .A1(n3577), .A2(n3576), .A3(n3575), .A4(n3574), .ZN(n3578)
         );
  NAND2_X1 U4502 ( .A1(n3730), .A2(n3629), .ZN(n3581) );
  NAND2_X1 U4503 ( .A1(n3695), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3580) );
  NAND2_X1 U4504 ( .A1(n3946), .A2(n3694), .ZN(n3586) );
  NAND2_X1 U4505 ( .A1(n3583), .A2(n3582), .ZN(n3632) );
  XNOR2_X1 U4506 ( .A(n3632), .B(n3629), .ZN(n3584) );
  NAND2_X1 U4507 ( .A1(n3584), .A2(n3512), .ZN(n3585) );
  NAND2_X1 U4508 ( .A1(n3586), .A2(n3585), .ZN(n3587) );
  INV_X1 U4509 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6419) );
  XNOR2_X1 U4510 ( .A(n3587), .B(n6419), .ZN(n4886) );
  NAND2_X1 U4511 ( .A1(n4887), .A2(n4886), .ZN(n4885) );
  NAND2_X1 U4512 ( .A1(n3587), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3588)
         );
  NAND2_X1 U4513 ( .A1(n4885), .A2(n3588), .ZN(n6360) );
  AOI22_X1 U4514 ( .A1(n4229), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3592) );
  AOI22_X1 U4515 ( .A1(n4351), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4516 ( .A1(n3982), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3590) );
  AOI22_X1 U4517 ( .A1(n4694), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3589) );
  NAND4_X1 U4518 ( .A1(n3592), .A2(n3591), .A3(n3590), .A4(n3589), .ZN(n3598)
         );
  AOI22_X1 U4519 ( .A1(n3460), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4520 ( .A1(n3461), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4521 ( .A1(n4234), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4522 ( .A1(n4356), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3593) );
  NAND4_X1 U4523 ( .A1(n3596), .A2(n3595), .A3(n3594), .A4(n3593), .ZN(n3597)
         );
  NAND2_X1 U4524 ( .A1(n3730), .A2(n3630), .ZN(n3600) );
  NAND2_X1 U4525 ( .A1(n3695), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3599) );
  NAND2_X1 U4526 ( .A1(n3600), .A2(n3599), .ZN(n3610) );
  NAND2_X1 U4527 ( .A1(n3905), .A2(n3694), .ZN(n3606) );
  INV_X1 U4528 ( .A(n3629), .ZN(n3602) );
  OR2_X1 U4529 ( .A1(n3632), .A2(n3602), .ZN(n3603) );
  XNOR2_X1 U4530 ( .A(n3603), .B(n3630), .ZN(n3604) );
  NAND2_X1 U4531 ( .A1(n3604), .A2(n3512), .ZN(n3605) );
  NAND2_X1 U4532 ( .A1(n3606), .A2(n3605), .ZN(n3607) );
  INV_X1 U4533 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3790) );
  XNOR2_X1 U4534 ( .A(n3607), .B(n3790), .ZN(n6359) );
  NAND2_X1 U4535 ( .A1(n6360), .A2(n6359), .ZN(n6358) );
  NAND2_X1 U4536 ( .A1(n3607), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3608)
         );
  INV_X1 U4537 ( .A(n3609), .ZN(n3612) );
  AOI22_X1 U4538 ( .A1(n4229), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4539 ( .A1(n4351), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4540 ( .A1(n3982), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4541 ( .A1(n4694), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3613) );
  NAND4_X1 U4542 ( .A1(n3616), .A2(n3615), .A3(n3614), .A4(n3613), .ZN(n3622)
         );
  AOI22_X1 U4543 ( .A1(n3460), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4544 ( .A1(n3461), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4545 ( .A1(n4234), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4546 ( .A1(n4356), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3617) );
  NAND4_X1 U4547 ( .A1(n3620), .A2(n3619), .A3(n3618), .A4(n3617), .ZN(n3621)
         );
  NAND2_X1 U4548 ( .A1(n3730), .A2(n3642), .ZN(n3624) );
  NAND2_X1 U4549 ( .A1(n3695), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3623) );
  NAND2_X1 U4550 ( .A1(n3624), .A2(n3623), .ZN(n3626) );
  INV_X1 U4551 ( .A(n3626), .ZN(n3627) );
  NAND2_X1 U4552 ( .A1(n3628), .A2(n3627), .ZN(n3912) );
  NAND3_X1 U4553 ( .A1(n3640), .A2(n3694), .A3(n3912), .ZN(n3635) );
  NAND2_X1 U4554 ( .A1(n3630), .A2(n3629), .ZN(n3631) );
  OR2_X1 U4555 ( .A1(n3632), .A2(n3631), .ZN(n3641) );
  XNOR2_X1 U4556 ( .A(n3641), .B(n3642), .ZN(n3633) );
  NAND2_X1 U4557 ( .A1(n3633), .A2(n3512), .ZN(n3634) );
  NAND2_X1 U4558 ( .A1(n3635), .A2(n3634), .ZN(n3636) );
  INV_X1 U4559 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4949) );
  XNOR2_X1 U4560 ( .A(n3636), .B(n4949), .ZN(n4939) );
  INV_X1 U4561 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3638) );
  NAND2_X1 U4562 ( .A1(n3730), .A2(n3652), .ZN(n3637) );
  OAI21_X1 U4563 ( .B1(n3638), .B2(n3726), .A(n3637), .ZN(n3639) );
  NAND2_X1 U4564 ( .A1(n3965), .A2(n3694), .ZN(n3646) );
  INV_X1 U4565 ( .A(n3641), .ZN(n3643) );
  NAND2_X1 U4566 ( .A1(n3643), .A2(n3642), .ZN(n3654) );
  XNOR2_X1 U4567 ( .A(n3654), .B(n3652), .ZN(n3644) );
  NAND2_X1 U4568 ( .A1(n3644), .A2(n3512), .ZN(n3645) );
  NAND2_X1 U4569 ( .A1(n3646), .A2(n3645), .ZN(n3647) );
  INV_X1 U4570 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6418) );
  XNOR2_X1 U4571 ( .A(n3647), .B(n6418), .ZN(n6351) );
  NAND2_X1 U4572 ( .A1(n3647), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3648)
         );
  NAND2_X1 U4573 ( .A1(n6350), .A2(n3648), .ZN(n5070) );
  NAND2_X1 U4574 ( .A1(n3652), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3649) );
  NOR2_X1 U4575 ( .A1(n3650), .A2(n3649), .ZN(n3651) );
  INV_X1 U4576 ( .A(n3652), .ZN(n3653) );
  OR3_X1 U4577 ( .A1(n3654), .A2(n3653), .A3(n6745), .ZN(n3655) );
  NAND2_X1 U4578 ( .A1(n3658), .A2(n3655), .ZN(n3656) );
  INV_X1 U4579 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6410) );
  XNOR2_X1 U4580 ( .A(n3656), .B(n6410), .ZN(n5069) );
  NAND2_X1 U4581 ( .A1(n5070), .A2(n5069), .ZN(n5068) );
  NAND2_X1 U4582 ( .A1(n3656), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3657)
         );
  NAND2_X1 U4583 ( .A1(n5068), .A2(n3657), .ZN(n5213) );
  INV_X1 U4584 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U4585 ( .A1(n6101), .A2(n6399), .ZN(n5214) );
  NAND2_X1 U4586 ( .A1(n5213), .A2(n5214), .ZN(n3659) );
  OR2_X1 U4587 ( .A1(n3155), .A2(n6399), .ZN(n5215) );
  INV_X1 U4588 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3660) );
  NAND2_X1 U4589 ( .A1(n3155), .A2(n3660), .ZN(n5297) );
  INV_X1 U4590 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5357) );
  AND2_X1 U4591 ( .A1(n3658), .A2(n5357), .ZN(n3663) );
  OR2_X1 U4592 ( .A1(n3658), .A2(n3660), .ZN(n5355) );
  INV_X1 U4593 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5534) );
  NOR2_X1 U4594 ( .A1(n3155), .A2(n5534), .ZN(n5521) );
  XNOR2_X1 U4595 ( .A(n6101), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5819)
         );
  NAND2_X1 U4596 ( .A1(n5818), .A2(n5819), .ZN(n3665) );
  NAND2_X1 U4597 ( .A1(n6101), .A2(n3817), .ZN(n3664) );
  NAND2_X1 U4598 ( .A1(n3665), .A2(n3664), .ZN(n5812) );
  INV_X1 U4599 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5813) );
  AND2_X1 U4600 ( .A1(n6101), .A2(n5813), .ZN(n3666) );
  INV_X1 U4601 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5942) );
  NAND2_X1 U4602 ( .A1(n6101), .A2(n5942), .ZN(n3667) );
  INV_X1 U4603 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U4604 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3869) );
  OR2_X1 U4605 ( .A1(n6101), .A2(n6099), .ZN(n5797) );
  NOR2_X1 U4606 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3668) );
  OR2_X1 U4607 ( .A1(n6101), .A2(n3668), .ZN(n3669) );
  NAND2_X1 U4608 ( .A1(n3674), .A2(n3670), .ZN(n6091) );
  INV_X1 U4609 ( .A(n6091), .ZN(n3671) );
  NAND2_X1 U4610 ( .A1(n3671), .A2(n6093), .ZN(n6092) );
  INV_X1 U4611 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6093) );
  OAI21_X1 U4612 ( .B1(n3674), .B2(n6093), .A(n3155), .ZN(n3672) );
  XNOR2_X1 U4613 ( .A(n3155), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5784)
         );
  INV_X1 U4614 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3841) );
  NOR2_X1 U4615 ( .A1(n3155), .A2(n3841), .ZN(n3673) );
  XNOR2_X1 U4616 ( .A(n3658), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5778)
         );
  AND2_X1 U4617 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5918) );
  AND2_X1 U4618 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3886) );
  NAND2_X1 U4619 ( .A1(n5918), .A2(n3886), .ZN(n3894) );
  OR3_X1 U4620 ( .A1(n3674), .A2(n6100), .A3(n3894), .ZN(n3675) );
  NAND2_X1 U4621 ( .A1(n3730), .A2(n4783), .ZN(n3678) );
  NAND2_X1 U4622 ( .A1(n3678), .A2(n3398), .ZN(n3689) );
  NAND2_X1 U4623 ( .A1(n5370), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3700) );
  NAND2_X1 U4624 ( .A1(n3370), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3679) );
  NAND2_X1 U4625 ( .A1(n3700), .A2(n3679), .ZN(n3680) );
  NAND2_X1 U4626 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n5407), .ZN(n3683) );
  NAND2_X1 U4627 ( .A1(n3680), .A2(n3683), .ZN(n3681) );
  NAND2_X1 U4628 ( .A1(n3701), .A2(n3681), .ZN(n3754) );
  NOR2_X1 U4629 ( .A1(n3754), .A2(n6656), .ZN(n3690) );
  INV_X1 U4630 ( .A(n3683), .ZN(n3684) );
  AOI21_X1 U4631 ( .B1(n3682), .B2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n3684), 
        .ZN(n3688) );
  AOI21_X1 U4632 ( .B1(n3768), .B2(n3688), .A(n3859), .ZN(n3687) );
  NAND2_X1 U4633 ( .A1(n3685), .A2(n3398), .ZN(n3686) );
  NAND2_X1 U4634 ( .A1(n4669), .A2(n3686), .ZN(n3713) );
  OAI22_X1 U4635 ( .A1(n3689), .A2(n3690), .B1(n3687), .B2(n3713), .ZN(n3697)
         );
  NAND2_X1 U4636 ( .A1(n3730), .A2(n3688), .ZN(n3693) );
  INV_X1 U4637 ( .A(n3689), .ZN(n3692) );
  INV_X1 U4638 ( .A(n3690), .ZN(n3691) );
  OAI22_X1 U4639 ( .A1(n3697), .A2(n3693), .B1(n3692), .B2(n3691), .ZN(n3699)
         );
  INV_X1 U4640 ( .A(n3754), .ZN(n3696) );
  AOI21_X1 U4641 ( .B1(n3697), .B2(n3696), .A(n3731), .ZN(n3698) );
  NAND2_X1 U4642 ( .A1(n6625), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3717) );
  NAND2_X1 U4643 ( .A1(n4601), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3702) );
  NAND2_X1 U4644 ( .A1(n3717), .A2(n3702), .ZN(n3704) );
  NAND2_X1 U4645 ( .A1(n3703), .A2(n3704), .ZN(n3707) );
  INV_X1 U4646 ( .A(n3704), .ZN(n3705) );
  NAND2_X1 U4647 ( .A1(n3707), .A2(n3718), .ZN(n3755) );
  INV_X1 U4648 ( .A(n3755), .ZN(n3709) );
  NAND2_X1 U4649 ( .A1(n3730), .A2(n3709), .ZN(n3712) );
  INV_X1 U4650 ( .A(n3713), .ZN(n3708) );
  OAI211_X1 U4651 ( .C1(n3709), .C2(n3726), .A(n3712), .B(n3708), .ZN(n3710)
         );
  NAND2_X1 U4652 ( .A1(n3711), .A2(n3710), .ZN(n3716) );
  INV_X1 U4653 ( .A(n3712), .ZN(n3714) );
  NAND2_X1 U4654 ( .A1(n3714), .A2(n3713), .ZN(n3715) );
  NAND2_X1 U4655 ( .A1(n3716), .A2(n3715), .ZN(n3728) );
  NAND2_X1 U4656 ( .A1(n3718), .A2(n3717), .ZN(n3721) );
  XNOR2_X1 U4657 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3720) );
  NAND2_X1 U4658 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3729), .ZN(n3719) );
  NOR2_X1 U4659 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n3719), .ZN(n3725)
         );
  NOR2_X1 U4660 ( .A1(n3721), .A2(n3720), .ZN(n3722) );
  OR2_X1 U4661 ( .A1(n3723), .A2(n3722), .ZN(n3724) );
  NAND2_X1 U4662 ( .A1(n3753), .A2(n3726), .ZN(n3727) );
  NAND2_X1 U4663 ( .A1(n3728), .A2(n3727), .ZN(n3734) );
  AOI222_X1 U4664 ( .A1(n3729), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B1(
        n3729), .B2(n3949), .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n3949), 
        .ZN(n3756) );
  NAND2_X1 U4665 ( .A1(n3756), .A2(n3730), .ZN(n3733) );
  AOI22_X1 U4666 ( .A1(n3753), .A2(n3735), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6656), .ZN(n3732) );
  NAND2_X1 U4667 ( .A1(n3756), .A2(n3735), .ZN(n3736) );
  NAND2_X1 U4668 ( .A1(n3385), .A2(n3383), .ZN(n3738) );
  OR3_X1 U4669 ( .A1(n5597), .A2(n3685), .A3(n6613), .ZN(n3749) );
  INV_X1 U4670 ( .A(n4429), .ZN(n5589) );
  AND2_X1 U4671 ( .A1(n4676), .A2(n3858), .ZN(n4675) );
  OR2_X1 U4672 ( .A1(n4675), .A2(n3740), .ZN(n3744) );
  NAND2_X1 U4673 ( .A1(n3741), .A2(n4874), .ZN(n3742) );
  NAND2_X1 U4674 ( .A1(n6745), .A2(n3742), .ZN(n3743) );
  NAND2_X1 U4675 ( .A1(n3744), .A2(n3743), .ZN(n3860) );
  INV_X1 U4676 ( .A(n3860), .ZN(n3747) );
  NOR2_X1 U4677 ( .A1(n3745), .A2(n4832), .ZN(n3857) );
  NAND2_X1 U4678 ( .A1(n6613), .A2(n3859), .ZN(n3746) );
  NAND2_X1 U4679 ( .A1(n3857), .A2(n3746), .ZN(n3769) );
  OR2_X1 U4680 ( .A1(n3747), .A2(n3769), .ZN(n3748) );
  NAND2_X1 U4681 ( .A1(n5589), .A2(n3748), .ZN(n3868) );
  NAND2_X1 U4682 ( .A1(n3749), .A2(n3868), .ZN(n4520) );
  INV_X1 U4683 ( .A(n3750), .ZN(n3752) );
  INV_X1 U4684 ( .A(STATE_REG_0__SCAN_IN), .ZN(n3751) );
  NAND2_X1 U4685 ( .A1(n3752), .A2(n3751), .ZN(n6673) );
  NAND2_X1 U4686 ( .A1(n4783), .A2(n6673), .ZN(n3760) );
  INV_X1 U4687 ( .A(n3753), .ZN(n3758) );
  NOR2_X1 U4688 ( .A1(n3755), .A2(n3754), .ZN(n3757) );
  AOI21_X1 U4689 ( .B1(n3758), .B2(n3757), .A(n3756), .ZN(n5590) );
  INV_X1 U4690 ( .A(n5590), .ZN(n3759) );
  NOR2_X1 U4691 ( .A1(n3759), .A2(READY_N), .ZN(n4521) );
  AND3_X1 U4692 ( .A1(n3760), .A2(n4832), .A3(n4521), .ZN(n3762) );
  OAI21_X1 U4693 ( .B1(n4520), .B2(n3762), .A(n6652), .ZN(n3767) );
  NAND2_X1 U4694 ( .A1(n3685), .A2(n6673), .ZN(n4435) );
  NAND3_X1 U4695 ( .A1(n4540), .A2(n5605), .A3(n4435), .ZN(n3763) );
  NAND3_X1 U4696 ( .A1(n3763), .A2(n4874), .A3(n3858), .ZN(n3764) );
  NAND2_X1 U4697 ( .A1(n3764), .A2(n3313), .ZN(n3765) );
  OR2_X1 U4698 ( .A1(n4563), .A2(n3765), .ZN(n3766) );
  NOR2_X1 U4699 ( .A1(n3769), .A2(n4669), .ZN(n5588) );
  INV_X1 U4700 ( .A(n5588), .ZN(n4593) );
  NAND2_X4 U4701 ( .A1(n4783), .A2(n3154), .ZN(n4666) );
  AOI22_X1 U4702 ( .A1(n3854), .A2(n3385), .B1(n4540), .B2(n4465), .ZN(n3770)
         );
  NAND4_X1 U4703 ( .A1(n4593), .A2(n3770), .A3(n4542), .A4(n6607), .ZN(n3771)
         );
  NAND2_X1 U4704 ( .A1(n4418), .A2(n6454), .ZN(n3893) );
  INV_X1 U4705 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U4706 ( .A1(n4462), .A2(n6064), .ZN(n3775) );
  NAND2_X1 U4707 ( .A1(n4465), .A2(n6064), .ZN(n3773) );
  INV_X1 U4708 ( .A(n4819), .ZN(n3772) );
  OAI211_X1 U4709 ( .C1(n3833), .C2(n3676), .A(n3773), .B(n4455), .ZN(n3774)
         );
  NAND2_X1 U4710 ( .A1(n3775), .A2(n3774), .ZN(n3853) );
  NAND2_X1 U4711 ( .A1(n4438), .A2(n4668), .ZN(n3777) );
  NAND2_X1 U4712 ( .A1(n3777), .A2(n3776), .ZN(n3781) );
  INV_X1 U4713 ( .A(n4455), .ZN(n3778) );
  NAND2_X1 U4714 ( .A1(n3778), .A2(n4666), .ZN(n4440) );
  NAND2_X1 U4715 ( .A1(n4666), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3779)
         );
  AND2_X1 U4716 ( .A1(n4440), .A2(n3779), .ZN(n3780) );
  NAND2_X1 U4717 ( .A1(n4455), .A2(EBX_REG_0__SCAN_IN), .ZN(n3782) );
  OAI21_X1 U4718 ( .B1(n3833), .B2(EBX_REG_0__SCAN_IN), .A(n3782), .ZN(n4579)
         );
  XNOR2_X1 U4719 ( .A(n3783), .B(n4579), .ZN(n4663) );
  NAND2_X1 U4720 ( .A1(n4663), .A2(n4465), .ZN(n4664) );
  NAND3_X1 U4721 ( .A1(n5685), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .A3(n4666), 
        .ZN(n3784) );
  AND2_X1 U4722 ( .A1(n4440), .A2(n3784), .ZN(n3785) );
  INV_X1 U4723 ( .A(n4768), .ZN(n3788) );
  MUX2_X1 U4724 ( .A(n4449), .B(n5685), .S(EBX_REG_3__SCAN_IN), .Z(n3787) );
  NAND2_X1 U4725 ( .A1(n4581), .A2(n6444), .ZN(n3786) );
  NAND2_X1 U4726 ( .A1(n3787), .A2(n3786), .ZN(n4769) );
  NOR2_X1 U4727 ( .A1(n3788), .A2(n4769), .ZN(n3789) );
  MUX2_X1 U4728 ( .A(n4449), .B(n5685), .S(EBX_REG_5__SCAN_IN), .Z(n3792) );
  NAND2_X1 U4729 ( .A1(n3790), .A2(n4581), .ZN(n3791) );
  AND2_X1 U4730 ( .A1(n3792), .A2(n3791), .ZN(n4791) );
  INV_X1 U4731 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4763) );
  NAND2_X1 U4732 ( .A1(n4453), .A2(n4763), .ZN(n3795) );
  NAND2_X1 U4733 ( .A1(n4455), .A2(n6419), .ZN(n3793) );
  OAI211_X1 U4734 ( .C1(EBX_REG_4__SCAN_IN), .C2(n4666), .A(n3793), .B(n5685), 
        .ZN(n3794) );
  NAND2_X1 U4735 ( .A1(n3795), .A2(n3794), .ZN(n4792) );
  NAND2_X1 U4736 ( .A1(n4791), .A2(n4792), .ZN(n3796) );
  INV_X1 U4737 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4879) );
  NAND2_X1 U4738 ( .A1(n4453), .A2(n4879), .ZN(n3800) );
  NAND2_X1 U4739 ( .A1(n4455), .A2(n4949), .ZN(n3798) );
  NAND2_X1 U4740 ( .A1(n4465), .A2(n4879), .ZN(n3797) );
  NAND3_X1 U4741 ( .A1(n3798), .A2(n5685), .A3(n3797), .ZN(n3799) );
  NAND2_X1 U4742 ( .A1(n3800), .A2(n3799), .ZN(n4842) );
  NAND2_X1 U4743 ( .A1(n6418), .A2(n4581), .ZN(n3802) );
  MUX2_X1 U4744 ( .A(n4449), .B(n5685), .S(EBX_REG_7__SCAN_IN), .Z(n3801) );
  NAND2_X1 U4745 ( .A1(n3802), .A2(n3801), .ZN(n4959) );
  INV_X1 U4746 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4985) );
  NAND2_X1 U4747 ( .A1(n4453), .A2(n4985), .ZN(n3807) );
  NAND2_X1 U4748 ( .A1(n4455), .A2(n6410), .ZN(n3805) );
  NAND2_X1 U4749 ( .A1(n4465), .A2(n4985), .ZN(n3804) );
  NAND3_X1 U4750 ( .A1(n3805), .A2(n5685), .A3(n3804), .ZN(n3806) );
  MUX2_X1 U4751 ( .A(n4449), .B(n5685), .S(EBX_REG_9__SCAN_IN), .Z(n3809) );
  NAND2_X1 U4752 ( .A1(n4581), .A2(n6399), .ZN(n3808) );
  NAND2_X1 U4753 ( .A1(n3809), .A2(n3808), .ZN(n5081) );
  MUX2_X1 U4754 ( .A(n4438), .B(n4455), .S(EBX_REG_10__SCAN_IN), .Z(n3812) );
  NAND2_X1 U4755 ( .A1(n4666), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3810) );
  AND2_X1 U4756 ( .A1(n4440), .A2(n3810), .ZN(n3811) );
  NAND2_X1 U4757 ( .A1(n3812), .A2(n3811), .ZN(n5225) );
  NAND2_X1 U4758 ( .A1(n5226), .A2(n5225), .ZN(n5244) );
  INV_X1 U4759 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5251) );
  NAND2_X1 U4760 ( .A1(n4462), .A2(n5251), .ZN(n3815) );
  NAND2_X1 U4761 ( .A1(n4465), .A2(n5251), .ZN(n3813) );
  OAI211_X1 U4762 ( .C1(n3833), .C2(n5357), .A(n3813), .B(n4455), .ZN(n3814)
         );
  NAND2_X1 U4763 ( .A1(n3815), .A2(n3814), .ZN(n5245) );
  INV_X1 U4764 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U4765 ( .A1(n4462), .A2(n5507), .ZN(n3819) );
  INV_X1 U4766 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3817) );
  NAND2_X1 U4767 ( .A1(n4465), .A2(n5507), .ZN(n3816) );
  OAI211_X1 U4768 ( .C1(n3833), .C2(n3817), .A(n3816), .B(n4455), .ZN(n3818)
         );
  MUX2_X1 U4769 ( .A(n4438), .B(n4455), .S(EBX_REG_12__SCAN_IN), .Z(n3822) );
  NAND2_X1 U4770 ( .A1(n4666), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3820) );
  AND2_X1 U4771 ( .A1(n4440), .A2(n3820), .ZN(n3821) );
  NAND2_X1 U4772 ( .A1(n3822), .A2(n3821), .ZN(n5504) );
  MUX2_X1 U4773 ( .A(n4438), .B(n4455), .S(EBX_REG_14__SCAN_IN), .Z(n3825) );
  NAND2_X1 U4774 ( .A1(n4666), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3823) );
  AND2_X1 U4775 ( .A1(n4440), .A2(n3823), .ZN(n3824) );
  NAND2_X1 U4776 ( .A1(n3825), .A2(n3824), .ZN(n5548) );
  INV_X1 U4777 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U4778 ( .A1(n4462), .A2(n5708), .ZN(n3828) );
  NAND2_X1 U4779 ( .A1(n4465), .A2(n5708), .ZN(n3826) );
  OAI211_X1 U4780 ( .C1(n3833), .C2(n5942), .A(n3826), .B(n4455), .ZN(n3827)
         );
  MUX2_X1 U4781 ( .A(n4438), .B(n4455), .S(EBX_REG_16__SCAN_IN), .Z(n3831) );
  NAND2_X1 U4782 ( .A1(n4666), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3829) );
  AND2_X1 U4783 ( .A1(n4440), .A2(n3829), .ZN(n3830) );
  INV_X1 U4784 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U4785 ( .A1(n4462), .A2(n6296), .ZN(n3835) );
  INV_X1 U4786 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U4787 ( .A1(n4465), .A2(n6296), .ZN(n3832) );
  OAI211_X1 U4788 ( .C1(n3833), .C2(n6129), .A(n3832), .B(n4455), .ZN(n3834)
         );
  NAND2_X1 U4789 ( .A1(n3835), .A2(n3834), .ZN(n6131) );
  INV_X1 U4790 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U4791 ( .A1(n4453), .A2(n6068), .ZN(n3839) );
  NAND2_X1 U4792 ( .A1(n4455), .A2(n6093), .ZN(n3837) );
  NAND2_X1 U4793 ( .A1(n4465), .A2(n6068), .ZN(n3836) );
  NAND3_X1 U4794 ( .A1(n3837), .A2(n5685), .A3(n3836), .ZN(n3838) );
  NAND2_X1 U4795 ( .A1(n3839), .A2(n3838), .ZN(n6058) );
  NOR2_X1 U4797 ( .A1(n4666), .A2(EBX_REG_20__SCAN_IN), .ZN(n3840) );
  AOI21_X1 U4798 ( .B1(n4581), .B2(n3841), .A(n3840), .ZN(n5686) );
  INV_X1 U4799 ( .A(n4581), .ZN(n4470) );
  OR2_X1 U4800 ( .A1(n4470), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3843)
         );
  INV_X1 U4801 ( .A(EBX_REG_18__SCAN_IN), .ZN(n3842) );
  NAND2_X1 U4802 ( .A1(n4465), .A2(n3842), .ZN(n5690) );
  NAND2_X1 U4803 ( .A1(n3843), .A2(n5690), .ZN(n5691) );
  NAND2_X1 U4804 ( .A1(n3833), .A2(EBX_REG_20__SCAN_IN), .ZN(n3845) );
  NAND2_X1 U4805 ( .A1(n5691), .A2(n5685), .ZN(n3844) );
  OAI211_X1 U4806 ( .C1(n5686), .C2(n5691), .A(n3845), .B(n3844), .ZN(n3846)
         );
  INV_X1 U4807 ( .A(n3846), .ZN(n3847) );
  INV_X1 U4808 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U4809 ( .A1(n5913), .A2(n4581), .ZN(n3849) );
  MUX2_X1 U4810 ( .A(n4449), .B(n5685), .S(EBX_REG_21__SCAN_IN), .Z(n3848) );
  NAND2_X1 U4811 ( .A1(n3849), .A2(n3848), .ZN(n5677) );
  MUX2_X1 U4812 ( .A(n4438), .B(n4455), .S(EBX_REG_22__SCAN_IN), .Z(n3852) );
  NAND2_X1 U4813 ( .A1(n4666), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3850) );
  AND2_X1 U4814 ( .A1(n4440), .A2(n3850), .ZN(n3851) );
  AOI21_X1 U4815 ( .B1(n3853), .B2(n5668), .A(n5661), .ZN(n6062) );
  INV_X1 U4816 ( .A(n6062), .ZN(n3890) );
  NAND2_X1 U4817 ( .A1(n3854), .A2(n4492), .ZN(n3855) );
  NAND2_X1 U4818 ( .A1(n4540), .A2(n3512), .ZN(n6642) );
  NAND2_X1 U4819 ( .A1(n3855), .A2(n6642), .ZN(n3856) );
  AND2_X2 U4820 ( .A1(n3872), .A2(n3856), .ZN(n6448) );
  NOR2_X1 U4821 ( .A1(n3857), .A2(n4581), .ZN(n3862) );
  INV_X1 U4822 ( .A(n3858), .ZN(n4678) );
  NAND2_X1 U4823 ( .A1(n3859), .A2(n4783), .ZN(n4963) );
  OR2_X1 U4824 ( .A1(n4963), .A2(n4832), .ZN(n4526) );
  OAI211_X1 U4825 ( .C1(n3313), .C2(n4678), .A(n3860), .B(n4526), .ZN(n3861)
         );
  NAND2_X1 U4826 ( .A1(n3172), .A2(n4698), .ZN(n3864) );
  NAND2_X1 U4827 ( .A1(n3872), .A2(n3864), .ZN(n5952) );
  OR2_X1 U4828 ( .A1(n5952), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3865)
         );
  INV_X2 U4829 ( .A(n6403), .ZN(n6457) );
  OR2_X1 U4830 ( .A1(n3872), .A2(n6457), .ZN(n4682) );
  NAND2_X1 U4831 ( .A1(n3865), .A2(n4682), .ZN(n5923) );
  NAND2_X1 U4832 ( .A1(n4526), .A2(n4783), .ZN(n3866) );
  NOR2_X1 U4833 ( .A1(n3866), .A2(n6613), .ZN(n3867) );
  NAND2_X1 U4834 ( .A1(n3868), .A2(n3867), .ZN(n4594) );
  INV_X1 U4835 ( .A(n4594), .ZN(n5593) );
  NAND2_X1 U4836 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6452) );
  NAND2_X1 U4837 ( .A1(n3534), .A2(n6452), .ZN(n6420) );
  NAND4_X1 U4838 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .A4(n6420), .ZN(n4948) );
  NOR2_X1 U4839 ( .A1(n4949), .A2(n4948), .ZN(n5307) );
  NOR2_X1 U4840 ( .A1(n6418), .A2(n6410), .ZN(n6402) );
  INV_X1 U4841 ( .A(n6402), .ZN(n5308) );
  NAND2_X1 U4842 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5309) );
  NOR2_X1 U4843 ( .A1(n5308), .A2(n5309), .ZN(n3874) );
  NAND2_X1 U4844 ( .A1(n5307), .A2(n3874), .ZN(n5532) );
  NAND3_X1 U4845 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5949) );
  NOR2_X1 U4846 ( .A1(n5813), .A2(n5949), .ZN(n5941) );
  NAND3_X1 U4847 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5941), .ZN(n5924) );
  NOR2_X1 U4848 ( .A1(n5532), .A2(n5924), .ZN(n5928) );
  INV_X1 U4849 ( .A(n3869), .ZN(n3884) );
  AND2_X1 U4850 ( .A1(n3884), .A2(n5918), .ZN(n3875) );
  AND2_X1 U4851 ( .A1(n5928), .A2(n3875), .ZN(n3870) );
  NOR2_X1 U4852 ( .A1(n6453), .A2(n3870), .ZN(n3871) );
  NOR2_X1 U4853 ( .A1(n5923), .A2(n3871), .ZN(n3881) );
  NAND2_X1 U4854 ( .A1(n3872), .A2(n6617), .ZN(n5947) );
  NAND3_X1 U4855 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n3873) );
  NOR2_X1 U4856 ( .A1(n4949), .A2(n3873), .ZN(n5304) );
  NAND4_X1 U4857 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n3874), .A4(n5304), .ZN(n5926) );
  INV_X1 U4858 ( .A(n5926), .ZN(n3878) );
  INV_X1 U4859 ( .A(n3875), .ZN(n3876) );
  NOR2_X1 U4860 ( .A1(n5924), .A2(n3876), .ZN(n3877) );
  NAND2_X1 U4861 ( .A1(n3878), .A2(n3877), .ZN(n3879) );
  NAND2_X1 U4862 ( .A1(n5925), .A2(n3879), .ZN(n3880) );
  AND2_X1 U4863 ( .A1(n3881), .A2(n3880), .ZN(n5910) );
  INV_X1 U4864 ( .A(n3886), .ZN(n5901) );
  NAND2_X1 U4865 ( .A1(n5847), .A2(n5901), .ZN(n3882) );
  AND2_X1 U4866 ( .A1(n5910), .A2(n3882), .ZN(n5827) );
  INV_X1 U4867 ( .A(n5827), .ZN(n3888) );
  INV_X1 U4868 ( .A(REIP_REG_23__SCAN_IN), .ZN(n3883) );
  NOR2_X1 U4869 ( .A1(n6403), .A2(n3883), .ZN(n4423) );
  NOR2_X1 U4870 ( .A1(n6453), .A2(n5532), .ZN(n5955) );
  INV_X1 U4871 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4589) );
  NAND2_X1 U4872 ( .A1(n4589), .A2(n5947), .ZN(n4683) );
  NAND2_X1 U4873 ( .A1(n5925), .A2(n4683), .ZN(n5922) );
  NOR2_X1 U4874 ( .A1(n5922), .A2(n5926), .ZN(n5533) );
  NAND2_X1 U4875 ( .A1(n3884), .A2(n6130), .ZN(n6125) );
  INV_X1 U4876 ( .A(n5918), .ZN(n3885) );
  NOR2_X1 U4877 ( .A1(n6125), .A2(n3885), .ZN(n5914) );
  NAND2_X1 U4878 ( .A1(n5914), .A2(n3886), .ZN(n5892) );
  NOR2_X1 U4879 ( .A1(n5892), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3887)
         );
  AOI211_X1 U4880 ( .C1(n3888), .C2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n4423), .B(n3887), .ZN(n3889) );
  INV_X1 U4881 ( .A(n3891), .ZN(n3892) );
  NAND2_X1 U4882 ( .A1(n3893), .A2(n3892), .ZN(U2995) );
  NAND2_X1 U4883 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5833) );
  OAI21_X1 U4884 ( .B1(n3894), .B2(n5833), .A(n3658), .ZN(n3895) );
  NAND2_X1 U4885 ( .A1(n6091), .A2(n3895), .ZN(n3898) );
  NOR2_X1 U4886 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5899) );
  NOR2_X1 U4887 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5891) );
  NOR2_X1 U4888 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5919) );
  AND3_X1 U4889 ( .A1(n5899), .A2(n5891), .A3(n5919), .ZN(n3896) );
  NAND2_X1 U4890 ( .A1(n3898), .A2(n3897), .ZN(n5565) );
  INV_X1 U4891 ( .A(n5565), .ZN(n3899) );
  INV_X1 U4892 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U4893 ( .A1(n3155), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5754) );
  NOR2_X2 U4894 ( .A1(n5727), .A2(n5754), .ZN(n5746) );
  AND2_X1 U4895 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U4896 ( .A1(n5746), .A2(n5834), .ZN(n5738) );
  NAND2_X1 U4897 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5835) );
  INV_X1 U4898 ( .A(n3901), .ZN(n3902) );
  INV_X1 U4899 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4454) );
  INV_X1 U4900 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5749) );
  NAND2_X1 U4901 ( .A1(n4454), .A2(n5749), .ZN(n5865) );
  NOR2_X1 U4902 ( .A1(n5739), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5726)
         );
  INV_X1 U4903 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5845) );
  NAND3_X1 U4904 ( .A1(n3902), .A2(n5726), .A3(n5845), .ZN(n3903) );
  XNOR2_X1 U4905 ( .A(n3904), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5843)
         );
  NAND2_X1 U4906 ( .A1(n3905), .A2(n4087), .ZN(n3911) );
  INV_X1 U4907 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3908) );
  OAI21_X1 U4908 ( .B1(n3951), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3960), 
        .ZN(n6365) );
  NAND2_X1 U4909 ( .A1(n6365), .A2(n4430), .ZN(n3907) );
  NAND2_X1 U4910 ( .A1(n4401), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3906)
         );
  OAI211_X1 U4911 ( .C1(n4161), .C2(n3908), .A(n3907), .B(n3906), .ZN(n3909)
         );
  INV_X1 U4912 ( .A(n3909), .ZN(n3910) );
  NAND2_X1 U4913 ( .A1(n3911), .A2(n3910), .ZN(n4767) );
  NAND2_X1 U4914 ( .A1(n3912), .A2(n4087), .ZN(n3918) );
  INV_X1 U4915 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3914) );
  INV_X1 U4916 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6163) );
  OAI21_X1 U4917 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6163), .A(n6655), 
        .ZN(n3913) );
  OAI21_X1 U4918 ( .B1(n4161), .B2(n3914), .A(n3913), .ZN(n3916) );
  XNOR2_X1 U4919 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n3960), .ZN(n4942) );
  NAND2_X1 U4920 ( .A1(n4942), .A2(n4430), .ZN(n3915) );
  NAND2_X1 U4921 ( .A1(n3916), .A2(n3915), .ZN(n3917) );
  NAND2_X1 U4922 ( .A1(n3918), .A2(n3917), .ZN(n4838) );
  INV_X1 U4923 ( .A(n4087), .ZN(n4027) );
  INV_X1 U4924 ( .A(n4401), .ZN(n3919) );
  NAND2_X1 U4925 ( .A1(n3920), .A2(n4087), .ZN(n3924) );
  INV_X1 U4926 ( .A(n4161), .ZN(n4402) );
  AOI22_X1 U4927 ( .A1(n4402), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6655), .ZN(n3922) );
  NAND2_X1 U4928 ( .A1(n3932), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3921) );
  AND2_X1 U4929 ( .A1(n3922), .A2(n3921), .ZN(n3923) );
  NAND2_X1 U4930 ( .A1(n3924), .A2(n3923), .ZN(n4661) );
  NAND2_X1 U4931 ( .A1(n6616), .A2(n4087), .ZN(n3930) );
  AOI22_X1 U4932 ( .A1(n3926), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6655), .ZN(n3928) );
  NAND2_X1 U4933 ( .A1(n3932), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3927) );
  AND2_X1 U4934 ( .A1(n3928), .A2(n3927), .ZN(n3929) );
  NAND2_X1 U4935 ( .A1(n3930), .A2(n3929), .ZN(n4583) );
  NAND2_X1 U4936 ( .A1(n4584), .A2(n4583), .ZN(n4582) );
  OR2_X1 U4937 ( .A1(n4583), .A2(n4395), .ZN(n3931) );
  NAND2_X1 U4938 ( .A1(n4582), .A2(n3931), .ZN(n4662) );
  AND2_X2 U4939 ( .A1(n4661), .A2(n4662), .ZN(n4659) );
  OAI21_X1 U4940 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3933), .ZN(n6383) );
  AOI22_X1 U4941 ( .A1(n4430), .A2(n6383), .B1(n4401), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3935) );
  NAND2_X1 U4942 ( .A1(n4402), .A2(EAX_REG_2__SCAN_IN), .ZN(n3934) );
  OAI211_X1 U4943 ( .C1(n3950), .C2(n4601), .A(n3935), .B(n3934), .ZN(n4753)
         );
  NAND2_X1 U4944 ( .A1(n3936), .A2(n4659), .ZN(n3937) );
  NAND2_X1 U4945 ( .A1(n4798), .A2(n4087), .ZN(n3945) );
  OAI21_X1 U4946 ( .B1(n3940), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n3952), 
        .ZN(n6373) );
  AOI22_X1 U4947 ( .A1(n6373), .A2(n4430), .B1(n4401), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3942) );
  NAND2_X1 U4948 ( .A1(n3926), .A2(EAX_REG_3__SCAN_IN), .ZN(n3941) );
  OAI211_X1 U4949 ( .C1(n3950), .C2(n3939), .A(n3942), .B(n3941), .ZN(n3943)
         );
  INV_X1 U4950 ( .A(n3943), .ZN(n3944) );
  NAND2_X1 U4951 ( .A1(n3946), .A2(n4087), .ZN(n3956) );
  INV_X1 U4952 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3949) );
  OAI21_X1 U4953 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6163), .A(n6655), 
        .ZN(n3948) );
  NAND2_X1 U4954 ( .A1(n3926), .A2(EAX_REG_4__SCAN_IN), .ZN(n3947) );
  OAI211_X1 U4955 ( .C1(n3950), .C2(n3949), .A(n3948), .B(n3947), .ZN(n3954)
         );
  AOI21_X1 U4956 ( .B1(n3952), .B2(n6263), .A(n3951), .ZN(n6268) );
  NAND2_X1 U4957 ( .A1(n6268), .A2(n4430), .ZN(n3953) );
  NAND2_X1 U4958 ( .A1(n3954), .A2(n3953), .ZN(n3955) );
  NAND3_X1 U4959 ( .A1(n4752), .A2(n4766), .A3(n4758), .ZN(n4756) );
  INV_X1 U4960 ( .A(n4756), .ZN(n3957) );
  NAND2_X1 U4961 ( .A1(n3958), .A2(n3957), .ZN(n4839) );
  OAI21_X1 U4962 ( .B1(n3961), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3979), 
        .ZN(n6357) );
  NAND2_X1 U4963 ( .A1(n6357), .A2(n4430), .ZN(n3963) );
  AOI22_X1 U4964 ( .A1(n3926), .A2(EAX_REG_7__SCAN_IN), .B1(n4401), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3962) );
  NAND2_X1 U4965 ( .A1(n3963), .A2(n3962), .ZN(n3964) );
  XNOR2_X1 U4966 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3979), .ZN(n5072) );
  AOI22_X1 U4967 ( .A1(n3459), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3969) );
  INV_X1 U4968 ( .A(n3425), .ZN(n3982) );
  AOI22_X1 U4969 ( .A1(n4694), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3982), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4970 ( .A1(n3547), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4971 ( .A1(n4351), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3966) );
  NAND4_X1 U4972 ( .A1(n3969), .A2(n3968), .A3(n3967), .A4(n3966), .ZN(n3975)
         );
  AOI22_X1 U4973 ( .A1(n4229), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4974 ( .A1(n4379), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4975 ( .A1(n3461), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U4976 ( .A1(n4234), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3970) );
  NAND4_X1 U4977 ( .A1(n3973), .A2(n3972), .A3(n3971), .A4(n3970), .ZN(n3974)
         );
  OR2_X1 U4978 ( .A1(n3975), .A2(n3974), .ZN(n3976) );
  AOI22_X1 U4979 ( .A1(n4087), .A2(n3976), .B1(n4401), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3978) );
  NAND2_X1 U4980 ( .A1(n3926), .A2(EAX_REG_8__SCAN_IN), .ZN(n3977) );
  OAI211_X1 U4981 ( .C1(n5072), .C2(n4395), .A(n3978), .B(n3977), .ZN(n4975)
         );
  NAND2_X1 U4982 ( .A1(n4972), .A2(n4975), .ZN(n4973) );
  INV_X1 U4983 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3981) );
  XNOR2_X1 U4984 ( .A(n3999), .B(n3981), .ZN(n5217) );
  AOI22_X1 U4985 ( .A1(n3459), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U4986 ( .A1(n4351), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4987 ( .A1(n3982), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4988 ( .A1(n3461), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3983) );
  NAND4_X1 U4989 ( .A1(n3986), .A2(n3985), .A3(n3984), .A4(n3983), .ZN(n3992)
         );
  AOI22_X1 U4990 ( .A1(n4229), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U4991 ( .A1(n4694), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U4992 ( .A1(n4356), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U4993 ( .A1(n4234), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3987) );
  NAND4_X1 U4994 ( .A1(n3990), .A2(n3989), .A3(n3988), .A4(n3987), .ZN(n3991)
         );
  OAI21_X1 U4995 ( .B1(n3992), .B2(n3991), .A(n4087), .ZN(n3995) );
  NAND2_X1 U4996 ( .A1(n4402), .A2(EAX_REG_9__SCAN_IN), .ZN(n3994) );
  NAND2_X1 U4997 ( .A1(n4401), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3993)
         );
  NAND3_X1 U4998 ( .A1(n3995), .A2(n3994), .A3(n3993), .ZN(n3996) );
  AOI21_X1 U4999 ( .B1(n5217), .B2(n4430), .A(n3996), .ZN(n5079) );
  XOR2_X1 U5000 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n4024), .Z(n6231) );
  INV_X1 U5001 ( .A(n6231), .ZN(n5301) );
  AOI22_X1 U5002 ( .A1(n4372), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U5003 ( .A1(n4379), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U5004 ( .A1(n4351), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U5005 ( .A1(n3982), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4000) );
  NAND4_X1 U5006 ( .A1(n4003), .A2(n4002), .A3(n4001), .A4(n4000), .ZN(n4009)
         );
  AOI22_X1 U5007 ( .A1(n3459), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U5008 ( .A1(n4229), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U5009 ( .A1(n4694), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U5010 ( .A1(n4234), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4004) );
  NAND4_X1 U5011 ( .A1(n4007), .A2(n4006), .A3(n4005), .A4(n4004), .ZN(n4008)
         );
  OAI21_X1 U5012 ( .B1(n4009), .B2(n4008), .A(n4087), .ZN(n4012) );
  NAND2_X1 U5013 ( .A1(n3926), .A2(EAX_REG_10__SCAN_IN), .ZN(n4011) );
  NAND2_X1 U5014 ( .A1(n4401), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4010)
         );
  NAND3_X1 U5015 ( .A1(n4012), .A2(n4011), .A3(n4010), .ZN(n4013) );
  AOI21_X1 U5016 ( .B1(n5301), .B2(n4430), .A(n4013), .ZN(n5223) );
  AOI22_X1 U5017 ( .A1(n3460), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U5018 ( .A1(n4372), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U5019 ( .A1(n3547), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U5020 ( .A1(n4229), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4014) );
  NAND4_X1 U5021 ( .A1(n4017), .A2(n4016), .A3(n4015), .A4(n4014), .ZN(n4023)
         );
  AOI22_X1 U5022 ( .A1(n4694), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U5023 ( .A1(n4351), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U5024 ( .A1(n4234), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U5025 ( .A1(n3982), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4018) );
  NAND4_X1 U5026 ( .A1(n4021), .A2(n4020), .A3(n4019), .A4(n4018), .ZN(n4022)
         );
  NOR2_X1 U5027 ( .A1(n4023), .A2(n4022), .ZN(n4028) );
  XNOR2_X1 U5028 ( .A(n4030), .B(n4029), .ZN(n5360) );
  NAND2_X1 U5029 ( .A1(n5360), .A2(n4430), .ZN(n4026) );
  AOI22_X1 U5030 ( .A1(n3926), .A2(EAX_REG_11__SCAN_IN), .B1(n4401), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4025) );
  OAI211_X1 U5031 ( .C1(n4028), .C2(n4027), .A(n4026), .B(n4025), .ZN(n5242)
         );
  XOR2_X1 U5032 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n4044), .Z(n6222) );
  AOI22_X1 U5033 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4694), .B1(n3982), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U5034 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4372), .B1(n3460), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U5035 ( .A1(n3547), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4234), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U5036 ( .A1(n4374), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4031) );
  NAND4_X1 U5037 ( .A1(n4034), .A2(n4033), .A3(n4032), .A4(n4031), .ZN(n4040)
         );
  AOI22_X1 U5038 ( .A1(n4351), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U5039 ( .A1(n4379), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U5040 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3461), .B1(n4382), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U5041 ( .A1(n4229), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4035) );
  NAND4_X1 U5042 ( .A1(n4038), .A2(n4037), .A3(n4036), .A4(n4035), .ZN(n4039)
         );
  OR2_X1 U5043 ( .A1(n4040), .A2(n4039), .ZN(n4041) );
  AOI22_X1 U5044 ( .A1(n4087), .A2(n4041), .B1(n4401), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4043) );
  NAND2_X1 U5045 ( .A1(n3926), .A2(EAX_REG_12__SCAN_IN), .ZN(n4042) );
  OAI211_X1 U5046 ( .C1(n6222), .C2(n4395), .A(n4043), .B(n4042), .ZN(n5258)
         );
  INV_X1 U5047 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4045) );
  XNOR2_X1 U5048 ( .A(n4061), .B(n4045), .ZN(n5820) );
  NAND2_X1 U5049 ( .A1(n5820), .A2(n4430), .ZN(n4047) );
  AOI22_X1 U5050 ( .A1(n3926), .A2(EAX_REG_13__SCAN_IN), .B1(n4401), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4046) );
  NAND2_X1 U5051 ( .A1(n4047), .A2(n4046), .ZN(n4059) );
  XNOR2_X2 U5052 ( .A(n5257), .B(n4059), .ZN(n5501) );
  AOI22_X1 U5053 ( .A1(n4229), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U5054 ( .A1(n4379), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4234), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4050) );
  AOI22_X1 U5055 ( .A1(n4356), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U5056 ( .A1(n4694), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4048) );
  NAND4_X1 U5057 ( .A1(n4051), .A2(n4050), .A3(n4049), .A4(n4048), .ZN(n4057)
         );
  AOI22_X1 U5058 ( .A1(n4351), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3982), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U5059 ( .A1(n3461), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U5060 ( .A1(n3459), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U5061 ( .A1(n3547), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4052) );
  NAND4_X1 U5062 ( .A1(n4055), .A2(n4054), .A3(n4053), .A4(n4052), .ZN(n4056)
         );
  OR2_X1 U5063 ( .A1(n4057), .A2(n4056), .ZN(n4058) );
  AND2_X1 U5064 ( .A1(n4087), .A2(n4058), .ZN(n5500) );
  NAND2_X1 U5065 ( .A1(n5501), .A2(n5500), .ZN(n5499) );
  INV_X1 U5066 ( .A(n4059), .ZN(n4060) );
  NAND2_X1 U5067 ( .A1(n5499), .A2(n5543), .ZN(n4077) );
  XNOR2_X1 U5068 ( .A(n4078), .B(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6212)
         );
  NAND2_X1 U5069 ( .A1(n6212), .A2(n4430), .ZN(n4076) );
  AOI22_X1 U5070 ( .A1(n3460), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U5071 ( .A1(n4356), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5072 ( .A1(n3547), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U5073 ( .A1(n4374), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4062) );
  NAND4_X1 U5074 ( .A1(n4065), .A2(n4064), .A3(n4063), .A4(n4062), .ZN(n4071)
         );
  AOI22_X1 U5075 ( .A1(n4229), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U5076 ( .A1(n4351), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4234), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U5077 ( .A1(n3982), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U5078 ( .A1(n4694), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4066) );
  NAND4_X1 U5079 ( .A1(n4069), .A2(n4068), .A3(n4067), .A4(n4066), .ZN(n4070)
         );
  OAI21_X1 U5080 ( .B1(n4071), .B2(n4070), .A(n4087), .ZN(n4074) );
  NAND2_X1 U5081 ( .A1(n4402), .A2(EAX_REG_14__SCAN_IN), .ZN(n4073) );
  NAND2_X1 U5082 ( .A1(n4401), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4072)
         );
  AND3_X1 U5083 ( .A1(n4074), .A2(n4073), .A3(n4072), .ZN(n4075) );
  NAND2_X1 U5084 ( .A1(n4076), .A2(n4075), .ZN(n5542) );
  NAND2_X1 U5085 ( .A1(n4077), .A2(n5542), .ZN(n5540) );
  INV_X1 U5086 ( .A(n5540), .ZN(n4096) );
  XNOR2_X1 U5087 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n4098), .ZN(n5807)
         );
  INV_X1 U5088 ( .A(n5807), .ZN(n4094) );
  AOI22_X1 U5089 ( .A1(n4694), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U5090 ( .A1(n3460), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4234), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U5091 ( .A1(n3461), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4080) );
  AOI22_X1 U5092 ( .A1(n4229), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4079) );
  NAND4_X1 U5093 ( .A1(n4082), .A2(n4081), .A3(n4080), .A4(n4079), .ZN(n4089)
         );
  AOI22_X1 U5094 ( .A1(n3982), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U5095 ( .A1(n4372), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U5096 ( .A1(n4356), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U5097 ( .A1(n4351), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4083) );
  NAND4_X1 U5098 ( .A1(n4086), .A2(n4085), .A3(n4084), .A4(n4083), .ZN(n4088)
         );
  OAI21_X1 U5099 ( .B1(n4089), .B2(n4088), .A(n4087), .ZN(n4092) );
  NAND2_X1 U5100 ( .A1(n4402), .A2(EAX_REG_15__SCAN_IN), .ZN(n4091) );
  NAND2_X1 U5101 ( .A1(n4401), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4090)
         );
  NAND3_X1 U5102 ( .A1(n4092), .A2(n4091), .A3(n4090), .ZN(n4093) );
  AOI21_X1 U5103 ( .B1(n4094), .B2(n4430), .A(n4093), .ZN(n5551) );
  XNOR2_X1 U5104 ( .A(n4127), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6202)
         );
  AOI22_X1 U5105 ( .A1(n4228), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5106 ( .A1(n4229), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U5107 ( .A1(n4351), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U5108 ( .A1(n3461), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4099) );
  NAND4_X1 U5109 ( .A1(n4102), .A2(n4101), .A3(n4100), .A4(n4099), .ZN(n4108)
         );
  AOI22_X1 U5110 ( .A1(n3459), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4234), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U5111 ( .A1(n4372), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U5112 ( .A1(n4356), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5113 ( .A1(n4694), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4103) );
  NAND4_X1 U5114 ( .A1(n4106), .A2(n4105), .A3(n4104), .A4(n4103), .ZN(n4107)
         );
  NOR2_X1 U5115 ( .A1(n4108), .A2(n4107), .ZN(n4110) );
  AOI22_X1 U5116 ( .A1(n3926), .A2(EAX_REG_16__SCAN_IN), .B1(n4401), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4109) );
  OAI21_X1 U5117 ( .B1(n4367), .B2(n4110), .A(n4109), .ZN(n4111) );
  AOI21_X1 U5118 ( .B1(n6202), .B2(n4430), .A(n4111), .ZN(n5704) );
  AOI22_X1 U5119 ( .A1(n4356), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4116) );
  AOI22_X1 U5120 ( .A1(n4229), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4115) );
  AOI22_X1 U5121 ( .A1(n4351), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4234), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4114) );
  AOI22_X1 U5122 ( .A1(n3982), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4113) );
  NAND4_X1 U5123 ( .A1(n4116), .A2(n4115), .A3(n4114), .A4(n4113), .ZN(n4122)
         );
  AOI22_X1 U5124 ( .A1(n3460), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U5125 ( .A1(n4694), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4119) );
  AOI22_X1 U5126 ( .A1(n3461), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U5127 ( .A1(n4381), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4117) );
  NAND4_X1 U5128 ( .A1(n4120), .A2(n4119), .A3(n4118), .A4(n4117), .ZN(n4121)
         );
  NOR2_X1 U5129 ( .A1(n4122), .A2(n4121), .ZN(n4126) );
  NAND2_X1 U5130 ( .A1(n6655), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4123)
         );
  NAND2_X1 U5131 ( .A1(n4395), .A2(n4123), .ZN(n4124) );
  AOI21_X1 U5132 ( .B1(n4402), .B2(EAX_REG_17__SCAN_IN), .A(n4124), .ZN(n4125)
         );
  OAI21_X1 U5133 ( .B1(n4367), .B2(n4126), .A(n4125), .ZN(n4130) );
  OAI21_X1 U5134 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4128), .A(n4146), 
        .ZN(n6196) );
  OR2_X1 U5135 ( .A1(n4395), .A2(n6196), .ZN(n4129) );
  NAND2_X1 U5136 ( .A1(n4130), .A2(n4129), .ZN(n6106) );
  AOI22_X1 U5137 ( .A1(n4229), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U5138 ( .A1(n4351), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U5139 ( .A1(n4228), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U5140 ( .A1(n4694), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4131) );
  NAND4_X1 U5141 ( .A1(n4134), .A2(n4133), .A3(n4132), .A4(n4131), .ZN(n4140)
         );
  AOI22_X1 U5142 ( .A1(n3460), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U5143 ( .A1(n3461), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4137) );
  AOI22_X1 U5144 ( .A1(n4234), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U5145 ( .A1(n4356), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4135) );
  NAND4_X1 U5146 ( .A1(n4138), .A2(n4137), .A3(n4136), .A4(n4135), .ZN(n4139)
         );
  NOR2_X1 U5147 ( .A1(n4140), .A2(n4139), .ZN(n4143) );
  INV_X1 U5148 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5794) );
  AOI21_X1 U5149 ( .B1(n5794), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4141) );
  AOI21_X1 U5150 ( .B1(n4402), .B2(EAX_REG_18__SCAN_IN), .A(n4141), .ZN(n4142)
         );
  OAI21_X1 U5151 ( .B1(n4367), .B2(n4143), .A(n4142), .ZN(n4145) );
  XNOR2_X1 U5152 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4146), .ZN(n6183)
         );
  NAND2_X1 U5153 ( .A1(n4430), .A2(n6183), .ZN(n4144) );
  NAND2_X1 U5154 ( .A1(n5695), .A2(n5698), .ZN(n5697) );
  INV_X1 U5155 ( .A(n5697), .ZN(n4165) );
  OR2_X1 U5156 ( .A1(n4147), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4148)
         );
  NAND2_X1 U5157 ( .A1(n4148), .A2(n4196), .ZN(n6098) );
  AOI22_X1 U5158 ( .A1(n4229), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4152) );
  AOI22_X1 U5159 ( .A1(n4694), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4151) );
  AOI22_X1 U5160 ( .A1(n4351), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U5161 ( .A1(n4234), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4149) );
  NAND4_X1 U5162 ( .A1(n4152), .A2(n4151), .A3(n4150), .A4(n4149), .ZN(n4158)
         );
  AOI22_X1 U5163 ( .A1(n3460), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4156) );
  AOI22_X1 U5164 ( .A1(n3547), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U5165 ( .A1(n4372), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5166 ( .A1(n4356), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4153) );
  NAND4_X1 U5167 ( .A1(n4156), .A2(n4155), .A3(n4154), .A4(n4153), .ZN(n4157)
         );
  NOR2_X1 U5168 ( .A1(n4158), .A2(n4157), .ZN(n4159) );
  NOR2_X1 U5169 ( .A1(n4367), .A2(n4159), .ZN(n4163) );
  INV_X1 U5170 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4519) );
  NAND2_X1 U5171 ( .A1(n6655), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4160)
         );
  OAI211_X1 U5172 ( .C1(n4161), .C2(n4519), .A(n4395), .B(n4160), .ZN(n4162)
         );
  OAI22_X1 U5173 ( .A1(n6098), .A2(n4395), .B1(n4163), .B2(n4162), .ZN(n6057)
         );
  NAND2_X1 U5174 ( .A1(n4165), .A2(n4164), .ZN(n5680) );
  AOI22_X1 U5175 ( .A1(n4229), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U5176 ( .A1(n4351), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U5177 ( .A1(n3982), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4167) );
  AOI22_X1 U5178 ( .A1(n4694), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4166) );
  NAND4_X1 U5179 ( .A1(n4169), .A2(n4168), .A3(n4167), .A4(n4166), .ZN(n4175)
         );
  AOI22_X1 U5180 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n3460), .B1(n4372), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4173) );
  AOI22_X1 U5181 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n3481), .B1(n4381), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4172) );
  AOI22_X1 U5182 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4234), .B1(n4374), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4171) );
  AOI22_X1 U5183 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4356), .B1(n4382), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4170) );
  NAND4_X1 U5184 ( .A1(n4173), .A2(n4172), .A3(n4171), .A4(n4170), .ZN(n4174)
         );
  NOR2_X1 U5185 ( .A1(n4175), .A2(n4174), .ZN(n4179) );
  INV_X1 U5186 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4176) );
  AOI21_X1 U5187 ( .B1(n4176), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4177) );
  AOI21_X1 U5188 ( .B1(n4402), .B2(EAX_REG_20__SCAN_IN), .A(n4177), .ZN(n4178)
         );
  OAI21_X1 U5189 ( .B1(n4367), .B2(n4179), .A(n4178), .ZN(n4181) );
  XNOR2_X1 U5190 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n4196), .ZN(n6044)
         );
  NAND2_X1 U5191 ( .A1(n6044), .A2(n4430), .ZN(n4180) );
  NAND2_X1 U5192 ( .A1(n4181), .A2(n4180), .ZN(n5682) );
  NOR2_X2 U5193 ( .A1(n5680), .A2(n5682), .ZN(n5674) );
  AOI22_X1 U5194 ( .A1(n3982), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4185) );
  AOI22_X1 U5195 ( .A1(n4356), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4234), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4184) );
  AOI22_X1 U5196 ( .A1(n4694), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4183) );
  AOI22_X1 U5197 ( .A1(n4372), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4182) );
  NAND4_X1 U5198 ( .A1(n4185), .A2(n4184), .A3(n4183), .A4(n4182), .ZN(n4191)
         );
  AOI22_X1 U5199 ( .A1(n4351), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4189) );
  AOI22_X1 U5200 ( .A1(n3460), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4188) );
  AOI22_X1 U5201 ( .A1(n4229), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4187) );
  AOI22_X1 U5202 ( .A1(n3481), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4186) );
  NAND4_X1 U5203 ( .A1(n4189), .A2(n4188), .A3(n4187), .A4(n4186), .ZN(n4190)
         );
  NOR2_X1 U5204 ( .A1(n4191), .A2(n4190), .ZN(n4195) );
  NAND2_X1 U5205 ( .A1(n6655), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4192)
         );
  NAND2_X1 U5206 ( .A1(n4395), .A2(n4192), .ZN(n4193) );
  AOI21_X1 U5207 ( .B1(n4402), .B2(EAX_REG_21__SCAN_IN), .A(n4193), .ZN(n4194)
         );
  OAI21_X1 U5208 ( .B1(n4367), .B2(n4195), .A(n4194), .ZN(n4200) );
  OAI21_X1 U5209 ( .B1(n4198), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n4245), 
        .ZN(n6034) );
  OR2_X1 U5210 ( .A1(n6034), .A2(n4395), .ZN(n4199) );
  NAND2_X1 U5211 ( .A1(n5674), .A2(n5673), .ZN(n5669) );
  AOI22_X1 U5212 ( .A1(n3460), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4204) );
  AOI22_X1 U5213 ( .A1(n4356), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4203) );
  AOI22_X1 U5214 ( .A1(n3982), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4202) );
  AOI22_X1 U5215 ( .A1(n4372), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4201) );
  NAND4_X1 U5216 ( .A1(n4204), .A2(n4203), .A3(n4202), .A4(n4201), .ZN(n4210)
         );
  AOI22_X1 U5217 ( .A1(n4384), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3481), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4208) );
  AOI22_X1 U5218 ( .A1(n4380), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4207) );
  AOI22_X1 U5219 ( .A1(n4694), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4206) );
  AOI22_X1 U5220 ( .A1(n4234), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4205) );
  NAND4_X1 U5221 ( .A1(n4208), .A2(n4207), .A3(n4206), .A4(n4205), .ZN(n4209)
         );
  NOR2_X1 U5222 ( .A1(n4210), .A2(n4209), .ZN(n4213) );
  OAI21_X1 U5223 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5772), .A(n4395), .ZN(
        n4211) );
  AOI21_X1 U5224 ( .B1(n4402), .B2(EAX_REG_22__SCAN_IN), .A(n4211), .ZN(n4212)
         );
  OAI21_X1 U5225 ( .B1(n4367), .B2(n4213), .A(n4212), .ZN(n4215) );
  XNOR2_X1 U5226 ( .A(n4245), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6024)
         );
  NAND2_X1 U5227 ( .A1(n6024), .A2(n4430), .ZN(n4214) );
  NAND2_X1 U5228 ( .A1(n4215), .A2(n4214), .ZN(n5670) );
  AOI22_X1 U5229 ( .A1(n3460), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4221) );
  AOI22_X1 U5230 ( .A1(n4694), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4234), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U5231 ( .A1(n4351), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4219) );
  AOI22_X1 U5232 ( .A1(n4372), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4218) );
  NAND4_X1 U5233 ( .A1(n4221), .A2(n4220), .A3(n4219), .A4(n4218), .ZN(n4227)
         );
  AOI22_X1 U5234 ( .A1(n4379), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4225) );
  AOI22_X1 U5235 ( .A1(n3461), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4224) );
  AOI22_X1 U5236 ( .A1(n4356), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4223) );
  AOI22_X1 U5237 ( .A1(n4229), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4222) );
  NAND4_X1 U5238 ( .A1(n4225), .A2(n4224), .A3(n4223), .A4(n4222), .ZN(n4226)
         );
  NOR2_X1 U5239 ( .A1(n4227), .A2(n4226), .ZN(n4250) );
  AOI22_X1 U5240 ( .A1(n4228), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4233) );
  AOI22_X1 U5241 ( .A1(n4229), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4232) );
  AOI22_X1 U5242 ( .A1(n4694), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4231) );
  AOI22_X1 U5243 ( .A1(n4351), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4230) );
  NAND4_X1 U5244 ( .A1(n4233), .A2(n4232), .A3(n4231), .A4(n4230), .ZN(n4240)
         );
  AOI22_X1 U5245 ( .A1(n3460), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4238) );
  AOI22_X1 U5246 ( .A1(n4234), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4237) );
  AOI22_X1 U5247 ( .A1(n4356), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4236) );
  AOI22_X1 U5248 ( .A1(n3461), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4235) );
  NAND4_X1 U5249 ( .A1(n4238), .A2(n4237), .A3(n4236), .A4(n4235), .ZN(n4239)
         );
  NOR2_X1 U5250 ( .A1(n4240), .A2(n4239), .ZN(n4251) );
  XNOR2_X1 U5251 ( .A(n4250), .B(n4251), .ZN(n4244) );
  NAND2_X1 U5252 ( .A1(n6655), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4241)
         );
  NAND2_X1 U5253 ( .A1(n4395), .A2(n4241), .ZN(n4242) );
  AOI21_X1 U5254 ( .B1(n4402), .B2(EAX_REG_23__SCAN_IN), .A(n4242), .ZN(n4243)
         );
  OAI21_X1 U5255 ( .B1(n4367), .B2(n4244), .A(n4243), .ZN(n4249) );
  OR2_X1 U5256 ( .A1(n4246), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4247)
         );
  NAND2_X1 U5257 ( .A1(n4285), .A2(n4247), .ZN(n6017) );
  NAND2_X1 U5258 ( .A1(n4249), .A2(n4248), .ZN(n4420) );
  NOR2_X1 U5259 ( .A1(n4251), .A2(n4250), .ZN(n4269) );
  AOI22_X1 U5260 ( .A1(n4229), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4255) );
  AOI22_X1 U5261 ( .A1(n4351), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4254) );
  AOI22_X1 U5262 ( .A1(n3982), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4253) );
  AOI22_X1 U5263 ( .A1(n4694), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4252) );
  NAND4_X1 U5264 ( .A1(n4255), .A2(n4254), .A3(n4253), .A4(n4252), .ZN(n4261)
         );
  AOI22_X1 U5265 ( .A1(n3459), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4259) );
  AOI22_X1 U5266 ( .A1(n3461), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4258) );
  AOI22_X1 U5267 ( .A1(n4234), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4257) );
  AOI22_X1 U5268 ( .A1(n4356), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4256) );
  NAND4_X1 U5269 ( .A1(n4259), .A2(n4258), .A3(n4257), .A4(n4256), .ZN(n4260)
         );
  INV_X1 U5270 ( .A(n4268), .ZN(n4262) );
  XNOR2_X1 U5271 ( .A(n4269), .B(n4262), .ZN(n4266) );
  XNOR2_X1 U5272 ( .A(n4285), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6009)
         );
  NAND2_X1 U5273 ( .A1(n4402), .A2(EAX_REG_24__SCAN_IN), .ZN(n4264) );
  NAND2_X1 U5274 ( .A1(n4401), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4263)
         );
  OAI211_X1 U5275 ( .C1(n6009), .C2(n4395), .A(n4264), .B(n4263), .ZN(n4265)
         );
  AOI21_X1 U5276 ( .B1(n4266), .B2(n4393), .A(n4265), .ZN(n5659) );
  NAND2_X1 U5277 ( .A1(n4269), .A2(n4268), .ZN(n4290) );
  AOI22_X1 U5278 ( .A1(n4351), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4273) );
  AOI22_X1 U5279 ( .A1(n3547), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4272) );
  AOI22_X1 U5280 ( .A1(n4372), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4271) );
  AOI22_X1 U5281 ( .A1(n4229), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4270) );
  NAND4_X1 U5282 ( .A1(n4273), .A2(n4272), .A3(n4271), .A4(n4270), .ZN(n4279)
         );
  AOI22_X1 U5283 ( .A1(n3982), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4277) );
  AOI22_X1 U5284 ( .A1(n4694), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4276) );
  AOI22_X1 U5285 ( .A1(n3461), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4234), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4275) );
  AOI22_X1 U5286 ( .A1(n4381), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4274) );
  NAND4_X1 U5287 ( .A1(n4277), .A2(n4276), .A3(n4275), .A4(n4274), .ZN(n4278)
         );
  NOR2_X1 U5288 ( .A1(n4279), .A2(n4278), .ZN(n4291) );
  XNOR2_X1 U5289 ( .A(n4290), .B(n4291), .ZN(n4283) );
  NAND2_X1 U5290 ( .A1(n6655), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4280)
         );
  NAND2_X1 U5291 ( .A1(n4395), .A2(n4280), .ZN(n4281) );
  AOI21_X1 U5292 ( .B1(n4402), .B2(EAX_REG_25__SCAN_IN), .A(n4281), .ZN(n4282)
         );
  OAI21_X1 U5293 ( .B1(n4283), .B2(n4367), .A(n4282), .ZN(n4289) );
  INV_X1 U5294 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4284) );
  OR2_X1 U5295 ( .A1(n4286), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4287)
         );
  NAND2_X1 U5296 ( .A1(n4287), .A2(n4325), .ZN(n6090) );
  NOR2_X1 U5297 ( .A1(n4291), .A2(n4290), .ZN(n4320) );
  AOI22_X1 U5298 ( .A1(n4229), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4295) );
  AOI22_X1 U5299 ( .A1(n4351), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4294) );
  AOI22_X1 U5300 ( .A1(n3982), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4293) );
  AOI22_X1 U5301 ( .A1(n4694), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4292) );
  NAND4_X1 U5302 ( .A1(n4295), .A2(n4294), .A3(n4293), .A4(n4292), .ZN(n4301)
         );
  AOI22_X1 U5303 ( .A1(n3460), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4299) );
  AOI22_X1 U5304 ( .A1(n3481), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4298) );
  AOI22_X1 U5305 ( .A1(n4234), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4297) );
  AOI22_X1 U5306 ( .A1(n4356), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4296) );
  NAND4_X1 U5307 ( .A1(n4299), .A2(n4298), .A3(n4297), .A4(n4296), .ZN(n4300)
         );
  OR2_X1 U5308 ( .A1(n4301), .A2(n4300), .ZN(n4319) );
  INV_X1 U5309 ( .A(n4319), .ZN(n4302) );
  XNOR2_X1 U5310 ( .A(n4320), .B(n4302), .ZN(n4303) );
  NAND2_X1 U5311 ( .A1(n4303), .A2(n4393), .ZN(n4308) );
  NAND2_X1 U5312 ( .A1(n6655), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4304)
         );
  NAND2_X1 U5313 ( .A1(n4395), .A2(n4304), .ZN(n4305) );
  AOI21_X1 U5314 ( .B1(n4402), .B2(EAX_REG_26__SCAN_IN), .A(n4305), .ZN(n4307)
         );
  XNOR2_X1 U5315 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .B(n4325), .ZN(n6000)
         );
  AOI22_X1 U5316 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4229), .B1(n3460), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4312) );
  AOI22_X1 U5317 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4694), .B1(n4234), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4311) );
  AOI22_X1 U5318 ( .A1(n4379), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4310) );
  AOI22_X1 U5319 ( .A1(n3476), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4309) );
  NAND4_X1 U5320 ( .A1(n4312), .A2(n4311), .A3(n4310), .A4(n4309), .ZN(n4318)
         );
  AOI22_X1 U5321 ( .A1(n4351), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3481), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4316) );
  AOI22_X1 U5322 ( .A1(n4372), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4315) );
  AOI22_X1 U5323 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4356), .B1(n4382), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4314) );
  AOI22_X1 U5324 ( .A1(n3982), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4313) );
  NAND4_X1 U5325 ( .A1(n4316), .A2(n4315), .A3(n4314), .A4(n4313), .ZN(n4317)
         );
  NOR2_X1 U5326 ( .A1(n4318), .A2(n4317), .ZN(n4341) );
  NAND2_X1 U5327 ( .A1(n4320), .A2(n4319), .ZN(n4340) );
  XNOR2_X1 U5328 ( .A(n4341), .B(n4340), .ZN(n4324) );
  NAND2_X1 U5329 ( .A1(n6655), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4321)
         );
  NAND2_X1 U5330 ( .A1(n4395), .A2(n4321), .ZN(n4322) );
  AOI21_X1 U5331 ( .B1(n4402), .B2(EAX_REG_27__SCAN_IN), .A(n4322), .ZN(n4323)
         );
  OAI21_X1 U5332 ( .B1(n4324), .B2(n4367), .A(n4323), .ZN(n4329) );
  INV_X1 U5333 ( .A(n4325), .ZN(n4326) );
  OAI21_X1 U5334 ( .B1(n4327), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n4346), 
        .ZN(n5993) );
  OR2_X1 U5335 ( .A1(n5993), .A2(n4395), .ZN(n4328) );
  NAND2_X1 U5336 ( .A1(n4329), .A2(n4328), .ZN(n5648) );
  AOI22_X1 U5337 ( .A1(n4229), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4333) );
  AOI22_X1 U5338 ( .A1(n4351), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4332) );
  AOI22_X1 U5339 ( .A1(n3982), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4331) );
  AOI22_X1 U5340 ( .A1(n4694), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4330) );
  NAND4_X1 U5341 ( .A1(n4333), .A2(n4332), .A3(n4331), .A4(n4330), .ZN(n4339)
         );
  AOI22_X1 U5342 ( .A1(n3460), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4337) );
  AOI22_X1 U5343 ( .A1(n3481), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4336) );
  AOI22_X1 U5344 ( .A1(n4234), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4335) );
  AOI22_X1 U5345 ( .A1(n4356), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4334) );
  NAND4_X1 U5346 ( .A1(n4337), .A2(n4336), .A3(n4335), .A4(n4334), .ZN(n4338)
         );
  OR2_X1 U5347 ( .A1(n4339), .A2(n4338), .ZN(n4363) );
  NOR2_X1 U5348 ( .A1(n4341), .A2(n4340), .ZN(n4364) );
  XOR2_X1 U5349 ( .A(n4363), .B(n4364), .Z(n4342) );
  NAND2_X1 U5350 ( .A1(n4342), .A2(n4393), .ZN(n4345) );
  INV_X1 U5351 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5568) );
  AOI21_X1 U5352 ( .B1(n5568), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4343) );
  AOI21_X1 U5353 ( .B1(n4402), .B2(EAX_REG_28__SCAN_IN), .A(n4343), .ZN(n4344)
         );
  XNOR2_X1 U5354 ( .A(n4346), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5983)
         );
  INV_X1 U5355 ( .A(n4347), .ZN(n4349) );
  INV_X1 U5356 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4348) );
  NAND2_X1 U5357 ( .A1(n4349), .A2(n4348), .ZN(n4350) );
  NAND2_X1 U5358 ( .A1(n4411), .A2(n4350), .ZN(n5742) );
  AOI22_X1 U5359 ( .A1(n4351), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4355) );
  AOI22_X1 U5360 ( .A1(n3481), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4354) );
  AOI22_X1 U5361 ( .A1(n4372), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4353) );
  AOI22_X1 U5362 ( .A1(n3982), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4352) );
  NAND4_X1 U5363 ( .A1(n4355), .A2(n4354), .A3(n4353), .A4(n4352), .ZN(n4362)
         );
  AOI22_X1 U5364 ( .A1(n4229), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4360) );
  AOI22_X1 U5365 ( .A1(n4694), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4234), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4359) );
  AOI22_X1 U5366 ( .A1(n4379), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4358) );
  AOI22_X1 U5367 ( .A1(n3476), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4357) );
  NAND4_X1 U5368 ( .A1(n4360), .A2(n4359), .A3(n4358), .A4(n4357), .ZN(n4361)
         );
  NOR2_X1 U5369 ( .A1(n4362), .A2(n4361), .ZN(n4371) );
  NAND2_X1 U5370 ( .A1(n4364), .A2(n4363), .ZN(n4370) );
  XNOR2_X1 U5371 ( .A(n4371), .B(n4370), .ZN(n4368) );
  AOI21_X1 U5372 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6655), .A(n4430), 
        .ZN(n4366) );
  NAND2_X1 U5373 ( .A1(n4402), .A2(EAX_REG_29__SCAN_IN), .ZN(n4365) );
  OAI211_X1 U5374 ( .C1(n4368), .C2(n4367), .A(n4366), .B(n4365), .ZN(n4369)
         );
  OAI21_X1 U5375 ( .B1(n4395), .B2(n5742), .A(n4369), .ZN(n5620) );
  NOR2_X1 U5376 ( .A1(n4371), .A2(n4370), .ZN(n4392) );
  AOI22_X1 U5377 ( .A1(n3459), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4378) );
  AOI22_X1 U5378 ( .A1(n3982), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3481), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4377) );
  AOI22_X1 U5379 ( .A1(n3476), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4373), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4376) );
  AOI22_X1 U5380 ( .A1(n4234), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4374), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4375) );
  NAND4_X1 U5381 ( .A1(n4378), .A2(n4377), .A3(n4376), .A4(n4375), .ZN(n4390)
         );
  AOI22_X1 U5382 ( .A1(n4380), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4379), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4388) );
  AOI22_X1 U5383 ( .A1(n4694), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4387) );
  AOI22_X1 U5384 ( .A1(n4356), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4382), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4386) );
  AOI22_X1 U5385 ( .A1(n4384), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4385) );
  NAND4_X1 U5386 ( .A1(n4388), .A2(n4387), .A3(n4386), .A4(n4385), .ZN(n4389)
         );
  NOR2_X1 U5387 ( .A1(n4390), .A2(n4389), .ZN(n4391) );
  XNOR2_X1 U5388 ( .A(n4392), .B(n4391), .ZN(n4394) );
  NAND2_X1 U5389 ( .A1(n4394), .A2(n4393), .ZN(n4400) );
  INV_X1 U5390 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5733) );
  OAI21_X1 U5391 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5733), .A(n4395), .ZN(
        n4396) );
  AOI21_X1 U5392 ( .B1(n4402), .B2(EAX_REG_30__SCAN_IN), .A(n4396), .ZN(n4399)
         );
  XNOR2_X1 U5393 ( .A(n4411), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5731)
         );
  AND2_X1 U5394 ( .A1(n5731), .A2(n4397), .ZN(n4398) );
  AOI22_X1 U5395 ( .A1(n4402), .A2(EAX_REG_31__SCAN_IN), .B1(n4401), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4403) );
  INV_X1 U5396 ( .A(n4403), .ZN(n4404) );
  AND2_X1 U5397 ( .A1(n6656), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4431) );
  NAND2_X1 U5398 ( .A1(n4431), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6663) );
  NAND2_X1 U5399 ( .A1(n5584), .A2(n6378), .ZN(n4417) );
  NAND2_X1 U5400 ( .A1(n4406), .A2(n6543), .ZN(n6742) );
  NAND2_X1 U5401 ( .A1(n6742), .A2(n6656), .ZN(n4407) );
  NAND2_X1 U5402 ( .A1(n6656), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4409) );
  NAND2_X1 U5403 ( .A1(n6163), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4408) );
  AND2_X1 U5404 ( .A1(n4409), .A2(n4408), .ZN(n4653) );
  INV_X1 U5405 ( .A(n4653), .ZN(n4410) );
  INV_X1 U5406 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4412) );
  NAND2_X1 U5407 ( .A1(n6457), .A2(REIP_REG_31__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U5408 ( .A1(n6374), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4414)
         );
  OAI211_X1 U5409 ( .C1(n6384), .C2(n4870), .A(n5832), .B(n4414), .ZN(n4415)
         );
  INV_X1 U5410 ( .A(n4415), .ZN(n4416) );
  OAI211_X1 U5411 ( .C1(n5843), .C2(n6164), .A(n4417), .B(n4416), .ZN(U2955)
         );
  NAND2_X1 U5412 ( .A1(n4418), .A2(n6380), .ZN(n4427) );
  NAND2_X1 U5413 ( .A1(n4419), .A2(n4420), .ZN(n4421) );
  NAND2_X1 U5414 ( .A1(n3164), .A2(n4421), .ZN(n6019) );
  NOR2_X1 U5415 ( .A1(n6384), .A2(n6017), .ZN(n4422) );
  AOI211_X1 U5416 ( .C1(n6374), .C2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n4423), 
        .B(n4422), .ZN(n4424) );
  NAND2_X1 U5417 ( .A1(n4427), .A2(n4426), .ZN(U2963) );
  AND2_X1 U5418 ( .A1(n4431), .A2(n4430), .ZN(n6654) );
  OR2_X1 U5419 ( .A1(n6457), .A2(n6654), .ZN(n4432) );
  NAND2_X1 U5420 ( .A1(n4712), .A2(n6655), .ZN(n6647) );
  NOR3_X1 U5421 ( .A1(n6656), .A2(n6722), .A3(n6647), .ZN(n6645) );
  NOR2_X1 U5422 ( .A1(n4870), .A2(n4712), .ZN(n4434) );
  INV_X1 U5423 ( .A(REIP_REG_28__SCAN_IN), .ZN(n7067) );
  INV_X1 U5424 ( .A(REIP_REG_27__SCAN_IN), .ZN(n7051) );
  NAND2_X1 U5425 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5633) );
  INV_X1 U5426 ( .A(REIP_REG_20__SCAN_IN), .ZN(n7078) );
  INV_X1 U5427 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6702) );
  INV_X1 U5428 ( .A(REIP_REG_18__SCAN_IN), .ZN(n7045) );
  NOR3_X1 U5429 ( .A1(n7078), .A2(n6702), .A3(n7045), .ZN(n4481) );
  NAND2_X1 U5430 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n6197) );
  NOR2_X1 U5431 ( .A1(STATEBS16_REG_SCAN_IN), .A2(READY_N), .ZN(n4475) );
  AND3_X1 U5432 ( .A1(n4435), .A2(n4475), .A3(n4874), .ZN(n4436) );
  INV_X1 U5433 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6694) );
  INV_X1 U5434 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6689) );
  INV_X1 U5435 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6688) );
  INV_X1 U5436 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6684) );
  NAND3_X1 U5437 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6270) );
  NOR2_X1 U5438 ( .A1(n6684), .A2(n6270), .ZN(n6253) );
  AND2_X1 U5439 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6253), .ZN(n4881) );
  NAND2_X1 U5440 ( .A1(REIP_REG_6__SCAN_IN), .A2(n4881), .ZN(n6239) );
  OR2_X1 U5441 ( .A1(n6688), .A2(n6239), .ZN(n4982) );
  NOR2_X1 U5442 ( .A1(n6689), .A2(n4982), .ZN(n5086) );
  NAND4_X1 U5443 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5086), .A3(
        REIP_REG_10__SCAN_IN), .A4(REIP_REG_9__SCAN_IN), .ZN(n5512) );
  NOR2_X1 U5444 ( .A1(n6694), .A2(n5512), .ZN(n5514) );
  NAND2_X1 U5445 ( .A1(REIP_REG_13__SCAN_IN), .A2(n5514), .ZN(n4480) );
  NAND2_X1 U5446 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6207), .ZN(n6200) );
  NAND2_X1 U5447 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6188), .ZN(n6180) );
  NAND4_X1 U5448 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n6036), .ZN(n6011) );
  NOR2_X1 U5449 ( .A1(n5633), .A2(n6011), .ZN(n6004) );
  NAND2_X1 U5450 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6004), .ZN(n5999) );
  NOR3_X1 U5451 ( .A1(n7067), .A2(n7051), .A3(n5999), .ZN(n4488) );
  INV_X1 U5452 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6913) );
  INV_X1 U5453 ( .A(REIP_REG_29__SCAN_IN), .ZN(n7097) );
  NOR3_X1 U5454 ( .A1(n6913), .A2(n7097), .A3(REIP_REG_31__SCAN_IN), .ZN(n4478) );
  AND2_X1 U5455 ( .A1(n4666), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4437)
         );
  AOI21_X1 U5456 ( .B1(n4470), .B2(EBX_REG_30__SCAN_IN), .A(n4437), .ZN(n4501)
         );
  MUX2_X1 U5457 ( .A(n4438), .B(n4455), .S(EBX_REG_24__SCAN_IN), .Z(n4442) );
  NAND2_X1 U5458 ( .A1(n4666), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4439) );
  AND2_X1 U5459 ( .A1(n4440), .A2(n4439), .ZN(n4441) );
  NAND2_X1 U5460 ( .A1(n4442), .A2(n4441), .ZN(n5660) );
  MUX2_X1 U5461 ( .A(n4449), .B(n5685), .S(EBX_REG_25__SCAN_IN), .Z(n4444) );
  NAND2_X1 U5462 ( .A1(n4581), .A2(n6115), .ZN(n4443) );
  NAND2_X1 U5463 ( .A1(n4444), .A2(n4443), .ZN(n5636) );
  INV_X1 U5464 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U5465 ( .A1(n4453), .A2(n6008), .ZN(n4448) );
  INV_X1 U5466 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U5467 ( .A1(n4455), .A2(n5885), .ZN(n4446) );
  NAND2_X1 U5468 ( .A1(n4465), .A2(n6008), .ZN(n4445) );
  NAND3_X1 U5469 ( .A1(n4446), .A2(n5685), .A3(n4445), .ZN(n4447) );
  MUX2_X1 U5470 ( .A(n4449), .B(n5685), .S(EBX_REG_27__SCAN_IN), .Z(n4451) );
  NAND2_X1 U5471 ( .A1(n4581), .A2(n5749), .ZN(n4450) );
  NAND2_X1 U5472 ( .A1(n4451), .A2(n4450), .ZN(n5651) );
  INV_X1 U5473 ( .A(n5651), .ZN(n4452) );
  INV_X1 U5474 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U5475 ( .A1(n4453), .A2(n5985), .ZN(n4459) );
  NAND2_X1 U5476 ( .A1(n4455), .A2(n4454), .ZN(n4457) );
  NAND2_X1 U5477 ( .A1(n4465), .A2(n5985), .ZN(n4456) );
  NAND3_X1 U5478 ( .A1(n4457), .A2(n5685), .A3(n4456), .ZN(n4458) );
  NAND2_X1 U5479 ( .A1(n4459), .A2(n4458), .ZN(n5577) );
  OR2_X1 U5480 ( .A1(n4470), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4467)
         );
  INV_X1 U5481 ( .A(n4467), .ZN(n4460) );
  MUX2_X1 U5482 ( .A(EBX_REG_29__SCAN_IN), .B(n4460), .S(n5685), .Z(n4461) );
  INV_X1 U5483 ( .A(n4461), .ZN(n4464) );
  INV_X1 U5484 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U5485 ( .A1(n4462), .A2(n5644), .ZN(n4463) );
  NAND2_X1 U5486 ( .A1(n4464), .A2(n4463), .ZN(n5615) );
  NOR2_X1 U5487 ( .A1(n4469), .A2(n5615), .ZN(n5617) );
  NAND2_X1 U5488 ( .A1(n4465), .A2(n5644), .ZN(n4466) );
  NAND2_X1 U5489 ( .A1(n4467), .A2(n4466), .ZN(n4468) );
  OAI22_X1 U5490 ( .A1(n4470), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4666), .ZN(n4471) );
  INV_X1 U5491 ( .A(n4471), .ZN(n4472) );
  NOR2_X1 U5492 ( .A1(n4666), .A2(n4475), .ZN(n4474) );
  INV_X1 U5493 ( .A(n4475), .ZN(n4873) );
  OR2_X1 U5494 ( .A1(n6673), .A2(n4873), .ZN(n6641) );
  AND2_X1 U5495 ( .A1(n3512), .A2(n6641), .ZN(n4872) );
  AOI22_X1 U5496 ( .A1(n4476), .A2(n4872), .B1(PHYADDRPOINTER_REG_31__SCAN_IN), 
        .B2(n6230), .ZN(n4477) );
  INV_X1 U5497 ( .A(n4488), .ZN(n4479) );
  NOR3_X1 U5498 ( .A1(n4479), .A2(REIP_REG_30__SCAN_IN), .A3(n7097), .ZN(n5611) );
  NAND2_X1 U5499 ( .A1(n6271), .A2(n5248), .ZN(n6261) );
  NAND3_X1 U5500 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4482) );
  INV_X1 U5501 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6701) );
  INV_X1 U5502 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6697) );
  NOR3_X1 U5503 ( .A1(n6701), .A2(n5557), .A3(n6197), .ZN(n6049) );
  INV_X1 U5504 ( .A(n6261), .ZN(n6050) );
  AOI21_X1 U5505 ( .B1(n6049), .B2(n4481), .A(n6050), .ZN(n6042) );
  AOI21_X1 U5506 ( .B1(n6261), .B2(n4482), .A(n6042), .ZN(n6023) );
  INV_X1 U5507 ( .A(n5633), .ZN(n4483) );
  NAND2_X1 U5508 ( .A1(n4483), .A2(REIP_REG_26__SCAN_IN), .ZN(n4484) );
  NAND2_X1 U5509 ( .A1(n6261), .A2(n4484), .ZN(n4485) );
  NAND2_X1 U5510 ( .A1(n6023), .A2(n4485), .ZN(n6005) );
  AND2_X1 U5511 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4486) );
  NOR2_X1 U5512 ( .A1(n6271), .A2(n4486), .ZN(n4487) );
  NOR2_X1 U5513 ( .A1(n6005), .A2(n4487), .ZN(n5986) );
  NAND2_X1 U5514 ( .A1(n4488), .A2(n7097), .ZN(n5621) );
  NAND2_X1 U5515 ( .A1(n5986), .A2(n5621), .ZN(n5613) );
  OAI21_X1 U5516 ( .B1(n5611), .B2(n5613), .A(REIP_REG_31__SCAN_IN), .ZN(n4489) );
  XNOR2_X1 U5517 ( .A(n5619), .B(n4491), .ZN(n5735) );
  NAND3_X1 U5518 ( .A1(n4493), .A2(n4492), .A3(n5582), .ZN(n4494) );
  OR2_X1 U5519 ( .A1(n4494), .A2(n3382), .ZN(n4670) );
  OAI22_X1 U5520 ( .A1(n4594), .A2(n5597), .B1(n4666), .B2(n4670), .ZN(n4495)
         );
  INV_X2 U5521 ( .A(n6066), .ZN(n5709) );
  NAND2_X1 U5522 ( .A1(n5735), .A2(n6066), .ZN(n4509) );
  INV_X1 U5523 ( .A(n4496), .ZN(n4502) );
  INV_X1 U5524 ( .A(n4469), .ZN(n4497) );
  NAND2_X1 U5525 ( .A1(n4502), .A2(n4497), .ZN(n4499) );
  INV_X1 U5526 ( .A(n4501), .ZN(n4498) );
  NAND2_X1 U5527 ( .A1(n4499), .A2(n4498), .ZN(n4504) );
  NAND2_X1 U5528 ( .A1(n4469), .A2(n3833), .ZN(n4500) );
  NAND3_X1 U5529 ( .A1(n4502), .A2(n4501), .A3(n4500), .ZN(n4503) );
  OAI21_X2 U5530 ( .B1(n4505), .B2(n4504), .A(n4503), .ZN(n5844) );
  INV_X1 U5531 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U5532 ( .A1(n4506), .A2(EBX_REG_30__SCAN_IN), .ZN(n4507) );
  NAND2_X1 U5533 ( .A1(n4509), .A2(n3234), .ZN(U2829) );
  NAND2_X1 U5534 ( .A1(n4669), .A2(n4666), .ZN(n5604) );
  INV_X1 U5535 ( .A(n5604), .ZN(n4512) );
  INV_X1 U5536 ( .A(n6741), .ZN(n4510) );
  OAI21_X1 U5537 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n6543), .A(n4515), .ZN(
        n5980) );
  OAI22_X1 U5538 ( .A1(n4510), .A2(n5604), .B1(n5980), .B2(
        READREQUEST_REG_SCAN_IN), .ZN(n4511) );
  OAI21_X1 U5539 ( .B1(n4512), .B2(n5981), .A(n4511), .ZN(U3474) );
  OR2_X1 U5540 ( .A1(n4515), .A2(n4783), .ZN(n4554) );
  INV_X1 U5541 ( .A(EAX_REG_15__SCAN_IN), .ZN(n4517) );
  INV_X1 U5542 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4516) );
  INV_X1 U5543 ( .A(n4515), .ZN(n4513) );
  INV_X1 U5544 ( .A(n4559), .ZN(n4610) );
  NAND2_X1 U5545 ( .A1(n4783), .A2(n5605), .ZN(n4514) );
  INV_X1 U5546 ( .A(DATAI_15_), .ZN(n7082) );
  OAI222_X1 U5547 ( .A1(n4554), .A2(n4517), .B1(n4516), .B2(n4610), .C1(n4674), 
        .C2(n7082), .ZN(U2954) );
  NAND2_X1 U5548 ( .A1(n4637), .A2(DATAI_3_), .ZN(n4627) );
  NAND2_X1 U5549 ( .A1(n4559), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4518) );
  OAI211_X1 U5550 ( .C1(n4554), .C2(n4519), .A(n4627), .B(n4518), .ZN(U2927)
         );
  NAND2_X1 U5551 ( .A1(n6656), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6719) );
  INV_X1 U5552 ( .A(n4520), .ZN(n4530) );
  NAND2_X1 U5553 ( .A1(n5597), .A2(n5588), .ZN(n4524) );
  INV_X1 U5554 ( .A(n4542), .ZN(n4522) );
  NAND2_X1 U5555 ( .A1(n4522), .A2(n4521), .ZN(n4523) );
  NAND2_X1 U5556 ( .A1(n4524), .A2(n4523), .ZN(n4672) );
  INV_X1 U5557 ( .A(n4672), .ZN(n4529) );
  AOI21_X1 U5558 ( .B1(n4666), .B2(n6673), .A(READY_N), .ZN(n4525) );
  OAI211_X1 U5559 ( .C1(n4540), .C2(n6617), .A(n5597), .B(n4525), .ZN(n4527)
         );
  AND2_X1 U5560 ( .A1(n4527), .A2(n4526), .ZN(n4528) );
  INV_X1 U5561 ( .A(n6652), .ZN(n6650) );
  INV_X1 U5562 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7094) );
  NAND2_X1 U5563 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4725) );
  NOR2_X1 U5564 ( .A1(n6656), .A2(n4725), .ZN(n4720) );
  INV_X1 U5565 ( .A(n4720), .ZN(n6718) );
  OAI22_X1 U5566 ( .A1(n4708), .A2(n6650), .B1(n7094), .B2(n6718), .ZN(n4533)
         );
  INV_X1 U5567 ( .A(n4533), .ZN(n4531) );
  NAND2_X1 U5568 ( .A1(n6719), .A2(n4531), .ZN(n6727) );
  INV_X1 U5569 ( .A(n4990), .ZN(n5372) );
  OR2_X1 U5570 ( .A1(n3538), .A2(n5372), .ZN(n4532) );
  XNOR2_X1 U5571 ( .A(n4532), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6259)
         );
  NOR2_X1 U5572 ( .A1(n4542), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4707) );
  AND2_X1 U5573 ( .A1(n6722), .A2(n4533), .ZN(n4534) );
  NAND3_X1 U5574 ( .A1(n6259), .A2(n4707), .A3(n4534), .ZN(n4535) );
  OAI21_X1 U5575 ( .B1(n6727), .B2(n3949), .A(n4535), .ZN(U3455) );
  INV_X1 U5576 ( .A(n6727), .ZN(n6729) );
  INV_X1 U5577 ( .A(n4538), .ZN(n4539) );
  NOR2_X1 U5578 ( .A1(n4540), .A2(n4539), .ZN(n4541) );
  AND2_X1 U5579 ( .A1(n4542), .A2(n4541), .ZN(n4543) );
  NAND2_X1 U5580 ( .A1(n3172), .A2(n4543), .ZN(n6615) );
  INV_X1 U5581 ( .A(n6615), .ZN(n4592) );
  OR2_X1 U5582 ( .A1(n4537), .A2(n4592), .ZN(n4549) );
  NOR2_X1 U5583 ( .A1(n4544), .A2(n4545), .ZN(n4547) );
  AOI22_X1 U5584 ( .A1(n6617), .A2(n3370), .B1(n4547), .B2(n4546), .ZN(n4548)
         );
  NAND2_X1 U5585 ( .A1(n4549), .A2(n4548), .ZN(n6619) );
  INV_X1 U5586 ( .A(n6732), .ZN(n4606) );
  INV_X1 U5587 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4550) );
  AOI22_X1 U5588 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4550), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4684), .ZN(n4603) );
  NAND2_X1 U5589 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4604) );
  INV_X1 U5590 ( .A(n4604), .ZN(n6726) );
  INV_X1 U5591 ( .A(n4544), .ZN(n4551) );
  INV_X1 U5592 ( .A(n4722), .ZN(n6724) );
  NOR2_X1 U5593 ( .A1(n6724), .A2(n4545), .ZN(n4607) );
  AOI222_X1 U5594 ( .A1(n6619), .A2(n4606), .B1(n4603), .B2(n6726), .C1(n4551), 
        .C2(n4607), .ZN(n4553) );
  NAND2_X1 U5595 ( .A1(n6729), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4552) );
  OAI21_X1 U5596 ( .B1(n6729), .B2(n4553), .A(n4552), .ZN(U3460) );
  INV_X2 U5597 ( .A(n4554), .ZN(n4649) );
  AOI22_X1 U5598 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n4559), .B1(n4649), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n4555) );
  NAND2_X1 U5599 ( .A1(n4637), .A2(DATAI_12_), .ZN(n4621) );
  NAND2_X1 U5600 ( .A1(n4555), .A2(n4621), .ZN(U2936) );
  AOI22_X1 U5601 ( .A1(UWORD_REG_11__SCAN_IN), .A2(n4559), .B1(n4649), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n4556) );
  NAND2_X1 U5602 ( .A1(n4637), .A2(DATAI_11_), .ZN(n4625) );
  NAND2_X1 U5603 ( .A1(n4556), .A2(n4625), .ZN(U2935) );
  AOI22_X1 U5604 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n4559), .B1(n4649), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n4557) );
  NAND2_X1 U5605 ( .A1(n4637), .A2(DATAI_2_), .ZN(n4612) );
  NAND2_X1 U5606 ( .A1(n4557), .A2(n4612), .ZN(U2926) );
  AOI22_X1 U5607 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n4559), .B1(n4649), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n4558) );
  NAND2_X1 U5608 ( .A1(n4637), .A2(DATAI_1_), .ZN(n4614) );
  NAND2_X1 U5609 ( .A1(n4558), .A2(n4614), .ZN(U2925) );
  AOI22_X1 U5610 ( .A1(UWORD_REG_10__SCAN_IN), .A2(n4559), .B1(n4649), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n4560) );
  INV_X1 U5611 ( .A(DATAI_10_), .ZN(n5228) );
  OR2_X1 U5612 ( .A1(n4674), .A2(n5228), .ZN(n4623) );
  NAND2_X1 U5613 ( .A1(n4560), .A2(n4623), .ZN(U2934) );
  INV_X1 U5614 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4566) );
  INV_X1 U5615 ( .A(n6642), .ZN(n4561) );
  INV_X1 U5616 ( .A(n6673), .ZN(n5603) );
  OAI21_X1 U5617 ( .B1(n6617), .B2(n4561), .A(n5603), .ZN(n4562) );
  NAND2_X1 U5618 ( .A1(n4564), .A2(n4874), .ZN(n4745) );
  NOR2_X1 U5619 ( .A1(n4725), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6743) );
  AOI22_X1 U5620 ( .A1(n6743), .A2(UWORD_REG_8__SCAN_IN), .B1(n6346), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4565) );
  OAI21_X1 U5621 ( .B1(n4566), .B2(n4745), .A(n4565), .ZN(U2899) );
  INV_X1 U5622 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5623 ( .A1(n6743), .A2(UWORD_REG_9__SCAN_IN), .B1(n6346), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4567) );
  OAI21_X1 U5624 ( .B1(n4568), .B2(n4745), .A(n4567), .ZN(U2898) );
  INV_X1 U5625 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4570) );
  AOI22_X1 U5626 ( .A1(n6743), .A2(UWORD_REG_11__SCAN_IN), .B1(n6346), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4569) );
  OAI21_X1 U5627 ( .B1(n4570), .B2(n4745), .A(n4569), .ZN(U2896) );
  INV_X1 U5628 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4572) );
  AOI22_X1 U5629 ( .A1(n6743), .A2(UWORD_REG_12__SCAN_IN), .B1(n6346), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4571) );
  OAI21_X1 U5630 ( .B1(n4572), .B2(n4745), .A(n4571), .ZN(U2895) );
  INV_X1 U5631 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4574) );
  AOI22_X1 U5632 ( .A1(n6743), .A2(UWORD_REG_13__SCAN_IN), .B1(n6346), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4573) );
  OAI21_X1 U5633 ( .B1(n4574), .B2(n4745), .A(n4573), .ZN(U2894) );
  INV_X1 U5634 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4576) );
  AOI22_X1 U5635 ( .A1(n6743), .A2(UWORD_REG_10__SCAN_IN), .B1(n6346), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4575) );
  OAI21_X1 U5636 ( .B1(n4576), .B2(n4745), .A(n4575), .ZN(U2897) );
  INV_X1 U5637 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4578) );
  AOI22_X1 U5638 ( .A1(n6743), .A2(UWORD_REG_14__SCAN_IN), .B1(n6346), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4577) );
  OAI21_X1 U5639 ( .B1(n4578), .B2(n4745), .A(n4577), .ZN(U2893) );
  INV_X1 U5640 ( .A(n4579), .ZN(n4580) );
  AOI21_X1 U5641 ( .B1(n4581), .B2(n4589), .A(n4580), .ZN(n4962) );
  INV_X1 U5642 ( .A(n4962), .ZN(n4586) );
  INV_X1 U5643 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4585) );
  OAI21_X1 U5644 ( .B1(n4584), .B2(n4583), .A(n4582), .ZN(n6317) );
  OAI222_X1 U5645 ( .A1(n4586), .A2(n6293), .B1(n4585), .B2(n6297), .C1(n6317), 
        .C2(n5709), .ZN(U2859) );
  XNOR2_X1 U5646 ( .A(n4587), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4658)
         );
  AND2_X1 U5647 ( .A1(n6457), .A2(REIP_REG_0__SCAN_IN), .ZN(n4655) );
  AOI21_X1 U5648 ( .B1(n4682), .B2(n5947), .A(n4589), .ZN(n4588) );
  AOI211_X1 U5649 ( .C1(n6448), .C2(n4962), .A(n4655), .B(n4588), .ZN(n4590)
         );
  NAND2_X1 U5650 ( .A1(n6453), .A2(n5952), .ZN(n5948) );
  NAND2_X1 U5651 ( .A1(n5948), .A2(n4589), .ZN(n4681) );
  OAI211_X1 U5652 ( .C1(n4658), .C2(n6138), .A(n4590), .B(n4681), .ZN(U3018)
         );
  OR2_X1 U5653 ( .A1(n4591), .A2(n4592), .ZN(n4600) );
  NAND2_X1 U5654 ( .A1(n4594), .A2(n4593), .ZN(n4701) );
  XNOR2_X1 U5655 ( .A(n4545), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4598)
         );
  XNOR2_X1 U5656 ( .A(n3370), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4595)
         );
  NAND2_X1 U5657 ( .A1(n6617), .A2(n4595), .ZN(n4596) );
  OAI21_X1 U5658 ( .B1(n4598), .B2(n4698), .A(n4596), .ZN(n4597) );
  AOI21_X1 U5659 ( .B1(n4701), .B2(n4598), .A(n4597), .ZN(n4599) );
  NAND2_X1 U5660 ( .A1(n4600), .A2(n4599), .ZN(n4704) );
  NAND3_X1 U5661 ( .A1(n4722), .A2(n4545), .A3(n4601), .ZN(n4602) );
  OAI21_X1 U5662 ( .B1(n4604), .B2(n4603), .A(n4602), .ZN(n4605) );
  AOI21_X1 U5663 ( .B1(n4704), .B2(n4606), .A(n4605), .ZN(n4609) );
  OAI21_X1 U5664 ( .B1(n6729), .B2(n4607), .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .ZN(n4608) );
  OAI21_X1 U5665 ( .B1(n4609), .B2(n6729), .A(n4608), .ZN(U3459) );
  AOI22_X1 U5666 ( .A1(UWORD_REG_14__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n4611) );
  NAND2_X1 U5667 ( .A1(n4637), .A2(DATAI_14_), .ZN(n4630) );
  NAND2_X1 U5668 ( .A1(n4611), .A2(n4630), .ZN(U2938) );
  AOI22_X1 U5669 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n4613) );
  NAND2_X1 U5670 ( .A1(n4613), .A2(n4612), .ZN(U2941) );
  AOI22_X1 U5671 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n4615) );
  NAND2_X1 U5672 ( .A1(n4615), .A2(n4614), .ZN(U2940) );
  AOI22_X1 U5673 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n4616) );
  NAND2_X1 U5674 ( .A1(n4637), .A2(DATAI_4_), .ZN(n4639) );
  NAND2_X1 U5675 ( .A1(n4616), .A2(n4639), .ZN(U2928) );
  AOI22_X1 U5676 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n4617) );
  NAND2_X1 U5677 ( .A1(n4637), .A2(DATAI_5_), .ZN(n4641) );
  NAND2_X1 U5678 ( .A1(n4617), .A2(n4641), .ZN(U2929) );
  AOI22_X1 U5679 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n4618) );
  NAND2_X1 U5680 ( .A1(n4637), .A2(DATAI_6_), .ZN(n4643) );
  NAND2_X1 U5681 ( .A1(n4618), .A2(n4643), .ZN(U2930) );
  AOI22_X1 U5682 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n4619) );
  NAND2_X1 U5683 ( .A1(n4637), .A2(DATAI_7_), .ZN(n4633) );
  NAND2_X1 U5684 ( .A1(n4619), .A2(n4633), .ZN(U2931) );
  AOI22_X1 U5685 ( .A1(UWORD_REG_8__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n4620) );
  NAND2_X1 U5686 ( .A1(n4637), .A2(DATAI_8_), .ZN(n4635) );
  NAND2_X1 U5687 ( .A1(n4620), .A2(n4635), .ZN(U2932) );
  AOI22_X1 U5688 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n4622) );
  NAND2_X1 U5689 ( .A1(n4622), .A2(n4621), .ZN(U2951) );
  AOI22_X1 U5690 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n4624) );
  NAND2_X1 U5691 ( .A1(n4624), .A2(n4623), .ZN(U2949) );
  AOI22_X1 U5692 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n4626) );
  NAND2_X1 U5693 ( .A1(n4626), .A2(n4625), .ZN(U2950) );
  AOI22_X1 U5694 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n4628) );
  NAND2_X1 U5695 ( .A1(n4628), .A2(n4627), .ZN(U2942) );
  AOI22_X1 U5696 ( .A1(UWORD_REG_13__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n4629) );
  NAND2_X1 U5697 ( .A1(n4637), .A2(DATAI_13_), .ZN(n4645) );
  NAND2_X1 U5698 ( .A1(n4629), .A2(n4645), .ZN(U2937) );
  AOI22_X1 U5699 ( .A1(LWORD_REG_14__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n4631) );
  NAND2_X1 U5700 ( .A1(n4631), .A2(n4630), .ZN(U2953) );
  AOI22_X1 U5701 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_0__SCAN_IN), .ZN(n4632) );
  NAND2_X1 U5702 ( .A1(n4637), .A2(DATAI_0_), .ZN(n4651) );
  NAND2_X1 U5703 ( .A1(n4632), .A2(n4651), .ZN(U2939) );
  AOI22_X1 U5704 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4634) );
  NAND2_X1 U5705 ( .A1(n4634), .A2(n4633), .ZN(U2946) );
  AOI22_X1 U5706 ( .A1(LWORD_REG_8__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4636) );
  NAND2_X1 U5707 ( .A1(n4636), .A2(n4635), .ZN(U2947) );
  AOI22_X1 U5708 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4638) );
  NAND2_X1 U5709 ( .A1(n4637), .A2(DATAI_9_), .ZN(n4647) );
  NAND2_X1 U5710 ( .A1(n4638), .A2(n4647), .ZN(U2948) );
  AOI22_X1 U5711 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n4640) );
  NAND2_X1 U5712 ( .A1(n4640), .A2(n4639), .ZN(U2943) );
  AOI22_X1 U5713 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n4642) );
  NAND2_X1 U5714 ( .A1(n4642), .A2(n4641), .ZN(U2944) );
  AOI22_X1 U5715 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n4644) );
  NAND2_X1 U5716 ( .A1(n4644), .A2(n4643), .ZN(U2945) );
  AOI22_X1 U5717 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n4646) );
  NAND2_X1 U5718 ( .A1(n4646), .A2(n4645), .ZN(U2952) );
  AOI22_X1 U5719 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n4648) );
  NAND2_X1 U5720 ( .A1(n4648), .A2(n4647), .ZN(U2933) );
  AOI22_X1 U5721 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n4650), .B1(n4649), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n4652) );
  NAND2_X1 U5722 ( .A1(n4652), .A2(n4651), .ZN(U2924) );
  NAND2_X1 U5723 ( .A1(n4653), .A2(n6111), .ZN(n4656) );
  NOR2_X1 U5724 ( .A1(n6317), .A2(n6108), .ZN(n4654) );
  AOI211_X1 U5725 ( .C1(PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n4656), .A(n4655), 
        .B(n4654), .ZN(n4657) );
  OAI21_X1 U5726 ( .B1(n4658), .B2(n6164), .A(n4657), .ZN(U2986) );
  INV_X1 U5727 ( .A(n4659), .ZN(n4660) );
  OAI21_X1 U5728 ( .B1(n4662), .B2(n4661), .A(n4660), .ZN(n5174) );
  INV_X1 U5729 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4668) );
  INV_X1 U5730 ( .A(n4663), .ZN(n4667) );
  INV_X1 U5731 ( .A(n4664), .ZN(n4665) );
  AOI21_X1 U5732 ( .B1(n4667), .B2(n4666), .A(n4665), .ZN(n4689) );
  OAI222_X1 U5733 ( .A1(n5709), .A2(n5174), .B1(n6297), .B2(n4668), .C1(n6293), 
        .C2(n4689), .ZN(U2858) );
  NOR2_X1 U5734 ( .A1(n4670), .A2(n4669), .ZN(n4671) );
  NAND2_X2 U5735 ( .A1(n6314), .A2(n4675), .ZN(n6316) );
  INV_X1 U5736 ( .A(n4676), .ZN(n4677) );
  NOR2_X2 U5737 ( .A1(n6310), .A2(n6307), .ZN(n6315) );
  INV_X1 U5738 ( .A(DATAI_1_), .ZN(n7029) );
  INV_X1 U5739 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6345) );
  OAI222_X1 U5740 ( .A1(n5174), .A2(n6316), .B1(n6315), .B2(n7029), .C1(n6314), 
        .C2(n6345), .ZN(U2890) );
  XOR2_X1 U5741 ( .A(n4680), .B(n4679), .Z(n4747) );
  NAND2_X1 U5742 ( .A1(n4747), .A2(n6454), .ZN(n4688) );
  INV_X1 U5743 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6733) );
  NOR2_X1 U5744 ( .A1(n6403), .A2(n6733), .ZN(n4749) );
  AOI21_X1 U5745 ( .B1(n4682), .B2(n4681), .A(n4684), .ZN(n4686) );
  AND3_X1 U5746 ( .A1(n4684), .A2(n4683), .A3(n5847), .ZN(n4685) );
  NOR3_X1 U5747 ( .A1(n4749), .A2(n4686), .A3(n4685), .ZN(n4687) );
  OAI211_X1 U5748 ( .C1(n4689), .C2(n6405), .A(n4688), .B(n4687), .ZN(U3017)
         );
  NAND2_X1 U5749 ( .A1(n4690), .A2(n6615), .ZN(n4703) );
  MUX2_X1 U5750 ( .A(n4691), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4545), 
        .Z(n4693) );
  NOR2_X1 U5751 ( .A1(n4693), .A2(n4692), .ZN(n4700) );
  OAI21_X1 U5752 ( .B1(n4694), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n3447), 
        .ZN(n5977) );
  XNOR2_X1 U5753 ( .A(n4695), .B(n3939), .ZN(n4696) );
  NAND2_X1 U5754 ( .A1(n6617), .A2(n4696), .ZN(n4697) );
  OAI21_X1 U5755 ( .B1(n5977), .B2(n4698), .A(n4697), .ZN(n4699) );
  AOI21_X1 U5756 ( .B1(n4701), .B2(n4700), .A(n4699), .ZN(n4702) );
  NAND2_X1 U5757 ( .A1(n4703), .A2(n4702), .ZN(n5976) );
  INV_X1 U5758 ( .A(n4708), .ZN(n6620) );
  MUX2_X1 U5759 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5976), .S(n6620), 
        .Z(n6631) );
  NAND2_X1 U5760 ( .A1(n4704), .A2(n6620), .ZN(n4706) );
  NAND2_X1 U5761 ( .A1(n4708), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4705) );
  NAND2_X1 U5762 ( .A1(n4706), .A2(n4705), .ZN(n6626) );
  NAND3_X1 U5763 ( .A1(n6631), .A2(n4712), .A3(n6626), .ZN(n4716) );
  NAND2_X1 U5764 ( .A1(n6259), .A2(n4707), .ZN(n4711) );
  MUX2_X1 U5765 ( .A(n4708), .B(n7094), .S(STATE2_REG_1__SCAN_IN), .Z(n4709)
         );
  NAND2_X1 U5766 ( .A1(n4709), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U5767 ( .A1(n4711), .A2(n4710), .ZN(n4717) );
  NOR2_X1 U5768 ( .A1(FLUSH_REG_SCAN_IN), .A2(n4712), .ZN(n4713) );
  AND2_X1 U5769 ( .A1(n4692), .A2(n4713), .ZN(n4714) );
  NOR2_X1 U5770 ( .A1(n4717), .A2(n4714), .ZN(n4715) );
  NAND2_X1 U5771 ( .A1(n4716), .A2(n4715), .ZN(n6612) );
  INV_X1 U5772 ( .A(n4717), .ZN(n4718) );
  NAND2_X1 U5773 ( .A1(n4718), .A2(n4544), .ZN(n4719) );
  NAND2_X1 U5774 ( .A1(n6612), .A2(n4719), .ZN(n4724) );
  NAND2_X1 U5775 ( .A1(n4724), .A2(n7094), .ZN(n4721) );
  NAND2_X1 U5776 ( .A1(n4721), .A2(n4720), .ZN(n4723) );
  INV_X1 U5777 ( .A(n6463), .ZN(n4730) );
  INV_X1 U5778 ( .A(n4724), .ZN(n4726) );
  NOR2_X1 U5779 ( .A1(n4726), .A2(n4725), .ZN(n6646) );
  INV_X1 U5780 ( .A(n6616), .ZN(n5405) );
  AND2_X1 U5781 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6722), .ZN(n5974) );
  OAI22_X1 U5782 ( .A1(n4727), .A2(n6543), .B1(n5405), .B2(n5974), .ZN(n4728)
         );
  OAI21_X1 U5783 ( .B1(n6646), .B2(n4728), .A(n4730), .ZN(n4729) );
  OAI21_X1 U5784 ( .B1(n4730), .B2(n5407), .A(n4729), .ZN(U3465) );
  INV_X1 U5785 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4732) );
  AOI22_X1 U5786 ( .A1(n6638), .A2(UWORD_REG_0__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4731) );
  OAI21_X1 U5787 ( .B1(n4732), .B2(n4745), .A(n4731), .ZN(U2907) );
  INV_X1 U5788 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4734) );
  AOI22_X1 U5789 ( .A1(n6638), .A2(UWORD_REG_5__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4733) );
  OAI21_X1 U5790 ( .B1(n4734), .B2(n4745), .A(n4733), .ZN(U2902) );
  INV_X1 U5791 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4736) );
  AOI22_X1 U5792 ( .A1(n6638), .A2(UWORD_REG_2__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4735) );
  OAI21_X1 U5793 ( .B1(n4736), .B2(n4745), .A(n4735), .ZN(U2905) );
  AOI22_X1 U5794 ( .A1(n6638), .A2(UWORD_REG_3__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4737) );
  OAI21_X1 U5795 ( .B1(n4519), .B2(n4745), .A(n4737), .ZN(U2904) );
  INV_X1 U5796 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4739) );
  AOI22_X1 U5797 ( .A1(n6638), .A2(UWORD_REG_4__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4738) );
  OAI21_X1 U5798 ( .B1(n4739), .B2(n4745), .A(n4738), .ZN(U2903) );
  INV_X1 U5799 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4741) );
  AOI22_X1 U5800 ( .A1(n6638), .A2(UWORD_REG_1__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4740) );
  OAI21_X1 U5801 ( .B1(n4741), .B2(n4745), .A(n4740), .ZN(U2906) );
  INV_X1 U5802 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4743) );
  AOI22_X1 U5803 ( .A1(n6743), .A2(UWORD_REG_7__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4742) );
  OAI21_X1 U5804 ( .B1(n4743), .B2(n4745), .A(n4742), .ZN(U2900) );
  INV_X1 U5805 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4746) );
  AOI22_X1 U5806 ( .A1(n6743), .A2(UWORD_REG_6__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4744) );
  OAI21_X1 U5807 ( .B1(n4746), .B2(n4745), .A(n4744), .ZN(U2901) );
  NAND2_X1 U5808 ( .A1(n4747), .A2(n6380), .ZN(n4751) );
  NOR2_X1 U5809 ( .A1(n6384), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4748)
         );
  AOI211_X1 U5810 ( .C1(n6374), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4749), 
        .B(n4748), .ZN(n4750) );
  OAI211_X1 U5811 ( .C1(n6108), .C2(n5174), .A(n4751), .B(n4750), .ZN(U2985)
         );
  NOR2_X1 U5812 ( .A1(n4754), .A2(n4753), .ZN(n4755) );
  NOR2_X1 U5813 ( .A1(n4752), .A2(n4755), .ZN(n6379) );
  INV_X1 U5814 ( .A(n6379), .ZN(n5239) );
  INV_X1 U5815 ( .A(DATAI_2_), .ZN(n7036) );
  INV_X1 U5816 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6343) );
  OAI222_X1 U5817 ( .A1(n5239), .A2(n6316), .B1(n6315), .B2(n7036), .C1(n6314), 
        .C2(n6343), .ZN(U2889) );
  NAND2_X1 U5818 ( .A1(n4752), .A2(n4766), .ZN(n4760) );
  INV_X1 U5819 ( .A(n4758), .ZN(n4759) );
  NAND2_X1 U5820 ( .A1(n4760), .A2(n4759), .ZN(n4761) );
  NAND2_X1 U5821 ( .A1(n4757), .A2(n4761), .ZN(n6266) );
  INV_X1 U5822 ( .A(n6430), .ZN(n4762) );
  OAI222_X1 U5823 ( .A1(n6266), .A2(n5709), .B1(n4763), .B2(n6297), .C1(n6293), 
        .C2(n4762), .ZN(U2855) );
  INV_X1 U5824 ( .A(DATAI_4_), .ZN(n7095) );
  INV_X1 U5825 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6339) );
  OAI222_X1 U5826 ( .A1(n6266), .A2(n6316), .B1(n6315), .B2(n7095), .C1(n6314), 
        .C2(n6339), .ZN(U2887) );
  INV_X1 U5827 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4765) );
  XNOR2_X1 U5828 ( .A(n4764), .B(n4768), .ZN(n6446) );
  OAI222_X1 U5829 ( .A1(n5709), .A2(n5239), .B1(n4765), .B2(n6297), .C1(n6293), 
        .C2(n6446), .ZN(U2857) );
  XOR2_X1 U5830 ( .A(n4752), .B(n4766), .Z(n6370) );
  INV_X1 U5831 ( .A(n6370), .ZN(n4772) );
  INV_X1 U5832 ( .A(DATAI_3_), .ZN(n6862) );
  INV_X1 U5833 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6341) );
  OAI222_X1 U5834 ( .A1(n4772), .A2(n6316), .B1(n6315), .B2(n6862), .C1(n6314), 
        .C2(n6341), .ZN(U2888) );
  XNOR2_X1 U5835 ( .A(n4767), .B(n4757), .ZN(n6362) );
  INV_X1 U5836 ( .A(n6362), .ZN(n4796) );
  INV_X1 U5837 ( .A(DATAI_5_), .ZN(n7085) );
  OAI222_X1 U5838 ( .A1(n6316), .A2(n4796), .B1(n6314), .B2(n3908), .C1(n7085), 
        .C2(n6315), .ZN(U2886) );
  NAND2_X1 U5839 ( .A1(n4764), .A2(n4768), .ZN(n4770) );
  NAND2_X1 U5840 ( .A1(n4770), .A2(n4769), .ZN(n4771) );
  INV_X1 U5841 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4773) );
  OAI222_X1 U5842 ( .A1(n6438), .A2(n6293), .B1(n4773), .B2(n6297), .C1(n4772), 
        .C2(n5709), .ZN(U2856) );
  OR2_X1 U5843 ( .A1(n4591), .A2(n4537), .ZN(n5455) );
  NOR2_X1 U5844 ( .A1(n5455), .A2(n4990), .ZN(n6470) );
  INV_X1 U5845 ( .A(n6525), .ZN(n4774) );
  AOI21_X1 U5846 ( .B1(n6470), .B2(n6616), .A(n4774), .ZN(n4777) );
  OR2_X1 U5847 ( .A1(n6543), .A2(n4777), .ZN(n4775) );
  OAI21_X1 U5848 ( .B1(n6468), .B2(n6655), .A(n4775), .ZN(n6528) );
  INV_X1 U5849 ( .A(n6528), .ZN(n4894) );
  INV_X1 U5850 ( .A(n6543), .ZN(n6537) );
  NAND2_X1 U5851 ( .A1(n5964), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6538) );
  NOR2_X1 U5852 ( .A1(n5365), .A2(n6538), .ZN(n5969) );
  INV_X1 U5853 ( .A(n5969), .ZN(n4778) );
  NAND3_X1 U5854 ( .A1(n4778), .A2(n6537), .A3(n4777), .ZN(n4779) );
  OAI21_X1 U5855 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6722), .A(n5264), 
        .ZN(n6542) );
  OAI211_X1 U5856 ( .C1(n6537), .C2(n4780), .A(n4779), .B(n5180), .ZN(n6529)
         );
  NAND2_X1 U5857 ( .A1(n6529), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4786) );
  INV_X1 U5858 ( .A(n5365), .ZN(n4781) );
  INV_X1 U5859 ( .A(n6532), .ZN(n4788) );
  NAND2_X1 U5860 ( .A1(n6378), .A2(DATAI_25_), .ZN(n6559) );
  INV_X1 U5861 ( .A(n6559), .ZN(n6482) );
  NAND2_X1 U5862 ( .A1(n6378), .A2(DATAI_17_), .ZN(n6554) );
  NAND2_X1 U5863 ( .A1(n4833), .A2(n4783), .ZN(n6553) );
  OAI22_X1 U5864 ( .A1(n6526), .A2(n6554), .B1(n6525), .B2(n6553), .ZN(n4784)
         );
  AOI21_X1 U5865 ( .B1(n4788), .B2(n6482), .A(n4784), .ZN(n4785) );
  OAI211_X1 U5866 ( .C1(n4894), .C2(n5432), .A(n4786), .B(n4785), .ZN(U3077)
         );
  NAND2_X1 U5867 ( .A1(n6529), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4790) );
  NAND2_X1 U5868 ( .A1(n6378), .A2(DATAI_28_), .ZN(n6580) );
  INV_X1 U5869 ( .A(n6580), .ZN(n6494) );
  NAND2_X1 U5870 ( .A1(n6378), .A2(DATAI_20_), .ZN(n6575) );
  NAND2_X1 U5871 ( .A1(n4833), .A2(n3385), .ZN(n6574) );
  OAI22_X1 U5872 ( .A1(n6526), .A2(n6575), .B1(n6525), .B2(n6574), .ZN(n4787)
         );
  AOI21_X1 U5873 ( .B1(n4788), .B2(n6494), .A(n4787), .ZN(n4789) );
  OAI211_X1 U5874 ( .C1(n4894), .C2(n5428), .A(n4790), .B(n4789), .ZN(U3080)
         );
  AOI21_X1 U5875 ( .B1(n4793), .B2(n4792), .A(n4791), .ZN(n4794) );
  OR2_X1 U5876 ( .A1(n4794), .A2(n4843), .ZN(n6248) );
  INV_X1 U5877 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4795) );
  OAI222_X1 U5878 ( .A1(n6248), .A2(n6293), .B1(n5709), .B2(n4796), .C1(n4795), 
        .C2(n6297), .ZN(U2854) );
  AND2_X1 U5879 ( .A1(n4690), .A2(n6616), .ZN(n5179) );
  NAND2_X1 U5880 ( .A1(n4591), .A2(n4537), .ZN(n5130) );
  INV_X1 U5881 ( .A(n5130), .ZN(n4797) );
  NAND3_X1 U5882 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6625), .A3(n5370), .ZN(n5132) );
  NOR2_X1 U5883 ( .A1(n5407), .A2(n5132), .ZN(n4806) );
  AOI21_X1 U5884 ( .B1(n5179), .B2(n4797), .A(n4806), .ZN(n4803) );
  OR3_X1 U5885 ( .A1(n6539), .A2(n5964), .A3(n6163), .ZN(n4799) );
  AOI22_X1 U5886 ( .A1(n4803), .A2(n4801), .B1(n6543), .B2(n5132), .ZN(n4800)
         );
  NAND2_X1 U5887 ( .A1(n5180), .A2(n4800), .ZN(n4831) );
  INV_X1 U5888 ( .A(DATAI_6_), .ZN(n4869) );
  INV_X1 U5889 ( .A(n4801), .ZN(n4802) );
  OAI22_X1 U5890 ( .A1(n4803), .A2(n4802), .B1(n6655), .B2(n5132), .ZN(n4830)
         );
  AOI22_X1 U5891 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4831), .B1(n6591), 
        .B2(n4830), .ZN(n4809) );
  NAND2_X1 U5892 ( .A1(n6378), .A2(DATAI_30_), .ZN(n6594) );
  INV_X1 U5893 ( .A(n6594), .ZN(n6502) );
  NAND2_X1 U5894 ( .A1(n6378), .A2(DATAI_22_), .ZN(n6589) );
  NAND2_X1 U5895 ( .A1(n4833), .A2(n4805), .ZN(n6588) );
  INV_X1 U5896 ( .A(n4806), .ZN(n4834) );
  OAI22_X1 U5897 ( .A1(n5039), .A2(n6589), .B1(n6588), .B2(n4834), .ZN(n4807)
         );
  AOI21_X1 U5898 ( .B1(n6502), .B2(n5129), .A(n4807), .ZN(n4808) );
  NAND2_X1 U5899 ( .A1(n4809), .A2(n4808), .ZN(U3098) );
  INV_X1 U5900 ( .A(DATAI_0_), .ZN(n6847) );
  AOI22_X1 U5901 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4831), .B1(n6549), 
        .B2(n4830), .ZN(n4812) );
  NAND2_X1 U5902 ( .A1(n6378), .A2(DATAI_24_), .ZN(n6552) );
  INV_X1 U5903 ( .A(n6552), .ZN(n6478) );
  NAND2_X1 U5904 ( .A1(n6378), .A2(DATAI_16_), .ZN(n6535) );
  NAND2_X1 U5905 ( .A1(n4833), .A2(n4874), .ZN(n6534) );
  OAI22_X1 U5906 ( .A1(n5039), .A2(n6535), .B1(n6534), .B2(n4834), .ZN(n4810)
         );
  AOI21_X1 U5907 ( .B1(n6478), .B2(n5129), .A(n4810), .ZN(n4811) );
  NAND2_X1 U5908 ( .A1(n4812), .A2(n4811), .ZN(U3092) );
  AOI22_X1 U5909 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4831), .B1(n6577), 
        .B2(n4830), .ZN(n4815) );
  OAI22_X1 U5910 ( .A1(n5039), .A2(n6575), .B1(n6574), .B2(n4834), .ZN(n4813)
         );
  AOI21_X1 U5911 ( .B1(n6494), .B2(n5129), .A(n4813), .ZN(n4814) );
  NAND2_X1 U5912 ( .A1(n4815), .A2(n4814), .ZN(U3096) );
  AOI22_X1 U5913 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4831), .B1(n6584), 
        .B2(n4830), .ZN(n4818) );
  NAND2_X1 U5914 ( .A1(n6378), .A2(DATAI_29_), .ZN(n6582) );
  INV_X1 U5915 ( .A(n6582), .ZN(n6498) );
  NAND2_X1 U5916 ( .A1(n6378), .A2(DATAI_21_), .ZN(n6587) );
  NAND2_X1 U5917 ( .A1(n4833), .A2(n3398), .ZN(n6581) );
  OAI22_X1 U5918 ( .A1(n5039), .A2(n6587), .B1(n6581), .B2(n4834), .ZN(n4816)
         );
  AOI21_X1 U5919 ( .B1(n6498), .B2(n5129), .A(n4816), .ZN(n4817) );
  NAND2_X1 U5920 ( .A1(n4818), .A2(n4817), .ZN(U3097) );
  AOI22_X1 U5921 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4831), .B1(n6570), 
        .B2(n4830), .ZN(n4822) );
  NAND2_X1 U5922 ( .A1(n6378), .A2(DATAI_27_), .ZN(n6573) );
  INV_X1 U5923 ( .A(n6573), .ZN(n6490) );
  NAND2_X1 U5924 ( .A1(n6378), .A2(DATAI_19_), .ZN(n6568) );
  NAND2_X1 U5925 ( .A1(n4833), .A2(n4819), .ZN(n6567) );
  OAI22_X1 U5926 ( .A1(n5039), .A2(n6568), .B1(n6567), .B2(n4834), .ZN(n4820)
         );
  AOI21_X1 U5927 ( .B1(n6490), .B2(n5129), .A(n4820), .ZN(n4821) );
  NAND2_X1 U5928 ( .A1(n4822), .A2(n4821), .ZN(U3095) );
  AOI22_X1 U5929 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4831), .B1(n6556), 
        .B2(n4830), .ZN(n4825) );
  OAI22_X1 U5930 ( .A1(n5039), .A2(n6554), .B1(n6553), .B2(n4834), .ZN(n4823)
         );
  AOI21_X1 U5931 ( .B1(n6482), .B2(n5129), .A(n4823), .ZN(n4824) );
  NAND2_X1 U5932 ( .A1(n4825), .A2(n4824), .ZN(U3093) );
  INV_X1 U5933 ( .A(DATAI_7_), .ZN(n7042) );
  AOI22_X1 U5934 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4831), .B1(n6601), 
        .B2(n4830), .ZN(n4829) );
  INV_X1 U5935 ( .A(DATAI_31_), .ZN(n4826) );
  NOR2_X1 U5936 ( .A1(n6108), .A2(n4826), .ZN(n6509) );
  NAND2_X1 U5937 ( .A1(n6378), .A2(DATAI_23_), .ZN(n6606) );
  NAND2_X1 U5938 ( .A1(n4833), .A2(n3383), .ZN(n6596) );
  OAI22_X1 U5939 ( .A1(n5039), .A2(n6606), .B1(n6596), .B2(n4834), .ZN(n4827)
         );
  AOI21_X1 U5940 ( .B1(n6509), .B2(n5129), .A(n4827), .ZN(n4828) );
  NAND2_X1 U5941 ( .A1(n4829), .A2(n4828), .ZN(U3099) );
  AOI22_X1 U5942 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4831), .B1(n6563), 
        .B2(n4830), .ZN(n4837) );
  NAND2_X1 U5943 ( .A1(n6378), .A2(DATAI_26_), .ZN(n6566) );
  INV_X1 U5944 ( .A(n6566), .ZN(n6486) );
  NAND2_X1 U5945 ( .A1(n6378), .A2(DATAI_18_), .ZN(n6561) );
  NAND2_X1 U5946 ( .A1(n4833), .A2(n4832), .ZN(n6560) );
  OAI22_X1 U5947 ( .A1(n5039), .A2(n6561), .B1(n6560), .B2(n4834), .ZN(n4835)
         );
  AOI21_X1 U5948 ( .B1(n6486), .B2(n5129), .A(n4835), .ZN(n4836) );
  NAND2_X1 U5949 ( .A1(n4837), .A2(n4836), .ZN(U3094) );
  AOI21_X1 U5950 ( .B1(n3957), .B2(n4767), .A(n4838), .ZN(n4840) );
  INV_X1 U5951 ( .A(n4839), .ZN(n4957) );
  NOR2_X1 U5952 ( .A1(n4840), .A2(n4957), .ZN(n4943) );
  INV_X1 U5953 ( .A(n4943), .ZN(n4884) );
  OAI21_X1 U5954 ( .B1(n4843), .B2(n4842), .A(n4841), .ZN(n4844) );
  INV_X1 U5955 ( .A(n4844), .ZN(n4953) );
  AOI22_X1 U5956 ( .A1(n6065), .A2(n4953), .B1(EBX_REG_6__SCAN_IN), .B2(n4506), 
        .ZN(n4845) );
  OAI21_X1 U5957 ( .B1(n4884), .B2(n5709), .A(n4845), .ZN(U2853) );
  NOR2_X1 U5958 ( .A1(n4690), .A2(n5130), .ZN(n5267) );
  NAND3_X1 U5959 ( .A1(n6630), .A2(n6625), .A3(n5370), .ZN(n5262) );
  NOR2_X1 U5960 ( .A1(n5407), .A2(n5262), .ZN(n4866) );
  AOI21_X1 U5961 ( .B1(n5267), .B2(n6616), .A(n4866), .ZN(n4848) );
  AOI21_X1 U5962 ( .B1(n3236), .B2(STATEBS16_REG_SCAN_IN), .A(n6543), .ZN(
        n4847) );
  AOI22_X1 U5963 ( .A1(n4848), .A2(n4847), .B1(n6543), .B2(n5262), .ZN(n4846)
         );
  NAND2_X1 U5964 ( .A1(n5180), .A2(n4846), .ZN(n4865) );
  INV_X1 U5965 ( .A(n4847), .ZN(n4849) );
  OAI22_X1 U5966 ( .A1(n4849), .A2(n4848), .B1(n6655), .B2(n5262), .ZN(n4864)
         );
  AOI22_X1 U5967 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4865), .B1(n6563), 
        .B2(n4864), .ZN(n4851) );
  INV_X1 U5968 ( .A(n6561), .ZN(n5470) );
  INV_X1 U5969 ( .A(n6560), .ZN(n6485) );
  AOI22_X1 U5970 ( .A1(n5317), .A2(n5470), .B1(n6485), .B2(n4866), .ZN(n4850)
         );
  OAI211_X1 U5971 ( .C1(n6566), .C2(n5296), .A(n4851), .B(n4850), .ZN(U3030)
         );
  AOI22_X1 U5972 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4865), .B1(n6570), 
        .B2(n4864), .ZN(n4853) );
  INV_X1 U5973 ( .A(n6568), .ZN(n5486) );
  INV_X1 U5974 ( .A(n6567), .ZN(n6489) );
  AOI22_X1 U5975 ( .A1(n5317), .A2(n5486), .B1(n6489), .B2(n4866), .ZN(n4852)
         );
  OAI211_X1 U5976 ( .C1(n6573), .C2(n5296), .A(n4853), .B(n4852), .ZN(U3031)
         );
  AOI22_X1 U5977 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4865), .B1(n6591), 
        .B2(n4864), .ZN(n4855) );
  INV_X1 U5978 ( .A(n6589), .ZN(n5478) );
  INV_X1 U5979 ( .A(n6588), .ZN(n6501) );
  AOI22_X1 U5980 ( .A1(n5317), .A2(n5478), .B1(n6501), .B2(n4866), .ZN(n4854)
         );
  OAI211_X1 U5981 ( .C1(n6594), .C2(n5296), .A(n4855), .B(n4854), .ZN(U3034)
         );
  AOI22_X1 U5982 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4865), .B1(n6577), 
        .B2(n4864), .ZN(n4857) );
  INV_X1 U5983 ( .A(n6575), .ZN(n5466) );
  INV_X1 U5984 ( .A(n6574), .ZN(n6493) );
  AOI22_X1 U5985 ( .A1(n5317), .A2(n5466), .B1(n6493), .B2(n4866), .ZN(n4856)
         );
  OAI211_X1 U5986 ( .C1(n6580), .C2(n5296), .A(n4857), .B(n4856), .ZN(U3032)
         );
  AOI22_X1 U5987 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4865), .B1(n6549), 
        .B2(n4864), .ZN(n4859) );
  INV_X1 U5988 ( .A(n6535), .ZN(n5492) );
  INV_X1 U5989 ( .A(n6534), .ZN(n6469) );
  AOI22_X1 U5990 ( .A1(n5317), .A2(n5492), .B1(n6469), .B2(n4866), .ZN(n4858)
         );
  OAI211_X1 U5991 ( .C1(n6552), .C2(n5296), .A(n4859), .B(n4858), .ZN(U3028)
         );
  AOI22_X1 U5992 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4865), .B1(n6556), 
        .B2(n4864), .ZN(n4861) );
  INV_X1 U5993 ( .A(n6554), .ZN(n5474) );
  INV_X1 U5994 ( .A(n6553), .ZN(n6481) );
  AOI22_X1 U5995 ( .A1(n5317), .A2(n5474), .B1(n6481), .B2(n4866), .ZN(n4860)
         );
  OAI211_X1 U5996 ( .C1(n6559), .C2(n5296), .A(n4861), .B(n4860), .ZN(U3029)
         );
  AOI22_X1 U5997 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4865), .B1(n6584), 
        .B2(n4864), .ZN(n4863) );
  INV_X1 U5998 ( .A(n6587), .ZN(n5462) );
  INV_X1 U5999 ( .A(n6581), .ZN(n6497) );
  AOI22_X1 U6000 ( .A1(n5317), .A2(n5462), .B1(n6497), .B2(n4866), .ZN(n4862)
         );
  OAI211_X1 U6001 ( .C1(n6582), .C2(n5296), .A(n4863), .B(n4862), .ZN(U3033)
         );
  INV_X1 U6002 ( .A(n6509), .ZN(n6597) );
  AOI22_X1 U6003 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4865), .B1(n6601), 
        .B2(n4864), .ZN(n4868) );
  INV_X1 U6004 ( .A(n6606), .ZN(n5482) );
  INV_X1 U6005 ( .A(n6596), .ZN(n6506) );
  AOI22_X1 U6006 ( .A1(n5317), .A2(n5482), .B1(n6506), .B2(n4866), .ZN(n4867)
         );
  OAI211_X1 U6007 ( .C1(n6597), .C2(n5296), .A(n4868), .B(n4867), .ZN(U3035)
         );
  OAI222_X1 U6008 ( .A1(n4884), .A2(n6316), .B1(n6315), .B2(n4869), .C1(n6314), 
        .C2(n3914), .ZN(U2885) );
  INV_X1 U6009 ( .A(n4872), .ZN(n4876) );
  INV_X1 U6010 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5643) );
  NAND3_X1 U6011 ( .A1(n4874), .A2(n5643), .A3(n4873), .ZN(n4875) );
  NAND2_X1 U6012 ( .A1(n4876), .A2(n4875), .ZN(n4877) );
  OAI21_X1 U6013 ( .B1(n6271), .B2(n4881), .A(n5248), .ZN(n6255) );
  AOI22_X1 U6014 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6230), .B1(
        REIP_REG_6__SCAN_IN), .B2(n6255), .ZN(n4878) );
  OAI211_X1 U6015 ( .C1(n6054), .C2(n4879), .A(n4878), .B(n6249), .ZN(n4880)
         );
  AOI21_X1 U6016 ( .B1(n4942), .B2(n6267), .A(n4880), .ZN(n4883) );
  NOR2_X1 U6017 ( .A1(n6271), .A2(REIP_REG_6__SCAN_IN), .ZN(n6245) );
  AOI22_X1 U6018 ( .A1(n6245), .A2(n4881), .B1(n6260), .B2(n4953), .ZN(n4882)
         );
  OAI211_X1 U6019 ( .C1(n6192), .C2(n4884), .A(n4883), .B(n4882), .ZN(U2821)
         );
  OAI21_X1 U6020 ( .B1(n4887), .B2(n4886), .A(n4885), .ZN(n6431) );
  NAND2_X1 U6021 ( .A1(n6457), .A2(REIP_REG_4__SCAN_IN), .ZN(n6428) );
  OAI21_X1 U6022 ( .B1(n6111), .B2(n6263), .A(n6428), .ZN(n4889) );
  NOR2_X1 U6023 ( .A1(n6266), .A2(n6108), .ZN(n4888) );
  AOI211_X1 U6024 ( .C1(n5808), .C2(n6268), .A(n4889), .B(n4888), .ZN(n4890)
         );
  OAI21_X1 U6025 ( .B1(n6164), .B2(n6431), .A(n4890), .ZN(U2982) );
  OAI22_X1 U6026 ( .A1(n6526), .A2(n6606), .B1(n6525), .B2(n6596), .ZN(n4892)
         );
  NOR2_X1 U6027 ( .A1(n6532), .A2(n6597), .ZN(n4891) );
  AOI211_X1 U6028 ( .C1(n6529), .C2(INSTQUEUE_REG_7__7__SCAN_IN), .A(n4892), 
        .B(n4891), .ZN(n4893) );
  OAI21_X1 U6029 ( .B1(n4894), .B2(n5420), .A(n4893), .ZN(U3083) );
  INV_X1 U6030 ( .A(n4895), .ZN(n4896) );
  OR2_X1 U6031 ( .A1(n4776), .A2(n4896), .ZN(n5176) );
  INV_X1 U6032 ( .A(n4537), .ZN(n5034) );
  NOR2_X1 U6033 ( .A1(n4591), .A2(n5034), .ZN(n5373) );
  NAND3_X1 U6034 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n5370), .ZN(n4991) );
  NOR2_X1 U6035 ( .A1(n5407), .A2(n4991), .ZN(n4897) );
  AOI21_X1 U6036 ( .B1(n5179), .B2(n5373), .A(n4897), .ZN(n4898) );
  OAI22_X1 U6037 ( .A1(n4898), .A2(n6543), .B1(n4991), .B2(n6655), .ZN(n4935)
         );
  INV_X1 U6038 ( .A(n4897), .ZN(n4933) );
  NAND2_X1 U6039 ( .A1(n4904), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5092) );
  NAND2_X1 U6040 ( .A1(n4898), .A2(n5092), .ZN(n4899) );
  OR2_X1 U6041 ( .A1(n6543), .A2(n4899), .ZN(n4901) );
  NAND2_X1 U6042 ( .A1(n6543), .A2(n4991), .ZN(n4900) );
  INV_X1 U6043 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4902) );
  OAI22_X1 U6044 ( .A1(n6567), .A2(n4933), .B1(n4932), .B2(n4902), .ZN(n4903)
         );
  AOI21_X1 U6045 ( .B1(n6570), .B2(n4935), .A(n4903), .ZN(n4906) );
  NAND2_X1 U6046 ( .A1(n5494), .A2(n5486), .ZN(n4905) );
  OAI211_X1 U6047 ( .C1(n5027), .C2(n6573), .A(n4906), .B(n4905), .ZN(U3127)
         );
  INV_X1 U6048 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4907) );
  OAI22_X1 U6049 ( .A1(n6560), .A2(n4933), .B1(n4932), .B2(n4907), .ZN(n4908)
         );
  AOI21_X1 U6050 ( .B1(n6563), .B2(n4935), .A(n4908), .ZN(n4910) );
  NAND2_X1 U6051 ( .A1(n5494), .A2(n5470), .ZN(n4909) );
  OAI211_X1 U6052 ( .C1(n5027), .C2(n6566), .A(n4910), .B(n4909), .ZN(U3126)
         );
  INV_X1 U6053 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4911) );
  OAI22_X1 U6054 ( .A1(n6588), .A2(n4933), .B1(n4932), .B2(n4911), .ZN(n4912)
         );
  AOI21_X1 U6055 ( .B1(n6591), .B2(n4935), .A(n4912), .ZN(n4914) );
  NAND2_X1 U6056 ( .A1(n5494), .A2(n5478), .ZN(n4913) );
  OAI211_X1 U6057 ( .C1(n5027), .C2(n6594), .A(n4914), .B(n4913), .ZN(U3130)
         );
  INV_X1 U6058 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4915) );
  OAI22_X1 U6059 ( .A1(n6596), .A2(n4933), .B1(n4932), .B2(n4915), .ZN(n4916)
         );
  AOI21_X1 U6060 ( .B1(n6601), .B2(n4935), .A(n4916), .ZN(n4918) );
  NAND2_X1 U6061 ( .A1(n5494), .A2(n5482), .ZN(n4917) );
  OAI211_X1 U6062 ( .C1(n5027), .C2(n6597), .A(n4918), .B(n4917), .ZN(U3131)
         );
  INV_X1 U6063 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4919) );
  OAI22_X1 U6064 ( .A1(n6553), .A2(n4933), .B1(n4932), .B2(n4919), .ZN(n4920)
         );
  AOI21_X1 U6065 ( .B1(n6556), .B2(n4935), .A(n4920), .ZN(n4922) );
  NAND2_X1 U6066 ( .A1(n5494), .A2(n5474), .ZN(n4921) );
  OAI211_X1 U6067 ( .C1(n5027), .C2(n6559), .A(n4922), .B(n4921), .ZN(U3125)
         );
  INV_X1 U6068 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4923) );
  OAI22_X1 U6069 ( .A1(n6574), .A2(n4933), .B1(n4932), .B2(n4923), .ZN(n4924)
         );
  AOI21_X1 U6070 ( .B1(n6577), .B2(n4935), .A(n4924), .ZN(n4926) );
  NAND2_X1 U6071 ( .A1(n5494), .A2(n5466), .ZN(n4925) );
  OAI211_X1 U6072 ( .C1(n5027), .C2(n6580), .A(n4926), .B(n4925), .ZN(U3128)
         );
  INV_X1 U6073 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4927) );
  OAI22_X1 U6074 ( .A1(n6534), .A2(n4933), .B1(n4932), .B2(n4927), .ZN(n4928)
         );
  AOI21_X1 U6075 ( .B1(n6549), .B2(n4935), .A(n4928), .ZN(n4930) );
  NAND2_X1 U6076 ( .A1(n5494), .A2(n5492), .ZN(n4929) );
  OAI211_X1 U6077 ( .C1(n5027), .C2(n6552), .A(n4930), .B(n4929), .ZN(U3124)
         );
  INV_X1 U6078 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4931) );
  OAI22_X1 U6079 ( .A1(n6581), .A2(n4933), .B1(n4932), .B2(n4931), .ZN(n4934)
         );
  AOI21_X1 U6080 ( .B1(n6584), .B2(n4935), .A(n4934), .ZN(n4937) );
  NAND2_X1 U6081 ( .A1(n5494), .A2(n5462), .ZN(n4936) );
  OAI211_X1 U6082 ( .C1(n5027), .C2(n6582), .A(n4937), .B(n4936), .ZN(U3129)
         );
  OAI21_X1 U6083 ( .B1(n4940), .B2(n4939), .A(n4938), .ZN(n4955) );
  AND2_X1 U6084 ( .A1(n6457), .A2(REIP_REG_6__SCAN_IN), .ZN(n4952) );
  NOR2_X1 U6085 ( .A1(n6111), .A2(n3959), .ZN(n4941) );
  AOI211_X1 U6086 ( .C1(n5808), .C2(n4942), .A(n4952), .B(n4941), .ZN(n4945)
         );
  NAND2_X1 U6087 ( .A1(n4943), .A2(n6378), .ZN(n4944) );
  OAI211_X1 U6088 ( .C1(n4955), .C2(n6164), .A(n4945), .B(n4944), .ZN(U2980)
         );
  NAND2_X1 U6090 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4947) );
  AOI21_X1 U6091 ( .B1(n5925), .B2(n4947), .A(n5923), .ZN(n6451) );
  INV_X1 U6092 ( .A(n6451), .ZN(n4946) );
  AOI21_X1 U6093 ( .B1(n4948), .B2(n5847), .A(n4946), .ZN(n6427) );
  OAI21_X1 U6094 ( .B1(n5922), .B2(n4947), .A(n6453), .ZN(n5306) );
  INV_X1 U6095 ( .A(n5306), .ZN(n6421) );
  OAI33_X1 U6096 ( .A1(1'b0), .A2(n6427), .A3(n4949), .B1(
        INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6421), .B3(n4948), .ZN(n4951) );
  AOI211_X1 U6097 ( .C1(n6448), .C2(n4953), .A(n4952), .B(n4951), .ZN(n4954)
         );
  OAI21_X1 U6098 ( .B1(n6138), .B2(n4955), .A(n4954), .ZN(U3012) );
  XNOR2_X1 U6099 ( .A(n4957), .B(n4956), .ZN(n6354) );
  INV_X1 U6100 ( .A(n6354), .ZN(n4971) );
  INV_X1 U6101 ( .A(n4977), .ZN(n4958) );
  AOI21_X1 U6102 ( .B1(n4959), .B2(n4841), .A(n4958), .ZN(n6411) );
  AOI22_X1 U6103 ( .A1(n6411), .A2(n6065), .B1(EBX_REG_7__SCAN_IN), .B2(n4506), 
        .ZN(n4960) );
  OAI21_X1 U6104 ( .B1(n4971), .B2(n5709), .A(n4960), .ZN(U2852) );
  NAND2_X1 U6105 ( .A1(n4965), .A2(n5596), .ZN(n4961) );
  NAND2_X1 U6106 ( .A1(n4961), .A2(n6192), .ZN(n6288) );
  INV_X1 U6107 ( .A(n6288), .ZN(n5238) );
  AOI22_X1 U6108 ( .A1(n6260), .A2(n4962), .B1(REIP_REG_0__SCAN_IN), .B2(n6261), .ZN(n4969) );
  INV_X1 U6109 ( .A(n4963), .ZN(n4964) );
  AND2_X1 U6110 ( .A1(n4965), .A2(n4964), .ZN(n6283) );
  NAND2_X1 U6111 ( .A1(n6283), .A2(n6616), .ZN(n4968) );
  NAND2_X1 U6112 ( .A1(n6282), .A2(EBX_REG_0__SCAN_IN), .ZN(n4967) );
  OAI21_X1 U6113 ( .B1(n6230), .B2(n6267), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4966) );
  AND4_X1 U6114 ( .A1(n4969), .A2(n4968), .A3(n4967), .A4(n4966), .ZN(n4970)
         );
  OAI21_X1 U6115 ( .B1(n5238), .B2(n6317), .A(n4970), .ZN(U2827) );
  INV_X1 U6116 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6334) );
  OAI222_X1 U6117 ( .A1(n6316), .A2(n4971), .B1(n6314), .B2(n6334), .C1(n7042), 
        .C2(n6315), .ZN(U2884) );
  OAI21_X1 U6118 ( .B1(n4972), .B2(n4975), .A(n4974), .ZN(n5071) );
  NAND2_X1 U6119 ( .A1(n4977), .A2(n4976), .ZN(n4978) );
  NAND2_X1 U6120 ( .A1(n5082), .A2(n4978), .ZN(n6404) );
  INV_X1 U6121 ( .A(n6404), .ZN(n4979) );
  AOI22_X1 U6122 ( .A1(n4979), .A2(n6065), .B1(EBX_REG_8__SCAN_IN), .B2(n4506), 
        .ZN(n4980) );
  OAI21_X1 U6123 ( .B1(n5071), .B2(n5709), .A(n4980), .ZN(U2851) );
  INV_X1 U6124 ( .A(n6271), .ZN(n6254) );
  INV_X1 U6125 ( .A(n5086), .ZN(n4981) );
  NAND2_X1 U6126 ( .A1(n6254), .A2(n4981), .ZN(n4983) );
  OAI22_X1 U6127 ( .A1(n6286), .A2(n6404), .B1(n4982), .B2(n4983), .ZN(n4987)
         );
  NAND2_X1 U6128 ( .A1(n4983), .A2(n5248), .ZN(n6233) );
  AOI22_X1 U6129 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n6230), .B1(
        REIP_REG_8__SCAN_IN), .B2(n6233), .ZN(n4984) );
  OAI211_X1 U6130 ( .C1(n6054), .C2(n4985), .A(n4984), .B(n6249), .ZN(n4986)
         );
  AOI211_X1 U6131 ( .C1(n5072), .C2(n6267), .A(n4987), .B(n4986), .ZN(n4988)
         );
  OAI21_X1 U6132 ( .B1(n6192), .B2(n5071), .A(n4988), .ZN(U2819) );
  INV_X1 U6133 ( .A(DATAI_8_), .ZN(n7033) );
  INV_X1 U6134 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6332) );
  OAI222_X1 U6135 ( .A1(n5071), .A2(n6316), .B1(n6315), .B2(n7033), .C1(n6314), 
        .C2(n6332), .ZN(U2883) );
  AOI21_X1 U6136 ( .B1(n5027), .B2(n6605), .A(n6163), .ZN(n4989) );
  AOI211_X1 U6137 ( .C1(n5373), .C2(n4990), .A(n6543), .B(n4989), .ZN(n4995)
         );
  NOR2_X1 U6138 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4991), .ZN(n5024)
         );
  AND2_X1 U6139 ( .A1(n4996), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5456) );
  INV_X1 U6140 ( .A(n5456), .ZN(n6473) );
  INV_X1 U6141 ( .A(n4992), .ZN(n5263) );
  NAND2_X1 U6142 ( .A1(n5263), .A2(n5322), .ZN(n5138) );
  AOI21_X1 U6143 ( .B1(n5138), .B2(STATE2_REG_2__SCAN_IN), .A(n4993), .ZN(
        n5133) );
  OAI211_X1 U6144 ( .C1(n6722), .C2(n5024), .A(n6473), .B(n5133), .ZN(n4994)
         );
  INV_X1 U6145 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5000) );
  NAND2_X1 U6146 ( .A1(n5373), .A2(n6537), .ZN(n5367) );
  INV_X1 U6147 ( .A(n4690), .ZN(n5973) );
  NOR2_X1 U6148 ( .A1(n4996), .A2(n6655), .ZN(n6465) );
  INV_X1 U6149 ( .A(n6465), .ZN(n5134) );
  OAI22_X1 U6150 ( .A1(n5367), .A2(n5973), .B1(n5134), .B2(n5138), .ZN(n5025)
         );
  AOI22_X1 U6151 ( .A1(n6549), .A2(n5025), .B1(n6469), .B2(n5024), .ZN(n4997)
         );
  OAI21_X1 U6152 ( .B1(n6535), .B2(n5027), .A(n4997), .ZN(n4998) );
  AOI21_X1 U6153 ( .B1(n6478), .B2(n5029), .A(n4998), .ZN(n4999) );
  OAI21_X1 U6154 ( .B1(n5032), .B2(n5000), .A(n4999), .ZN(U3116) );
  INV_X1 U6155 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5004) );
  AOI22_X1 U6156 ( .A1(n6570), .A2(n5025), .B1(n6489), .B2(n5024), .ZN(n5001)
         );
  OAI21_X1 U6157 ( .B1(n6568), .B2(n5027), .A(n5001), .ZN(n5002) );
  AOI21_X1 U6158 ( .B1(n6490), .B2(n5029), .A(n5002), .ZN(n5003) );
  OAI21_X1 U6159 ( .B1(n5032), .B2(n5004), .A(n5003), .ZN(U3119) );
  INV_X1 U6160 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5008) );
  AOI22_X1 U6161 ( .A1(n6601), .A2(n5025), .B1(n6506), .B2(n5024), .ZN(n5005)
         );
  OAI21_X1 U6162 ( .B1(n6606), .B2(n5027), .A(n5005), .ZN(n5006) );
  AOI21_X1 U6163 ( .B1(n6509), .B2(n5029), .A(n5006), .ZN(n5007) );
  OAI21_X1 U6164 ( .B1(n5032), .B2(n5008), .A(n5007), .ZN(U3123) );
  AOI22_X1 U6165 ( .A1(n6563), .A2(n5025), .B1(n6485), .B2(n5024), .ZN(n5009)
         );
  OAI21_X1 U6166 ( .B1(n6561), .B2(n5027), .A(n5009), .ZN(n5010) );
  AOI21_X1 U6167 ( .B1(n6486), .B2(n5029), .A(n5010), .ZN(n5011) );
  OAI21_X1 U6168 ( .B1(n5032), .B2(n3294), .A(n5011), .ZN(U3118) );
  INV_X1 U6169 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5015) );
  AOI22_X1 U6170 ( .A1(n6591), .A2(n5025), .B1(n6501), .B2(n5024), .ZN(n5012)
         );
  OAI21_X1 U6171 ( .B1(n6589), .B2(n5027), .A(n5012), .ZN(n5013) );
  AOI21_X1 U6172 ( .B1(n6502), .B2(n5029), .A(n5013), .ZN(n5014) );
  OAI21_X1 U6173 ( .B1(n5032), .B2(n5015), .A(n5014), .ZN(U3122) );
  INV_X1 U6174 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5019) );
  AOI22_X1 U6175 ( .A1(n6556), .A2(n5025), .B1(n6481), .B2(n5024), .ZN(n5016)
         );
  OAI21_X1 U6176 ( .B1(n6554), .B2(n5027), .A(n5016), .ZN(n5017) );
  AOI21_X1 U6177 ( .B1(n6482), .B2(n5029), .A(n5017), .ZN(n5018) );
  OAI21_X1 U6178 ( .B1(n5032), .B2(n5019), .A(n5018), .ZN(U3117) );
  INV_X1 U6179 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5023) );
  AOI22_X1 U6180 ( .A1(n6577), .A2(n5025), .B1(n6493), .B2(n5024), .ZN(n5020)
         );
  OAI21_X1 U6181 ( .B1(n6575), .B2(n5027), .A(n5020), .ZN(n5021) );
  AOI21_X1 U6182 ( .B1(n6494), .B2(n5029), .A(n5021), .ZN(n5022) );
  OAI21_X1 U6183 ( .B1(n5032), .B2(n5023), .A(n5022), .ZN(U3120) );
  INV_X1 U6184 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5031) );
  AOI22_X1 U6185 ( .A1(n6584), .A2(n5025), .B1(n6497), .B2(n5024), .ZN(n5026)
         );
  OAI21_X1 U6186 ( .B1(n6587), .B2(n5027), .A(n5026), .ZN(n5028) );
  AOI21_X1 U6187 ( .B1(n6498), .B2(n5029), .A(n5028), .ZN(n5030) );
  OAI21_X1 U6188 ( .B1(n5032), .B2(n5031), .A(n5030), .ZN(U3121) );
  NAND2_X1 U6189 ( .A1(n5039), .A2(n6598), .ZN(n5033) );
  AOI21_X1 U6190 ( .B1(n5033), .B2(STATEBS16_REG_SCAN_IN), .A(n6543), .ZN(
        n5037) );
  AND2_X1 U6191 ( .A1(n4591), .A2(n5034), .ZN(n5094) );
  AND2_X1 U6192 ( .A1(n5094), .A2(n4690), .ZN(n6541) );
  NOR3_X1 U6193 ( .A1(n6473), .A2(n5322), .A3(n6630), .ZN(n5035) );
  INV_X1 U6194 ( .A(n5322), .ZN(n6464) );
  OAI21_X1 U6195 ( .B1(n6464), .B2(n6655), .A(n5264), .ZN(n6475) );
  NOR2_X1 U6196 ( .A1(n6465), .A2(n6475), .ZN(n5320) );
  INV_X1 U6197 ( .A(n6541), .ZN(n5036) );
  NAND3_X1 U6198 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6625), .ZN(n6546) );
  OR2_X1 U6199 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6546), .ZN(n5062)
         );
  AOI22_X1 U6200 ( .A1(n5037), .A2(n5036), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5062), .ZN(n5038) );
  NAND2_X1 U6201 ( .A1(n5061), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5042)
         );
  OAI22_X1 U6202 ( .A1(n6598), .A2(n6575), .B1(n5062), .B2(n6574), .ZN(n5040)
         );
  AOI21_X1 U6203 ( .B1(n5064), .B2(n6494), .A(n5040), .ZN(n5041) );
  OAI211_X1 U6204 ( .C1(n5067), .C2(n5428), .A(n5042), .B(n5041), .ZN(U3104)
         );
  INV_X1 U6205 ( .A(n6570), .ZN(n5436) );
  NAND2_X1 U6206 ( .A1(n5061), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5045)
         );
  OAI22_X1 U6207 ( .A1(n6598), .A2(n6568), .B1(n5062), .B2(n6567), .ZN(n5043)
         );
  AOI21_X1 U6208 ( .B1(n5064), .B2(n6490), .A(n5043), .ZN(n5044) );
  OAI211_X1 U6209 ( .C1(n5067), .C2(n5436), .A(n5045), .B(n5044), .ZN(U3103)
         );
  NAND2_X1 U6210 ( .A1(n5061), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5048)
         );
  OAI22_X1 U6211 ( .A1(n6598), .A2(n6589), .B1(n5062), .B2(n6588), .ZN(n5046)
         );
  AOI21_X1 U6212 ( .B1(n5064), .B2(n6502), .A(n5046), .ZN(n5047) );
  OAI211_X1 U6213 ( .C1(n5067), .C2(n5444), .A(n5048), .B(n5047), .ZN(U3106)
         );
  NAND2_X1 U6214 ( .A1(n5061), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5051)
         );
  OAI22_X1 U6215 ( .A1(n6598), .A2(n6554), .B1(n5062), .B2(n6553), .ZN(n5049)
         );
  AOI21_X1 U6216 ( .B1(n5064), .B2(n6482), .A(n5049), .ZN(n5050) );
  OAI211_X1 U6217 ( .C1(n5067), .C2(n5432), .A(n5051), .B(n5050), .ZN(U3101)
         );
  NAND2_X1 U6218 ( .A1(n5061), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5054)
         );
  OAI22_X1 U6219 ( .A1(n6598), .A2(n6535), .B1(n6534), .B2(n5062), .ZN(n5052)
         );
  AOI21_X1 U6220 ( .B1(n5064), .B2(n6478), .A(n5052), .ZN(n5053) );
  OAI211_X1 U6221 ( .C1(n5067), .C2(n5451), .A(n5054), .B(n5053), .ZN(U3100)
         );
  NAND2_X1 U6222 ( .A1(n5061), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5057)
         );
  OAI22_X1 U6223 ( .A1(n6598), .A2(n6561), .B1(n5062), .B2(n6560), .ZN(n5055)
         );
  AOI21_X1 U6224 ( .B1(n5064), .B2(n6486), .A(n5055), .ZN(n5056) );
  OAI211_X1 U6225 ( .C1(n5067), .C2(n5424), .A(n5057), .B(n5056), .ZN(U3102)
         );
  NAND2_X1 U6226 ( .A1(n5061), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5060)
         );
  OAI22_X1 U6227 ( .A1(n6598), .A2(n6606), .B1(n5062), .B2(n6596), .ZN(n5058)
         );
  AOI21_X1 U6228 ( .B1(n5064), .B2(n6509), .A(n5058), .ZN(n5059) );
  OAI211_X1 U6229 ( .C1(n5067), .C2(n5420), .A(n5060), .B(n5059), .ZN(U3107)
         );
  NAND2_X1 U6230 ( .A1(n5061), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5066)
         );
  OAI22_X1 U6231 ( .A1(n6598), .A2(n6587), .B1(n5062), .B2(n6581), .ZN(n5063)
         );
  AOI21_X1 U6232 ( .B1(n5064), .B2(n6498), .A(n5063), .ZN(n5065) );
  OAI211_X1 U6233 ( .C1(n5067), .C2(n5440), .A(n5066), .B(n5065), .ZN(U3105)
         );
  OAI21_X1 U6234 ( .B1(n5070), .B2(n5069), .A(n5068), .ZN(n6401) );
  INV_X1 U6235 ( .A(n5071), .ZN(n5076) );
  INV_X1 U6236 ( .A(n5072), .ZN(n5074) );
  AOI22_X1 U6237 ( .A1(n6374), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6457), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5073) );
  OAI21_X1 U6238 ( .B1(n5074), .B2(n6384), .A(n5073), .ZN(n5075) );
  AOI21_X1 U6239 ( .B1(n5076), .B2(n6378), .A(n5075), .ZN(n5077) );
  OAI21_X1 U6240 ( .B1(n6401), .B2(n6164), .A(n5077), .ZN(U2978) );
  NAND2_X1 U6241 ( .A1(n4974), .A2(n5079), .ZN(n5080) );
  NAND2_X1 U6242 ( .A1(n5078), .A2(n5080), .ZN(n5221) );
  INV_X1 U6243 ( .A(DATAI_9_), .ZN(n7075) );
  INV_X1 U6244 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6330) );
  OAI222_X1 U6245 ( .A1(n5221), .A2(n6316), .B1(n6315), .B2(n7075), .C1(n6314), 
        .C2(n6330), .ZN(U2882) );
  INV_X1 U6246 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5084) );
  AND2_X1 U6247 ( .A1(n5082), .A2(n5081), .ZN(n5083) );
  OR2_X1 U6248 ( .A1(n5083), .A2(n5226), .ZN(n5085) );
  OAI222_X1 U6249 ( .A1(n5221), .A2(n5709), .B1(n5084), .B2(n6297), .C1(n6293), 
        .C2(n5085), .ZN(U2850) );
  INV_X1 U6250 ( .A(n5085), .ZN(n6394) );
  NAND2_X1 U6251 ( .A1(n6254), .A2(n5086), .ZN(n6228) );
  NOR2_X1 U6252 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6228), .ZN(n6234) );
  INV_X1 U6253 ( .A(n6234), .ZN(n5087) );
  OAI21_X1 U6254 ( .B1(n6280), .B2(n5217), .A(n5087), .ZN(n5090) );
  AOI22_X1 U6255 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6282), .B1(
        REIP_REG_9__SCAN_IN), .B2(n6233), .ZN(n5088) );
  OAI211_X1 U6256 ( .C1(n6279), .C2(n3981), .A(n5088), .B(n6249), .ZN(n5089)
         );
  AOI211_X1 U6257 ( .C1(n6394), .C2(n6260), .A(n5090), .B(n5089), .ZN(n5091)
         );
  OAI21_X1 U6258 ( .B1(n6192), .B2(n5221), .A(n5091), .ZN(U2818) );
  NAND2_X1 U6259 ( .A1(n5092), .A2(n6539), .ZN(n5970) );
  NOR3_X1 U6260 ( .A1(n5970), .A2(n3502), .A3(n6538), .ZN(n5093) );
  NOR2_X1 U6261 ( .A1(n5093), .A2(n6543), .ZN(n5100) );
  NOR2_X1 U6262 ( .A1(n6533), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5097)
         );
  AOI21_X1 U6263 ( .B1(n5324), .B2(n6616), .A(n5097), .ZN(n5099) );
  INV_X1 U6264 ( .A(n5099), .ZN(n5095) );
  NAND3_X1 U6265 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6630), .A3(n6625), .ZN(n5316) );
  INV_X1 U6266 ( .A(n5316), .ZN(n5102) );
  AOI22_X1 U6267 ( .A1(n5100), .A2(n5095), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5102), .ZN(n5128) );
  INV_X1 U6268 ( .A(n4798), .ZN(n5972) );
  NAND3_X1 U6269 ( .A1(n5972), .A2(n4776), .A3(n5964), .ZN(n5096) );
  NOR2_X2 U6270 ( .A1(n5096), .A2(n5415), .ZN(n5351) );
  INV_X1 U6271 ( .A(n5097), .ZN(n5123) );
  OAI22_X1 U6272 ( .A1(n5404), .A2(n6606), .B1(n6596), .B2(n5123), .ZN(n5098)
         );
  AOI21_X1 U6273 ( .B1(n6509), .B2(n5351), .A(n5098), .ZN(n5104) );
  NAND2_X1 U6274 ( .A1(n5100), .A2(n5099), .ZN(n5101) );
  NAND2_X1 U6275 ( .A1(n5125), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5103) );
  OAI211_X1 U6276 ( .C1(n5128), .C2(n5420), .A(n5104), .B(n5103), .ZN(U3051)
         );
  OAI22_X1 U6277 ( .A1(n5404), .A2(n6561), .B1(n6560), .B2(n5123), .ZN(n5105)
         );
  AOI21_X1 U6278 ( .B1(n6486), .B2(n5351), .A(n5105), .ZN(n5107) );
  NAND2_X1 U6279 ( .A1(n5125), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5106) );
  OAI211_X1 U6280 ( .C1(n5128), .C2(n5424), .A(n5107), .B(n5106), .ZN(U3046)
         );
  OAI22_X1 U6281 ( .A1(n5404), .A2(n6587), .B1(n6581), .B2(n5123), .ZN(n5108)
         );
  AOI21_X1 U6282 ( .B1(n6498), .B2(n5351), .A(n5108), .ZN(n5110) );
  NAND2_X1 U6283 ( .A1(n5125), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5109) );
  OAI211_X1 U6284 ( .C1(n5128), .C2(n5440), .A(n5110), .B(n5109), .ZN(U3049)
         );
  OAI22_X1 U6285 ( .A1(n5404), .A2(n6568), .B1(n6567), .B2(n5123), .ZN(n5111)
         );
  AOI21_X1 U6286 ( .B1(n6490), .B2(n5351), .A(n5111), .ZN(n5113) );
  NAND2_X1 U6287 ( .A1(n5125), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5112) );
  OAI211_X1 U6288 ( .C1(n5128), .C2(n5436), .A(n5113), .B(n5112), .ZN(U3047)
         );
  OAI22_X1 U6289 ( .A1(n5404), .A2(n6589), .B1(n6588), .B2(n5123), .ZN(n5114)
         );
  AOI21_X1 U6290 ( .B1(n6502), .B2(n5351), .A(n5114), .ZN(n5116) );
  NAND2_X1 U6291 ( .A1(n5125), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5115) );
  OAI211_X1 U6292 ( .C1(n5128), .C2(n5444), .A(n5116), .B(n5115), .ZN(U3050)
         );
  OAI22_X1 U6293 ( .A1(n5404), .A2(n6575), .B1(n6574), .B2(n5123), .ZN(n5117)
         );
  AOI21_X1 U6294 ( .B1(n6494), .B2(n5351), .A(n5117), .ZN(n5119) );
  NAND2_X1 U6295 ( .A1(n5125), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5118) );
  OAI211_X1 U6296 ( .C1(n5128), .C2(n5428), .A(n5119), .B(n5118), .ZN(U3048)
         );
  OAI22_X1 U6297 ( .A1(n5404), .A2(n6554), .B1(n6553), .B2(n5123), .ZN(n5120)
         );
  AOI21_X1 U6298 ( .B1(n6482), .B2(n5351), .A(n5120), .ZN(n5122) );
  NAND2_X1 U6299 ( .A1(n5125), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n5121) );
  OAI211_X1 U6300 ( .C1(n5128), .C2(n5432), .A(n5122), .B(n5121), .ZN(U3045)
         );
  OAI22_X1 U6301 ( .A1(n5404), .A2(n6535), .B1(n6534), .B2(n5123), .ZN(n5124)
         );
  AOI21_X1 U6302 ( .B1(n6478), .B2(n5351), .A(n5124), .ZN(n5127) );
  NAND2_X1 U6303 ( .A1(n5125), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n5126) );
  OAI211_X1 U6304 ( .C1(n5128), .C2(n5451), .A(n5127), .B(n5126), .ZN(U3044)
         );
  NAND3_X1 U6305 ( .A1(n5168), .A2(n6537), .A3(n6526), .ZN(n5131) );
  NOR2_X1 U6306 ( .A1(n6543), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5374) );
  INV_X1 U6307 ( .A(n5374), .ZN(n6471) );
  NOR2_X1 U6308 ( .A1(n5973), .A2(n5130), .ZN(n5137) );
  AOI21_X1 U6309 ( .B1(n5131), .B2(n6471), .A(n5137), .ZN(n5136) );
  NOR2_X1 U6310 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5132), .ZN(n5140)
         );
  OAI211_X1 U6311 ( .C1(n6722), .C2(n5140), .A(n5134), .B(n5133), .ZN(n5135)
         );
  NAND2_X1 U6312 ( .A1(n5162), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5143) );
  INV_X1 U6313 ( .A(n5137), .ZN(n5139) );
  OAI22_X1 U6314 ( .A1(n5139), .A2(n6543), .B1(n6473), .B2(n5138), .ZN(n5165)
         );
  INV_X1 U6315 ( .A(n5140), .ZN(n5163) );
  OAI22_X1 U6316 ( .A1(n6526), .A2(n6559), .B1(n6553), .B2(n5163), .ZN(n5141)
         );
  AOI21_X1 U6317 ( .B1(n6556), .B2(n5165), .A(n5141), .ZN(n5142) );
  OAI211_X1 U6318 ( .C1(n5168), .C2(n6554), .A(n5143), .B(n5142), .ZN(U3085)
         );
  NAND2_X1 U6319 ( .A1(n5162), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5146) );
  OAI22_X1 U6320 ( .A1(n6526), .A2(n6582), .B1(n6581), .B2(n5163), .ZN(n5144)
         );
  AOI21_X1 U6321 ( .B1(n6584), .B2(n5165), .A(n5144), .ZN(n5145) );
  OAI211_X1 U6322 ( .C1(n5168), .C2(n6587), .A(n5146), .B(n5145), .ZN(U3089)
         );
  NAND2_X1 U6323 ( .A1(n5162), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5149) );
  OAI22_X1 U6324 ( .A1(n6526), .A2(n6580), .B1(n6574), .B2(n5163), .ZN(n5147)
         );
  AOI21_X1 U6325 ( .B1(n6577), .B2(n5165), .A(n5147), .ZN(n5148) );
  OAI211_X1 U6326 ( .C1(n5168), .C2(n6575), .A(n5149), .B(n5148), .ZN(U3088)
         );
  NAND2_X1 U6327 ( .A1(n5162), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5152) );
  OAI22_X1 U6328 ( .A1(n6526), .A2(n6573), .B1(n6567), .B2(n5163), .ZN(n5150)
         );
  AOI21_X1 U6329 ( .B1(n6570), .B2(n5165), .A(n5150), .ZN(n5151) );
  OAI211_X1 U6330 ( .C1(n5168), .C2(n6568), .A(n5152), .B(n5151), .ZN(U3087)
         );
  NAND2_X1 U6331 ( .A1(n5162), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5155) );
  OAI22_X1 U6332 ( .A1(n6526), .A2(n6597), .B1(n6596), .B2(n5163), .ZN(n5153)
         );
  AOI21_X1 U6333 ( .B1(n6601), .B2(n5165), .A(n5153), .ZN(n5154) );
  OAI211_X1 U6334 ( .C1(n5168), .C2(n6606), .A(n5155), .B(n5154), .ZN(U3091)
         );
  NAND2_X1 U6335 ( .A1(n5162), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5158) );
  OAI22_X1 U6336 ( .A1(n6526), .A2(n6594), .B1(n6588), .B2(n5163), .ZN(n5156)
         );
  AOI21_X1 U6337 ( .B1(n6591), .B2(n5165), .A(n5156), .ZN(n5157) );
  OAI211_X1 U6338 ( .C1(n5168), .C2(n6589), .A(n5158), .B(n5157), .ZN(U3090)
         );
  NAND2_X1 U6339 ( .A1(n5162), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5161) );
  OAI22_X1 U6340 ( .A1(n6526), .A2(n6552), .B1(n6534), .B2(n5163), .ZN(n5159)
         );
  AOI21_X1 U6341 ( .B1(n6549), .B2(n5165), .A(n5159), .ZN(n5160) );
  OAI211_X1 U6342 ( .C1(n5168), .C2(n6535), .A(n5161), .B(n5160), .ZN(U3084)
         );
  NAND2_X1 U6343 ( .A1(n5162), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5167) );
  OAI22_X1 U6344 ( .A1(n6526), .A2(n6566), .B1(n6560), .B2(n5163), .ZN(n5164)
         );
  AOI21_X1 U6345 ( .B1(n6563), .B2(n5165), .A(n5164), .ZN(n5166) );
  OAI211_X1 U6346 ( .C1(n5168), .C2(n6561), .A(n5167), .B(n5166), .ZN(U3086)
         );
  OR2_X1 U6347 ( .A1(n6271), .A2(REIP_REG_1__SCAN_IN), .ZN(n5230) );
  AOI22_X1 U6348 ( .A1(n6230), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6262), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5169) );
  OAI211_X1 U6349 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6280), .A(n5230), 
        .B(n5169), .ZN(n5172) );
  INV_X1 U6350 ( .A(n6283), .ZN(n5170) );
  OAI22_X1 U6351 ( .A1(n4537), .A2(n5170), .B1(n6054), .B2(n4668), .ZN(n5171)
         );
  AOI211_X1 U6352 ( .C1(n6260), .C2(n4663), .A(n5172), .B(n5171), .ZN(n5173)
         );
  OAI21_X1 U6353 ( .B1(n5174), .B2(n5238), .A(n5173), .ZN(U2826) );
  INV_X1 U6354 ( .A(n5185), .ZN(n5177) );
  OAI21_X1 U6355 ( .B1(n5177), .B2(n6108), .A(n6471), .ZN(n5183) );
  INV_X1 U6356 ( .A(n5455), .ZN(n5460) );
  INV_X1 U6357 ( .A(n5178), .ZN(n5207) );
  AOI21_X1 U6358 ( .B1(n5179), .B2(n5460), .A(n5207), .ZN(n5184) );
  OAI21_X1 U6359 ( .B1(n6537), .B2(n5181), .A(n5180), .ZN(n5182) );
  INV_X1 U6360 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5188) );
  OAI22_X1 U6361 ( .A1(n5184), .A2(n6543), .B1(n5453), .B2(n6655), .ZN(n5208)
         );
  AOI22_X1 U6362 ( .A1(n6556), .A2(n5208), .B1(n5207), .B2(n6481), .ZN(n5187)
         );
  AOI22_X1 U6363 ( .A1(n6482), .A2(n5493), .B1(n3152), .B2(n5474), .ZN(n5186)
         );
  OAI211_X1 U6364 ( .C1(n5212), .C2(n5188), .A(n5187), .B(n5186), .ZN(U3141)
         );
  INV_X1 U6365 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5191) );
  AOI22_X1 U6366 ( .A1(n6584), .A2(n5208), .B1(n5207), .B2(n6497), .ZN(n5190)
         );
  AOI22_X1 U6367 ( .A1(n6498), .A2(n5493), .B1(n3152), .B2(n5462), .ZN(n5189)
         );
  OAI211_X1 U6368 ( .C1(n5212), .C2(n5191), .A(n5190), .B(n5189), .ZN(U3145)
         );
  INV_X1 U6369 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5194) );
  AOI22_X1 U6370 ( .A1(n6577), .A2(n5208), .B1(n5207), .B2(n6493), .ZN(n5193)
         );
  AOI22_X1 U6371 ( .A1(n6494), .A2(n5493), .B1(n3152), .B2(n5466), .ZN(n5192)
         );
  OAI211_X1 U6372 ( .C1(n5212), .C2(n5194), .A(n5193), .B(n5192), .ZN(U3144)
         );
  INV_X1 U6373 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5197) );
  AOI22_X1 U6374 ( .A1(n6570), .A2(n5208), .B1(n5207), .B2(n6489), .ZN(n5196)
         );
  AOI22_X1 U6375 ( .A1(n6490), .A2(n5493), .B1(n3152), .B2(n5486), .ZN(n5195)
         );
  OAI211_X1 U6376 ( .C1(n5212), .C2(n5197), .A(n5196), .B(n5195), .ZN(U3143)
         );
  INV_X1 U6377 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5200) );
  AOI22_X1 U6378 ( .A1(n6601), .A2(n5208), .B1(n5207), .B2(n6506), .ZN(n5199)
         );
  AOI22_X1 U6379 ( .A1(n6509), .A2(n5493), .B1(n3152), .B2(n5482), .ZN(n5198)
         );
  OAI211_X1 U6380 ( .C1(n5212), .C2(n5200), .A(n5199), .B(n5198), .ZN(U3147)
         );
  INV_X1 U6381 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5203) );
  AOI22_X1 U6382 ( .A1(n6591), .A2(n5208), .B1(n5207), .B2(n6501), .ZN(n5202)
         );
  AOI22_X1 U6383 ( .A1(n6502), .A2(n5493), .B1(n3152), .B2(n5478), .ZN(n5201)
         );
  OAI211_X1 U6384 ( .C1(n5212), .C2(n5203), .A(n5202), .B(n5201), .ZN(U3146)
         );
  INV_X1 U6385 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n5206) );
  AOI22_X1 U6386 ( .A1(n6549), .A2(n5208), .B1(n5207), .B2(n6469), .ZN(n5205)
         );
  AOI22_X1 U6387 ( .A1(n6478), .A2(n5493), .B1(n3152), .B2(n5492), .ZN(n5204)
         );
  OAI211_X1 U6388 ( .C1(n5212), .C2(n5206), .A(n5205), .B(n5204), .ZN(U3140)
         );
  INV_X1 U6389 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5211) );
  AOI22_X1 U6390 ( .A1(n6563), .A2(n5208), .B1(n5207), .B2(n6485), .ZN(n5210)
         );
  AOI22_X1 U6391 ( .A1(n6486), .A2(n5493), .B1(n3152), .B2(n5470), .ZN(n5209)
         );
  OAI211_X1 U6392 ( .C1(n5212), .C2(n5211), .A(n5210), .B(n5209), .ZN(U3142)
         );
  NAND2_X1 U6393 ( .A1(n5215), .A2(n5214), .ZN(n5216) );
  XNOR2_X1 U6394 ( .A(n5213), .B(n5216), .ZN(n6396) );
  NAND2_X1 U6395 ( .A1(n6396), .A2(n6380), .ZN(n5220) );
  AND2_X1 U6396 ( .A1(n6457), .A2(REIP_REG_9__SCAN_IN), .ZN(n6393) );
  NOR2_X1 U6397 ( .A1(n6384), .A2(n5217), .ZN(n5218) );
  AOI211_X1 U6398 ( .C1(n6374), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6393), 
        .B(n5218), .ZN(n5219) );
  OAI211_X1 U6399 ( .C1(n6108), .C2(n5221), .A(n5220), .B(n5219), .ZN(U2977)
         );
  AND2_X1 U6400 ( .A1(n5078), .A2(n5223), .ZN(n5224) );
  NOR2_X1 U6401 ( .A1(n5222), .A2(n5224), .ZN(n6232) );
  INV_X1 U6402 ( .A(n6232), .ZN(n5229) );
  INV_X1 U6403 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5227) );
  OAI21_X1 U6404 ( .B1(n5226), .B2(n5225), .A(n5244), .ZN(n5310) );
  OAI222_X1 U6405 ( .A1(n5229), .A2(n5709), .B1(n5227), .B2(n6297), .C1(n6293), 
        .C2(n5310), .ZN(U2849) );
  INV_X1 U6406 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6328) );
  OAI222_X1 U6407 ( .A1(n5229), .A2(n6316), .B1(n6315), .B2(n5228), .C1(n6314), 
        .C2(n6328), .ZN(U2881) );
  NAND2_X1 U6408 ( .A1(n5230), .A2(n5248), .ZN(n6276) );
  NOR2_X1 U6409 ( .A1(n6280), .A2(n6383), .ZN(n5232) );
  NOR3_X1 U6410 ( .A1(n6271), .A2(REIP_REG_2__SCAN_IN), .A3(n6733), .ZN(n5231)
         );
  AOI211_X1 U6411 ( .C1(n6230), .C2(PHYADDRPOINTER_REG_2__SCAN_IN), .A(n5232), 
        .B(n5231), .ZN(n5235) );
  INV_X1 U6412 ( .A(n4591), .ZN(n5233) );
  AOI22_X1 U6413 ( .A1(n5233), .A2(n6283), .B1(n6282), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n5234) );
  OAI211_X1 U6414 ( .C1(n6446), .C2(n6286), .A(n5235), .B(n5234), .ZN(n5236)
         );
  AOI21_X1 U6415 ( .B1(REIP_REG_2__SCAN_IN), .B2(n6276), .A(n5236), .ZN(n5237)
         );
  OAI21_X1 U6416 ( .B1(n5239), .B2(n5238), .A(n5237), .ZN(U2825) );
  INV_X1 U6417 ( .A(n5240), .ZN(n5241) );
  OAI21_X1 U6418 ( .B1(n5222), .B2(n5242), .A(n5241), .ZN(n5364) );
  AOI21_X1 U6419 ( .B1(n5245), .B2(n5244), .A(n5243), .ZN(n6386) );
  AOI22_X1 U6420 ( .A1(n6386), .A2(n6065), .B1(EBX_REG_11__SCAN_IN), .B2(n4506), .ZN(n5246) );
  OAI21_X1 U6421 ( .B1(n5364), .B2(n5709), .A(n5246), .ZN(U2848) );
  INV_X1 U6422 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6692) );
  INV_X1 U6423 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6690) );
  NOR4_X1 U6424 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6692), .A3(n6690), .A4(n6228), .ZN(n5255) );
  INV_X1 U6425 ( .A(n5512), .ZN(n5247) );
  NAND2_X1 U6426 ( .A1(n5248), .A2(n5247), .ZN(n5249) );
  NAND2_X1 U6427 ( .A1(n6261), .A2(n5249), .ZN(n6219) );
  INV_X1 U6428 ( .A(n6219), .ZN(n5513) );
  AOI22_X1 U6429 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6230), .B1(
        REIP_REG_11__SCAN_IN), .B2(n5513), .ZN(n5250) );
  OAI211_X1 U6430 ( .C1(n6054), .C2(n5251), .A(n5250), .B(n6249), .ZN(n5254)
         );
  INV_X1 U6431 ( .A(n6386), .ZN(n5252) );
  OAI22_X1 U6432 ( .A1(n5252), .A2(n6286), .B1(n5360), .B2(n6280), .ZN(n5253)
         );
  NOR3_X1 U6433 ( .A1(n5255), .A2(n5254), .A3(n5253), .ZN(n5256) );
  OAI21_X1 U6434 ( .B1(n5364), .B2(n6192), .A(n5256), .ZN(U2816) );
  OAI21_X1 U6435 ( .B1(n5240), .B2(n5258), .A(n5257), .ZN(n5523) );
  XNOR2_X1 U6436 ( .A(n5259), .B(n5504), .ZN(n6218) );
  AOI22_X1 U6437 ( .A1(n6218), .A2(n6065), .B1(EBX_REG_12__SCAN_IN), .B2(n4506), .ZN(n5260) );
  OAI21_X1 U6438 ( .B1(n5523), .B2(n5709), .A(n5260), .ZN(U2847) );
  INV_X1 U6439 ( .A(DATAI_12_), .ZN(n6875) );
  INV_X1 U6440 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6324) );
  OAI222_X1 U6441 ( .A1(n5523), .A2(n6316), .B1(n6315), .B2(n6875), .C1(n6314), 
        .C2(n6324), .ZN(U2879) );
  INV_X1 U6442 ( .A(DATAI_11_), .ZN(n7020) );
  INV_X1 U6443 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6326) );
  OAI222_X1 U6444 ( .A1(n5364), .A2(n6316), .B1(n6315), .B2(n7020), .C1(n6314), 
        .C2(n6326), .ZN(U2880) );
  NOR2_X1 U6445 ( .A1(n3152), .A2(n6543), .ZN(n5261) );
  AOI21_X1 U6446 ( .B1(n5261), .B2(n5296), .A(n5374), .ZN(n5266) );
  OR2_X1 U6447 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5262), .ZN(n5290)
         );
  NOR2_X1 U6448 ( .A1(n5263), .A2(n6464), .ZN(n5368) );
  OAI21_X1 U6449 ( .B1(n5368), .B2(n6655), .A(n5264), .ZN(n5375) );
  AOI211_X1 U6450 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5290), .A(n6465), .B(
        n5375), .ZN(n5265) );
  NAND2_X1 U6451 ( .A1(n5289), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5270) );
  AOI22_X1 U6452 ( .A1(n5267), .A2(n6537), .B1(n5456), .B2(n5368), .ZN(n5291)
         );
  OAI22_X1 U6453 ( .A1(n5436), .A2(n5291), .B1(n6567), .B2(n5290), .ZN(n5268)
         );
  AOI21_X1 U6454 ( .B1(n6490), .B2(n3152), .A(n5268), .ZN(n5269) );
  OAI211_X1 U6455 ( .C1(n5296), .C2(n6568), .A(n5270), .B(n5269), .ZN(U3023)
         );
  NAND2_X1 U6456 ( .A1(n5289), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5273) );
  OAI22_X1 U6457 ( .A1(n5420), .A2(n5291), .B1(n6596), .B2(n5290), .ZN(n5271)
         );
  AOI21_X1 U6458 ( .B1(n6509), .B2(n3152), .A(n5271), .ZN(n5272) );
  OAI211_X1 U6459 ( .C1(n5296), .C2(n6606), .A(n5273), .B(n5272), .ZN(U3027)
         );
  NAND2_X1 U6460 ( .A1(n5289), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5276) );
  OAI22_X1 U6461 ( .A1(n5451), .A2(n5291), .B1(n6534), .B2(n5290), .ZN(n5274)
         );
  AOI21_X1 U6462 ( .B1(n6478), .B2(n3152), .A(n5274), .ZN(n5275) );
  OAI211_X1 U6463 ( .C1(n5296), .C2(n6535), .A(n5276), .B(n5275), .ZN(U3020)
         );
  NAND2_X1 U6464 ( .A1(n5289), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5279) );
  OAI22_X1 U6465 ( .A1(n5428), .A2(n5291), .B1(n6574), .B2(n5290), .ZN(n5277)
         );
  AOI21_X1 U6466 ( .B1(n6494), .B2(n3152), .A(n5277), .ZN(n5278) );
  OAI211_X1 U6467 ( .C1(n5296), .C2(n6575), .A(n5279), .B(n5278), .ZN(U3024)
         );
  NAND2_X1 U6468 ( .A1(n5289), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5282) );
  OAI22_X1 U6469 ( .A1(n5432), .A2(n5291), .B1(n6553), .B2(n5290), .ZN(n5280)
         );
  AOI21_X1 U6470 ( .B1(n6482), .B2(n3152), .A(n5280), .ZN(n5281) );
  OAI211_X1 U6471 ( .C1(n5296), .C2(n6554), .A(n5282), .B(n5281), .ZN(U3021)
         );
  NAND2_X1 U6472 ( .A1(n5289), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5285) );
  OAI22_X1 U6473 ( .A1(n5424), .A2(n5291), .B1(n6560), .B2(n5290), .ZN(n5283)
         );
  AOI21_X1 U6474 ( .B1(n6486), .B2(n3152), .A(n5283), .ZN(n5284) );
  OAI211_X1 U6475 ( .C1(n5296), .C2(n6561), .A(n5285), .B(n5284), .ZN(U3022)
         );
  NAND2_X1 U6476 ( .A1(n5289), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5288) );
  OAI22_X1 U6477 ( .A1(n5444), .A2(n5291), .B1(n6588), .B2(n5290), .ZN(n5286)
         );
  AOI21_X1 U6478 ( .B1(n6502), .B2(n3152), .A(n5286), .ZN(n5287) );
  OAI211_X1 U6479 ( .C1(n5296), .C2(n6589), .A(n5288), .B(n5287), .ZN(U3026)
         );
  NAND2_X1 U6480 ( .A1(n5289), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5295) );
  OAI22_X1 U6481 ( .A1(n5440), .A2(n5291), .B1(n6581), .B2(n5290), .ZN(n5292)
         );
  AOI21_X1 U6482 ( .B1(n6498), .B2(n3152), .A(n5292), .ZN(n5294) );
  OAI211_X1 U6483 ( .C1(n5296), .C2(n6587), .A(n5295), .B(n5294), .ZN(U3025)
         );
  NAND2_X1 U6484 ( .A1(n5355), .A2(n5297), .ZN(n5299) );
  XOR2_X1 U6485 ( .A(n5299), .B(n5298), .Z(n5315) );
  AOI22_X1 U6486 ( .A1(n6374), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6457), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5300) );
  OAI21_X1 U6487 ( .B1(n6384), .B2(n5301), .A(n5300), .ZN(n5302) );
  AOI21_X1 U6488 ( .B1(n6232), .B2(n6378), .A(n5302), .ZN(n5303) );
  OAI21_X1 U6489 ( .B1(n5315), .B2(n6164), .A(n5303), .ZN(U2976) );
  OAI21_X1 U6490 ( .B1(n6453), .B2(n6420), .A(n6451), .ZN(n6432) );
  INV_X1 U6491 ( .A(n6432), .ZN(n6445) );
  AOI22_X1 U6492 ( .A1(n5304), .A2(n6445), .B1(n5939), .B2(n6451), .ZN(n5305)
         );
  INV_X1 U6493 ( .A(n5305), .ZN(n6417) );
  OAI21_X1 U6494 ( .B1(n6402), .B2(n5939), .A(n6417), .ZN(n6392) );
  NAND2_X1 U6495 ( .A1(n5307), .A2(n5306), .ZN(n6412) );
  NOR2_X1 U6496 ( .A1(n5308), .A2(n6412), .ZN(n6395) );
  OAI211_X1 U6497 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6395), .B(n5309), .ZN(n5312) );
  INV_X1 U6498 ( .A(n5310), .ZN(n6227) );
  NAND2_X1 U6499 ( .A1(n6227), .A2(n6448), .ZN(n5311) );
  OAI211_X1 U6500 ( .C1(n6692), .C2(n6403), .A(n5312), .B(n5311), .ZN(n5313)
         );
  AOI21_X1 U6501 ( .B1(n6392), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5313), 
        .ZN(n5314) );
  OAI21_X1 U6502 ( .B1(n5315), .B2(n6138), .A(n5314), .ZN(U3008) );
  NOR2_X1 U6503 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5316), .ZN(n5325)
         );
  OAI21_X1 U6504 ( .B1(n5351), .B2(n5317), .A(n6471), .ZN(n5319) );
  INV_X1 U6505 ( .A(n5324), .ZN(n5318) );
  NAND2_X1 U6506 ( .A1(n5319), .A2(n5318), .ZN(n5321) );
  NAND2_X1 U6507 ( .A1(n5347), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5328) );
  NOR3_X1 U6508 ( .A1(n6473), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n5322), 
        .ZN(n5323) );
  AOI21_X1 U6509 ( .B1(n5324), .B2(n6537), .A(n5323), .ZN(n5349) );
  INV_X1 U6510 ( .A(n5325), .ZN(n5348) );
  OAI22_X1 U6511 ( .A1(n5420), .A2(n5349), .B1(n6596), .B2(n5348), .ZN(n5326)
         );
  AOI21_X1 U6512 ( .B1(n5482), .B2(n5351), .A(n5326), .ZN(n5327) );
  OAI211_X1 U6513 ( .C1(n5354), .C2(n6597), .A(n5328), .B(n5327), .ZN(U3043)
         );
  NAND2_X1 U6514 ( .A1(n5347), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5331) );
  OAI22_X1 U6515 ( .A1(n5428), .A2(n5349), .B1(n6574), .B2(n5348), .ZN(n5329)
         );
  AOI21_X1 U6516 ( .B1(n5466), .B2(n5351), .A(n5329), .ZN(n5330) );
  OAI211_X1 U6517 ( .C1(n5354), .C2(n6580), .A(n5331), .B(n5330), .ZN(U3040)
         );
  NAND2_X1 U6518 ( .A1(n5347), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5334) );
  OAI22_X1 U6519 ( .A1(n5424), .A2(n5349), .B1(n6560), .B2(n5348), .ZN(n5332)
         );
  AOI21_X1 U6520 ( .B1(n5470), .B2(n5351), .A(n5332), .ZN(n5333) );
  OAI211_X1 U6521 ( .C1(n5354), .C2(n6566), .A(n5334), .B(n5333), .ZN(U3038)
         );
  NAND2_X1 U6522 ( .A1(n5347), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5337) );
  OAI22_X1 U6523 ( .A1(n5440), .A2(n5349), .B1(n6581), .B2(n5348), .ZN(n5335)
         );
  AOI21_X1 U6524 ( .B1(n5462), .B2(n5351), .A(n5335), .ZN(n5336) );
  OAI211_X1 U6525 ( .C1(n5354), .C2(n6582), .A(n5337), .B(n5336), .ZN(U3041)
         );
  NAND2_X1 U6526 ( .A1(n5347), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5340) );
  OAI22_X1 U6527 ( .A1(n5444), .A2(n5349), .B1(n6588), .B2(n5348), .ZN(n5338)
         );
  AOI21_X1 U6528 ( .B1(n5478), .B2(n5351), .A(n5338), .ZN(n5339) );
  OAI211_X1 U6529 ( .C1(n5354), .C2(n6594), .A(n5340), .B(n5339), .ZN(U3042)
         );
  NAND2_X1 U6530 ( .A1(n5347), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5343) );
  OAI22_X1 U6531 ( .A1(n5451), .A2(n5349), .B1(n6534), .B2(n5348), .ZN(n5341)
         );
  AOI21_X1 U6532 ( .B1(n5492), .B2(n5351), .A(n5341), .ZN(n5342) );
  OAI211_X1 U6533 ( .C1(n6552), .C2(n5354), .A(n5343), .B(n5342), .ZN(U3036)
         );
  NAND2_X1 U6534 ( .A1(n5347), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5346) );
  OAI22_X1 U6535 ( .A1(n5436), .A2(n5349), .B1(n6567), .B2(n5348), .ZN(n5344)
         );
  AOI21_X1 U6536 ( .B1(n5486), .B2(n5351), .A(n5344), .ZN(n5345) );
  OAI211_X1 U6537 ( .C1(n5354), .C2(n6573), .A(n5346), .B(n5345), .ZN(U3039)
         );
  NAND2_X1 U6538 ( .A1(n5347), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5353) );
  OAI22_X1 U6539 ( .A1(n5432), .A2(n5349), .B1(n6553), .B2(n5348), .ZN(n5350)
         );
  AOI21_X1 U6540 ( .B1(n5474), .B2(n5351), .A(n5350), .ZN(n5352) );
  OAI211_X1 U6541 ( .C1(n5354), .C2(n6559), .A(n5353), .B(n5352), .ZN(U3037)
         );
  NAND2_X1 U6542 ( .A1(n5356), .A2(n5355), .ZN(n5359) );
  XNOR2_X1 U6543 ( .A(n3658), .B(n5357), .ZN(n5358) );
  XNOR2_X1 U6544 ( .A(n5359), .B(n5358), .ZN(n6388) );
  NAND2_X1 U6545 ( .A1(n6388), .A2(n6380), .ZN(n5363) );
  AND2_X1 U6546 ( .A1(n6457), .A2(REIP_REG_11__SCAN_IN), .ZN(n6385) );
  NOR2_X1 U6547 ( .A1(n6384), .A2(n5360), .ZN(n5361) );
  AOI211_X1 U6548 ( .C1(n6374), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6385), 
        .B(n5361), .ZN(n5362) );
  OAI211_X1 U6549 ( .C1(n6108), .C2(n5364), .A(n5363), .B(n5362), .ZN(U2975)
         );
  INV_X1 U6550 ( .A(n5416), .ZN(n5366) );
  NOR2_X2 U6551 ( .A1(n5366), .A2(n5415), .ZN(n5448) );
  INV_X1 U6552 ( .A(n5367), .ZN(n5369) );
  AOI22_X1 U6553 ( .A1(n5369), .A2(n5973), .B1(n6465), .B2(n5368), .ZN(n5399)
         );
  NAND3_X1 U6554 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6630), .A3(n5370), .ZN(n5411) );
  OR2_X1 U6555 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5411), .ZN(n5398)
         );
  OAI22_X1 U6556 ( .A1(n5420), .A2(n5399), .B1(n6596), .B2(n5398), .ZN(n5371)
         );
  AOI21_X1 U6557 ( .B1(n5482), .B2(n5448), .A(n5371), .ZN(n5379) );
  AOI21_X1 U6558 ( .B1(n5416), .B2(STATEBS16_REG_SCAN_IN), .A(n6543), .ZN(
        n5410) );
  NAND2_X1 U6559 ( .A1(n5373), .A2(n5372), .ZN(n5406) );
  OAI211_X1 U6560 ( .C1(n5404), .C2(n5374), .A(n5410), .B(n5406), .ZN(n5377)
         );
  AOI211_X1 U6561 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5398), .A(n5456), .B(
        n5375), .ZN(n5376) );
  NAND2_X1 U6562 ( .A1(n5377), .A2(n5376), .ZN(n5401) );
  NAND2_X1 U6563 ( .A1(n5401), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5378) );
  OAI211_X1 U6564 ( .C1(n5404), .C2(n6597), .A(n5379), .B(n5378), .ZN(U3059)
         );
  OAI22_X1 U6565 ( .A1(n5440), .A2(n5399), .B1(n6581), .B2(n5398), .ZN(n5380)
         );
  AOI21_X1 U6566 ( .B1(n5462), .B2(n5448), .A(n5380), .ZN(n5382) );
  NAND2_X1 U6567 ( .A1(n5401), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5381) );
  OAI211_X1 U6568 ( .C1(n5404), .C2(n6582), .A(n5382), .B(n5381), .ZN(U3057)
         );
  OAI22_X1 U6569 ( .A1(n5444), .A2(n5399), .B1(n6588), .B2(n5398), .ZN(n5383)
         );
  AOI21_X1 U6570 ( .B1(n5478), .B2(n5448), .A(n5383), .ZN(n5385) );
  NAND2_X1 U6571 ( .A1(n5401), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5384) );
  OAI211_X1 U6572 ( .C1(n5404), .C2(n6594), .A(n5385), .B(n5384), .ZN(U3058)
         );
  OAI22_X1 U6573 ( .A1(n5432), .A2(n5399), .B1(n6553), .B2(n5398), .ZN(n5386)
         );
  AOI21_X1 U6574 ( .B1(n5474), .B2(n5448), .A(n5386), .ZN(n5388) );
  NAND2_X1 U6575 ( .A1(n5401), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5387) );
  OAI211_X1 U6576 ( .C1(n5404), .C2(n6559), .A(n5388), .B(n5387), .ZN(U3053)
         );
  OAI22_X1 U6577 ( .A1(n5424), .A2(n5399), .B1(n6560), .B2(n5398), .ZN(n5389)
         );
  AOI21_X1 U6578 ( .B1(n5470), .B2(n5448), .A(n5389), .ZN(n5391) );
  NAND2_X1 U6579 ( .A1(n5401), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5390) );
  OAI211_X1 U6580 ( .C1(n5404), .C2(n6566), .A(n5391), .B(n5390), .ZN(U3054)
         );
  OAI22_X1 U6581 ( .A1(n5428), .A2(n5399), .B1(n6574), .B2(n5398), .ZN(n5392)
         );
  AOI21_X1 U6582 ( .B1(n5466), .B2(n5448), .A(n5392), .ZN(n5394) );
  NAND2_X1 U6583 ( .A1(n5401), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5393) );
  OAI211_X1 U6584 ( .C1(n5404), .C2(n6580), .A(n5394), .B(n5393), .ZN(U3056)
         );
  OAI22_X1 U6585 ( .A1(n5436), .A2(n5399), .B1(n6567), .B2(n5398), .ZN(n5395)
         );
  AOI21_X1 U6586 ( .B1(n5486), .B2(n5448), .A(n5395), .ZN(n5397) );
  NAND2_X1 U6587 ( .A1(n5401), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5396) );
  OAI211_X1 U6588 ( .C1(n5404), .C2(n6573), .A(n5397), .B(n5396), .ZN(U3055)
         );
  OAI22_X1 U6589 ( .A1(n5451), .A2(n5399), .B1(n6534), .B2(n5398), .ZN(n5400)
         );
  AOI21_X1 U6590 ( .B1(n5492), .B2(n5448), .A(n5400), .ZN(n5403) );
  NAND2_X1 U6591 ( .A1(n5401), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5402) );
  OAI211_X1 U6592 ( .C1(n5404), .C2(n6552), .A(n5403), .B(n5402), .ZN(U3052)
         );
  OR2_X1 U6593 ( .A1(n5406), .A2(n5405), .ZN(n5408) );
  OR2_X1 U6594 ( .A1(n5407), .A2(n5411), .ZN(n5446) );
  NAND2_X1 U6595 ( .A1(n5408), .A2(n5446), .ZN(n5413) );
  INV_X1 U6596 ( .A(n5411), .ZN(n5409) );
  AOI22_X1 U6597 ( .A1(n5410), .A2(n5413), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5409), .ZN(n5452) );
  INV_X1 U6598 ( .A(n5410), .ZN(n5414) );
  AOI21_X1 U6599 ( .B1(n6543), .B2(n5411), .A(n6542), .ZN(n5412) );
  NAND2_X1 U6600 ( .A1(n5445), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U6601 ( .A1(n5416), .A2(n5415), .ZN(n6477) );
  OAI22_X1 U6602 ( .A1(n6477), .A2(n6606), .B1(n6596), .B2(n5446), .ZN(n5417)
         );
  AOI21_X1 U6603 ( .B1(n6509), .B2(n5448), .A(n5417), .ZN(n5418) );
  OAI211_X1 U6604 ( .C1(n5452), .C2(n5420), .A(n5419), .B(n5418), .ZN(U3067)
         );
  NAND2_X1 U6605 ( .A1(n5445), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5423) );
  OAI22_X1 U6606 ( .A1(n6477), .A2(n6561), .B1(n6560), .B2(n5446), .ZN(n5421)
         );
  AOI21_X1 U6607 ( .B1(n6486), .B2(n5448), .A(n5421), .ZN(n5422) );
  OAI211_X1 U6608 ( .C1(n5452), .C2(n5424), .A(n5423), .B(n5422), .ZN(U3062)
         );
  NAND2_X1 U6609 ( .A1(n5445), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5427) );
  OAI22_X1 U6610 ( .A1(n6477), .A2(n6575), .B1(n6574), .B2(n5446), .ZN(n5425)
         );
  AOI21_X1 U6611 ( .B1(n6494), .B2(n5448), .A(n5425), .ZN(n5426) );
  OAI211_X1 U6612 ( .C1(n5452), .C2(n5428), .A(n5427), .B(n5426), .ZN(U3064)
         );
  NAND2_X1 U6613 ( .A1(n5445), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n5431) );
  OAI22_X1 U6614 ( .A1(n6477), .A2(n6554), .B1(n6553), .B2(n5446), .ZN(n5429)
         );
  AOI21_X1 U6615 ( .B1(n6482), .B2(n5448), .A(n5429), .ZN(n5430) );
  OAI211_X1 U6616 ( .C1(n5452), .C2(n5432), .A(n5431), .B(n5430), .ZN(U3061)
         );
  NAND2_X1 U6617 ( .A1(n5445), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5435) );
  OAI22_X1 U6618 ( .A1(n6477), .A2(n6568), .B1(n6567), .B2(n5446), .ZN(n5433)
         );
  AOI21_X1 U6619 ( .B1(n6490), .B2(n5448), .A(n5433), .ZN(n5434) );
  OAI211_X1 U6620 ( .C1(n5452), .C2(n5436), .A(n5435), .B(n5434), .ZN(U3063)
         );
  NAND2_X1 U6621 ( .A1(n5445), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n5439) );
  OAI22_X1 U6622 ( .A1(n6477), .A2(n6587), .B1(n6581), .B2(n5446), .ZN(n5437)
         );
  AOI21_X1 U6623 ( .B1(n6498), .B2(n5448), .A(n5437), .ZN(n5438) );
  OAI211_X1 U6624 ( .C1(n5452), .C2(n5440), .A(n5439), .B(n5438), .ZN(U3065)
         );
  NAND2_X1 U6625 ( .A1(n5445), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5443) );
  OAI22_X1 U6626 ( .A1(n6477), .A2(n6589), .B1(n6588), .B2(n5446), .ZN(n5441)
         );
  AOI21_X1 U6627 ( .B1(n6502), .B2(n5448), .A(n5441), .ZN(n5442) );
  OAI211_X1 U6628 ( .C1(n5452), .C2(n5444), .A(n5443), .B(n5442), .ZN(U3066)
         );
  NAND2_X1 U6629 ( .A1(n5445), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n5450) );
  OAI22_X1 U6630 ( .A1(n6477), .A2(n6535), .B1(n6534), .B2(n5446), .ZN(n5447)
         );
  AOI21_X1 U6631 ( .B1(n6478), .B2(n5448), .A(n5447), .ZN(n5449) );
  OAI211_X1 U6632 ( .C1(n5452), .C2(n5451), .A(n5450), .B(n5449), .ZN(U3060)
         );
  NOR2_X1 U6633 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5453), .ZN(n5490)
         );
  OAI21_X1 U6634 ( .B1(n5494), .B2(n5493), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5454) );
  NAND3_X1 U6635 ( .A1(n5455), .A2(n6537), .A3(n5454), .ZN(n5458) );
  NOR3_X1 U6636 ( .A1(n6475), .A2(n6630), .A3(n5456), .ZN(n5457) );
  OAI211_X1 U6637 ( .C1(n5490), .C2(n6722), .A(n5458), .B(n5457), .ZN(n5459)
         );
  INV_X1 U6638 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U6639 ( .A1(n5460), .A2(n6537), .ZN(n6467) );
  NAND3_X1 U6640 ( .A1(n6465), .A2(n6464), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5461) );
  OAI21_X1 U6641 ( .B1(n6467), .B2(n5973), .A(n5461), .ZN(n5491) );
  AOI22_X1 U6642 ( .A1(n6584), .A2(n5491), .B1(n6497), .B2(n5490), .ZN(n5464)
         );
  AOI22_X1 U6643 ( .A1(n6498), .A2(n5494), .B1(n5493), .B2(n5462), .ZN(n5463)
         );
  OAI211_X1 U6644 ( .C1(n5498), .C2(n5465), .A(n5464), .B(n5463), .ZN(U3137)
         );
  INV_X1 U6645 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5469) );
  AOI22_X1 U6646 ( .A1(n6577), .A2(n5491), .B1(n6493), .B2(n5490), .ZN(n5468)
         );
  AOI22_X1 U6647 ( .A1(n6494), .A2(n5494), .B1(n5493), .B2(n5466), .ZN(n5467)
         );
  OAI211_X1 U6648 ( .C1(n5498), .C2(n5469), .A(n5468), .B(n5467), .ZN(U3136)
         );
  INV_X1 U6649 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5473) );
  AOI22_X1 U6650 ( .A1(n6563), .A2(n5491), .B1(n6485), .B2(n5490), .ZN(n5472)
         );
  AOI22_X1 U6651 ( .A1(n6486), .A2(n5494), .B1(n5493), .B2(n5470), .ZN(n5471)
         );
  OAI211_X1 U6652 ( .C1(n5498), .C2(n5473), .A(n5472), .B(n5471), .ZN(U3134)
         );
  INV_X1 U6653 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5477) );
  AOI22_X1 U6654 ( .A1(n6556), .A2(n5491), .B1(n6481), .B2(n5490), .ZN(n5476)
         );
  AOI22_X1 U6655 ( .A1(n6482), .A2(n5494), .B1(n5493), .B2(n5474), .ZN(n5475)
         );
  OAI211_X1 U6656 ( .C1(n5498), .C2(n5477), .A(n5476), .B(n5475), .ZN(U3133)
         );
  INV_X1 U6657 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5481) );
  AOI22_X1 U6658 ( .A1(n6591), .A2(n5491), .B1(n6501), .B2(n5490), .ZN(n5480)
         );
  AOI22_X1 U6659 ( .A1(n6502), .A2(n5494), .B1(n5493), .B2(n5478), .ZN(n5479)
         );
  OAI211_X1 U6660 ( .C1(n5498), .C2(n5481), .A(n5480), .B(n5479), .ZN(U3138)
         );
  INV_X1 U6661 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5485) );
  AOI22_X1 U6662 ( .A1(n6601), .A2(n5491), .B1(n6506), .B2(n5490), .ZN(n5484)
         );
  AOI22_X1 U6663 ( .A1(n6509), .A2(n5494), .B1(n5493), .B2(n5482), .ZN(n5483)
         );
  OAI211_X1 U6664 ( .C1(n5498), .C2(n5485), .A(n5484), .B(n5483), .ZN(U3139)
         );
  INV_X1 U6665 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5489) );
  AOI22_X1 U6666 ( .A1(n6570), .A2(n5491), .B1(n6489), .B2(n5490), .ZN(n5488)
         );
  AOI22_X1 U6667 ( .A1(n6490), .A2(n5494), .B1(n5493), .B2(n5486), .ZN(n5487)
         );
  OAI211_X1 U6668 ( .C1(n5498), .C2(n5489), .A(n5488), .B(n5487), .ZN(U3135)
         );
  INV_X1 U6669 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5497) );
  AOI22_X1 U6670 ( .A1(n6549), .A2(n5491), .B1(n6469), .B2(n5490), .ZN(n5496)
         );
  AOI22_X1 U6671 ( .A1(n6478), .A2(n5494), .B1(n5493), .B2(n5492), .ZN(n5495)
         );
  OAI211_X1 U6672 ( .C1(n5498), .C2(n5497), .A(n5496), .B(n5495), .ZN(U3132)
         );
  OR2_X1 U6673 ( .A1(n5501), .A2(n5500), .ZN(n5502) );
  NAND2_X1 U6674 ( .A1(n5499), .A2(n5502), .ZN(n5824) );
  AOI21_X1 U6675 ( .B1(n5243), .B2(n5504), .A(n5503), .ZN(n5506) );
  OR2_X1 U6676 ( .A1(n5506), .A2(n5505), .ZN(n5510) );
  OAI22_X1 U6677 ( .A1(n5510), .A2(n6293), .B1(n5507), .B2(n6297), .ZN(n5508)
         );
  INV_X1 U6678 ( .A(n5508), .ZN(n5509) );
  OAI21_X1 U6679 ( .B1(n5824), .B2(n5709), .A(n5509), .ZN(U2846) );
  INV_X1 U6680 ( .A(n5510), .ZN(n6150) );
  AOI22_X1 U6681 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6282), .B1(n6260), .B2(n6150), .ZN(n5511) );
  OAI211_X1 U6682 ( .C1(n6279), .C2(n4045), .A(n5511), .B(n6249), .ZN(n5518)
         );
  NOR3_X1 U6683 ( .A1(n6271), .A2(REIP_REG_12__SCAN_IN), .A3(n5512), .ZN(n6221) );
  OAI21_X1 U6684 ( .B1(n6221), .B2(n5513), .A(REIP_REG_13__SCAN_IN), .ZN(n5516) );
  INV_X1 U6685 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6696) );
  NAND3_X1 U6686 ( .A1(n6254), .A2(n6696), .A3(n5514), .ZN(n5515) );
  OAI211_X1 U6687 ( .C1(n5820), .C2(n6280), .A(n5516), .B(n5515), .ZN(n5517)
         );
  NOR2_X1 U6688 ( .A1(n5518), .A2(n5517), .ZN(n5519) );
  OAI21_X1 U6689 ( .B1(n5824), .B2(n6192), .A(n5519), .ZN(U2814) );
  NOR2_X1 U6690 ( .A1(n5521), .A2(n3168), .ZN(n5522) );
  XNOR2_X1 U6691 ( .A(n5520), .B(n5522), .ZN(n5539) );
  INV_X1 U6692 ( .A(n5523), .ZN(n6223) );
  INV_X1 U6693 ( .A(n6222), .ZN(n5525) );
  AOI22_X1 U6694 ( .A1(n6374), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n6457), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n5524) );
  OAI21_X1 U6695 ( .B1(n6384), .B2(n5525), .A(n5524), .ZN(n5526) );
  AOI21_X1 U6696 ( .B1(n6223), .B2(n6378), .A(n5526), .ZN(n5527) );
  OAI21_X1 U6697 ( .B1(n5539), .B2(n6164), .A(n5527), .ZN(U2974) );
  INV_X1 U6698 ( .A(n6156), .ZN(n6387) );
  NAND3_X1 U6699 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n5534), .A3(n6387), .ZN(n5529) );
  NAND2_X1 U6700 ( .A1(n6218), .A2(n6448), .ZN(n5528) );
  OAI211_X1 U6701 ( .C1(n6694), .C2(n6403), .A(n5529), .B(n5528), .ZN(n5537)
         );
  AOI21_X1 U6702 ( .B1(n5925), .B2(n5926), .A(n5923), .ZN(n5530) );
  INV_X1 U6703 ( .A(n5530), .ZN(n5531) );
  AOI21_X1 U6704 ( .B1(n6450), .B2(n5532), .A(n5531), .ZN(n6391) );
  OAI21_X1 U6705 ( .B1(n6450), .B2(n5533), .A(n5357), .ZN(n5535) );
  AOI21_X1 U6706 ( .B1(n6391), .B2(n5535), .A(n5534), .ZN(n5536) );
  NOR2_X1 U6707 ( .A1(n5537), .A2(n5536), .ZN(n5538) );
  OAI21_X1 U6708 ( .B1(n5539), .B2(n6138), .A(n5538), .ZN(U3006) );
  INV_X1 U6709 ( .A(DATAI_13_), .ZN(n7001) );
  INV_X1 U6710 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6322) );
  OAI222_X1 U6711 ( .A1(n5824), .A2(n6316), .B1(n6315), .B2(n7001), .C1(n6314), 
        .C2(n6322), .ZN(U2878) );
  INV_X1 U6712 ( .A(n5542), .ZN(n5544) );
  NAND3_X1 U6713 ( .A1(n5499), .A2(n5544), .A3(n5543), .ZN(n5545) );
  AND2_X1 U6714 ( .A1(n5541), .A2(n5545), .ZN(n6214) );
  INV_X1 U6715 ( .A(n6214), .ZN(n5550) );
  INV_X1 U6716 ( .A(n6315), .ZN(n5562) );
  AOI22_X1 U6717 ( .A1(n5562), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n6311), .ZN(n5546) );
  OAI21_X1 U6718 ( .B1(n5550), .B2(n6316), .A(n5546), .ZN(U2877) );
  INV_X1 U6719 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5549) );
  INV_X1 U6720 ( .A(n5555), .ZN(n5547) );
  OAI21_X1 U6721 ( .B1(n5505), .B2(n5548), .A(n5547), .ZN(n6217) );
  OAI222_X1 U6722 ( .A1(n5550), .A2(n5709), .B1(n6297), .B2(n5549), .C1(n6217), 
        .C2(n6293), .ZN(U2845) );
  INV_X1 U6723 ( .A(n5541), .ZN(n5553) );
  OAI21_X1 U6724 ( .B1(n5553), .B2(n4095), .A(n5552), .ZN(n5811) );
  OAI21_X1 U6725 ( .B1(n5555), .B2(n5554), .A(n5700), .ZN(n5707) );
  INV_X1 U6726 ( .A(n5707), .ZN(n6142) );
  NAND2_X1 U6727 ( .A1(n6267), .A2(n5807), .ZN(n5556) );
  OAI211_X1 U6728 ( .C1(n6279), .C2(n4097), .A(n5556), .B(n6249), .ZN(n5560)
         );
  AND2_X1 U6729 ( .A1(n6261), .A2(n5557), .ZN(n6211) );
  AOI22_X1 U6730 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6282), .B1(
        REIP_REG_15__SCAN_IN), .B2(n6211), .ZN(n5558) );
  OAI21_X1 U6731 ( .B1(REIP_REG_15__SCAN_IN), .B2(n6200), .A(n5558), .ZN(n5559) );
  AOI211_X1 U6732 ( .C1(n6142), .C2(n6260), .A(n5560), .B(n5559), .ZN(n5561)
         );
  OAI21_X1 U6733 ( .B1(n5811), .B2(n6192), .A(n5561), .ZN(U2812) );
  AOI22_X1 U6734 ( .A1(n5562), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6311), .ZN(n5563) );
  OAI21_X1 U6735 ( .B1(n5811), .B2(n6316), .A(n5563), .ZN(U2876) );
  INV_X1 U6736 ( .A(n5727), .ZN(n5737) );
  NAND2_X1 U6737 ( .A1(n5737), .A2(n5564), .ZN(n5566) );
  XNOR2_X1 U6738 ( .A(n5567), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5873)
         );
  INV_X1 U6739 ( .A(n5983), .ZN(n5573) );
  NAND2_X1 U6740 ( .A1(n6457), .A2(REIP_REG_28__SCAN_IN), .ZN(n5867) );
  OAI21_X1 U6741 ( .B1(n6111), .B2(n5568), .A(n5867), .ZN(n5569) );
  INV_X1 U6742 ( .A(n5569), .ZN(n5572) );
  INV_X1 U6743 ( .A(n5574), .ZN(n5575) );
  OAI21_X1 U6744 ( .B1(n6164), .B2(n5873), .A(n5575), .ZN(U2958) );
  OR2_X1 U6745 ( .A1(n5649), .A2(n5577), .ZN(n5578) );
  NAND2_X1 U6746 ( .A1(n4469), .A2(n5578), .ZN(n5984) );
  INV_X1 U6747 ( .A(n5984), .ZN(n5871) );
  AOI22_X1 U6748 ( .A1(n5871), .A2(n6065), .B1(EBX_REG_28__SCAN_IN), .B2(n4506), .ZN(n5579) );
  OAI21_X1 U6749 ( .B1(n5576), .B2(n5709), .A(n5579), .ZN(U2831) );
  AOI22_X1 U6750 ( .A1(n6307), .A2(DATAI_28_), .B1(n6311), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U6751 ( .A1(n6310), .A2(DATAI_12_), .ZN(n5580) );
  OAI211_X1 U6752 ( .C1(n5576), .C2(n6316), .A(n5581), .B(n5580), .ZN(U2863)
         );
  AND2_X1 U6753 ( .A1(n6314), .A2(n5582), .ZN(n5583) );
  NAND2_X1 U6754 ( .A1(n5584), .A2(n5583), .ZN(n5586) );
  AOI22_X1 U6755 ( .A1(n6307), .A2(DATAI_31_), .B1(n6311), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U6756 ( .A1(n5586), .A2(n5585), .ZN(U2860) );
  NAND2_X1 U6757 ( .A1(n6607), .A2(n5599), .ZN(n5587) );
  NOR2_X1 U6758 ( .A1(n5588), .A2(n5587), .ZN(n5591) );
  OAI22_X1 U6759 ( .A1(n5597), .A2(n5591), .B1(n5590), .B2(n5589), .ZN(n5592)
         );
  INV_X1 U6760 ( .A(n5592), .ZN(n5595) );
  NAND2_X1 U6761 ( .A1(n5593), .A2(n5597), .ZN(n5594) );
  AND2_X1 U6762 ( .A1(n5595), .A2(n5594), .ZN(n6608) );
  INV_X1 U6763 ( .A(n6608), .ZN(n5607) );
  OR2_X1 U6764 ( .A1(n5597), .A2(n5596), .ZN(n5602) );
  INV_X1 U6765 ( .A(n5598), .ZN(n5600) );
  NAND2_X1 U6766 ( .A1(n5600), .A2(n5599), .ZN(n5601) );
  NAND2_X1 U6767 ( .A1(n5602), .A2(n5601), .ZN(n6158) );
  OR2_X1 U6768 ( .A1(n5604), .A2(n5603), .ZN(n5606) );
  INV_X1 U6769 ( .A(READY_N), .ZN(n5605) );
  AND2_X1 U6770 ( .A1(n5606), .A2(n5605), .ZN(n6744) );
  OR2_X1 U6771 ( .A1(n6158), .A2(n6744), .ZN(n6610) );
  AND2_X1 U6772 ( .A1(n6610), .A2(n6652), .ZN(n6165) );
  MUX2_X1 U6773 ( .A(MORE_REG_SCAN_IN), .B(n5607), .S(n6165), .Z(U3471) );
  INV_X1 U6774 ( .A(n5735), .ZN(n5712) );
  OAI22_X1 U6775 ( .A1(n5608), .A2(n6054), .B1(n5733), .B2(n6279), .ZN(n5609)
         );
  AOI21_X1 U6776 ( .B1(n6267), .B2(n5731), .A(n5609), .ZN(n5610) );
  OAI21_X1 U6777 ( .B1(n5844), .B2(n6286), .A(n5610), .ZN(n5612) );
  AOI211_X1 U6778 ( .C1(REIP_REG_30__SCAN_IN), .C2(n5613), .A(n5612), .B(n5611), .ZN(n5614) );
  OAI21_X1 U6779 ( .B1(n5712), .B2(n6192), .A(n5614), .ZN(U2797) );
  AND2_X1 U6780 ( .A1(n4469), .A2(n5615), .ZN(n5616) );
  AOI21_X1 U6781 ( .B1(n5620), .B2(n5618), .A(n5619), .ZN(n5744) );
  NAND2_X1 U6782 ( .A1(n5744), .A2(n6244), .ZN(n5626) );
  OAI22_X1 U6783 ( .A1(n5644), .A2(n6054), .B1(n4348), .B2(n6279), .ZN(n5624)
         );
  OAI22_X1 U6784 ( .A1(n5986), .A2(n7097), .B1(n5742), .B2(n6280), .ZN(n5623)
         );
  INV_X1 U6785 ( .A(n5621), .ZN(n5622) );
  NOR3_X1 U6786 ( .A1(n5624), .A2(n5623), .A3(n5622), .ZN(n5625) );
  OAI211_X1 U6787 ( .C1(n6286), .C2(n5861), .A(n5626), .B(n5625), .ZN(U2798)
         );
  INV_X1 U6788 ( .A(n5627), .ZN(n5632) );
  INV_X1 U6789 ( .A(n5629), .ZN(n5631) );
  AOI21_X1 U6790 ( .B1(n5632), .B2(n5631), .A(n5630), .ZN(n6087) );
  INV_X1 U6791 ( .A(n6087), .ZN(n5723) );
  INV_X1 U6792 ( .A(n6011), .ZN(n5634) );
  OAI211_X1 U6793 ( .C1(REIP_REG_24__SCAN_IN), .C2(REIP_REG_25__SCAN_IN), .A(
        n5634), .B(n5633), .ZN(n5635) );
  INV_X1 U6794 ( .A(n5635), .ZN(n5641) );
  INV_X1 U6795 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6860) );
  OAI22_X1 U6796 ( .A1(n6023), .A2(n6860), .B1(n6090), .B2(n6280), .ZN(n5640)
         );
  NAND2_X1 U6797 ( .A1(n5663), .A2(n5636), .ZN(n5637) );
  NAND2_X1 U6798 ( .A1(n3158), .A2(n5637), .ZN(n6112) );
  AOI22_X1 U6799 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6282), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6230), .ZN(n5638) );
  OAI21_X1 U6800 ( .B1(n6112), .B2(n6286), .A(n5638), .ZN(n5639) );
  NOR3_X1 U6801 ( .A1(n5641), .A2(n5640), .A3(n5639), .ZN(n5642) );
  OAI21_X1 U6802 ( .B1(n5723), .B2(n6192), .A(n5642), .ZN(U2802) );
  OAI22_X1 U6803 ( .A1(n5839), .A2(n6293), .B1(n6297), .B2(n5643), .ZN(U2828)
         );
  INV_X1 U6804 ( .A(n5744), .ZN(n5715) );
  OAI22_X1 U6805 ( .A1(n5861), .A2(n6293), .B1(n5644), .B2(n6297), .ZN(n5645)
         );
  INV_X1 U6806 ( .A(n5645), .ZN(n5646) );
  OAI21_X1 U6807 ( .B1(n5715), .B2(n5709), .A(n5646), .ZN(U2830) );
  AOI21_X1 U6808 ( .B1(n5648), .B2(n5647), .A(n5570), .ZN(n5996) );
  INV_X1 U6809 ( .A(n5996), .ZN(n5718) );
  INV_X1 U6810 ( .A(n5655), .ZN(n5650) );
  AOI21_X1 U6811 ( .B1(n5651), .B2(n5650), .A(n5649), .ZN(n5995) );
  AOI22_X1 U6812 ( .A1(n5995), .A2(n6065), .B1(EBX_REG_27__SCAN_IN), .B2(n4506), .ZN(n5652) );
  OAI21_X1 U6813 ( .B1(n5718), .B2(n5709), .A(n5652), .ZN(U2832) );
  AND2_X1 U6814 ( .A1(n3158), .A2(n5654), .ZN(n5656) );
  OR2_X1 U6815 ( .A1(n5656), .A2(n5655), .ZN(n6001) );
  INV_X1 U6816 ( .A(n6001), .ZN(n5887) );
  AOI22_X1 U6817 ( .A1(n5887), .A2(n6065), .B1(EBX_REG_26__SCAN_IN), .B2(n4506), .ZN(n5657) );
  OAI21_X1 U6818 ( .B1(n6002), .B2(n5709), .A(n5657), .ZN(U2833) );
  INV_X1 U6819 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5658) );
  OAI222_X1 U6820 ( .A1(n5723), .A2(n5709), .B1(n5658), .B2(n6297), .C1(n6293), 
        .C2(n6112), .ZN(U2834) );
  AOI21_X1 U6821 ( .B1(n5659), .B2(n3164), .A(n5629), .ZN(n5767) );
  INV_X1 U6822 ( .A(n5767), .ZN(n6012) );
  INV_X1 U6823 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5664) );
  OR2_X1 U6824 ( .A1(n5661), .A2(n5660), .ZN(n5662) );
  NAND2_X1 U6825 ( .A1(n5663), .A2(n5662), .ZN(n6016) );
  OAI222_X1 U6826 ( .A1(n5709), .A2(n6012), .B1(n6297), .B2(n5664), .C1(n6016), 
        .C2(n6293), .ZN(U2835) );
  NAND2_X1 U6827 ( .A1(n5666), .A2(n5665), .ZN(n5667) );
  AND2_X1 U6828 ( .A1(n5668), .A2(n5667), .ZN(n5906) );
  INV_X1 U6829 ( .A(n5906), .ZN(n6025) );
  INV_X1 U6830 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5672) );
  NAND2_X1 U6831 ( .A1(n5676), .A2(n5670), .ZN(n5671) );
  NAND2_X1 U6832 ( .A1(n4419), .A2(n5671), .ZN(n6073) );
  OAI222_X1 U6833 ( .A1(n6293), .A2(n6025), .B1(n6297), .B2(n5672), .C1(n6073), 
        .C2(n5709), .ZN(U2837) );
  OR2_X1 U6834 ( .A1(n5674), .A2(n5673), .ZN(n5675) );
  NAND2_X1 U6835 ( .A1(n5676), .A2(n5675), .ZN(n6078) );
  INV_X1 U6836 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5679) );
  XNOR2_X1 U6837 ( .A(n5678), .B(n5677), .ZN(n6040) );
  OAI222_X1 U6838 ( .A1(n6078), .A2(n5709), .B1(n5679), .B2(n6297), .C1(n6293), 
        .C2(n6040), .ZN(U2838) );
  INV_X1 U6839 ( .A(n5682), .ZN(n5683) );
  XNOR2_X1 U6840 ( .A(n5681), .B(n5683), .ZN(n6082) );
  INV_X1 U6841 ( .A(n6082), .ZN(n5689) );
  MUX2_X1 U6842 ( .A(n5685), .B(n5691), .S(n5684), .Z(n5687) );
  XNOR2_X1 U6843 ( .A(n5687), .B(n5686), .ZN(n6041) );
  AOI22_X1 U6844 ( .A1(n6041), .A2(n6065), .B1(EBX_REG_20__SCAN_IN), .B2(n4506), .ZN(n5688) );
  OAI21_X1 U6845 ( .B1(n5689), .B2(n5709), .A(n5688), .ZN(U2839) );
  MUX2_X1 U6846 ( .A(n5691), .B(n5690), .S(n3833), .Z(n5692) );
  INV_X1 U6847 ( .A(n5692), .ZN(n5693) );
  NAND2_X1 U6848 ( .A1(n6133), .A2(n5693), .ZN(n6059) );
  OR2_X1 U6849 ( .A1(n6133), .A2(n5693), .ZN(n5694) );
  NAND2_X1 U6850 ( .A1(n6059), .A2(n5694), .ZN(n6186) );
  OAI21_X1 U6851 ( .B1(n5696), .B2(n5698), .A(n5697), .ZN(n6182) );
  OAI222_X1 U6852 ( .A1(n6186), .A2(n6293), .B1(n6297), .B2(n3842), .C1(n6182), 
        .C2(n5709), .ZN(U2841) );
  NAND2_X1 U6853 ( .A1(n5700), .A2(n5699), .ZN(n5701) );
  NAND2_X1 U6854 ( .A1(n6132), .A2(n5701), .ZN(n6206) );
  INV_X1 U6855 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5706) );
  INV_X1 U6856 ( .A(n5702), .ZN(n5703) );
  AOI21_X1 U6857 ( .B1(n5704), .B2(n5552), .A(n5703), .ZN(n6309) );
  INV_X1 U6858 ( .A(n6309), .ZN(n5705) );
  OAI222_X1 U6859 ( .A1(n6206), .A2(n6293), .B1(n6297), .B2(n5706), .C1(n5705), 
        .C2(n5709), .ZN(U2843) );
  OAI222_X1 U6860 ( .A1(n5811), .A2(n5709), .B1(n5708), .B2(n6297), .C1(n6293), 
        .C2(n5707), .ZN(U2844) );
  AOI22_X1 U6861 ( .A1(n6307), .A2(DATAI_30_), .B1(n6311), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U6862 ( .A1(n6310), .A2(DATAI_14_), .ZN(n5710) );
  OAI211_X1 U6863 ( .C1(n5712), .C2(n6316), .A(n5711), .B(n5710), .ZN(U2861)
         );
  AOI22_X1 U6864 ( .A1(n6307), .A2(DATAI_29_), .B1(n6311), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U6865 ( .A1(n6310), .A2(DATAI_13_), .ZN(n5713) );
  OAI211_X1 U6866 ( .C1(n5715), .C2(n6316), .A(n5714), .B(n5713), .ZN(U2862)
         );
  AOI22_X1 U6867 ( .A1(n6307), .A2(DATAI_27_), .B1(n6311), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5717) );
  NAND2_X1 U6868 ( .A1(n6310), .A2(DATAI_11_), .ZN(n5716) );
  OAI211_X1 U6869 ( .C1(n5718), .C2(n6316), .A(n5717), .B(n5716), .ZN(U2864)
         );
  AOI22_X1 U6870 ( .A1(n6307), .A2(DATAI_26_), .B1(n6311), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U6871 ( .A1(n6310), .A2(DATAI_10_), .ZN(n5719) );
  OAI211_X1 U6872 ( .C1(n6002), .C2(n6316), .A(n5720), .B(n5719), .ZN(U2865)
         );
  AOI22_X1 U6873 ( .A1(n6307), .A2(DATAI_25_), .B1(n6311), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5722) );
  NAND2_X1 U6874 ( .A1(n6310), .A2(DATAI_9_), .ZN(n5721) );
  OAI211_X1 U6875 ( .C1(n5723), .C2(n6316), .A(n5722), .B(n5721), .ZN(U2866)
         );
  AOI22_X1 U6876 ( .A1(n6307), .A2(DATAI_24_), .B1(n6311), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U6877 ( .A1(n6310), .A2(DATAI_8_), .ZN(n5724) );
  OAI211_X1 U6878 ( .C1(n6012), .C2(n6316), .A(n5725), .B(n5724), .ZN(U2867)
         );
  INV_X1 U6879 ( .A(n5738), .ZN(n5729) );
  AND2_X1 U6880 ( .A1(n5727), .A2(n5726), .ZN(n5728) );
  XNOR2_X1 U6881 ( .A(n5730), .B(n5845), .ZN(n5854) );
  NAND2_X1 U6882 ( .A1(n5808), .A2(n5731), .ZN(n5732) );
  NAND2_X1 U6883 ( .A1(n6457), .A2(REIP_REG_30__SCAN_IN), .ZN(n5848) );
  OAI211_X1 U6884 ( .C1(n5733), .C2(n6111), .A(n5732), .B(n5848), .ZN(n5734)
         );
  AOI21_X1 U6885 ( .B1(n5735), .B2(n6378), .A(n5734), .ZN(n5736) );
  OAI21_X1 U6886 ( .B1(n5854), .B2(n6164), .A(n5736), .ZN(U2956) );
  OAI21_X1 U6887 ( .B1(n5737), .B2(n5739), .A(n5738), .ZN(n5740) );
  XNOR2_X1 U6888 ( .A(n5740), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5864)
         );
  NAND2_X1 U6889 ( .A1(n6457), .A2(REIP_REG_29__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U6890 ( .A1(n6374), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5741)
         );
  OAI211_X1 U6891 ( .C1(n6384), .C2(n5742), .A(n5857), .B(n5741), .ZN(n5743)
         );
  AOI21_X1 U6892 ( .B1(n5744), .B2(n6378), .A(n5743), .ZN(n5745) );
  OAI21_X1 U6893 ( .B1(n5864), .B2(n6164), .A(n5745), .ZN(U2957) );
  INV_X1 U6894 ( .A(n5747), .ZN(n5748) );
  NOR2_X1 U6895 ( .A1(n5746), .A2(n5748), .ZN(n5750) );
  XNOR2_X1 U6896 ( .A(n5750), .B(n5749), .ZN(n5880) );
  NAND2_X1 U6897 ( .A1(n6457), .A2(REIP_REG_27__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U6898 ( .A1(n6374), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5751)
         );
  OAI211_X1 U6899 ( .C1(n6384), .C2(n5993), .A(n5875), .B(n5751), .ZN(n5752)
         );
  AOI21_X1 U6900 ( .B1(n5996), .B2(n6378), .A(n5752), .ZN(n5753) );
  OAI21_X1 U6901 ( .B1(n5880), .B2(n6164), .A(n5753), .ZN(U2959) );
  NAND2_X1 U6902 ( .A1(n5755), .A2(n5754), .ZN(n5756) );
  XNOR2_X1 U6903 ( .A(n5737), .B(n5756), .ZN(n5889) );
  INV_X1 U6904 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U6905 ( .A1(n6457), .A2(REIP_REG_26__SCAN_IN), .ZN(n5884) );
  OAI21_X1 U6906 ( .B1(n6111), .B2(n5757), .A(n5884), .ZN(n5759) );
  NOR2_X1 U6907 ( .A1(n6002), .A2(n6108), .ZN(n5758) );
  AOI211_X1 U6908 ( .C1(n5808), .C2(n6000), .A(n5759), .B(n5758), .ZN(n5760)
         );
  OAI21_X1 U6909 ( .B1(n5889), .B2(n6164), .A(n5760), .ZN(U2960) );
  NAND3_X1 U6910 ( .A1(n3658), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5761) );
  XNOR2_X1 U6911 ( .A(n5763), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5898)
         );
  INV_X1 U6912 ( .A(n6009), .ZN(n5765) );
  AND2_X1 U6913 ( .A1(n6457), .A2(REIP_REG_24__SCAN_IN), .ZN(n5895) );
  AOI21_X1 U6914 ( .B1(n6374), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5895), 
        .ZN(n5764) );
  OAI21_X1 U6915 ( .B1(n5765), .B2(n6384), .A(n5764), .ZN(n5766) );
  AOI21_X1 U6916 ( .B1(n5767), .B2(n6378), .A(n5766), .ZN(n5768) );
  OAI21_X1 U6917 ( .B1(n5898), .B2(n6164), .A(n5768), .ZN(U2962) );
  AOI21_X1 U6918 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n3155), .A(n5769), 
        .ZN(n5770) );
  XNOR2_X1 U6919 ( .A(n5771), .B(n5770), .ZN(n5908) );
  NAND2_X1 U6920 ( .A1(n6457), .A2(REIP_REG_22__SCAN_IN), .ZN(n5903) );
  OAI21_X1 U6921 ( .B1(n6111), .B2(n5772), .A(n5903), .ZN(n5774) );
  NOR2_X1 U6922 ( .A1(n6073), .A2(n6108), .ZN(n5773) );
  AOI211_X1 U6923 ( .C1(n5808), .C2(n6024), .A(n5774), .B(n5773), .ZN(n5775)
         );
  OAI21_X1 U6924 ( .B1(n5908), .B2(n6164), .A(n5775), .ZN(U2964) );
  OAI21_X1 U6925 ( .B1(n5778), .B2(n5777), .A(n5776), .ZN(n5909) );
  NAND2_X1 U6926 ( .A1(n5909), .A2(n6380), .ZN(n5782) );
  INV_X1 U6927 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5779) );
  NOR2_X1 U6928 ( .A1(n6403), .A2(n5779), .ZN(n5912) );
  NOR2_X1 U6929 ( .A1(n6384), .A2(n6034), .ZN(n5780) );
  AOI211_X1 U6930 ( .C1(n6374), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5912), 
        .B(n5780), .ZN(n5781) );
  OAI211_X1 U6931 ( .C1(n6108), .C2(n6078), .A(n5782), .B(n5781), .ZN(U2965)
         );
  XNOR2_X1 U6932 ( .A(n5783), .B(n5784), .ZN(n5931) );
  INV_X1 U6933 ( .A(n6044), .ZN(n5786) );
  NAND2_X1 U6934 ( .A1(n6374), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5785)
         );
  NAND2_X1 U6935 ( .A1(n6457), .A2(REIP_REG_20__SCAN_IN), .ZN(n5917) );
  OAI211_X1 U6936 ( .C1(n6384), .C2(n5786), .A(n5785), .B(n5917), .ZN(n5787)
         );
  AOI21_X1 U6937 ( .B1(n6082), .B2(n6378), .A(n5787), .ZN(n5788) );
  OAI21_X1 U6938 ( .B1(n5931), .B2(n6164), .A(n5788), .ZN(U2966) );
  INV_X1 U6939 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U6940 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n3658), .ZN(n5791) );
  NAND4_X1 U6941 ( .A1(n6100), .A2(n6099), .A3(n6129), .A4(n5789), .ZN(n5790)
         );
  OAI21_X1 U6942 ( .B1(n5791), .B2(n3165), .A(n5790), .ZN(n5792) );
  XNOR2_X1 U6943 ( .A(n5933), .B(n5792), .ZN(n5934) );
  AOI22_X1 U6944 ( .A1(n6380), .A2(n5934), .B1(n6457), .B2(
        REIP_REG_18__SCAN_IN), .ZN(n5793) );
  OAI21_X1 U6945 ( .B1(n5794), .B2(n6111), .A(n5793), .ZN(n5795) );
  AOI21_X1 U6946 ( .B1(n5808), .B2(n6183), .A(n5795), .ZN(n5796) );
  OAI21_X1 U6947 ( .B1(n6182), .B2(n6108), .A(n5796), .ZN(U2968) );
  INV_X1 U6948 ( .A(n5797), .ZN(n5800) );
  OAI21_X1 U6949 ( .B1(n5798), .B2(n5800), .A(n5789), .ZN(n5799) );
  OAI21_X1 U6950 ( .B1(n3165), .B2(n5800), .A(n5799), .ZN(n5946) );
  NAND2_X1 U6951 ( .A1(n6457), .A2(REIP_REG_16__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U6952 ( .A1(n6374), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5801)
         );
  OAI211_X1 U6953 ( .C1(n6384), .C2(n6202), .A(n5940), .B(n5801), .ZN(n5802)
         );
  AOI21_X1 U6954 ( .B1(n6309), .B2(n6378), .A(n5802), .ZN(n5803) );
  OAI21_X1 U6955 ( .B1(n5946), .B2(n6164), .A(n5803), .ZN(U2970) );
  XNOR2_X1 U6956 ( .A(n3155), .B(n5942), .ZN(n5805) );
  XNOR2_X1 U6957 ( .A(n5804), .B(n5805), .ZN(n6144) );
  NAND2_X1 U6958 ( .A1(n6144), .A2(n6380), .ZN(n5810) );
  NAND2_X1 U6959 ( .A1(n6457), .A2(REIP_REG_15__SCAN_IN), .ZN(n6140) );
  OAI21_X1 U6960 ( .B1(n6111), .B2(n4097), .A(n6140), .ZN(n5806) );
  AOI21_X1 U6961 ( .B1(n5808), .B2(n5807), .A(n5806), .ZN(n5809) );
  OAI211_X1 U6962 ( .C1(n6108), .C2(n5811), .A(n5810), .B(n5809), .ZN(U2971)
         );
  XNOR2_X1 U6963 ( .A(n3155), .B(n5813), .ZN(n5814) );
  XNOR2_X1 U6964 ( .A(n5812), .B(n5814), .ZN(n5963) );
  NAND2_X1 U6965 ( .A1(n6457), .A2(REIP_REG_14__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U6966 ( .A1(n6374), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5815)
         );
  OAI211_X1 U6967 ( .C1(n6384), .C2(n6212), .A(n5958), .B(n5815), .ZN(n5816)
         );
  AOI21_X1 U6968 ( .B1(n6214), .B2(n6378), .A(n5816), .ZN(n5817) );
  OAI21_X1 U6969 ( .B1(n5963), .B2(n6164), .A(n5817), .ZN(U2972) );
  XNOR2_X1 U6970 ( .A(n5818), .B(n5819), .ZN(n6152) );
  NAND2_X1 U6971 ( .A1(n6152), .A2(n6380), .ZN(n5823) );
  AND2_X1 U6972 ( .A1(n6457), .A2(REIP_REG_13__SCAN_IN), .ZN(n6149) );
  NOR2_X1 U6973 ( .A1(n6384), .A2(n5820), .ZN(n5821) );
  AOI211_X1 U6974 ( .C1(n6374), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6149), 
        .B(n5821), .ZN(n5822) );
  OAI211_X1 U6975 ( .C1(n6108), .C2(n5824), .A(n5823), .B(n5822), .ZN(U2973)
         );
  INV_X1 U6976 ( .A(n5835), .ZN(n5831) );
  NAND2_X1 U6977 ( .A1(n5922), .A2(n6453), .ZN(n5825) );
  NAND2_X1 U6978 ( .A1(n5825), .A2(n5833), .ZN(n5826) );
  NAND2_X1 U6979 ( .A1(n5827), .A2(n5826), .ZN(n6117) );
  NAND2_X1 U6980 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n5834), .ZN(n5828) );
  OAI21_X1 U6981 ( .B1(n5828), .B2(n6115), .A(n5847), .ZN(n5829) );
  INV_X1 U6982 ( .A(n5829), .ZN(n5830) );
  NOR2_X1 U6983 ( .A1(n6117), .A2(n5830), .ZN(n5846) );
  OAI21_X1 U6984 ( .B1(n5831), .B2(n5939), .A(n5846), .ZN(n5838) );
  INV_X1 U6985 ( .A(n5832), .ZN(n5837) );
  NOR2_X1 U6986 ( .A1(n5892), .A2(n5833), .ZN(n6116) );
  AND2_X1 U6987 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U6988 ( .A1(n6116), .A2(n5881), .ZN(n5877) );
  INV_X1 U6989 ( .A(n5834), .ZN(n5866) );
  NOR3_X1 U6990 ( .A1(n5856), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5835), 
        .ZN(n5836) );
  AOI211_X1 U6991 ( .C1(n5838), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5837), .B(n5836), .ZN(n5842) );
  INV_X1 U6992 ( .A(n5839), .ZN(n5840) );
  NAND2_X1 U6993 ( .A1(n5840), .A2(n6448), .ZN(n5841) );
  OAI211_X1 U6994 ( .C1(n5843), .C2(n6138), .A(n5842), .B(n5841), .ZN(U2987)
         );
  INV_X1 U6995 ( .A(n5844), .ZN(n5852) );
  NAND2_X1 U6996 ( .A1(n5845), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U6997 ( .A1(n5846), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5860) );
  OAI211_X1 U6998 ( .C1(n5847), .C2(n6117), .A(n5860), .B(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5849) );
  OAI211_X1 U6999 ( .C1(n5856), .C2(n5850), .A(n5849), .B(n5848), .ZN(n5851)
         );
  AOI21_X1 U7000 ( .B1(n5852), .B2(n6448), .A(n5851), .ZN(n5853) );
  OAI21_X1 U7001 ( .B1(n5854), .B2(n6138), .A(n5853), .ZN(U2988) );
  INV_X1 U7002 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U7003 ( .A1(n5856), .A2(n5855), .ZN(n5859) );
  INV_X1 U7004 ( .A(n5857), .ZN(n5858) );
  AOI21_X1 U7005 ( .B1(n5860), .B2(n5859), .A(n5858), .ZN(n5863) );
  OR2_X1 U7006 ( .A1(n5861), .A2(n6405), .ZN(n5862) );
  OAI211_X1 U7007 ( .C1(n5864), .C2(n6138), .A(n5863), .B(n5862), .ZN(U2989)
         );
  NAND2_X1 U7008 ( .A1(n5866), .A2(n5865), .ZN(n5869) );
  INV_X1 U7009 ( .A(n6117), .ZN(n5890) );
  OAI21_X1 U7010 ( .B1(n5939), .B2(n5881), .A(n5890), .ZN(n5874) );
  NAND2_X1 U7011 ( .A1(n5874), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5868) );
  OAI211_X1 U7012 ( .C1(n5877), .C2(n5869), .A(n5868), .B(n5867), .ZN(n5870)
         );
  AOI21_X1 U7013 ( .B1(n5871), .B2(n6448), .A(n5870), .ZN(n5872) );
  OAI21_X1 U7014 ( .B1(n5873), .B2(n6138), .A(n5872), .ZN(U2990) );
  NAND2_X1 U7015 ( .A1(n5874), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5876) );
  OAI211_X1 U7016 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5877), .A(n5876), .B(n5875), .ZN(n5878) );
  AOI21_X1 U7017 ( .B1(n5995), .B2(n6448), .A(n5878), .ZN(n5879) );
  OAI21_X1 U7018 ( .B1(n5880), .B2(n6138), .A(n5879), .ZN(U2991) );
  AOI21_X1 U7019 ( .B1(n5885), .B2(n6115), .A(n5881), .ZN(n5882) );
  NAND2_X1 U7020 ( .A1(n6116), .A2(n5882), .ZN(n5883) );
  OAI211_X1 U7021 ( .C1(n5890), .C2(n5885), .A(n5884), .B(n5883), .ZN(n5886)
         );
  AOI21_X1 U7022 ( .B1(n5887), .B2(n6448), .A(n5886), .ZN(n5888) );
  OAI21_X1 U7023 ( .B1(n5889), .B2(n6138), .A(n5888), .ZN(U2992) );
  INV_X1 U7024 ( .A(n6016), .ZN(n5896) );
  INV_X1 U7025 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5893) );
  AOI211_X1 U7026 ( .C1(n5893), .C2(n5892), .A(n5891), .B(n5890), .ZN(n5894)
         );
  AOI211_X1 U7027 ( .C1(n5896), .C2(n6448), .A(n5895), .B(n5894), .ZN(n5897)
         );
  OAI21_X1 U7028 ( .B1(n5898), .B2(n6138), .A(n5897), .ZN(U2994) );
  INV_X1 U7029 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5904) );
  INV_X1 U7030 ( .A(n5899), .ZN(n5900) );
  NAND3_X1 U7031 ( .A1(n5914), .A2(n5901), .A3(n5900), .ZN(n5902) );
  OAI211_X1 U7032 ( .C1(n5910), .C2(n5904), .A(n5903), .B(n5902), .ZN(n5905)
         );
  AOI21_X1 U7033 ( .B1(n5906), .B2(n6448), .A(n5905), .ZN(n5907) );
  OAI21_X1 U7034 ( .B1(n5908), .B2(n6138), .A(n5907), .ZN(U2996) );
  NAND2_X1 U7035 ( .A1(n5909), .A2(n6454), .ZN(n5916) );
  NOR2_X1 U7036 ( .A1(n5910), .A2(n5913), .ZN(n5911) );
  AOI211_X1 U7037 ( .C1(n5914), .C2(n5913), .A(n5912), .B(n5911), .ZN(n5915)
         );
  OAI211_X1 U7038 ( .C1(n6405), .C2(n6040), .A(n5916), .B(n5915), .ZN(U2997)
         );
  INV_X1 U7039 ( .A(n5917), .ZN(n5921) );
  NOR3_X1 U7040 ( .A1(n6125), .A2(n5919), .A3(n5918), .ZN(n5920) );
  AOI211_X1 U7041 ( .C1(n6041), .C2(n6448), .A(n5921), .B(n5920), .ZN(n5930)
         );
  INV_X1 U7042 ( .A(n5922), .ZN(n6458) );
  AOI221_X1 U7043 ( .B1(n5926), .B2(n5925), .C1(n5924), .C2(n5925), .A(n5923), 
        .ZN(n5927) );
  OAI221_X1 U7044 ( .B1(n6453), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .C1(
        n6453), .C2(n5928), .A(n5927), .ZN(n6128) );
  AOI21_X1 U7045 ( .B1(n6458), .B2(n6129), .A(n6128), .ZN(n5932) );
  OAI21_X1 U7046 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5939), .A(n5932), 
        .ZN(n6120) );
  NAND2_X1 U7047 ( .A1(n6120), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5929) );
  OAI211_X1 U7048 ( .C1(n5931), .C2(n6138), .A(n5930), .B(n5929), .ZN(U2998)
         );
  OAI22_X1 U7049 ( .A1(n5932), .A2(n5933), .B1(n6403), .B2(n7045), .ZN(n5938)
         );
  NAND3_X1 U7050 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6130), .A3(n5933), .ZN(n5936) );
  NAND2_X1 U7051 ( .A1(n6454), .A2(n5934), .ZN(n5935) );
  OAI211_X1 U7052 ( .C1(n6186), .C2(n6405), .A(n5936), .B(n5935), .ZN(n5937)
         );
  OR2_X1 U7053 ( .A1(n5938), .A2(n5937), .ZN(U3000) );
  OAI21_X1 U7054 ( .B1(n5941), .B2(n5939), .A(n6391), .ZN(n6143) );
  OAI21_X1 U7055 ( .B1(n6206), .B2(n6405), .A(n5940), .ZN(n5944) );
  NAND2_X1 U7056 ( .A1(n5941), .A2(n6387), .ZN(n6147) );
  AOI221_X1 U7057 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n5942), .C2(n6099), .A(n6147), 
        .ZN(n5943) );
  AOI211_X1 U7058 ( .C1(INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n6143), .A(n5944), .B(n5943), .ZN(n5945) );
  OAI21_X1 U7059 ( .B1(n5946), .B2(n6138), .A(n5945), .ZN(U3002) );
  NOR3_X1 U7060 ( .A1(n6156), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n5949), 
        .ZN(n5961) );
  INV_X1 U7061 ( .A(n5947), .ZN(n5950) );
  NAND2_X1 U7062 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5953) );
  AOI22_X1 U7063 ( .A1(n5950), .A2(n5949), .B1(n5953), .B2(n5948), .ZN(n5951)
         );
  NAND2_X1 U7064 ( .A1(n6391), .A2(n5951), .ZN(n6151) );
  INV_X1 U7065 ( .A(n6151), .ZN(n5957) );
  INV_X1 U7066 ( .A(n5952), .ZN(n5954) );
  NOR2_X1 U7067 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5953), .ZN(n6148)
         );
  OAI21_X1 U7068 ( .B1(n5955), .B2(n5954), .A(n6148), .ZN(n5956) );
  AOI21_X1 U7069 ( .B1(n5957), .B2(n5956), .A(n5813), .ZN(n5960) );
  OAI21_X1 U7070 ( .B1(n6217), .B2(n6405), .A(n5958), .ZN(n5959) );
  NOR3_X1 U7071 ( .A1(n5961), .A2(n5960), .A3(n5959), .ZN(n5962) );
  OAI21_X1 U7072 ( .B1(n5963), .B2(n6138), .A(n5962), .ZN(U3004) );
  OAI211_X1 U7073 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n5964), .A(n6538), .B(
        n6537), .ZN(n5965) );
  OAI21_X1 U7074 ( .B1(n5974), .B2(n4537), .A(n5965), .ZN(n5966) );
  MUX2_X1 U7075 ( .A(n5966), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(n6463), 
        .Z(U3464) );
  XNOR2_X1 U7076 ( .A(n4776), .B(n6538), .ZN(n5967) );
  OAI22_X1 U7077 ( .A1(n5967), .A2(n6543), .B1(n4591), .B2(n5974), .ZN(n5968)
         );
  MUX2_X1 U7078 ( .A(n5968), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(n6463), 
        .Z(U3463) );
  NOR2_X1 U7079 ( .A1(n5970), .A2(n5969), .ZN(n5971) );
  OAI222_X1 U7080 ( .A1(n5974), .A2(n5973), .B1(n6471), .B2(n5972), .C1(n6543), 
        .C2(n5971), .ZN(n5975) );
  MUX2_X1 U7081 ( .A(n5975), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(n6463), 
        .Z(U3462) );
  INV_X1 U7082 ( .A(n5976), .ZN(n5978) );
  OAI22_X1 U7083 ( .A1(n5978), .A2(n6732), .B1(n5977), .B2(n6724), .ZN(n5979)
         );
  MUX2_X1 U7084 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5979), .S(n6727), 
        .Z(U3456) );
  AND2_X1 U7085 ( .A1(n6337), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI21_X1 U7086 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n5981), .A(n5980), .ZN(
        n5982) );
  INV_X1 U7087 ( .A(n5982), .ZN(U2788) );
  AOI22_X1 U7088 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n6230), .B1(n5983), 
        .B2(n6267), .ZN(n5991) );
  OAI22_X1 U7089 ( .A1(n5576), .A2(n6192), .B1(n5984), .B2(n6286), .ZN(n5989)
         );
  NOR3_X1 U7090 ( .A1(REIP_REG_28__SCAN_IN), .A2(n7051), .A3(n5999), .ZN(n5988) );
  OAI22_X1 U7091 ( .A1(n5986), .A2(n7067), .B1(n5985), .B2(n6054), .ZN(n5987)
         );
  NAND2_X1 U7092 ( .A1(n5991), .A2(n5990), .ZN(U2799) );
  AOI22_X1 U7093 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6282), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6230), .ZN(n5992) );
  OAI21_X1 U7094 ( .B1(n5993), .B2(n6280), .A(n5992), .ZN(n5994) );
  AOI21_X1 U7095 ( .B1(REIP_REG_27__SCAN_IN), .B2(n6005), .A(n5994), .ZN(n5998) );
  AOI22_X1 U7096 ( .A1(n5996), .A2(n6244), .B1(n5995), .B2(n6260), .ZN(n5997)
         );
  OAI211_X1 U7097 ( .C1(REIP_REG_27__SCAN_IN), .C2(n5999), .A(n5998), .B(n5997), .ZN(U2800) );
  AOI22_X1 U7098 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6230), .B1(n6000), 
        .B2(n6267), .ZN(n6007) );
  OAI22_X1 U7099 ( .A1(n6002), .A2(n6192), .B1(n6001), .B2(n6286), .ZN(n6003)
         );
  OAI211_X1 U7100 ( .C1(n6008), .C2(n6054), .A(n6007), .B(n6006), .ZN(U2801)
         );
  INV_X1 U7101 ( .A(REIP_REG_24__SCAN_IN), .ZN(n7019) );
  AOI22_X1 U7102 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n6230), .B1(n6009), 
        .B2(n6267), .ZN(n6010) );
  OAI21_X1 U7103 ( .B1(n6023), .B2(n7019), .A(n6010), .ZN(n6014) );
  OAI22_X1 U7104 ( .A1(n6012), .A2(n6192), .B1(REIP_REG_24__SCAN_IN), .B2(
        n6011), .ZN(n6013) );
  AOI211_X1 U7105 ( .C1(EBX_REG_24__SCAN_IN), .C2(n6282), .A(n6014), .B(n6013), 
        .ZN(n6015) );
  OAI21_X1 U7106 ( .B1(n6016), .B2(n6286), .A(n6015), .ZN(U2803) );
  INV_X1 U7107 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6705) );
  NOR2_X1 U7108 ( .A1(n6705), .A2(n5779), .ZN(n6027) );
  AOI21_X1 U7109 ( .B1(n6027), .B2(n6036), .A(REIP_REG_23__SCAN_IN), .ZN(n6022) );
  OAI22_X1 U7110 ( .A1(n6064), .A2(n6054), .B1(n6017), .B2(n6280), .ZN(n6018)
         );
  AOI21_X1 U7111 ( .B1(PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6230), .A(n6018), 
        .ZN(n6021) );
  INV_X1 U7112 ( .A(n6019), .ZN(n6069) );
  AOI22_X1 U7113 ( .A1(n6069), .A2(n6244), .B1(n6062), .B2(n6260), .ZN(n6020)
         );
  OAI211_X1 U7114 ( .C1(n6023), .C2(n6022), .A(n6021), .B(n6020), .ZN(U2804)
         );
  AOI22_X1 U7115 ( .A1(EBX_REG_22__SCAN_IN), .A2(n6282), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6230), .ZN(n6032) );
  AOI22_X1 U7116 ( .A1(n6024), .A2(n6267), .B1(REIP_REG_22__SCAN_IN), .B2(
        n6042), .ZN(n6031) );
  OAI22_X1 U7117 ( .A1(n6073), .A2(n6192), .B1(n6025), .B2(n6286), .ZN(n6026)
         );
  INV_X1 U7118 ( .A(n6026), .ZN(n6030) );
  INV_X1 U7119 ( .A(n6027), .ZN(n6028) );
  OAI211_X1 U7120 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n6036), .B(n6028), .ZN(n6029) );
  NAND4_X1 U7121 ( .A1(n6032), .A2(n6031), .A3(n6030), .A4(n6029), .ZN(U2805)
         );
  AOI22_X1 U7122 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6282), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6230), .ZN(n6033) );
  OAI21_X1 U7123 ( .B1(n6034), .B2(n6280), .A(n6033), .ZN(n6035) );
  AOI221_X1 U7124 ( .B1(n6042), .B2(REIP_REG_21__SCAN_IN), .C1(n6036), .C2(
        n5779), .A(n6035), .ZN(n6039) );
  INV_X1 U7125 ( .A(n6078), .ZN(n6037) );
  NAND2_X1 U7126 ( .A1(n6037), .A2(n6244), .ZN(n6038) );
  OAI211_X1 U7127 ( .C1(n6286), .C2(n6040), .A(n6039), .B(n6038), .ZN(U2806)
         );
  AOI22_X1 U7128 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6282), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6230), .ZN(n6048) );
  AOI22_X1 U7129 ( .A1(n6082), .A2(n6244), .B1(n6260), .B2(n6041), .ZN(n6047)
         );
  NOR2_X1 U7130 ( .A1(n6702), .A2(n7045), .ZN(n6051) );
  OAI221_X1 U7131 ( .B1(REIP_REG_20__SCAN_IN), .B2(n6051), .C1(
        REIP_REG_20__SCAN_IN), .C2(n6043), .A(n6042), .ZN(n6046) );
  NAND2_X1 U7132 ( .A1(n6044), .A2(n6267), .ZN(n6045) );
  NAND4_X1 U7133 ( .A1(n6048), .A2(n6047), .A3(n6046), .A4(n6045), .ZN(U2807)
         );
  NOR2_X1 U7134 ( .A1(n6050), .A2(n6049), .ZN(n6187) );
  AOI211_X1 U7135 ( .C1(n6702), .C2(n7045), .A(n6051), .B(n6180), .ZN(n6052)
         );
  AOI211_X1 U7136 ( .C1(n6230), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6052), 
        .B(n6265), .ZN(n6053) );
  OAI21_X1 U7137 ( .B1(n6068), .B2(n6054), .A(n6053), .ZN(n6055) );
  AOI21_X1 U7138 ( .B1(REIP_REG_19__SCAN_IN), .B2(n6187), .A(n6055), .ZN(n6061) );
  INV_X1 U7139 ( .A(n5681), .ZN(n6056) );
  AOI21_X1 U7140 ( .B1(n6057), .B2(n5697), .A(n6056), .ZN(n6095) );
  XNOR2_X1 U7141 ( .A(n6059), .B(n6058), .ZN(n6121) );
  AOI22_X1 U7142 ( .A1(n6095), .A2(n6244), .B1(n6260), .B2(n6121), .ZN(n6060)
         );
  OAI211_X1 U7143 ( .C1(n6098), .C2(n6280), .A(n6061), .B(n6060), .ZN(U2808)
         );
  AOI22_X1 U7144 ( .A1(n6069), .A2(n6066), .B1(n6062), .B2(n6065), .ZN(n6063)
         );
  OAI21_X1 U7145 ( .B1(n6297), .B2(n6064), .A(n6063), .ZN(U2836) );
  AOI22_X1 U7146 ( .A1(n6095), .A2(n6066), .B1(n6065), .B2(n6121), .ZN(n6067)
         );
  OAI21_X1 U7147 ( .B1(n6297), .B2(n6068), .A(n6067), .ZN(U2840) );
  INV_X1 U7148 ( .A(n6316), .ZN(n6308) );
  AOI22_X1 U7149 ( .A1(n6069), .A2(n6308), .B1(n6307), .B2(DATAI_23_), .ZN(
        n6071) );
  AOI22_X1 U7150 ( .A1(EAX_REG_23__SCAN_IN), .A2(n6311), .B1(n6310), .B2(
        DATAI_7_), .ZN(n6070) );
  NAND2_X1 U7151 ( .A1(n6071), .A2(n6070), .ZN(U2868) );
  INV_X1 U7152 ( .A(n6307), .ZN(n6302) );
  INV_X1 U7153 ( .A(DATAI_22_), .ZN(n6072) );
  OAI22_X1 U7154 ( .A1(n6073), .A2(n6316), .B1(n6302), .B2(n6072), .ZN(n6074)
         );
  INV_X1 U7155 ( .A(n6074), .ZN(n6076) );
  AOI22_X1 U7156 ( .A1(EAX_REG_22__SCAN_IN), .A2(n6311), .B1(n6310), .B2(
        DATAI_6_), .ZN(n6075) );
  NAND2_X1 U7157 ( .A1(n6076), .A2(n6075), .ZN(U2869) );
  INV_X1 U7158 ( .A(DATAI_21_), .ZN(n6077) );
  OAI22_X1 U7159 ( .A1(n6078), .A2(n6316), .B1(n6302), .B2(n6077), .ZN(n6079)
         );
  INV_X1 U7160 ( .A(n6079), .ZN(n6081) );
  AOI22_X1 U7161 ( .A1(EAX_REG_21__SCAN_IN), .A2(n6311), .B1(n6310), .B2(
        DATAI_5_), .ZN(n6080) );
  NAND2_X1 U7162 ( .A1(n6081), .A2(n6080), .ZN(U2870) );
  AOI22_X1 U7163 ( .A1(n6082), .A2(n6308), .B1(n6307), .B2(DATAI_20_), .ZN(
        n6084) );
  AOI22_X1 U7164 ( .A1(EAX_REG_20__SCAN_IN), .A2(n6311), .B1(n6310), .B2(
        DATAI_4_), .ZN(n6083) );
  NAND2_X1 U7165 ( .A1(n6084), .A2(n6083), .ZN(U2871) );
  AOI22_X1 U7166 ( .A1(n6095), .A2(n6308), .B1(n6307), .B2(DATAI_19_), .ZN(
        n6086) );
  AOI22_X1 U7167 ( .A1(EAX_REG_19__SCAN_IN), .A2(n6311), .B1(n6310), .B2(
        DATAI_3_), .ZN(n6085) );
  NAND2_X1 U7168 ( .A1(n6086), .A2(n6085), .ZN(U2872) );
  AOI22_X1 U7169 ( .A1(n6457), .A2(REIP_REG_25__SCAN_IN), .B1(n6374), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6089) );
  OAI21_X1 U7170 ( .B1(n3899), .B2(n3239), .A(n3901), .ZN(n6114) );
  AOI22_X1 U7171 ( .A1(n6087), .A2(n6378), .B1(n6380), .B2(n6114), .ZN(n6088)
         );
  OAI211_X1 U7172 ( .C1(n6384), .C2(n6090), .A(n6089), .B(n6088), .ZN(U2961)
         );
  AOI22_X1 U7173 ( .A1(n6457), .A2(REIP_REG_19__SCAN_IN), .B1(n6374), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6097) );
  OAI21_X1 U7174 ( .B1(n3671), .B2(n6093), .A(n6092), .ZN(n6094) );
  XNOR2_X1 U7175 ( .A(n6094), .B(n6100), .ZN(n6122) );
  AOI22_X1 U7176 ( .A1(n6122), .A2(n6380), .B1(n6378), .B2(n6095), .ZN(n6096)
         );
  OAI211_X1 U7177 ( .C1(n6384), .C2(n6098), .A(n6097), .B(n6096), .ZN(U2967)
         );
  INV_X1 U7178 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6190) );
  OR3_X1 U7179 ( .A1(n5789), .A2(n6100), .A3(n6099), .ZN(n6104) );
  NOR2_X1 U7180 ( .A1(n3155), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6102)
         );
  NAND2_X1 U7181 ( .A1(n5789), .A2(n6102), .ZN(n6103) );
  NAND2_X1 U7182 ( .A1(n6104), .A2(n6103), .ZN(n6105) );
  XNOR2_X1 U7183 ( .A(n6105), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6139)
         );
  AND2_X1 U7184 ( .A1(n5702), .A2(n6106), .ZN(n6107) );
  OR2_X1 U7185 ( .A1(n6107), .A2(n5696), .ZN(n6303) );
  OAI222_X1 U7186 ( .A1(n6384), .A2(n6196), .B1(n6164), .B2(n6139), .C1(n6108), 
        .C2(n6303), .ZN(n6109) );
  INV_X1 U7187 ( .A(n6109), .ZN(n6110) );
  NAND2_X1 U7188 ( .A1(n6457), .A2(REIP_REG_17__SCAN_IN), .ZN(n6126) );
  OAI211_X1 U7189 ( .C1(n6190), .C2(n6111), .A(n6110), .B(n6126), .ZN(U2969)
         );
  INV_X1 U7190 ( .A(n6112), .ZN(n6113) );
  AOI22_X1 U7191 ( .A1(n6114), .A2(n6454), .B1(n6448), .B2(n6113), .ZN(n6119)
         );
  AOI22_X1 U7192 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n6117), .B1(n6116), .B2(n6115), .ZN(n6118) );
  OAI211_X1 U7193 ( .C1(n6860), .C2(n6403), .A(n6119), .B(n6118), .ZN(U2993)
         );
  AOI22_X1 U7194 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n6120), .B1(n6457), .B2(REIP_REG_19__SCAN_IN), .ZN(n6124) );
  AOI22_X1 U7195 ( .A1(n6122), .A2(n6454), .B1(n6448), .B2(n6121), .ZN(n6123)
         );
  OAI211_X1 U7196 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n6125), .A(n6124), .B(n6123), .ZN(U2999) );
  INV_X1 U7197 ( .A(n6126), .ZN(n6127) );
  AOI221_X1 U7198 ( .B1(n6130), .B2(n6129), .C1(n6128), .C2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n6127), .ZN(n6137) );
  AND2_X1 U7199 ( .A1(n6132), .A2(n6131), .ZN(n6134) );
  OR2_X1 U7200 ( .A1(n6134), .A2(n6133), .ZN(n6292) );
  INV_X1 U7201 ( .A(n6292), .ZN(n6135) );
  NAND2_X1 U7202 ( .A1(n6135), .A2(n6448), .ZN(n6136) );
  OAI211_X1 U7203 ( .C1(n6139), .C2(n6138), .A(n6137), .B(n6136), .ZN(U3001)
         );
  INV_X1 U7204 ( .A(n6140), .ZN(n6141) );
  AOI21_X1 U7205 ( .B1(n6142), .B2(n6448), .A(n6141), .ZN(n6146) );
  AOI22_X1 U7206 ( .A1(n6144), .A2(n6454), .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n6143), .ZN(n6145) );
  OAI211_X1 U7207 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n6147), .A(n6146), .B(n6145), .ZN(U3003) );
  INV_X1 U7208 ( .A(n6148), .ZN(n6155) );
  AOI21_X1 U7209 ( .B1(n6150), .B2(n6448), .A(n6149), .ZN(n6154) );
  AOI22_X1 U7210 ( .A1(n6152), .A2(n6454), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n6151), .ZN(n6153) );
  OAI211_X1 U7211 ( .C1(n6156), .C2(n6155), .A(n6154), .B(n6153), .ZN(U3005)
         );
  INV_X1 U7212 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6157) );
  INV_X2 U7213 ( .A(n7142), .ZN(n6713) );
  INV_X1 U7214 ( .A(ADS_N_REG_SCAN_IN), .ZN(n7032) );
  AOI221_X4 U7215 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_0__SCAN_IN), .C1(
        n6157), .C2(STATE_REG_0__SCAN_IN), .A(n6713), .ZN(n6717) );
  INV_X1 U7216 ( .A(n6717), .ZN(n6715) );
  OAI21_X1 U7217 ( .B1(n6713), .B2(n7032), .A(n6715), .ZN(U2789) );
  INV_X1 U7218 ( .A(n6647), .ZN(n6746) );
  NAND2_X1 U7219 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6746), .ZN(n6160) );
  OAI21_X1 U7220 ( .B1(n6158), .B2(n6650), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6159) );
  OAI21_X1 U7221 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6160), .A(n6159), .ZN(
        U2790) );
  NOR2_X1 U7222 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6162) );
  OAI21_X1 U7223 ( .B1(n6162), .B2(D_C_N_REG_SCAN_IN), .A(n7142), .ZN(n6161)
         );
  OAI21_X1 U7224 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n7142), .A(n6161), .ZN(
        U2791) );
  OAI21_X1 U7225 ( .B1(BS16_N), .B2(n6162), .A(n6717), .ZN(n6716) );
  OAI21_X1 U7226 ( .B1(n6717), .B2(n6163), .A(n6716), .ZN(U2792) );
  OAI21_X1 U7227 ( .B1(n6165), .B2(n7094), .A(n6164), .ZN(U2793) );
  NOR4_X1 U7228 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(
        DATAWIDTH_REG_5__SCAN_IN), .ZN(n6169) );
  NOR4_X1 U7229 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_7__SCAN_IN), .ZN(n6168) );
  NOR4_X1 U7230 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6167) );
  NOR4_X1 U7231 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6166) );
  NAND4_X1 U7232 ( .A1(n6169), .A2(n6168), .A3(n6167), .A4(n6166), .ZN(n6175)
         );
  NOR4_X1 U7233 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(
        DATAWIDTH_REG_13__SCAN_IN), .ZN(n6173) );
  AOI211_X1 U7234 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_8__SCAN_IN), .B(
        DATAWIDTH_REG_11__SCAN_IN), .ZN(n6172) );
  NOR4_X1 U7235 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6171)
         );
  NOR4_X1 U7236 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n6170) );
  NAND4_X1 U7237 ( .A1(n6173), .A2(n6172), .A3(n6171), .A4(n6170), .ZN(n6174)
         );
  NOR2_X1 U7238 ( .A1(n6175), .A2(n6174), .ZN(n6739) );
  INV_X1 U7239 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6711) );
  NOR3_X1 U7240 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6177) );
  OAI21_X1 U7241 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6177), .A(n6739), .ZN(n6176)
         );
  OAI21_X1 U7242 ( .B1(n6739), .B2(n6711), .A(n6176), .ZN(U2794) );
  INV_X1 U7243 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6888) );
  AOI21_X1 U7244 ( .B1(n6733), .B2(n6888), .A(n6177), .ZN(n6178) );
  INV_X1 U7245 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6863) );
  INV_X1 U7246 ( .A(n6739), .ZN(n6735) );
  AOI22_X1 U7247 ( .A1(n6739), .A2(n6178), .B1(n6863), .B2(n6735), .ZN(U2795)
         );
  AOI22_X1 U7248 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6282), .B1(
        REIP_REG_18__SCAN_IN), .B2(n6187), .ZN(n6179) );
  OAI21_X1 U7249 ( .B1(REIP_REG_18__SCAN_IN), .B2(n6180), .A(n6179), .ZN(n6181) );
  AOI211_X1 U7250 ( .C1(n6230), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6265), 
        .B(n6181), .ZN(n6185) );
  INV_X1 U7251 ( .A(n6182), .ZN(n6298) );
  AOI22_X1 U7252 ( .A1(n6298), .A2(n6244), .B1(n6267), .B2(n6183), .ZN(n6184)
         );
  OAI211_X1 U7253 ( .C1(n6286), .C2(n6186), .A(n6185), .B(n6184), .ZN(U2809)
         );
  OAI21_X1 U7254 ( .B1(REIP_REG_17__SCAN_IN), .B2(n6188), .A(n6187), .ZN(n6189) );
  OAI21_X1 U7255 ( .B1(n6279), .B2(n6190), .A(n6189), .ZN(n6191) );
  AOI211_X1 U7256 ( .C1(n6282), .C2(EBX_REG_17__SCAN_IN), .A(n6265), .B(n6191), 
        .ZN(n6195) );
  OAI22_X1 U7257 ( .A1(n6303), .A2(n6192), .B1(n6286), .B2(n6292), .ZN(n6193)
         );
  INV_X1 U7258 ( .A(n6193), .ZN(n6194) );
  OAI211_X1 U7259 ( .C1(n6196), .C2(n6280), .A(n6195), .B(n6194), .ZN(U2810)
         );
  OAI21_X1 U7260 ( .B1(REIP_REG_16__SCAN_IN), .B2(REIP_REG_15__SCAN_IN), .A(
        n6197), .ZN(n6199) );
  AOI22_X1 U7261 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6282), .B1(
        REIP_REG_16__SCAN_IN), .B2(n6211), .ZN(n6198) );
  OAI21_X1 U7262 ( .B1(n6200), .B2(n6199), .A(n6198), .ZN(n6201) );
  AOI211_X1 U7263 ( .C1(n6230), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6265), 
        .B(n6201), .ZN(n6205) );
  INV_X1 U7264 ( .A(n6202), .ZN(n6203) );
  AOI22_X1 U7265 ( .A1(n6309), .A2(n6244), .B1(n6203), .B2(n6267), .ZN(n6204)
         );
  OAI211_X1 U7266 ( .C1(n6286), .C2(n6206), .A(n6205), .B(n6204), .ZN(U2811)
         );
  INV_X1 U7267 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6209) );
  AOI22_X1 U7268 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6282), .B1(n6207), .B2(n6697), .ZN(n6208) );
  OAI211_X1 U7269 ( .C1(n6279), .C2(n6209), .A(n6208), .B(n6249), .ZN(n6210)
         );
  AOI21_X1 U7270 ( .B1(REIP_REG_14__SCAN_IN), .B2(n6211), .A(n6210), .ZN(n6216) );
  INV_X1 U7271 ( .A(n6212), .ZN(n6213) );
  AOI22_X1 U7272 ( .A1(n6214), .A2(n6244), .B1(n6213), .B2(n6267), .ZN(n6215)
         );
  OAI211_X1 U7273 ( .C1(n6286), .C2(n6217), .A(n6216), .B(n6215), .ZN(U2813)
         );
  AOI22_X1 U7274 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n6230), .B1(n6260), 
        .B2(n6218), .ZN(n6226) );
  NOR2_X1 U7275 ( .A1(n6694), .A2(n6219), .ZN(n6220) );
  AOI211_X1 U7276 ( .C1(n6282), .C2(EBX_REG_12__SCAN_IN), .A(n6221), .B(n6220), 
        .ZN(n6225) );
  AOI22_X1 U7277 ( .A1(n6223), .A2(n6244), .B1(n6267), .B2(n6222), .ZN(n6224)
         );
  NAND4_X1 U7278 ( .A1(n6226), .A2(n6225), .A3(n6224), .A4(n6249), .ZN(U2815)
         );
  AOI22_X1 U7279 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6282), .B1(n6260), .B2(n6227), .ZN(n6238) );
  NOR3_X1 U7280 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6690), .A3(n6228), .ZN(n6229) );
  AOI211_X1 U7281 ( .C1(n6230), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6265), 
        .B(n6229), .ZN(n6237) );
  AOI22_X1 U7282 ( .A1(n6232), .A2(n6244), .B1(n6267), .B2(n6231), .ZN(n6236)
         );
  OAI21_X1 U7283 ( .B1(n6234), .B2(n6233), .A(REIP_REG_10__SCAN_IN), .ZN(n6235) );
  NAND4_X1 U7284 ( .A1(n6238), .A2(n6237), .A3(n6236), .A4(n6235), .ZN(U2817)
         );
  NOR3_X1 U7285 ( .A1(n6271), .A2(REIP_REG_7__SCAN_IN), .A3(n6239), .ZN(n6243)
         );
  INV_X1 U7286 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6241) );
  AOI22_X1 U7287 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6282), .B1(n6260), .B2(n6411), 
        .ZN(n6240) );
  OAI211_X1 U7288 ( .C1(n6279), .C2(n6241), .A(n6240), .B(n6249), .ZN(n6242)
         );
  AOI211_X1 U7289 ( .C1(n6354), .C2(n6244), .A(n6243), .B(n6242), .ZN(n6247)
         );
  OAI21_X1 U7290 ( .B1(n6245), .B2(n6255), .A(REIP_REG_7__SCAN_IN), .ZN(n6246)
         );
  OAI211_X1 U7291 ( .C1(n6280), .C2(n6357), .A(n6247), .B(n6246), .ZN(U2820)
         );
  INV_X1 U7292 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6251) );
  INV_X1 U7293 ( .A(n6248), .ZN(n6422) );
  AOI22_X1 U7294 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6282), .B1(n6260), .B2(n6422), 
        .ZN(n6250) );
  OAI211_X1 U7295 ( .C1(n6279), .C2(n6251), .A(n6250), .B(n6249), .ZN(n6252)
         );
  AOI21_X1 U7296 ( .B1(n6362), .B2(n6288), .A(n6252), .ZN(n6258) );
  AND2_X1 U7297 ( .A1(n6254), .A2(n6253), .ZN(n6256) );
  OAI21_X1 U7298 ( .B1(n6256), .B2(REIP_REG_5__SCAN_IN), .A(n6255), .ZN(n6257)
         );
  OAI211_X1 U7299 ( .C1(n6280), .C2(n6365), .A(n6258), .B(n6257), .ZN(U2822)
         );
  AOI22_X1 U7300 ( .A1(n6260), .A2(n6430), .B1(n6259), .B2(n6283), .ZN(n6275)
         );
  OAI21_X1 U7301 ( .B1(n6262), .B2(n6270), .A(n6261), .ZN(n6291) );
  OAI22_X1 U7302 ( .A1(n6291), .A2(n6684), .B1(n6263), .B2(n6279), .ZN(n6264)
         );
  AOI211_X1 U7303 ( .C1(n6282), .C2(EBX_REG_4__SCAN_IN), .A(n6265), .B(n6264), 
        .ZN(n6274) );
  INV_X1 U7304 ( .A(n6266), .ZN(n6269) );
  AOI22_X1 U7305 ( .A1(n6269), .A2(n6288), .B1(n6268), .B2(n6267), .ZN(n6273)
         );
  OR3_X1 U7306 ( .A1(n6271), .A2(REIP_REG_4__SCAN_IN), .A3(n6270), .ZN(n6272)
         );
  NAND4_X1 U7307 ( .A1(n6275), .A2(n6274), .A3(n6273), .A4(n6272), .ZN(U2823)
         );
  INV_X1 U7308 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6683) );
  INV_X1 U7309 ( .A(n6276), .ZN(n6277) );
  NAND2_X1 U7310 ( .A1(n6277), .A2(REIP_REG_2__SCAN_IN), .ZN(n6290) );
  INV_X1 U7311 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6278) );
  OAI22_X1 U7312 ( .A1(n6373), .A2(n6280), .B1(n6279), .B2(n6278), .ZN(n6281)
         );
  AOI21_X1 U7313 ( .B1(n6282), .B2(EBX_REG_3__SCAN_IN), .A(n6281), .ZN(n6285)
         );
  NAND2_X1 U7314 ( .A1(n6283), .A2(n4690), .ZN(n6284) );
  OAI211_X1 U7315 ( .C1(n6286), .C2(n6438), .A(n6285), .B(n6284), .ZN(n6287)
         );
  AOI21_X1 U7316 ( .B1(n6370), .B2(n6288), .A(n6287), .ZN(n6289) );
  OAI221_X1 U7317 ( .B1(n6291), .B2(n6683), .C1(n6291), .C2(n6290), .A(n6289), 
        .ZN(U2824) );
  OAI22_X1 U7318 ( .A1(n6303), .A2(n5709), .B1(n6293), .B2(n6292), .ZN(n6294)
         );
  INV_X1 U7319 ( .A(n6294), .ZN(n6295) );
  OAI21_X1 U7320 ( .B1(n6297), .B2(n6296), .A(n6295), .ZN(U2842) );
  AOI22_X1 U7321 ( .A1(n6298), .A2(n6308), .B1(n6307), .B2(DATAI_18_), .ZN(
        n6300) );
  AOI22_X1 U7322 ( .A1(EAX_REG_18__SCAN_IN), .A2(n6311), .B1(n6310), .B2(
        DATAI_2_), .ZN(n6299) );
  NAND2_X1 U7323 ( .A1(n6300), .A2(n6299), .ZN(U2873) );
  INV_X1 U7324 ( .A(DATAI_17_), .ZN(n6301) );
  OAI22_X1 U7325 ( .A1(n6303), .A2(n6316), .B1(n6302), .B2(n6301), .ZN(n6304)
         );
  INV_X1 U7326 ( .A(n6304), .ZN(n6306) );
  AOI22_X1 U7327 ( .A1(EAX_REG_17__SCAN_IN), .A2(n6311), .B1(n6310), .B2(
        DATAI_1_), .ZN(n6305) );
  NAND2_X1 U7328 ( .A1(n6306), .A2(n6305), .ZN(U2874) );
  AOI22_X1 U7329 ( .A1(n6309), .A2(n6308), .B1(n6307), .B2(DATAI_16_), .ZN(
        n6313) );
  AOI22_X1 U7330 ( .A1(EAX_REG_16__SCAN_IN), .A2(n6311), .B1(n6310), .B2(
        DATAI_0_), .ZN(n6312) );
  NAND2_X1 U7331 ( .A1(n6313), .A2(n6312), .ZN(U2875) );
  INV_X1 U7332 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6349) );
  OAI222_X1 U7333 ( .A1(n6317), .A2(n6316), .B1(n6847), .B2(n6315), .C1(n6349), 
        .C2(n6314), .ZN(U2891) );
  AOI22_X1 U7334 ( .A1(n6638), .A2(LWORD_REG_15__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6318) );
  OAI21_X1 U7335 ( .B1(n4517), .B2(n6348), .A(n6318), .ZN(U2908) );
  INV_X1 U7336 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6320) );
  AOI22_X1 U7337 ( .A1(n6638), .A2(LWORD_REG_14__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6319) );
  OAI21_X1 U7338 ( .B1(n6320), .B2(n6348), .A(n6319), .ZN(U2909) );
  AOI22_X1 U7339 ( .A1(n6638), .A2(LWORD_REG_13__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6321) );
  OAI21_X1 U7340 ( .B1(n6322), .B2(n6348), .A(n6321), .ZN(U2910) );
  AOI22_X1 U7341 ( .A1(n6638), .A2(LWORD_REG_12__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6323) );
  OAI21_X1 U7342 ( .B1(n6324), .B2(n6348), .A(n6323), .ZN(U2911) );
  AOI22_X1 U7343 ( .A1(n6638), .A2(LWORD_REG_11__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6325) );
  OAI21_X1 U7344 ( .B1(n6326), .B2(n6348), .A(n6325), .ZN(U2912) );
  AOI22_X1 U7345 ( .A1(n6638), .A2(LWORD_REG_10__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6327) );
  OAI21_X1 U7346 ( .B1(n6328), .B2(n6348), .A(n6327), .ZN(U2913) );
  AOI22_X1 U7347 ( .A1(n6638), .A2(LWORD_REG_9__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6329) );
  OAI21_X1 U7348 ( .B1(n6330), .B2(n6348), .A(n6329), .ZN(U2914) );
  AOI22_X1 U7349 ( .A1(n6638), .A2(LWORD_REG_8__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6331) );
  OAI21_X1 U7350 ( .B1(n6332), .B2(n6348), .A(n6331), .ZN(U2915) );
  AOI22_X1 U7351 ( .A1(n6638), .A2(LWORD_REG_7__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6333) );
  OAI21_X1 U7352 ( .B1(n6334), .B2(n6348), .A(n6333), .ZN(U2916) );
  AOI22_X1 U7353 ( .A1(n6638), .A2(LWORD_REG_6__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6335) );
  OAI21_X1 U7354 ( .B1(n3914), .B2(n6348), .A(n6335), .ZN(U2917) );
  AOI22_X1 U7355 ( .A1(n6638), .A2(LWORD_REG_5__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6336) );
  OAI21_X1 U7356 ( .B1(n3908), .B2(n6348), .A(n6336), .ZN(U2918) );
  AOI22_X1 U7357 ( .A1(n6638), .A2(LWORD_REG_4__SCAN_IN), .B1(n6337), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6338) );
  OAI21_X1 U7358 ( .B1(n6339), .B2(n6348), .A(n6338), .ZN(U2919) );
  AOI22_X1 U7359 ( .A1(n6638), .A2(LWORD_REG_3__SCAN_IN), .B1(n6346), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6340) );
  OAI21_X1 U7360 ( .B1(n6341), .B2(n6348), .A(n6340), .ZN(U2920) );
  AOI22_X1 U7361 ( .A1(n6638), .A2(LWORD_REG_2__SCAN_IN), .B1(n6346), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6342) );
  OAI21_X1 U7362 ( .B1(n6343), .B2(n6348), .A(n6342), .ZN(U2921) );
  AOI22_X1 U7363 ( .A1(n6638), .A2(LWORD_REG_1__SCAN_IN), .B1(n6346), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6344) );
  OAI21_X1 U7364 ( .B1(n6345), .B2(n6348), .A(n6344), .ZN(U2922) );
  AOI22_X1 U7365 ( .A1(n6638), .A2(LWORD_REG_0__SCAN_IN), .B1(n6346), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6347) );
  OAI21_X1 U7366 ( .B1(n6349), .B2(n6348), .A(n6347), .ZN(U2923) );
  AOI22_X1 U7367 ( .A1(n6457), .A2(REIP_REG_7__SCAN_IN), .B1(n6374), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6356) );
  OAI21_X1 U7368 ( .B1(n6352), .B2(n6351), .A(n6350), .ZN(n6353) );
  INV_X1 U7369 ( .A(n6353), .ZN(n6414) );
  AOI22_X1 U7370 ( .A1(n6414), .A2(n6380), .B1(n6378), .B2(n6354), .ZN(n6355)
         );
  OAI211_X1 U7371 ( .C1(n6384), .C2(n6357), .A(n6356), .B(n6355), .ZN(U2979)
         );
  AOI22_X1 U7372 ( .A1(n6457), .A2(REIP_REG_5__SCAN_IN), .B1(n6374), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6364) );
  OAI21_X1 U7373 ( .B1(n6360), .B2(n6359), .A(n6358), .ZN(n6361) );
  INV_X1 U7374 ( .A(n6361), .ZN(n6423) );
  AOI22_X1 U7375 ( .A1(n6423), .A2(n6380), .B1(n6378), .B2(n6362), .ZN(n6363)
         );
  OAI211_X1 U7376 ( .C1(n6384), .C2(n6365), .A(n6364), .B(n6363), .ZN(U2981)
         );
  AOI22_X1 U7377 ( .A1(n6457), .A2(REIP_REG_3__SCAN_IN), .B1(n6374), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6372) );
  OAI21_X1 U7378 ( .B1(n6368), .B2(n6367), .A(n6366), .ZN(n6369) );
  INV_X1 U7379 ( .A(n6369), .ZN(n6440) );
  AOI22_X1 U7380 ( .A1(n6370), .A2(n6378), .B1(n6440), .B2(n6380), .ZN(n6371)
         );
  OAI211_X1 U7381 ( .C1(n6384), .C2(n6373), .A(n6372), .B(n6371), .ZN(U2983)
         );
  AOI22_X1 U7382 ( .A1(n6457), .A2(REIP_REG_2__SCAN_IN), .B1(n6374), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6382) );
  XOR2_X1 U7383 ( .A(n6375), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n6377) );
  XNOR2_X1 U7384 ( .A(n6377), .B(n6376), .ZN(n6455) );
  AOI22_X1 U7385 ( .A1(n6455), .A2(n6380), .B1(n6379), .B2(n6378), .ZN(n6381)
         );
  OAI211_X1 U7386 ( .C1(n6384), .C2(n6383), .A(n6382), .B(n6381), .ZN(U2984)
         );
  AOI21_X1 U7387 ( .B1(n6386), .B2(n6448), .A(n6385), .ZN(n6390) );
  AOI22_X1 U7388 ( .A1(n6454), .A2(n6388), .B1(n5357), .B2(n6387), .ZN(n6389)
         );
  OAI211_X1 U7389 ( .C1(n6391), .C2(n5357), .A(n6390), .B(n6389), .ZN(U3007)
         );
  INV_X1 U7390 ( .A(n6392), .ZN(n6400) );
  AOI21_X1 U7391 ( .B1(n6394), .B2(n6448), .A(n6393), .ZN(n6398) );
  AOI22_X1 U7392 ( .A1(n6396), .A2(n6454), .B1(n6395), .B2(n6399), .ZN(n6397)
         );
  OAI211_X1 U7393 ( .C1(n6400), .C2(n6399), .A(n6398), .B(n6397), .ZN(U3009)
         );
  INV_X1 U7394 ( .A(n6401), .ZN(n6408) );
  AOI211_X1 U7395 ( .C1(n6418), .C2(n6410), .A(n6402), .B(n6412), .ZN(n6407)
         );
  OAI22_X1 U7396 ( .A1(n6405), .A2(n6404), .B1(n6689), .B2(n6403), .ZN(n6406)
         );
  AOI211_X1 U7397 ( .C1(n6408), .C2(n6454), .A(n6407), .B(n6406), .ZN(n6409)
         );
  OAI21_X1 U7398 ( .B1(n6410), .B2(n6417), .A(n6409), .ZN(U3010) );
  AOI22_X1 U7399 ( .A1(n6411), .A2(n6448), .B1(n6457), .B2(REIP_REG_7__SCAN_IN), .ZN(n6416) );
  INV_X1 U7400 ( .A(n6412), .ZN(n6413) );
  AOI22_X1 U7401 ( .A1(n6414), .A2(n6454), .B1(n6413), .B2(n6418), .ZN(n6415)
         );
  OAI211_X1 U7402 ( .C1(n6418), .C2(n6417), .A(n6416), .B(n6415), .ZN(U3011)
         );
  NOR2_X1 U7403 ( .A1(n6444), .A2(n6419), .ZN(n6437) );
  INV_X1 U7404 ( .A(n6420), .ZN(n6449) );
  NOR2_X1 U7405 ( .A1(n6449), .A2(n6421), .ZN(n6441) );
  AOI21_X1 U7406 ( .B1(n6437), .B2(n6441), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6426) );
  AOI22_X1 U7407 ( .A1(n6423), .A2(n6454), .B1(n6448), .B2(n6422), .ZN(n6425)
         );
  NAND2_X1 U7408 ( .A1(n6457), .A2(REIP_REG_5__SCAN_IN), .ZN(n6424) );
  OAI211_X1 U7409 ( .C1(n6427), .C2(n6426), .A(n6425), .B(n6424), .ZN(U3013)
         );
  OAI21_X1 U7410 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6441), .ZN(n6436) );
  INV_X1 U7411 ( .A(n6428), .ZN(n6429) );
  AOI21_X1 U7412 ( .B1(n6448), .B2(n6430), .A(n6429), .ZN(n6435) );
  INV_X1 U7413 ( .A(n6431), .ZN(n6433) );
  AOI22_X1 U7414 ( .A1(n6433), .A2(n6454), .B1(INSTADDRPOINTER_REG_4__SCAN_IN), 
        .B2(n6432), .ZN(n6434) );
  OAI211_X1 U7415 ( .C1(n6437), .C2(n6436), .A(n6435), .B(n6434), .ZN(U3014)
         );
  INV_X1 U7416 ( .A(n6438), .ZN(n6439) );
  AOI22_X1 U7417 ( .A1(n6448), .A2(n6439), .B1(n6457), .B2(REIP_REG_3__SCAN_IN), .ZN(n6443) );
  AOI22_X1 U7418 ( .A1(n6441), .A2(n6444), .B1(n6440), .B2(n6454), .ZN(n6442)
         );
  OAI211_X1 U7419 ( .C1(n6445), .C2(n6444), .A(n6443), .B(n6442), .ZN(U3015)
         );
  INV_X1 U7420 ( .A(n6446), .ZN(n6447) );
  AOI22_X1 U7421 ( .A1(n6450), .A2(n6449), .B1(n6448), .B2(n6447), .ZN(n6462)
         );
  OAI21_X1 U7422 ( .B1(n6453), .B2(n6452), .A(n6451), .ZN(n6456) );
  AOI22_X1 U7423 ( .A1(n6456), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6455), 
        .B2(n6454), .ZN(n6461) );
  NAND2_X1 U7424 ( .A1(n6457), .A2(REIP_REG_2__SCAN_IN), .ZN(n6460) );
  NAND3_X1 U7425 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6458), .A3(n3534), 
        .ZN(n6459) );
  NAND4_X1 U7426 ( .A1(n6462), .A2(n6461), .A3(n6460), .A4(n6459), .ZN(U3016)
         );
  AND2_X1 U7427 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6463), .ZN(U3019)
         );
  NAND3_X1 U7428 ( .A1(n6465), .A2(n6464), .A3(n6630), .ZN(n6466) );
  OAI21_X1 U7429 ( .B1(n6467), .B2(n4690), .A(n6466), .ZN(n6507) );
  NOR2_X1 U7430 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6468), .ZN(n6505)
         );
  AOI22_X1 U7431 ( .A1(n6549), .A2(n6507), .B1(n6469), .B2(n6505), .ZN(n6480)
         );
  NAND3_X1 U7432 ( .A1(n6477), .A2(n6537), .A3(n6532), .ZN(n6472) );
  AOI21_X1 U7433 ( .B1(n6472), .B2(n6471), .A(n6470), .ZN(n6476) );
  OAI211_X1 U7434 ( .C1(n6505), .C2(n6722), .A(n6473), .B(n6630), .ZN(n6474)
         );
  AOI22_X1 U7435 ( .A1(n6510), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6478), 
        .B2(n6508), .ZN(n6479) );
  OAI211_X1 U7436 ( .C1(n6535), .C2(n6532), .A(n6480), .B(n6479), .ZN(U3068)
         );
  AOI22_X1 U7437 ( .A1(n6556), .A2(n6507), .B1(n6481), .B2(n6505), .ZN(n6484)
         );
  AOI22_X1 U7438 ( .A1(n6510), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6482), 
        .B2(n6508), .ZN(n6483) );
  OAI211_X1 U7439 ( .C1(n6554), .C2(n6532), .A(n6484), .B(n6483), .ZN(U3069)
         );
  AOI22_X1 U7440 ( .A1(n6563), .A2(n6507), .B1(n6485), .B2(n6505), .ZN(n6488)
         );
  AOI22_X1 U7441 ( .A1(n6510), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6486), 
        .B2(n6508), .ZN(n6487) );
  OAI211_X1 U7442 ( .C1(n6561), .C2(n6532), .A(n6488), .B(n6487), .ZN(U3070)
         );
  AOI22_X1 U7443 ( .A1(n6570), .A2(n6507), .B1(n6489), .B2(n6505), .ZN(n6492)
         );
  AOI22_X1 U7444 ( .A1(n6510), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6490), 
        .B2(n6508), .ZN(n6491) );
  OAI211_X1 U7445 ( .C1(n6568), .C2(n6532), .A(n6492), .B(n6491), .ZN(U3071)
         );
  AOI22_X1 U7446 ( .A1(n6577), .A2(n6507), .B1(n6493), .B2(n6505), .ZN(n6496)
         );
  AOI22_X1 U7447 ( .A1(n6510), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6494), 
        .B2(n6508), .ZN(n6495) );
  OAI211_X1 U7448 ( .C1(n6575), .C2(n6532), .A(n6496), .B(n6495), .ZN(U3072)
         );
  AOI22_X1 U7449 ( .A1(n6584), .A2(n6507), .B1(n6497), .B2(n6505), .ZN(n6500)
         );
  AOI22_X1 U7450 ( .A1(n6510), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6498), 
        .B2(n6508), .ZN(n6499) );
  OAI211_X1 U7451 ( .C1(n6587), .C2(n6532), .A(n6500), .B(n6499), .ZN(U3073)
         );
  AOI22_X1 U7452 ( .A1(n6591), .A2(n6507), .B1(n6501), .B2(n6505), .ZN(n6504)
         );
  AOI22_X1 U7453 ( .A1(n6510), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6502), 
        .B2(n6508), .ZN(n6503) );
  OAI211_X1 U7454 ( .C1(n6589), .C2(n6532), .A(n6504), .B(n6503), .ZN(U3074)
         );
  AOI22_X1 U7455 ( .A1(n6601), .A2(n6507), .B1(n6506), .B2(n6505), .ZN(n6512)
         );
  AOI22_X1 U7456 ( .A1(n6510), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6509), 
        .B2(n6508), .ZN(n6511) );
  OAI211_X1 U7457 ( .C1(n6606), .C2(n6532), .A(n6512), .B(n6511), .ZN(U3075)
         );
  OAI22_X1 U7458 ( .A1(n6526), .A2(n6535), .B1(n6525), .B2(n6534), .ZN(n6513)
         );
  INV_X1 U7459 ( .A(n6513), .ZN(n6515) );
  AOI22_X1 U7460 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6529), .B1(n6549), 
        .B2(n6528), .ZN(n6514) );
  OAI211_X1 U7461 ( .C1(n6552), .C2(n6532), .A(n6515), .B(n6514), .ZN(U3076)
         );
  OAI22_X1 U7462 ( .A1(n6526), .A2(n6561), .B1(n6525), .B2(n6560), .ZN(n6516)
         );
  INV_X1 U7463 ( .A(n6516), .ZN(n6518) );
  AOI22_X1 U7464 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6529), .B1(n6563), 
        .B2(n6528), .ZN(n6517) );
  OAI211_X1 U7465 ( .C1(n6566), .C2(n6532), .A(n6518), .B(n6517), .ZN(U3078)
         );
  OAI22_X1 U7466 ( .A1(n6526), .A2(n6568), .B1(n6525), .B2(n6567), .ZN(n6519)
         );
  INV_X1 U7467 ( .A(n6519), .ZN(n6521) );
  AOI22_X1 U7468 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6529), .B1(n6570), 
        .B2(n6528), .ZN(n6520) );
  OAI211_X1 U7469 ( .C1(n6573), .C2(n6532), .A(n6521), .B(n6520), .ZN(U3079)
         );
  OAI22_X1 U7470 ( .A1(n6526), .A2(n6587), .B1(n6525), .B2(n6581), .ZN(n6522)
         );
  INV_X1 U7471 ( .A(n6522), .ZN(n6524) );
  AOI22_X1 U7472 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6529), .B1(n6584), 
        .B2(n6528), .ZN(n6523) );
  OAI211_X1 U7473 ( .C1(n6582), .C2(n6532), .A(n6524), .B(n6523), .ZN(U3081)
         );
  OAI22_X1 U7474 ( .A1(n6526), .A2(n6589), .B1(n6525), .B2(n6588), .ZN(n6527)
         );
  INV_X1 U7475 ( .A(n6527), .ZN(n6531) );
  AOI22_X1 U7476 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6529), .B1(n6591), 
        .B2(n6528), .ZN(n6530) );
  OAI211_X1 U7477 ( .C1(n6594), .C2(n6532), .A(n6531), .B(n6530), .ZN(U3082)
         );
  NOR2_X1 U7478 ( .A1(n6533), .A2(n6630), .ZN(n6540) );
  INV_X1 U7479 ( .A(n6540), .ZN(n6595) );
  OAI22_X1 U7480 ( .A1(n6605), .A2(n6535), .B1(n6534), .B2(n6595), .ZN(n6536)
         );
  INV_X1 U7481 ( .A(n6536), .ZN(n6551) );
  OAI21_X1 U7482 ( .B1(n6539), .B2(n6538), .A(n6537), .ZN(n6548) );
  AOI21_X1 U7483 ( .B1(n6541), .B2(n6616), .A(n6540), .ZN(n6547) );
  INV_X1 U7484 ( .A(n6547), .ZN(n6545) );
  AOI21_X1 U7485 ( .B1(n6543), .B2(n6546), .A(n6542), .ZN(n6544) );
  OAI21_X1 U7486 ( .B1(n6548), .B2(n6545), .A(n6544), .ZN(n6602) );
  OAI22_X1 U7487 ( .A1(n6548), .A2(n6547), .B1(n6546), .B2(n6655), .ZN(n6600)
         );
  AOI22_X1 U7488 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6602), .B1(n6549), 
        .B2(n6600), .ZN(n6550) );
  OAI211_X1 U7489 ( .C1(n6552), .C2(n6598), .A(n6551), .B(n6550), .ZN(U3108)
         );
  OAI22_X1 U7490 ( .A1(n6605), .A2(n6554), .B1(n6553), .B2(n6595), .ZN(n6555)
         );
  INV_X1 U7491 ( .A(n6555), .ZN(n6558) );
  AOI22_X1 U7492 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6602), .B1(n6556), 
        .B2(n6600), .ZN(n6557) );
  OAI211_X1 U7493 ( .C1(n6559), .C2(n6598), .A(n6558), .B(n6557), .ZN(U3109)
         );
  OAI22_X1 U7494 ( .A1(n6605), .A2(n6561), .B1(n6560), .B2(n6595), .ZN(n6562)
         );
  INV_X1 U7495 ( .A(n6562), .ZN(n6565) );
  AOI22_X1 U7496 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6602), .B1(n6563), 
        .B2(n6600), .ZN(n6564) );
  OAI211_X1 U7497 ( .C1(n6566), .C2(n6598), .A(n6565), .B(n6564), .ZN(U3110)
         );
  OAI22_X1 U7498 ( .A1(n6605), .A2(n6568), .B1(n6567), .B2(n6595), .ZN(n6569)
         );
  INV_X1 U7499 ( .A(n6569), .ZN(n6572) );
  AOI22_X1 U7500 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6602), .B1(n6570), 
        .B2(n6600), .ZN(n6571) );
  OAI211_X1 U7501 ( .C1(n6573), .C2(n6598), .A(n6572), .B(n6571), .ZN(U3111)
         );
  OAI22_X1 U7502 ( .A1(n6605), .A2(n6575), .B1(n6574), .B2(n6595), .ZN(n6576)
         );
  INV_X1 U7503 ( .A(n6576), .ZN(n6579) );
  AOI22_X1 U7504 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6602), .B1(n6577), 
        .B2(n6600), .ZN(n6578) );
  OAI211_X1 U7505 ( .C1(n6580), .C2(n6598), .A(n6579), .B(n6578), .ZN(U3112)
         );
  OAI22_X1 U7506 ( .A1(n6598), .A2(n6582), .B1(n6581), .B2(n6595), .ZN(n6583)
         );
  INV_X1 U7507 ( .A(n6583), .ZN(n6586) );
  AOI22_X1 U7508 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6602), .B1(n6584), 
        .B2(n6600), .ZN(n6585) );
  OAI211_X1 U7509 ( .C1(n6587), .C2(n6605), .A(n6586), .B(n6585), .ZN(U3113)
         );
  OAI22_X1 U7510 ( .A1(n6605), .A2(n6589), .B1(n6588), .B2(n6595), .ZN(n6590)
         );
  INV_X1 U7511 ( .A(n6590), .ZN(n6593) );
  AOI22_X1 U7512 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6602), .B1(n6591), 
        .B2(n6600), .ZN(n6592) );
  OAI211_X1 U7513 ( .C1(n6594), .C2(n6598), .A(n6593), .B(n6592), .ZN(U3114)
         );
  OAI22_X1 U7514 ( .A1(n6598), .A2(n6597), .B1(n6596), .B2(n6595), .ZN(n6599)
         );
  INV_X1 U7515 ( .A(n6599), .ZN(n6604) );
  AOI22_X1 U7516 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6602), .B1(n6601), 
        .B2(n6600), .ZN(n6603) );
  OAI211_X1 U7517 ( .C1(n6606), .C2(n6605), .A(n6604), .B(n6603), .ZN(U3115)
         );
  NOR2_X1 U7518 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6609) );
  OAI211_X1 U7519 ( .C1(n6610), .C2(n6609), .A(n6608), .B(n6607), .ZN(n6611)
         );
  NOR2_X1 U7520 ( .A1(n6612), .A2(n6611), .ZN(n6637) );
  NOR2_X1 U7521 ( .A1(n6613), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6614)
         );
  AOI21_X1 U7522 ( .B1(n6616), .B2(n6615), .A(n6614), .ZN(n6721) );
  NAND2_X1 U7523 ( .A1(n6617), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6731) );
  AND2_X1 U7524 ( .A1(n6731), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6618)
         );
  AND2_X1 U7525 ( .A1(n6721), .A2(n6618), .ZN(n6622) );
  NAND2_X1 U7526 ( .A1(n6622), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6624) );
  NAND2_X1 U7527 ( .A1(n6620), .A2(n6619), .ZN(n6621) );
  OAI21_X1 U7528 ( .B1(n6622), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6621), 
        .ZN(n6623) );
  OAI211_X1 U7529 ( .C1(n6626), .C2(n6625), .A(n6624), .B(n6623), .ZN(n6628)
         );
  NAND2_X1 U7530 ( .A1(n6626), .A2(n6625), .ZN(n6627) );
  NAND2_X1 U7531 ( .A1(n6628), .A2(n6627), .ZN(n6629) );
  OAI21_X1 U7532 ( .B1(n6631), .B2(n6630), .A(n6629), .ZN(n6633) );
  NAND2_X1 U7533 ( .A1(n6631), .A2(n6630), .ZN(n6632) );
  NAND2_X1 U7534 ( .A1(n6633), .A2(n6632), .ZN(n6635) );
  INV_X1 U7535 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6634) );
  NAND2_X1 U7536 ( .A1(n6635), .A2(n6634), .ZN(n6636) );
  NAND2_X1 U7537 ( .A1(n6651), .A2(n6652), .ZN(n6640) );
  NAND2_X1 U7538 ( .A1(READY_N), .A2(n6638), .ZN(n6639) );
  NAND2_X1 U7539 ( .A1(n6640), .A2(n6639), .ZN(n6644) );
  OR2_X1 U7540 ( .A1(n6642), .A2(n6641), .ZN(n6643) );
  OAI21_X1 U7541 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5605), .A(n6720), .ZN(
        n6657) );
  AOI221_X1 U7542 ( .B1(n6646), .B2(STATE2_REG_0__SCAN_IN), .C1(n6657), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6645), .ZN(n6649) );
  OAI211_X1 U7543 ( .C1(n6647), .C2(n6724), .A(n6656), .B(n6720), .ZN(n6648)
         );
  OAI211_X1 U7544 ( .C1(n6651), .C2(n6650), .A(n6649), .B(n6648), .ZN(U3148)
         );
  AOI21_X1 U7545 ( .B1(n6653), .B2(n5605), .A(n6652), .ZN(n6660) );
  INV_X1 U7546 ( .A(n6654), .ZN(n6659) );
  NAND2_X1 U7547 ( .A1(n6656), .A2(n6655), .ZN(n6662) );
  NAND3_X1 U7548 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6662), .A3(n6657), .ZN(
        n6658) );
  OAI211_X1 U7549 ( .C1(n6661), .C2(n6660), .A(n6659), .B(n6658), .ZN(U3149)
         );
  OAI211_X1 U7550 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n5605), .A(n6718), .B(
        n6662), .ZN(n6664) );
  OAI21_X1 U7551 ( .B1(n6746), .B2(n6664), .A(n6663), .ZN(U3150) );
  AND2_X1 U7552 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6715), .ZN(U3151) );
  AND2_X1 U7553 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6715), .ZN(U3152) );
  AND2_X1 U7554 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6715), .ZN(U3153) );
  AND2_X1 U7555 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6715), .ZN(U3154) );
  AND2_X1 U7556 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6715), .ZN(U3155) );
  AND2_X1 U7557 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6715), .ZN(U3156) );
  AND2_X1 U7558 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6715), .ZN(U3157) );
  AND2_X1 U7559 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6715), .ZN(U3158) );
  AND2_X1 U7560 ( .A1(n6715), .A2(DATAWIDTH_REG_23__SCAN_IN), .ZN(U3159) );
  INV_X1 U7561 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6878) );
  NOR2_X1 U7562 ( .A1(n6717), .A2(n6878), .ZN(U3160) );
  AND2_X1 U7563 ( .A1(n6715), .A2(DATAWIDTH_REG_21__SCAN_IN), .ZN(U3161) );
  AND2_X1 U7564 ( .A1(n6715), .A2(DATAWIDTH_REG_20__SCAN_IN), .ZN(U3162) );
  INV_X1 U7565 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n7027) );
  NOR2_X1 U7566 ( .A1(n6717), .A2(n7027), .ZN(U3163) );
  INV_X1 U7567 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n7104) );
  NOR2_X1 U7568 ( .A1(n6717), .A2(n7104), .ZN(U3164) );
  INV_X1 U7569 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n7064) );
  NOR2_X1 U7570 ( .A1(n6717), .A2(n7064), .ZN(U3165) );
  AND2_X1 U7571 ( .A1(n6715), .A2(DATAWIDTH_REG_16__SCAN_IN), .ZN(U3166) );
  INV_X1 U7572 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6857) );
  NOR2_X1 U7573 ( .A1(n6717), .A2(n6857), .ZN(U3167) );
  INV_X1 U7574 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6845) );
  NOR2_X1 U7575 ( .A1(n6717), .A2(n6845), .ZN(U3168) );
  AND2_X1 U7576 ( .A1(n6715), .A2(DATAWIDTH_REG_13__SCAN_IN), .ZN(U3169) );
  INV_X1 U7577 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6915) );
  NOR2_X1 U7578 ( .A1(n6717), .A2(n6915), .ZN(U3170) );
  AND2_X1 U7579 ( .A1(n6715), .A2(DATAWIDTH_REG_11__SCAN_IN), .ZN(U3171) );
  INV_X1 U7580 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6911) );
  NOR2_X1 U7581 ( .A1(n6717), .A2(n6911), .ZN(U3172) );
  INV_X1 U7582 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6833) );
  NOR2_X1 U7583 ( .A1(n6717), .A2(n6833), .ZN(U3173) );
  AND2_X1 U7584 ( .A1(n6715), .A2(DATAWIDTH_REG_8__SCAN_IN), .ZN(U3174) );
  INV_X1 U7585 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6848) );
  NOR2_X1 U7586 ( .A1(n6717), .A2(n6848), .ZN(U3175) );
  AND2_X1 U7587 ( .A1(n6715), .A2(DATAWIDTH_REG_6__SCAN_IN), .ZN(U3176) );
  INV_X1 U7588 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n7081) );
  NOR2_X1 U7589 ( .A1(n6717), .A2(n7081), .ZN(U3177) );
  AND2_X1 U7590 ( .A1(n6715), .A2(DATAWIDTH_REG_4__SCAN_IN), .ZN(U3178) );
  INV_X1 U7591 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6877) );
  NOR2_X1 U7592 ( .A1(n6717), .A2(n6877), .ZN(U3179) );
  INV_X1 U7593 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6854) );
  NOR2_X1 U7594 ( .A1(n6717), .A2(n6854), .ZN(U3180) );
  NAND2_X1 U7595 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6668) );
  NAND2_X1 U7596 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6666) );
  NAND2_X1 U7597 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6669) );
  NAND2_X1 U7598 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6675) );
  NAND2_X1 U7599 ( .A1(n6669), .A2(n6675), .ZN(n6665) );
  INV_X1 U7600 ( .A(NA_N), .ZN(n7114) );
  AOI221_X1 U7601 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n7114), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6679) );
  AOI21_X1 U7602 ( .B1(n6666), .B2(n6665), .A(n6679), .ZN(n6667) );
  OAI221_X1 U7603 ( .B1(n6713), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n6713), 
        .C2(n6668), .A(n6667), .ZN(U3181) );
  INV_X1 U7604 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6676) );
  NOR2_X1 U7605 ( .A1(n3751), .A2(n6676), .ZN(n6671) );
  INV_X1 U7606 ( .A(n6668), .ZN(n6670) );
  OAI21_X1 U7607 ( .B1(n6671), .B2(n6670), .A(n6669), .ZN(n6672) );
  NAND3_X1 U7608 ( .A1(n6673), .A2(n6675), .A3(n6672), .ZN(U3182) );
  AOI221_X1 U7609 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n5605), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6674) );
  AOI221_X1 U7610 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6674), .C2(HOLD), .A(n3751), .ZN(n6680) );
  OR4_X1 U7611 ( .A1(n6676), .A2(n3751), .A3(n6675), .A4(NA_N), .ZN(n6678) );
  NAND3_X1 U7612 ( .A1(READY_N), .A2(STATE_REG_2__SCAN_IN), .A3(
        STATE_REG_1__SCAN_IN), .ZN(n6677) );
  OAI211_X1 U7613 ( .C1(n6680), .C2(n6679), .A(n6678), .B(n6677), .ZN(U3183)
         );
  INV_X1 U7614 ( .A(STATE_REG_2__SCAN_IN), .ZN(n7076) );
  NAND2_X1 U7615 ( .A1(n6713), .A2(n7076), .ZN(n6698) );
  INV_X1 U7616 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6682) );
  INV_X1 U7617 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6681) );
  OAI222_X1 U7618 ( .A1(n6698), .A2(n6682), .B1(n6681), .B2(n6713), .C1(n6733), 
        .C2(n6708), .ZN(U3184) );
  INV_X1 U7619 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n7002) );
  OAI222_X1 U7620 ( .A1(n6708), .A2(n6682), .B1(n7002), .B2(n6713), .C1(n6683), 
        .C2(n6709), .ZN(U3185) );
  INV_X1 U7621 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n7108) );
  OAI222_X1 U7622 ( .A1(n6708), .A2(n6683), .B1(n7108), .B2(n6713), .C1(n6684), 
        .C2(n6709), .ZN(U3186) );
  INV_X1 U7623 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n7061) );
  INV_X1 U7624 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6685) );
  OAI222_X1 U7625 ( .A1(n6708), .A2(n6684), .B1(n7061), .B2(n6713), .C1(n6685), 
        .C2(n6709), .ZN(U3187) );
  INV_X1 U7626 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n7047) );
  INV_X1 U7627 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6686) );
  OAI222_X1 U7628 ( .A1(n6708), .A2(n6685), .B1(n7047), .B2(n6713), .C1(n6686), 
        .C2(n6709), .ZN(U3188) );
  INV_X1 U7629 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n7030) );
  OAI222_X1 U7630 ( .A1(n6708), .A2(n6686), .B1(n7030), .B2(n6713), .C1(n6688), 
        .C2(n6709), .ZN(U3189) );
  INV_X1 U7631 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6687) );
  OAI222_X1 U7632 ( .A1(n6708), .A2(n6688), .B1(n6687), .B2(n6713), .C1(n6689), 
        .C2(n6698), .ZN(U3190) );
  INV_X1 U7633 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n7044) );
  OAI222_X1 U7634 ( .A1(n6698), .A2(n6690), .B1(n7044), .B2(n6713), .C1(n6689), 
        .C2(n6708), .ZN(U3191) );
  INV_X1 U7635 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n7070) );
  OAI222_X1 U7636 ( .A1(n6708), .A2(n6690), .B1(n7070), .B2(n6713), .C1(n6692), 
        .C2(n6698), .ZN(U3192) );
  INV_X1 U7637 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n6691) );
  INV_X1 U7638 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6693) );
  OAI222_X1 U7639 ( .A1(n6708), .A2(n6692), .B1(n6691), .B2(n6713), .C1(n6693), 
        .C2(n6698), .ZN(U3193) );
  INV_X1 U7640 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6836) );
  OAI222_X1 U7641 ( .A1(n6708), .A2(n6693), .B1(n6836), .B2(n6713), .C1(n6694), 
        .C2(n6698), .ZN(U3194) );
  INV_X1 U7642 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6903) );
  OAI222_X1 U7643 ( .A1(n6708), .A2(n6694), .B1(n6903), .B2(n6713), .C1(n6696), 
        .C2(n6698), .ZN(U3195) );
  INV_X1 U7644 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6695) );
  OAI222_X1 U7645 ( .A1(n6708), .A2(n6696), .B1(n6695), .B2(n6713), .C1(n6697), 
        .C2(n6698), .ZN(U3196) );
  INV_X1 U7646 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6699) );
  INV_X1 U7647 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n7079) );
  OAI222_X1 U7648 ( .A1(n6698), .A2(n6699), .B1(n7079), .B2(n6713), .C1(n6697), 
        .C2(n6708), .ZN(U3197) );
  INV_X1 U7649 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n7011) );
  INV_X1 U7650 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6916) );
  OAI222_X1 U7651 ( .A1(n6708), .A2(n6699), .B1(n7011), .B2(n6713), .C1(n6916), 
        .C2(n6698), .ZN(U3198) );
  INV_X1 U7652 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n6700) );
  OAI222_X1 U7653 ( .A1(n6708), .A2(n6916), .B1(n6700), .B2(n6713), .C1(n6701), 
        .C2(n6709), .ZN(U3199) );
  INV_X1 U7654 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6873) );
  OAI222_X1 U7655 ( .A1(n6709), .A2(n7045), .B1(n6873), .B2(n6713), .C1(n6701), 
        .C2(n6708), .ZN(U3200) );
  INV_X1 U7656 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6824) );
  OAI222_X1 U7657 ( .A1(n6708), .A2(n7045), .B1(n6824), .B2(n6713), .C1(n6702), 
        .C2(n6709), .ZN(U3201) );
  INV_X1 U7658 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n7026) );
  OAI222_X1 U7659 ( .A1(n6708), .A2(n6702), .B1(n7026), .B2(n6713), .C1(n7078), 
        .C2(n6709), .ZN(U3202) );
  INV_X1 U7660 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6703) );
  OAI222_X1 U7661 ( .A1(n6708), .A2(n7078), .B1(n6703), .B2(n6713), .C1(n5779), 
        .C2(n6709), .ZN(U3203) );
  INV_X1 U7662 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6704) );
  OAI222_X1 U7663 ( .A1(n6708), .A2(n5779), .B1(n6704), .B2(n6713), .C1(n6705), 
        .C2(n6709), .ZN(U3204) );
  INV_X1 U7664 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n7010) );
  OAI222_X1 U7665 ( .A1(n6708), .A2(n6705), .B1(n7010), .B2(n6713), .C1(n3883), 
        .C2(n6709), .ZN(U3205) );
  INV_X1 U7666 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n7111) );
  OAI222_X1 U7667 ( .A1(n6708), .A2(n3883), .B1(n7111), .B2(n6713), .C1(n7019), 
        .C2(n6709), .ZN(U3206) );
  INV_X1 U7668 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6887) );
  OAI222_X1 U7669 ( .A1(n6709), .A2(n6860), .B1(n6887), .B2(n6713), .C1(n7019), 
        .C2(n6708), .ZN(U3207) );
  INV_X1 U7670 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n7091) );
  INV_X1 U7671 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6706) );
  OAI222_X1 U7672 ( .A1(n6708), .A2(n6860), .B1(n7091), .B2(n6713), .C1(n6706), 
        .C2(n6709), .ZN(U3208) );
  INV_X1 U7673 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n7004) );
  OAI222_X1 U7674 ( .A1(n6708), .A2(n6706), .B1(n7004), .B2(n6713), .C1(n7051), 
        .C2(n6709), .ZN(U3209) );
  INV_X1 U7675 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6943) );
  OAI222_X1 U7676 ( .A1(n6708), .A2(n7051), .B1(n6943), .B2(n6713), .C1(n7067), 
        .C2(n6709), .ZN(U3210) );
  INV_X1 U7677 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n7007) );
  OAI222_X1 U7678 ( .A1(n6708), .A2(n7067), .B1(n7007), .B2(n6713), .C1(n7097), 
        .C2(n6709), .ZN(U3211) );
  INV_X1 U7679 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6707) );
  OAI222_X1 U7680 ( .A1(n6708), .A2(n7097), .B1(n6707), .B2(n6713), .C1(n6913), 
        .C2(n6709), .ZN(U3212) );
  INV_X1 U7681 ( .A(REIP_REG_31__SCAN_IN), .ZN(n7050) );
  INV_X1 U7682 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6831) );
  OAI222_X1 U7683 ( .A1(n6709), .A2(n7050), .B1(n6831), .B2(n6713), .C1(n6913), 
        .C2(n6708), .ZN(U3213) );
  INV_X1 U7684 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6736) );
  INV_X1 U7685 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n7110) );
  AOI22_X1 U7686 ( .A1(n6713), .A2(n6736), .B1(n7110), .B2(n7142), .ZN(U3446)
         );
  INV_X1 U7687 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6710) );
  AOI22_X1 U7688 ( .A1(n6713), .A2(n6711), .B1(n6710), .B2(n7142), .ZN(U3447)
         );
  INV_X1 U7689 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n7062) );
  INV_X1 U7690 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6712) );
  AOI22_X1 U7691 ( .A1(n6713), .A2(n7062), .B1(n6712), .B2(n7142), .ZN(U3448)
         );
  INV_X1 U7692 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n7005) );
  INV_X1 U7693 ( .A(n6716), .ZN(n6714) );
  AOI21_X1 U7694 ( .B1(n7005), .B2(n6715), .A(n6714), .ZN(U3451) );
  OAI21_X1 U7695 ( .B1(n6717), .B2(n6888), .A(n6716), .ZN(U3452) );
  OAI211_X1 U7696 ( .C1(n6722), .C2(n6720), .A(n6719), .B(n6718), .ZN(U3453)
         );
  INV_X1 U7697 ( .A(n6721), .ZN(n6723) );
  AOI21_X1 U7698 ( .B1(n6723), .B2(n6722), .A(STATE2_REG_1__SCAN_IN), .ZN(
        n6725) );
  OAI22_X1 U7699 ( .A1(n6726), .A2(n6725), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6724), .ZN(n6728) );
  AOI22_X1 U7700 ( .A1(n6729), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(n6728), .B2(n6727), .ZN(n6730) );
  OAI21_X1 U7701 ( .B1(n6732), .B2(n6731), .A(n6730), .ZN(U3461) );
  AOI21_X1 U7702 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6734) );
  AOI22_X1 U7703 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6734), .B2(n6733), .ZN(n6737) );
  AOI22_X1 U7704 ( .A1(n6739), .A2(n6737), .B1(n6736), .B2(n6735), .ZN(U3468)
         );
  OAI21_X1 U7705 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6739), .ZN(n6738) );
  OAI21_X1 U7706 ( .B1(n6739), .B2(n7062), .A(n6738), .ZN(U3469) );
  INV_X1 U7707 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6740) );
  AOI22_X1 U7708 ( .A1(n6713), .A2(READREQUEST_REG_SCAN_IN), .B1(n6740), .B2(
        n7142), .ZN(U3470) );
  AOI211_X1 U7709 ( .C1(n6743), .C2(n5605), .A(n6742), .B(n6741), .ZN(n6750)
         );
  OAI211_X1 U7710 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6745), .A(n6744), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6747) );
  AOI21_X1 U7711 ( .B1(n6747), .B2(STATE2_REG_0__SCAN_IN), .A(n6746), .ZN(
        n6749) );
  NAND2_X1 U7712 ( .A1(n6750), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6748) );
  OAI21_X1 U7713 ( .B1(n6750), .B2(n6749), .A(n6748), .ZN(U3472) );
  INV_X1 U7714 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n7105) );
  INV_X1 U7715 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6834) );
  AOI22_X1 U7716 ( .A1(n6713), .A2(n7105), .B1(n6834), .B2(n7142), .ZN(U3473)
         );
  OAI22_X1 U7717 ( .A1(BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_g48), .B1(
        DATAWIDTH_REG_8__SCAN_IN), .B2(keyinput_g112), .ZN(n6751) );
  AOI221_X1 U7718 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_g48), .C1(
        keyinput_g112), .C2(DATAWIDTH_REG_8__SCAN_IN), .A(n6751), .ZN(n6758)
         );
  OAI22_X1 U7719 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(keyinput_g124), .B1(
        keyinput_g125), .B2(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6752) );
  AOI221_X1 U7720 ( .B1(DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput_g124), .C1(
        DATAWIDTH_REG_21__SCAN_IN), .C2(keyinput_g125), .A(n6752), .ZN(n6757)
         );
  OAI22_X1 U7721 ( .A1(REIP_REG_28__SCAN_IN), .A2(keyinput_g54), .B1(
        keyinput_g5), .B2(DATAI_26_), .ZN(n6753) );
  AOI221_X1 U7722 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_g54), .C1(
        DATAI_26_), .C2(keyinput_g5), .A(n6753), .ZN(n6756) );
  OAI22_X1 U7723 ( .A1(REIP_REG_21__SCAN_IN), .A2(keyinput_g61), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(keyinput_g80), .ZN(n6754) );
  AOI221_X1 U7724 ( .B1(REIP_REG_21__SCAN_IN), .B2(keyinput_g61), .C1(
        keyinput_g80), .C2(ADDRESS_REG_20__SCAN_IN), .A(n6754), .ZN(n6755) );
  NAND4_X1 U7725 ( .A1(n6758), .A2(n6757), .A3(n6756), .A4(n6755), .ZN(n6786)
         );
  OAI22_X1 U7726 ( .A1(ADDRESS_REG_1__SCAN_IN), .A2(keyinput_g99), .B1(
        keyinput_g34), .B2(BS16_N), .ZN(n6759) );
  AOI221_X1 U7727 ( .B1(ADDRESS_REG_1__SCAN_IN), .B2(keyinput_g99), .C1(BS16_N), .C2(keyinput_g34), .A(n6759), .ZN(n6766) );
  OAI22_X1 U7728 ( .A1(REIP_REG_26__SCAN_IN), .A2(keyinput_g56), .B1(
        keyinput_g117), .B2(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6760) );
  AOI221_X1 U7729 ( .B1(REIP_REG_26__SCAN_IN), .B2(keyinput_g56), .C1(
        DATAWIDTH_REG_13__SCAN_IN), .C2(keyinput_g117), .A(n6760), .ZN(n6765)
         );
  OAI22_X1 U7730 ( .A1(REIP_REG_19__SCAN_IN), .A2(keyinput_g63), .B1(
        keyinput_g75), .B2(ADDRESS_REG_25__SCAN_IN), .ZN(n6761) );
  AOI221_X1 U7731 ( .B1(REIP_REG_19__SCAN_IN), .B2(keyinput_g63), .C1(
        ADDRESS_REG_25__SCAN_IN), .C2(keyinput_g75), .A(n6761), .ZN(n6764) );
  OAI22_X1 U7732 ( .A1(DATAI_27_), .A2(keyinput_g4), .B1(
        DATAWIDTH_REG_6__SCAN_IN), .B2(keyinput_g110), .ZN(n6762) );
  AOI221_X1 U7733 ( .B1(DATAI_27_), .B2(keyinput_g4), .C1(keyinput_g110), .C2(
        DATAWIDTH_REG_6__SCAN_IN), .A(n6762), .ZN(n6763) );
  NAND4_X1 U7734 ( .A1(n6766), .A2(n6765), .A3(n6764), .A4(n6763), .ZN(n6785)
         );
  OAI22_X1 U7735 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(keyinput_g123), .B1(
        keyinput_g109), .B2(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6767) );
  AOI221_X1 U7736 ( .B1(DATAWIDTH_REG_19__SCAN_IN), .B2(keyinput_g123), .C1(
        DATAWIDTH_REG_5__SCAN_IN), .C2(keyinput_g109), .A(n6767), .ZN(n6774)
         );
  OAI22_X1 U7737 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(keyinput_g127), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(keyinput_g86), .ZN(n6768) );
  AOI221_X1 U7738 ( .B1(DATAWIDTH_REG_23__SCAN_IN), .B2(keyinput_g127), .C1(
        keyinput_g86), .C2(ADDRESS_REG_14__SCAN_IN), .A(n6768), .ZN(n6773) );
  OAI22_X1 U7739 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput_g60), .B1(
        keyinput_g2), .B2(DATAI_29_), .ZN(n6769) );
  AOI221_X1 U7740 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_g60), .C1(
        DATAI_29_), .C2(keyinput_g2), .A(n6769), .ZN(n6772) );
  OAI22_X1 U7741 ( .A1(REIP_REG_18__SCAN_IN), .A2(keyinput_g64), .B1(
        keyinput_g49), .B2(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6770) );
  AOI221_X1 U7742 ( .B1(REIP_REG_18__SCAN_IN), .B2(keyinput_g64), .C1(
        BYTEENABLE_REG_2__SCAN_IN), .C2(keyinput_g49), .A(n6770), .ZN(n6771)
         );
  NAND4_X1 U7743 ( .A1(n6774), .A2(n6773), .A3(n6772), .A4(n6771), .ZN(n6784)
         );
  OAI22_X1 U7744 ( .A1(DATAI_10_), .A2(keyinput_g21), .B1(keyinput_g68), .B2(
        BE_N_REG_2__SCAN_IN), .ZN(n6775) );
  AOI221_X1 U7745 ( .B1(DATAI_10_), .B2(keyinput_g21), .C1(BE_N_REG_2__SCAN_IN), .C2(keyinput_g68), .A(n6775), .ZN(n6782) );
  OAI22_X1 U7746 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(keyinput_g115), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(keyinput_g88), .ZN(n6776) );
  AOI221_X1 U7747 ( .B1(DATAWIDTH_REG_11__SCAN_IN), .B2(keyinput_g115), .C1(
        keyinput_g88), .C2(ADDRESS_REG_12__SCAN_IN), .A(n6776), .ZN(n6781) );
  OAI22_X1 U7748 ( .A1(DATAI_7_), .A2(keyinput_g24), .B1(
        DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput_g104), .ZN(n6777) );
  AOI221_X1 U7749 ( .B1(DATAI_7_), .B2(keyinput_g24), .C1(keyinput_g104), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(n6777), .ZN(n6780) );
  OAI22_X1 U7750 ( .A1(D_C_N_REG_SCAN_IN), .A2(keyinput_g41), .B1(
        keyinput_g100), .B2(ADDRESS_REG_0__SCAN_IN), .ZN(n6778) );
  AOI221_X1 U7751 ( .B1(D_C_N_REG_SCAN_IN), .B2(keyinput_g41), .C1(
        ADDRESS_REG_0__SCAN_IN), .C2(keyinput_g100), .A(n6778), .ZN(n6779) );
  NAND4_X1 U7752 ( .A1(n6782), .A2(n6781), .A3(n6780), .A4(n6779), .ZN(n6783)
         );
  NOR4_X1 U7753 ( .A1(n6786), .A2(n6785), .A3(n6784), .A4(n6783), .ZN(n7141)
         );
  OAI22_X1 U7754 ( .A1(DATAI_14_), .A2(keyinput_g17), .B1(keyinput_g70), .B2(
        BE_N_REG_0__SCAN_IN), .ZN(n6787) );
  AOI221_X1 U7755 ( .B1(DATAI_14_), .B2(keyinput_g17), .C1(BE_N_REG_0__SCAN_IN), .C2(keyinput_g70), .A(n6787), .ZN(n6794) );
  OAI22_X1 U7756 ( .A1(REIP_REG_23__SCAN_IN), .A2(keyinput_g59), .B1(
        DATAWIDTH_REG_16__SCAN_IN), .B2(keyinput_g120), .ZN(n6788) );
  AOI221_X1 U7757 ( .B1(REIP_REG_23__SCAN_IN), .B2(keyinput_g59), .C1(
        keyinput_g120), .C2(DATAWIDTH_REG_16__SCAN_IN), .A(n6788), .ZN(n6793)
         );
  OAI22_X1 U7758 ( .A1(ADDRESS_REG_6__SCAN_IN), .A2(keyinput_g94), .B1(
        ADS_N_REG_SCAN_IN), .B2(keyinput_g38), .ZN(n6789) );
  AOI221_X1 U7759 ( .B1(ADDRESS_REG_6__SCAN_IN), .B2(keyinput_g94), .C1(
        keyinput_g38), .C2(ADS_N_REG_SCAN_IN), .A(n6789), .ZN(n6792) );
  OAI22_X1 U7760 ( .A1(DATAI_31_), .A2(keyinput_g0), .B1(DATAI_24_), .B2(
        keyinput_g7), .ZN(n6790) );
  AOI221_X1 U7761 ( .B1(DATAI_31_), .B2(keyinput_g0), .C1(keyinput_g7), .C2(
        DATAI_24_), .A(n6790), .ZN(n6791) );
  NAND4_X1 U7762 ( .A1(n6794), .A2(n6793), .A3(n6792), .A4(n6791), .ZN(n6928)
         );
  OAI22_X1 U7763 ( .A1(STATE_REG_0__SCAN_IN), .A2(keyinput_g103), .B1(
        REIP_REG_24__SCAN_IN), .B2(keyinput_g58), .ZN(n6795) );
  AOI221_X1 U7764 ( .B1(STATE_REG_0__SCAN_IN), .B2(keyinput_g103), .C1(
        keyinput_g58), .C2(REIP_REG_24__SCAN_IN), .A(n6795), .ZN(n6820) );
  OAI22_X1 U7765 ( .A1(DATAI_13_), .A2(keyinput_g18), .B1(DATAI_6_), .B2(
        keyinput_g25), .ZN(n6796) );
  AOI221_X1 U7766 ( .B1(DATAI_13_), .B2(keyinput_g18), .C1(keyinput_g25), .C2(
        DATAI_6_), .A(n6796), .ZN(n6799) );
  OAI22_X1 U7767 ( .A1(DATAI_1_), .A2(keyinput_g30), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(keyinput_g72), .ZN(n6797) );
  AOI221_X1 U7768 ( .B1(DATAI_1_), .B2(keyinput_g30), .C1(keyinput_g72), .C2(
        ADDRESS_REG_28__SCAN_IN), .A(n6797), .ZN(n6798) );
  OAI211_X1 U7769 ( .C1(n7061), .C2(keyinput_g97), .A(n6799), .B(n6798), .ZN(
        n6800) );
  AOI21_X1 U7770 ( .B1(n7061), .B2(keyinput_g97), .A(n6800), .ZN(n6819) );
  AOI22_X1 U7771 ( .A1(ADDRESS_REG_22__SCAN_IN), .A2(keyinput_g78), .B1(
        REIP_REG_17__SCAN_IN), .B2(keyinput_g65), .ZN(n6801) );
  OAI221_X1 U7772 ( .B1(ADDRESS_REG_22__SCAN_IN), .B2(keyinput_g78), .C1(
        REIP_REG_17__SCAN_IN), .C2(keyinput_g65), .A(n6801), .ZN(n6808) );
  AOI22_X1 U7773 ( .A1(ADDRESS_REG_26__SCAN_IN), .A2(keyinput_g74), .B1(
        REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_g42), .ZN(n6802) );
  OAI221_X1 U7774 ( .B1(ADDRESS_REG_26__SCAN_IN), .B2(keyinput_g74), .C1(
        REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_g42), .A(n6802), .ZN(n6807)
         );
  AOI22_X1 U7775 ( .A1(FLUSH_REG_SCAN_IN), .A2(keyinput_g45), .B1(
        STATE_REG_1__SCAN_IN), .B2(keyinput_g102), .ZN(n6803) );
  OAI221_X1 U7776 ( .B1(FLUSH_REG_SCAN_IN), .B2(keyinput_g45), .C1(
        STATE_REG_1__SCAN_IN), .C2(keyinput_g102), .A(n6803), .ZN(n6806) );
  AOI22_X1 U7777 ( .A1(DATAI_19_), .A2(keyinput_g12), .B1(DATAI_20_), .B2(
        keyinput_g11), .ZN(n6804) );
  OAI221_X1 U7778 ( .B1(DATAI_19_), .B2(keyinput_g12), .C1(DATAI_20_), .C2(
        keyinput_g11), .A(n6804), .ZN(n6805) );
  NOR4_X1 U7779 ( .A1(n6808), .A2(n6807), .A3(n6806), .A4(n6805), .ZN(n6818)
         );
  AOI22_X1 U7780 ( .A1(ADDRESS_REG_9__SCAN_IN), .A2(keyinput_g91), .B1(
        DATAI_5_), .B2(keyinput_g26), .ZN(n6809) );
  OAI221_X1 U7781 ( .B1(ADDRESS_REG_9__SCAN_IN), .B2(keyinput_g91), .C1(
        DATAI_5_), .C2(keyinput_g26), .A(n6809), .ZN(n6816) );
  AOI22_X1 U7782 ( .A1(ADDRESS_REG_15__SCAN_IN), .A2(keyinput_g85), .B1(
        STATEBS16_REG_SCAN_IN), .B2(keyinput_g43), .ZN(n6810) );
  OAI221_X1 U7783 ( .B1(ADDRESS_REG_15__SCAN_IN), .B2(keyinput_g85), .C1(
        STATEBS16_REG_SCAN_IN), .C2(keyinput_g43), .A(n6810), .ZN(n6815) );
  AOI22_X1 U7784 ( .A1(ADDRESS_REG_18__SCAN_IN), .A2(keyinput_g82), .B1(
        REIP_REG_31__SCAN_IN), .B2(keyinput_g51), .ZN(n6811) );
  OAI221_X1 U7785 ( .B1(ADDRESS_REG_18__SCAN_IN), .B2(keyinput_g82), .C1(
        REIP_REG_31__SCAN_IN), .C2(keyinput_g51), .A(n6811), .ZN(n6814) );
  AOI22_X1 U7786 ( .A1(NA_N), .A2(keyinput_g33), .B1(W_R_N_REG_SCAN_IN), .B2(
        keyinput_g46), .ZN(n6812) );
  OAI221_X1 U7787 ( .B1(NA_N), .B2(keyinput_g33), .C1(W_R_N_REG_SCAN_IN), .C2(
        keyinput_g46), .A(n6812), .ZN(n6813) );
  NOR4_X1 U7788 ( .A1(n6816), .A2(n6815), .A3(n6814), .A4(n6813), .ZN(n6817)
         );
  NAND4_X1 U7789 ( .A1(n6820), .A2(n6819), .A3(n6818), .A4(n6817), .ZN(n6927)
         );
  AOI22_X1 U7790 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(keyinput_g108), .B1(
        BE_N_REG_1__SCAN_IN), .B2(keyinput_g69), .ZN(n6821) );
  OAI221_X1 U7791 ( .B1(DATAWIDTH_REG_4__SCAN_IN), .B2(keyinput_g108), .C1(
        BE_N_REG_1__SCAN_IN), .C2(keyinput_g69), .A(n6821), .ZN(n6829) );
  AOI22_X1 U7792 ( .A1(ADDRESS_REG_21__SCAN_IN), .A2(keyinput_g79), .B1(
        DATAI_4_), .B2(keyinput_g27), .ZN(n6822) );
  OAI221_X1 U7793 ( .B1(ADDRESS_REG_21__SCAN_IN), .B2(keyinput_g79), .C1(
        DATAI_4_), .C2(keyinput_g27), .A(n6822), .ZN(n6828) );
  AOI22_X1 U7794 ( .A1(n6824), .A2(keyinput_g83), .B1(n7097), .B2(keyinput_g53), .ZN(n6823) );
  OAI221_X1 U7795 ( .B1(n6824), .B2(keyinput_g83), .C1(n7097), .C2(
        keyinput_g53), .A(n6823), .ZN(n6827) );
  AOI22_X1 U7796 ( .A1(n7062), .A2(keyinput_g47), .B1(n7064), .B2(
        keyinput_g121), .ZN(n6825) );
  OAI221_X1 U7797 ( .B1(n7062), .B2(keyinput_g47), .C1(n7064), .C2(
        keyinput_g121), .A(n6825), .ZN(n6826) );
  NOR4_X1 U7798 ( .A1(n6829), .A2(n6828), .A3(n6827), .A4(n6826), .ZN(n6871)
         );
  AOI22_X1 U7799 ( .A1(n7007), .A2(keyinput_g73), .B1(n6831), .B2(keyinput_g71), .ZN(n6830) );
  OAI221_X1 U7800 ( .B1(n7007), .B2(keyinput_g73), .C1(n6831), .C2(
        keyinput_g71), .A(n6830), .ZN(n6841) );
  AOI22_X1 U7801 ( .A1(n6834), .A2(keyinput_g40), .B1(keyinput_g113), .B2(
        n6833), .ZN(n6832) );
  OAI221_X1 U7802 ( .B1(n6834), .B2(keyinput_g40), .C1(n6833), .C2(
        keyinput_g113), .A(n6832), .ZN(n6840) );
  AOI22_X1 U7803 ( .A1(n7033), .A2(keyinput_g23), .B1(keyinput_g90), .B2(n6836), .ZN(n6835) );
  OAI221_X1 U7804 ( .B1(n7033), .B2(keyinput_g23), .C1(n6836), .C2(
        keyinput_g90), .A(n6835), .ZN(n6839) );
  AOI22_X1 U7805 ( .A1(n7044), .A2(keyinput_g93), .B1(n5605), .B2(keyinput_g35), .ZN(n6837) );
  OAI221_X1 U7806 ( .B1(n7044), .B2(keyinput_g93), .C1(n5605), .C2(
        keyinput_g35), .A(n6837), .ZN(n6838) );
  NOR4_X1 U7807 ( .A1(n6841), .A2(n6840), .A3(n6839), .A4(n6838), .ZN(n6870)
         );
  INV_X1 U7808 ( .A(DATAI_18_), .ZN(n7048) );
  AOI22_X1 U7809 ( .A1(n7048), .A2(keyinput_g13), .B1(keyinput_g122), .B2(
        n7104), .ZN(n6842) );
  OAI221_X1 U7810 ( .B1(n7048), .B2(keyinput_g13), .C1(n7104), .C2(
        keyinput_g122), .A(n6842), .ZN(n6852) );
  INV_X1 U7811 ( .A(DATAI_25_), .ZN(n7035) );
  AOI22_X1 U7812 ( .A1(n7030), .A2(keyinput_g95), .B1(n7035), .B2(keyinput_g6), 
        .ZN(n6843) );
  OAI221_X1 U7813 ( .B1(n7030), .B2(keyinput_g95), .C1(n7035), .C2(keyinput_g6), .A(n6843), .ZN(n6851) );
  AOI22_X1 U7814 ( .A1(n6072), .A2(keyinput_g9), .B1(keyinput_g118), .B2(n6845), .ZN(n6844) );
  OAI221_X1 U7815 ( .B1(n6072), .B2(keyinput_g9), .C1(n6845), .C2(
        keyinput_g118), .A(n6844), .ZN(n6850) );
  AOI22_X1 U7816 ( .A1(n6848), .A2(keyinput_g111), .B1(n6847), .B2(
        keyinput_g31), .ZN(n6846) );
  OAI221_X1 U7817 ( .B1(n6848), .B2(keyinput_g111), .C1(n6847), .C2(
        keyinput_g31), .A(n6846), .ZN(n6849) );
  NOR4_X1 U7818 ( .A1(n6852), .A2(n6851), .A3(n6850), .A4(n6849), .ZN(n6869)
         );
  INV_X1 U7819 ( .A(DATAI_30_), .ZN(n6855) );
  AOI22_X1 U7820 ( .A1(n6855), .A2(keyinput_g1), .B1(keyinput_g106), .B2(n6854), .ZN(n6853) );
  OAI221_X1 U7821 ( .B1(n6855), .B2(keyinput_g1), .C1(n6854), .C2(
        keyinput_g106), .A(n6853), .ZN(n6867) );
  INV_X1 U7822 ( .A(DATAI_16_), .ZN(n6858) );
  AOI22_X1 U7823 ( .A1(n6858), .A2(keyinput_g15), .B1(keyinput_g119), .B2(
        n6857), .ZN(n6856) );
  OAI221_X1 U7824 ( .B1(n6858), .B2(keyinput_g15), .C1(n6857), .C2(
        keyinput_g119), .A(n6856), .ZN(n6866) );
  AOI22_X1 U7825 ( .A1(n6860), .A2(keyinput_g57), .B1(keyinput_g76), .B2(n7091), .ZN(n6859) );
  OAI221_X1 U7826 ( .B1(n6860), .B2(keyinput_g57), .C1(n7091), .C2(
        keyinput_g76), .A(n6859), .ZN(n6865) );
  AOI22_X1 U7827 ( .A1(n6863), .A2(keyinput_g50), .B1(n6862), .B2(keyinput_g28), .ZN(n6861) );
  OAI221_X1 U7828 ( .B1(n6863), .B2(keyinput_g50), .C1(n6862), .C2(
        keyinput_g28), .A(n6861), .ZN(n6864) );
  NOR4_X1 U7829 ( .A1(n6867), .A2(n6866), .A3(n6865), .A4(n6864), .ZN(n6868)
         );
  NAND4_X1 U7830 ( .A1(n6871), .A2(n6870), .A3(n6869), .A4(n6868), .ZN(n6926)
         );
  AOI22_X1 U7831 ( .A1(n6873), .A2(keyinput_g84), .B1(keyinput_g92), .B2(n7070), .ZN(n6872) );
  OAI221_X1 U7832 ( .B1(n6873), .B2(keyinput_g84), .C1(n7070), .C2(
        keyinput_g92), .A(n6872), .ZN(n6883) );
  AOI22_X1 U7833 ( .A1(n6875), .A2(keyinput_g19), .B1(keyinput_g10), .B2(n6077), .ZN(n6874) );
  OAI221_X1 U7834 ( .B1(n6875), .B2(keyinput_g19), .C1(n6077), .C2(
        keyinput_g10), .A(n6874), .ZN(n6882) );
  AOI22_X1 U7835 ( .A1(n6878), .A2(keyinput_g126), .B1(n6877), .B2(
        keyinput_g107), .ZN(n6876) );
  OAI221_X1 U7836 ( .B1(n6878), .B2(keyinput_g126), .C1(n6877), .C2(
        keyinput_g107), .A(n6876), .ZN(n6881) );
  AOI22_X1 U7837 ( .A1(n7051), .A2(keyinput_g55), .B1(keyinput_g32), .B2(n7105), .ZN(n6879) );
  OAI221_X1 U7838 ( .B1(n7051), .B2(keyinput_g55), .C1(n7105), .C2(
        keyinput_g32), .A(n6879), .ZN(n6880) );
  NOR4_X1 U7839 ( .A1(n6883), .A2(n6882), .A3(n6881), .A4(n6880), .ZN(n6924)
         );
  INV_X1 U7840 ( .A(MORE_REG_SCAN_IN), .ZN(n6885) );
  AOI22_X1 U7841 ( .A1(n7036), .A2(keyinput_g29), .B1(keyinput_g44), .B2(n6885), .ZN(n6884) );
  OAI221_X1 U7842 ( .B1(n7036), .B2(keyinput_g29), .C1(n6885), .C2(
        keyinput_g44), .A(n6884), .ZN(n6897) );
  AOI22_X1 U7843 ( .A1(n6888), .A2(keyinput_g105), .B1(n6887), .B2(
        keyinput_g77), .ZN(n6886) );
  OAI221_X1 U7844 ( .B1(n6888), .B2(keyinput_g105), .C1(n6887), .C2(
        keyinput_g77), .A(n6886), .ZN(n6896) );
  INV_X1 U7845 ( .A(HOLD), .ZN(n6891) );
  INV_X1 U7846 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n6890) );
  AOI22_X1 U7847 ( .A1(n6891), .A2(keyinput_g36), .B1(keyinput_g67), .B2(n6890), .ZN(n6889) );
  OAI221_X1 U7848 ( .B1(n6891), .B2(keyinput_g36), .C1(n6890), .C2(
        keyinput_g67), .A(n6889), .ZN(n6895) );
  INV_X1 U7849 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n7098) );
  INV_X1 U7850 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6893) );
  AOI22_X1 U7851 ( .A1(n7098), .A2(keyinput_g39), .B1(keyinput_g37), .B2(n6893), .ZN(n6892) );
  OAI221_X1 U7852 ( .B1(n7098), .B2(keyinput_g39), .C1(n6893), .C2(
        keyinput_g37), .A(n6892), .ZN(n6894) );
  NOR4_X1 U7853 ( .A1(n6897), .A2(n6896), .A3(n6895), .A4(n6894), .ZN(n6923)
         );
  INV_X1 U7854 ( .A(DATAI_23_), .ZN(n6899) );
  AOI22_X1 U7855 ( .A1(n7082), .A2(keyinput_g16), .B1(n6899), .B2(keyinput_g8), 
        .ZN(n6898) );
  OAI221_X1 U7856 ( .B1(n7082), .B2(keyinput_g16), .C1(n6899), .C2(keyinput_g8), .A(n6898), .ZN(n6908) );
  AOI22_X1 U7857 ( .A1(n7078), .A2(keyinput_g62), .B1(keyinput_g98), .B2(n7108), .ZN(n6900) );
  OAI221_X1 U7858 ( .B1(n7078), .B2(keyinput_g62), .C1(n7108), .C2(
        keyinput_g98), .A(n6900), .ZN(n6907) );
  AOI22_X1 U7859 ( .A1(n7075), .A2(keyinput_g22), .B1(keyinput_g87), .B2(n7079), .ZN(n6901) );
  OAI221_X1 U7860 ( .B1(n7075), .B2(keyinput_g22), .C1(n7079), .C2(
        keyinput_g87), .A(n6901), .ZN(n6906) );
  INV_X1 U7861 ( .A(DATAI_28_), .ZN(n6904) );
  AOI22_X1 U7862 ( .A1(n6904), .A2(keyinput_g3), .B1(keyinput_g89), .B2(n6903), 
        .ZN(n6902) );
  OAI221_X1 U7863 ( .B1(n6904), .B2(keyinput_g3), .C1(n6903), .C2(keyinput_g89), .A(n6902), .ZN(n6905) );
  NOR4_X1 U7864 ( .A1(n6908), .A2(n6907), .A3(n6906), .A4(n6905), .ZN(n6922)
         );
  AOI22_X1 U7865 ( .A1(n6301), .A2(keyinput_g14), .B1(keyinput_g96), .B2(n7047), .ZN(n6909) );
  OAI221_X1 U7866 ( .B1(n6301), .B2(keyinput_g14), .C1(n7047), .C2(
        keyinput_g96), .A(n6909), .ZN(n6920) );
  AOI22_X1 U7867 ( .A1(n6911), .A2(keyinput_g114), .B1(n7076), .B2(
        keyinput_g101), .ZN(n6910) );
  OAI221_X1 U7868 ( .B1(n6911), .B2(keyinput_g114), .C1(n7076), .C2(
        keyinput_g101), .A(n6910), .ZN(n6919) );
  AOI22_X1 U7869 ( .A1(n7020), .A2(keyinput_g20), .B1(n6913), .B2(keyinput_g52), .ZN(n6912) );
  OAI221_X1 U7870 ( .B1(n7020), .B2(keyinput_g20), .C1(n6913), .C2(
        keyinput_g52), .A(n6912), .ZN(n6918) );
  AOI22_X1 U7871 ( .A1(n6916), .A2(keyinput_g66), .B1(keyinput_g116), .B2(
        n6915), .ZN(n6914) );
  OAI221_X1 U7872 ( .B1(n6916), .B2(keyinput_g66), .C1(n6915), .C2(
        keyinput_g116), .A(n6914), .ZN(n6917) );
  NOR4_X1 U7873 ( .A1(n6920), .A2(n6919), .A3(n6918), .A4(n6917), .ZN(n6921)
         );
  NAND4_X1 U7874 ( .A1(n6924), .A2(n6923), .A3(n6922), .A4(n6921), .ZN(n6925)
         );
  NOR4_X1 U7875 ( .A1(n6928), .A2(n6927), .A3(n6926), .A4(n6925), .ZN(n7140)
         );
  AOI22_X1 U7876 ( .A1(DATAI_20_), .A2(keyinput_f11), .B1(DATAI_10_), .B2(
        keyinput_f21), .ZN(n6929) );
  OAI221_X1 U7877 ( .B1(DATAI_20_), .B2(keyinput_f11), .C1(DATAI_10_), .C2(
        keyinput_f21), .A(n6929), .ZN(n6936) );
  AOI22_X1 U7878 ( .A1(keyinput_f89), .A2(ADDRESS_REG_11__SCAN_IN), .B1(
        keyinput_f80), .B2(ADDRESS_REG_20__SCAN_IN), .ZN(n6930) );
  OAI221_X1 U7879 ( .B1(keyinput_f89), .B2(ADDRESS_REG_11__SCAN_IN), .C1(
        keyinput_f80), .C2(ADDRESS_REG_20__SCAN_IN), .A(n6930), .ZN(n6935) );
  AOI22_X1 U7880 ( .A1(DATAI_12_), .A2(keyinput_f19), .B1(REIP_REG_21__SCAN_IN), .B2(keyinput_f61), .ZN(n6931) );
  OAI221_X1 U7881 ( .B1(DATAI_12_), .B2(keyinput_f19), .C1(
        REIP_REG_21__SCAN_IN), .C2(keyinput_f61), .A(n6931), .ZN(n6934) );
  AOI22_X1 U7882 ( .A1(keyinput_f41), .A2(D_C_N_REG_SCAN_IN), .B1(
        keyinput_f112), .B2(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6932) );
  OAI221_X1 U7883 ( .B1(keyinput_f41), .B2(D_C_N_REG_SCAN_IN), .C1(
        keyinput_f112), .C2(DATAWIDTH_REG_8__SCAN_IN), .A(n6932), .ZN(n6933)
         );
  NOR4_X1 U7884 ( .A1(n6936), .A2(n6935), .A3(n6934), .A4(n6933), .ZN(n7134)
         );
  AOI22_X1 U7885 ( .A1(keyinput_f91), .A2(ADDRESS_REG_9__SCAN_IN), .B1(
        DATAI_6_), .B2(keyinput_f25), .ZN(n6937) );
  OAI221_X1 U7886 ( .B1(keyinput_f91), .B2(ADDRESS_REG_9__SCAN_IN), .C1(
        DATAI_6_), .C2(keyinput_f25), .A(n6937), .ZN(n6963) );
  OAI22_X1 U7887 ( .A1(STATEBS16_REG_SCAN_IN), .A2(keyinput_f43), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(keyinput_f77), .ZN(n6938) );
  AOI221_X1 U7888 ( .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput_f43), .C1(
        keyinput_f77), .C2(ADDRESS_REG_23__SCAN_IN), .A(n6938), .ZN(n6942) );
  AOI22_X1 U7889 ( .A1(keyinput_f48), .A2(BYTEENABLE_REG_1__SCAN_IN), .B1(
        STATE_REG_0__SCAN_IN), .B2(keyinput_f103), .ZN(n6939) );
  OAI221_X1 U7890 ( .B1(keyinput_f48), .B2(BYTEENABLE_REG_1__SCAN_IN), .C1(
        STATE_REG_0__SCAN_IN), .C2(keyinput_f103), .A(n6939), .ZN(n6940) );
  AOI21_X1 U7891 ( .B1(keyinput_f74), .B2(n6943), .A(n6940), .ZN(n6941) );
  OAI211_X1 U7892 ( .C1(keyinput_f74), .C2(n6943), .A(n6942), .B(n6941), .ZN(
        n6962) );
  OAI22_X1 U7893 ( .A1(keyinput_f83), .A2(ADDRESS_REG_17__SCAN_IN), .B1(
        keyinput_f115), .B2(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6944) );
  AOI221_X1 U7894 ( .B1(keyinput_f83), .B2(ADDRESS_REG_17__SCAN_IN), .C1(
        DATAWIDTH_REG_11__SCAN_IN), .C2(keyinput_f115), .A(n6944), .ZN(n6951)
         );
  OAI22_X1 U7895 ( .A1(DATAI_26_), .A2(keyinput_f5), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(keyinput_f71), .ZN(n6945) );
  AOI221_X1 U7896 ( .B1(DATAI_26_), .B2(keyinput_f5), .C1(keyinput_f71), .C2(
        ADDRESS_REG_29__SCAN_IN), .A(n6945), .ZN(n6950) );
  OAI22_X1 U7897 ( .A1(DATAI_3_), .A2(keyinput_f28), .B1(keyinput_f124), .B2(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n6946) );
  AOI221_X1 U7898 ( .B1(DATAI_3_), .B2(keyinput_f28), .C1(
        DATAWIDTH_REG_20__SCAN_IN), .C2(keyinput_f124), .A(n6946), .ZN(n6949)
         );
  OAI22_X1 U7899 ( .A1(READY_N), .A2(keyinput_f35), .B1(M_IO_N_REG_SCAN_IN), 
        .B2(keyinput_f40), .ZN(n6947) );
  AOI221_X1 U7900 ( .B1(READY_N), .B2(keyinput_f35), .C1(keyinput_f40), .C2(
        M_IO_N_REG_SCAN_IN), .A(n6947), .ZN(n6948) );
  NAND4_X1 U7901 ( .A1(n6951), .A2(n6950), .A3(n6949), .A4(n6948), .ZN(n6961)
         );
  OAI22_X1 U7902 ( .A1(REIP_REG_30__SCAN_IN), .A2(keyinput_f52), .B1(
        REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_f42), .ZN(n6952) );
  AOI221_X1 U7903 ( .B1(REIP_REG_30__SCAN_IN), .B2(keyinput_f52), .C1(
        keyinput_f42), .C2(REQUESTPENDING_REG_SCAN_IN), .A(n6952), .ZN(n6959)
         );
  OAI22_X1 U7904 ( .A1(REIP_REG_26__SCAN_IN), .A2(keyinput_f56), .B1(
        keyinput_f84), .B2(ADDRESS_REG_16__SCAN_IN), .ZN(n6953) );
  AOI221_X1 U7905 ( .B1(REIP_REG_26__SCAN_IN), .B2(keyinput_f56), .C1(
        ADDRESS_REG_16__SCAN_IN), .C2(keyinput_f84), .A(n6953), .ZN(n6958) );
  OAI22_X1 U7906 ( .A1(DATAI_16_), .A2(keyinput_f15), .B1(
        DATAWIDTH_REG_21__SCAN_IN), .B2(keyinput_f125), .ZN(n6954) );
  AOI221_X1 U7907 ( .B1(DATAI_16_), .B2(keyinput_f15), .C1(keyinput_f125), 
        .C2(DATAWIDTH_REG_21__SCAN_IN), .A(n6954), .ZN(n6957) );
  OAI22_X1 U7908 ( .A1(REIP_REG_17__SCAN_IN), .A2(keyinput_f65), .B1(
        DATAWIDTH_REG_6__SCAN_IN), .B2(keyinput_f110), .ZN(n6955) );
  AOI221_X1 U7909 ( .B1(REIP_REG_17__SCAN_IN), .B2(keyinput_f65), .C1(
        keyinput_f110), .C2(DATAWIDTH_REG_6__SCAN_IN), .A(n6955), .ZN(n6956)
         );
  NAND4_X1 U7910 ( .A1(n6959), .A2(n6958), .A3(n6957), .A4(n6956), .ZN(n6960)
         );
  NOR4_X1 U7911 ( .A1(n6963), .A2(n6962), .A3(n6961), .A4(n6960), .ZN(n7133)
         );
  OAI22_X1 U7912 ( .A1(DATAI_29_), .A2(keyinput_f2), .B1(
        DATAWIDTH_REG_13__SCAN_IN), .B2(keyinput_f117), .ZN(n6964) );
  AOI221_X1 U7913 ( .B1(DATAI_29_), .B2(keyinput_f2), .C1(keyinput_f117), .C2(
        DATAWIDTH_REG_13__SCAN_IN), .A(n6964), .ZN(n6971) );
  OAI22_X1 U7914 ( .A1(REIP_REG_16__SCAN_IN), .A2(keyinput_f66), .B1(
        keyinput_f85), .B2(ADDRESS_REG_15__SCAN_IN), .ZN(n6965) );
  AOI221_X1 U7915 ( .B1(REIP_REG_16__SCAN_IN), .B2(keyinput_f66), .C1(
        ADDRESS_REG_15__SCAN_IN), .C2(keyinput_f85), .A(n6965), .ZN(n6970) );
  OAI22_X1 U7916 ( .A1(keyinput_f100), .A2(ADDRESS_REG_0__SCAN_IN), .B1(
        keyinput_f94), .B2(ADDRESS_REG_6__SCAN_IN), .ZN(n6966) );
  AOI221_X1 U7917 ( .B1(keyinput_f100), .B2(ADDRESS_REG_0__SCAN_IN), .C1(
        ADDRESS_REG_6__SCAN_IN), .C2(keyinput_f94), .A(n6966), .ZN(n6969) );
  OAI22_X1 U7918 ( .A1(keyinput_f88), .A2(ADDRESS_REG_12__SCAN_IN), .B1(
        keyinput_f50), .B2(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6967) );
  AOI221_X1 U7919 ( .B1(keyinput_f88), .B2(ADDRESS_REG_12__SCAN_IN), .C1(
        BYTEENABLE_REG_3__SCAN_IN), .C2(keyinput_f50), .A(n6967), .ZN(n6968)
         );
  NAND4_X1 U7920 ( .A1(n6971), .A2(n6970), .A3(n6969), .A4(n6968), .ZN(n6999)
         );
  OAI22_X1 U7921 ( .A1(keyinput_f69), .A2(BE_N_REG_1__SCAN_IN), .B1(
        keyinput_f116), .B2(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6972) );
  AOI221_X1 U7922 ( .B1(keyinput_f69), .B2(BE_N_REG_1__SCAN_IN), .C1(
        DATAWIDTH_REG_12__SCAN_IN), .C2(keyinput_f116), .A(n6972), .ZN(n6979)
         );
  OAI22_X1 U7923 ( .A1(keyinput_f118), .A2(DATAWIDTH_REG_14__SCAN_IN), .B1(
        keyinput_f113), .B2(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6973) );
  AOI221_X1 U7924 ( .B1(keyinput_f118), .B2(DATAWIDTH_REG_14__SCAN_IN), .C1(
        DATAWIDTH_REG_9__SCAN_IN), .C2(keyinput_f113), .A(n6973), .ZN(n6978)
         );
  OAI22_X1 U7925 ( .A1(MORE_REG_SCAN_IN), .A2(keyinput_f44), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(keyinput_f72), .ZN(n6974) );
  AOI221_X1 U7926 ( .B1(MORE_REG_SCAN_IN), .B2(keyinput_f44), .C1(keyinput_f72), .C2(ADDRESS_REG_28__SCAN_IN), .A(n6974), .ZN(n6977) );
  OAI22_X1 U7927 ( .A1(keyinput_f107), .A2(DATAWIDTH_REG_3__SCAN_IN), .B1(
        keyinput_f46), .B2(W_R_N_REG_SCAN_IN), .ZN(n6975) );
  AOI221_X1 U7928 ( .B1(keyinput_f107), .B2(DATAWIDTH_REG_3__SCAN_IN), .C1(
        W_R_N_REG_SCAN_IN), .C2(keyinput_f46), .A(n6975), .ZN(n6976) );
  NAND4_X1 U7929 ( .A1(n6979), .A2(n6978), .A3(n6977), .A4(n6976), .ZN(n6998)
         );
  OAI22_X1 U7930 ( .A1(REIP_REG_19__SCAN_IN), .A2(keyinput_f63), .B1(
        keyinput_f9), .B2(DATAI_22_), .ZN(n6980) );
  AOI221_X1 U7931 ( .B1(REIP_REG_19__SCAN_IN), .B2(keyinput_f63), .C1(
        DATAI_22_), .C2(keyinput_f9), .A(n6980), .ZN(n6987) );
  OAI22_X1 U7932 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput_f60), .B1(
        keyinput_f1), .B2(DATAI_30_), .ZN(n6981) );
  AOI221_X1 U7933 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_f60), .C1(
        DATAI_30_), .C2(keyinput_f1), .A(n6981), .ZN(n6986) );
  OAI22_X1 U7934 ( .A1(REIP_REG_25__SCAN_IN), .A2(keyinput_f57), .B1(
        DATAWIDTH_REG_23__SCAN_IN), .B2(keyinput_f127), .ZN(n6982) );
  AOI221_X1 U7935 ( .B1(REIP_REG_25__SCAN_IN), .B2(keyinput_f57), .C1(
        keyinput_f127), .C2(DATAWIDTH_REG_23__SCAN_IN), .A(n6982), .ZN(n6985)
         );
  OAI22_X1 U7936 ( .A1(DATAI_28_), .A2(keyinput_f3), .B1(keyinput_f108), .B2(
        DATAWIDTH_REG_4__SCAN_IN), .ZN(n6983) );
  AOI221_X1 U7937 ( .B1(DATAI_28_), .B2(keyinput_f3), .C1(
        DATAWIDTH_REG_4__SCAN_IN), .C2(keyinput_f108), .A(n6983), .ZN(n6984)
         );
  NAND4_X1 U7938 ( .A1(n6987), .A2(n6986), .A3(n6985), .A4(n6984), .ZN(n6997)
         );
  OAI22_X1 U7939 ( .A1(DATAI_0_), .A2(keyinput_f31), .B1(keyinput_f70), .B2(
        BE_N_REG_0__SCAN_IN), .ZN(n6988) );
  AOI221_X1 U7940 ( .B1(DATAI_0_), .B2(keyinput_f31), .C1(BE_N_REG_0__SCAN_IN), 
        .C2(keyinput_f70), .A(n6988), .ZN(n6995) );
  OAI22_X1 U7941 ( .A1(DATAI_17_), .A2(keyinput_f14), .B1(keyinput_f119), .B2(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n6989) );
  AOI221_X1 U7942 ( .B1(DATAI_17_), .B2(keyinput_f14), .C1(
        DATAWIDTH_REG_15__SCAN_IN), .C2(keyinput_f119), .A(n6989), .ZN(n6994)
         );
  OAI22_X1 U7943 ( .A1(DATAI_31_), .A2(keyinput_f0), .B1(keyinput_f10), .B2(
        DATAI_21_), .ZN(n6990) );
  AOI221_X1 U7944 ( .B1(DATAI_31_), .B2(keyinput_f0), .C1(DATAI_21_), .C2(
        keyinput_f10), .A(n6990), .ZN(n6993) );
  OAI22_X1 U7945 ( .A1(READREQUEST_REG_SCAN_IN), .A2(keyinput_f37), .B1(HOLD), 
        .B2(keyinput_f36), .ZN(n6991) );
  AOI221_X1 U7946 ( .B1(READREQUEST_REG_SCAN_IN), .B2(keyinput_f37), .C1(
        keyinput_f36), .C2(HOLD), .A(n6991), .ZN(n6992) );
  NAND4_X1 U7947 ( .A1(n6995), .A2(n6994), .A3(n6993), .A4(n6992), .ZN(n6996)
         );
  NOR4_X1 U7948 ( .A1(n6999), .A2(n6998), .A3(n6997), .A4(n6996), .ZN(n7132)
         );
  AOI22_X1 U7949 ( .A1(n7002), .A2(keyinput_f99), .B1(n7001), .B2(keyinput_f18), .ZN(n7000) );
  OAI221_X1 U7950 ( .B1(n7002), .B2(keyinput_f99), .C1(n7001), .C2(
        keyinput_f18), .A(n7000), .ZN(n7130) );
  OAI22_X1 U7951 ( .A1(keyinput_f104), .A2(n7005), .B1(n7004), .B2(
        keyinput_f75), .ZN(n7003) );
  AOI221_X1 U7952 ( .B1(n7005), .B2(keyinput_f104), .C1(n7004), .C2(
        keyinput_f75), .A(n7003), .ZN(n7014) );
  INV_X1 U7953 ( .A(DATAI_24_), .ZN(n7008) );
  OAI22_X1 U7954 ( .A1(n7008), .A2(keyinput_f7), .B1(n7007), .B2(keyinput_f73), 
        .ZN(n7006) );
  AOI221_X1 U7955 ( .B1(n7008), .B2(keyinput_f7), .C1(keyinput_f73), .C2(n7007), .A(n7006), .ZN(n7013) );
  OAI22_X1 U7956 ( .A1(n7011), .A2(keyinput_f86), .B1(n7010), .B2(keyinput_f79), .ZN(n7009) );
  AOI221_X1 U7957 ( .B1(n7011), .B2(keyinput_f86), .C1(keyinput_f79), .C2(
        n7010), .A(n7009), .ZN(n7012) );
  NAND3_X1 U7958 ( .A1(n7014), .A2(n7013), .A3(n7012), .ZN(n7129) );
  AOI22_X1 U7959 ( .A1(keyinput_f120), .A2(DATAWIDTH_REG_16__SCAN_IN), .B1(
        keyinput_f126), .B2(DATAWIDTH_REG_22__SCAN_IN), .ZN(n7015) );
  OAI221_X1 U7960 ( .B1(keyinput_f120), .B2(DATAWIDTH_REG_16__SCAN_IN), .C1(
        keyinput_f126), .C2(DATAWIDTH_REG_22__SCAN_IN), .A(n7015), .ZN(n7024)
         );
  AOI22_X1 U7961 ( .A1(DATAI_23_), .A2(keyinput_f8), .B1(STATE_REG_1__SCAN_IN), 
        .B2(keyinput_f102), .ZN(n7016) );
  OAI221_X1 U7962 ( .B1(DATAI_23_), .B2(keyinput_f8), .C1(STATE_REG_1__SCAN_IN), .C2(keyinput_f102), .A(n7016), .ZN(n7023) );
  AOI22_X1 U7963 ( .A1(keyinput_f114), .A2(DATAWIDTH_REG_10__SCAN_IN), .B1(
        keyinput_f90), .B2(ADDRESS_REG_10__SCAN_IN), .ZN(n7017) );
  OAI221_X1 U7964 ( .B1(keyinput_f114), .B2(DATAWIDTH_REG_10__SCAN_IN), .C1(
        keyinput_f90), .C2(ADDRESS_REG_10__SCAN_IN), .A(n7017), .ZN(n7022) );
  AOI22_X1 U7965 ( .A1(n7020), .A2(keyinput_f20), .B1(n7019), .B2(keyinput_f58), .ZN(n7018) );
  OAI221_X1 U7966 ( .B1(n7020), .B2(keyinput_f20), .C1(n7019), .C2(
        keyinput_f58), .A(n7018), .ZN(n7021) );
  NOR4_X1 U7967 ( .A1(n7024), .A2(n7023), .A3(n7022), .A4(n7021), .ZN(n7059)
         );
  OAI22_X1 U7968 ( .A1(keyinput_f123), .A2(n7027), .B1(n7026), .B2(
        keyinput_f82), .ZN(n7025) );
  AOI221_X1 U7969 ( .B1(n7027), .B2(keyinput_f123), .C1(n7026), .C2(
        keyinput_f82), .A(n7025), .ZN(n7058) );
  AOI22_X1 U7970 ( .A1(n7030), .A2(keyinput_f95), .B1(n7029), .B2(keyinput_f30), .ZN(n7028) );
  OAI221_X1 U7971 ( .B1(n7030), .B2(keyinput_f95), .C1(n7029), .C2(
        keyinput_f30), .A(n7028), .ZN(n7039) );
  AOI22_X1 U7972 ( .A1(n7033), .A2(keyinput_f23), .B1(keyinput_f38), .B2(n7032), .ZN(n7031) );
  OAI221_X1 U7973 ( .B1(n7033), .B2(keyinput_f23), .C1(n7032), .C2(
        keyinput_f38), .A(n7031), .ZN(n7038) );
  AOI22_X1 U7974 ( .A1(n7036), .A2(keyinput_f29), .B1(n7035), .B2(keyinput_f6), 
        .ZN(n7034) );
  OAI221_X1 U7975 ( .B1(n7036), .B2(keyinput_f29), .C1(n7035), .C2(keyinput_f6), .A(n7034), .ZN(n7037) );
  NOR3_X1 U7976 ( .A1(n7039), .A2(n7038), .A3(n7037), .ZN(n7057) );
  INV_X1 U7977 ( .A(keyinput_f111), .ZN(n7041) );
  AOI22_X1 U7978 ( .A1(n7042), .A2(keyinput_f24), .B1(DATAWIDTH_REG_7__SCAN_IN), .B2(n7041), .ZN(n7040) );
  OAI221_X1 U7979 ( .B1(n7042), .B2(keyinput_f24), .C1(n7041), .C2(
        DATAWIDTH_REG_7__SCAN_IN), .A(n7040), .ZN(n7055) );
  AOI22_X1 U7980 ( .A1(n7045), .A2(keyinput_f64), .B1(keyinput_f93), .B2(n7044), .ZN(n7043) );
  OAI221_X1 U7981 ( .B1(n7045), .B2(keyinput_f64), .C1(n7044), .C2(
        keyinput_f93), .A(n7043), .ZN(n7054) );
  AOI22_X1 U7982 ( .A1(n7048), .A2(keyinput_f13), .B1(keyinput_f96), .B2(n7047), .ZN(n7046) );
  OAI221_X1 U7983 ( .B1(n7048), .B2(keyinput_f13), .C1(n7047), .C2(
        keyinput_f96), .A(n7046), .ZN(n7053) );
  AOI22_X1 U7984 ( .A1(n7051), .A2(keyinput_f55), .B1(n7050), .B2(keyinput_f51), .ZN(n7049) );
  OAI221_X1 U7985 ( .B1(n7051), .B2(keyinput_f55), .C1(n7050), .C2(
        keyinput_f51), .A(n7049), .ZN(n7052) );
  NOR4_X1 U7986 ( .A1(n7055), .A2(n7054), .A3(n7053), .A4(n7052), .ZN(n7056)
         );
  NAND4_X1 U7987 ( .A1(n7059), .A2(n7058), .A3(n7057), .A4(n7056), .ZN(n7128)
         );
  OAI22_X1 U7988 ( .A1(keyinput_f47), .A2(n7062), .B1(n7061), .B2(keyinput_f97), .ZN(n7060) );
  AOI221_X1 U7989 ( .B1(n7062), .B2(keyinput_f47), .C1(n7061), .C2(
        keyinput_f97), .A(n7060), .ZN(n7126) );
  AOI22_X1 U7990 ( .A1(n3883), .A2(keyinput_f59), .B1(keyinput_f121), .B2(
        n7064), .ZN(n7063) );
  OAI221_X1 U7991 ( .B1(n3883), .B2(keyinput_f59), .C1(n7064), .C2(
        keyinput_f121), .A(n7063), .ZN(n7073) );
  INV_X1 U7992 ( .A(keyinput_f49), .ZN(n7066) );
  AOI22_X1 U7993 ( .A1(n7067), .A2(keyinput_f54), .B1(
        BYTEENABLE_REG_2__SCAN_IN), .B2(n7066), .ZN(n7065) );
  OAI221_X1 U7994 ( .B1(n7067), .B2(keyinput_f54), .C1(n7066), .C2(
        BYTEENABLE_REG_2__SCAN_IN), .A(n7065), .ZN(n7072) );
  INV_X1 U7995 ( .A(DATAI_27_), .ZN(n7069) );
  AOI22_X1 U7996 ( .A1(n7070), .A2(keyinput_f92), .B1(n7069), .B2(keyinput_f4), 
        .ZN(n7068) );
  OAI221_X1 U7997 ( .B1(n7070), .B2(keyinput_f92), .C1(n7069), .C2(keyinput_f4), .A(n7068), .ZN(n7071) );
  NOR3_X1 U7998 ( .A1(n7073), .A2(n7072), .A3(n7071), .ZN(n7125) );
  AOI22_X1 U7999 ( .A1(n7076), .A2(keyinput_f101), .B1(keyinput_f22), .B2(
        n7075), .ZN(n7074) );
  OAI221_X1 U8000 ( .B1(n7076), .B2(keyinput_f101), .C1(n7075), .C2(
        keyinput_f22), .A(n7074), .ZN(n7089) );
  AOI22_X1 U8001 ( .A1(n7079), .A2(keyinput_f87), .B1(n7078), .B2(keyinput_f62), .ZN(n7077) );
  OAI221_X1 U8002 ( .B1(n7079), .B2(keyinput_f87), .C1(n7078), .C2(
        keyinput_f62), .A(n7077), .ZN(n7088) );
  AOI22_X1 U8003 ( .A1(n7082), .A2(keyinput_f16), .B1(keyinput_f109), .B2(
        n7081), .ZN(n7080) );
  OAI221_X1 U8004 ( .B1(n7082), .B2(keyinput_f16), .C1(n7081), .C2(
        keyinput_f109), .A(n7080), .ZN(n7087) );
  INV_X1 U8005 ( .A(BS16_N), .ZN(n7084) );
  AOI22_X1 U8006 ( .A1(n7085), .A2(keyinput_f26), .B1(keyinput_f34), .B2(n7084), .ZN(n7083) );
  OAI221_X1 U8007 ( .B1(n7085), .B2(keyinput_f26), .C1(n7084), .C2(
        keyinput_f34), .A(n7083), .ZN(n7086) );
  NOR4_X1 U8008 ( .A1(n7089), .A2(n7088), .A3(n7087), .A4(n7086), .ZN(n7124)
         );
  INV_X1 U8009 ( .A(DATAI_19_), .ZN(n7092) );
  AOI22_X1 U8010 ( .A1(n7092), .A2(keyinput_f12), .B1(keyinput_f76), .B2(n7091), .ZN(n7090) );
  OAI221_X1 U8011 ( .B1(n7092), .B2(keyinput_f12), .C1(n7091), .C2(
        keyinput_f76), .A(n7090), .ZN(n7122) );
  AOI22_X1 U8012 ( .A1(n7095), .A2(keyinput_f27), .B1(keyinput_f45), .B2(n7094), .ZN(n7093) );
  OAI221_X1 U8013 ( .B1(n7095), .B2(keyinput_f27), .C1(n7094), .C2(
        keyinput_f45), .A(n7093), .ZN(n7121) );
  INV_X1 U8014 ( .A(DATAI_14_), .ZN(n7102) );
  XOR2_X1 U8015 ( .A(keyinput_f67), .B(BE_N_REG_3__SCAN_IN), .Z(n7100) );
  AOI22_X1 U8016 ( .A1(n7098), .A2(keyinput_f39), .B1(n7097), .B2(keyinput_f53), .ZN(n7096) );
  OAI221_X1 U8017 ( .B1(n7098), .B2(keyinput_f39), .C1(n7097), .C2(
        keyinput_f53), .A(n7096), .ZN(n7099) );
  AOI211_X1 U8018 ( .C1(n7102), .C2(keyinput_f17), .A(n7100), .B(n7099), .ZN(
        n7101) );
  OAI21_X1 U8019 ( .B1(n7102), .B2(keyinput_f17), .A(n7101), .ZN(n7120) );
  OAI22_X1 U8020 ( .A1(n7105), .A2(keyinput_f32), .B1(n7104), .B2(
        keyinput_f122), .ZN(n7103) );
  AOI221_X1 U8021 ( .B1(n7105), .B2(keyinput_f32), .C1(keyinput_f122), .C2(
        n7104), .A(n7103), .ZN(n7118) );
  INV_X1 U8022 ( .A(keyinput_f106), .ZN(n7107) );
  OAI22_X1 U8023 ( .A1(n7108), .A2(keyinput_f98), .B1(n7107), .B2(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n7106) );
  AOI221_X1 U8024 ( .B1(n7108), .B2(keyinput_f98), .C1(
        DATAWIDTH_REG_2__SCAN_IN), .C2(n7107), .A(n7106), .ZN(n7117) );
  OAI22_X1 U8025 ( .A1(n7111), .A2(keyinput_f78), .B1(n7110), .B2(keyinput_f68), .ZN(n7109) );
  AOI221_X1 U8026 ( .B1(n7111), .B2(keyinput_f78), .C1(keyinput_f68), .C2(
        n7110), .A(n7109), .ZN(n7116) );
  INV_X1 U8027 ( .A(keyinput_f105), .ZN(n7113) );
  OAI22_X1 U8028 ( .A1(keyinput_f33), .A2(n7114), .B1(n7113), .B2(
        DATAWIDTH_REG_1__SCAN_IN), .ZN(n7112) );
  AOI221_X1 U8029 ( .B1(n7114), .B2(keyinput_f33), .C1(n7113), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(n7112), .ZN(n7115) );
  NAND4_X1 U8030 ( .A1(n7118), .A2(n7117), .A3(n7116), .A4(n7115), .ZN(n7119)
         );
  NOR4_X1 U8031 ( .A1(n7122), .A2(n7121), .A3(n7120), .A4(n7119), .ZN(n7123)
         );
  NAND4_X1 U8032 ( .A1(n7126), .A2(n7125), .A3(n7124), .A4(n7123), .ZN(n7127)
         );
  NOR4_X1 U8033 ( .A1(n7130), .A2(n7129), .A3(n7128), .A4(n7127), .ZN(n7131)
         );
  NAND4_X1 U8034 ( .A1(n7134), .A2(n7133), .A3(n7132), .A4(n7131), .ZN(n7136)
         );
  AOI21_X1 U8035 ( .B1(keyinput_f81), .B2(n7136), .A(keyinput_g81), .ZN(n7138)
         );
  INV_X1 U8036 ( .A(keyinput_f81), .ZN(n7135) );
  AOI21_X1 U8037 ( .B1(n7136), .B2(n7135), .A(ADDRESS_REG_19__SCAN_IN), .ZN(
        n7137) );
  AOI22_X1 U8038 ( .A1(ADDRESS_REG_19__SCAN_IN), .A2(n7138), .B1(keyinput_g81), 
        .B2(n7137), .ZN(n7139) );
  AOI21_X1 U8039 ( .B1(n7141), .B2(n7140), .A(n7139), .ZN(n7144) );
  AOI22_X1 U8040 ( .A1(n6713), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n7142), .ZN(n7143) );
  XNOR2_X1 U8041 ( .A(n7144), .B(n7143), .ZN(U3445) );
  AND2_X1 U4796 ( .A1(n6133), .A2(n6058), .ZN(n5684) );
  CLKBUF_X1 U3604 ( .A(n3546), .Z(n3547) );
  CLKBUF_X1 U3607 ( .A(n3399), .Z(n4492) );
  CLKBUF_X1 U3621 ( .A(n3925), .Z(n6616) );
  CLKBUF_X1 U3627 ( .A(n4397), .Z(n4430) );
  CLKBUF_X1 U3931 ( .A(n6743), .Z(n6638) );
  OR2_X1 U3940 ( .A1(n5185), .A2(n4727), .ZN(n7145) );
endmodule

