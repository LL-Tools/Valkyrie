

module b17_C_SARLock_k_128_3 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192;

  MUX2_X1 U11191 ( .A(n14822), .B(n14821), .S(n15138), .Z(n14824) );
  NAND2_X1 U11192 ( .A1(n15570), .A2(n15566), .ZN(n16332) );
  NAND2_X1 U11194 ( .A1(n15568), .A2(n15565), .ZN(n15570) );
  OR2_X1 U11195 ( .A1(n15380), .A2(n15381), .ZN(n15383) );
  AOI21_X1 U11196 ( .B1(n12071), .B2(n12070), .A(n15138), .ZN(n10119) );
  OR2_X1 U11198 ( .A1(n11110), .A2(n11114), .ZN(n19585) );
  OR2_X1 U11199 ( .A1(n11096), .A2(n15847), .ZN(n19757) );
  OR2_X1 U11200 ( .A1(n11102), .A2(n13588), .ZN(n19829) );
  OR2_X1 U11201 ( .A1(n11096), .A2(n13588), .ZN(n15888) );
  INV_X1 U11202 ( .A(n11065), .ZN(n11433) );
  BUF_X2 U11204 ( .A(n13466), .Z(n17284) );
  BUF_X2 U11205 ( .A(n12749), .Z(n17279) );
  INV_X2 U11206 ( .A(n17019), .ZN(n9754) );
  NOR2_X2 U11207 ( .A1(n18778), .A2(n12662), .ZN(n12750) );
  AND2_X1 U11208 ( .A1(n10773), .A2(n10456), .ZN(n10897) );
  AND2_X1 U11209 ( .A1(n10636), .A2(n10456), .ZN(n10986) );
  AND2_X1 U11210 ( .A1(n10773), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10499) );
  AND2_X1 U11211 ( .A1(n10804), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10617) );
  AND2_X1 U11212 ( .A1(n9765), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10896) );
  CLKBUF_X2 U11214 ( .A(n11939), .Z(n9776) );
  AND2_X1 U11215 ( .A1(n11811), .A2(n12089), .ZN(n10015) );
  NAND2_X1 U11216 ( .A1(n15876), .A2(n10331), .ZN(n11431) );
  AND2_X1 U11217 ( .A1(n11663), .A2(n13681), .ZN(n11888) );
  NAND2_X2 U11218 ( .A1(n10259), .A2(n10258), .ZN(n11457) );
  AND2_X1 U11219 ( .A1(n11664), .A2(n13700), .ZN(n11847) );
  AND2_X1 U11220 ( .A1(n11663), .A2(n11664), .ZN(n11939) );
  AND2_X1 U11221 ( .A1(n11665), .A2(n11662), .ZN(n11830) );
  INV_X2 U11222 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11802) );
  INV_X1 U11223 ( .A(n10293), .ZN(n9751) );
  INV_X1 U11224 ( .A(n10293), .ZN(n10318) );
  NAND2_X2 U11225 ( .A1(n13833), .A2(n10237), .ZN(n10293) );
  INV_X1 U11226 ( .A(n10293), .ZN(n10797) );
  AND2_X1 U11227 ( .A1(n13209), .A2(n14360), .ZN(n11807) );
  AND2_X1 U11228 ( .A1(n11661), .A2(n13424), .ZN(n11836) );
  OR2_X1 U11229 ( .A1(n11110), .A2(n11108), .ZN(n15866) );
  INV_X1 U11230 ( .A(n15900), .ZN(n13504) );
  OR2_X1 U11231 ( .A1(n12667), .A2(n12665), .ZN(n17119) );
  AND2_X1 U11232 ( .A1(n11791), .A2(n11807), .ZN(n9929) );
  INV_X1 U11233 ( .A(n11547), .ZN(n11538) );
  BUF_X1 U11234 ( .A(n10910), .Z(n9747) );
  OR2_X1 U11235 ( .A1(n11110), .A2(n11109), .ZN(n19556) );
  INV_X1 U11237 ( .A(n13547), .ZN(n11788) );
  OR2_X1 U11239 ( .A1(n19010), .A2(n10058), .ZN(n10056) );
  AND2_X1 U11240 ( .A1(n10071), .A2(n19173), .ZN(n19011) );
  AND2_X1 U11241 ( .A1(n10363), .A2(n10370), .ZN(n11466) );
  INV_X1 U11242 ( .A(n17029), .ZN(n10031) );
  AND3_X1 U11243 ( .A1(n10214), .A2(n12713), .A3(n10215), .ZN(n12757) );
  INV_X4 U11244 ( .A(n17218), .ZN(n17302) );
  XNOR2_X1 U11245 ( .A(n14809), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14966) );
  INV_X1 U11248 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n20119) );
  NAND2_X1 U11249 ( .A1(n17961), .A2(n17922), .ZN(n17956) );
  AND2_X1 U11250 ( .A1(n13565), .A2(n13564), .ZN(n20227) );
  AOI211_X1 U11251 ( .C1(n14491), .C2(n19382), .A(n14486), .B(n14485), .ZN(
        n14487) );
  NOR2_X1 U11252 ( .A1(n12723), .A2(n12722), .ZN(n12919) );
  INV_X1 U11253 ( .A(n11888), .ZN(n9757) );
  XOR2_X1 U11254 ( .A(n15547), .B(n15749), .Z(n9746) );
  NAND2_X2 U11255 ( .A1(n9928), .A2(n9938), .ZN(n14883) );
  NAND2_X1 U11256 ( .A1(n9908), .A2(n9907), .ZN(n10910) );
  INV_X2 U11257 ( .A(n11461), .ZN(n10345) );
  NOR2_X2 U11258 ( .A1(n13573), .A2(n13574), .ZN(n13891) );
  AND2_X2 U11259 ( .A1(n10328), .A2(n10316), .ZN(n9763) );
  NAND2_X2 U11260 ( .A1(n10756), .A2(n10755), .ZN(n10142) );
  NAND2_X2 U11261 ( .A1(n15266), .A2(n10730), .ZN(n10756) );
  NAND2_X2 U11263 ( .A1(n10383), .A2(n10382), .ZN(n10385) );
  XNOR2_X2 U11264 ( .A(n11960), .B(n13789), .ZN(n13784) );
  NAND2_X2 U11265 ( .A1(n13709), .A2(n11930), .ZN(n11960) );
  INV_X1 U11266 ( .A(n17119), .ZN(n9749) );
  INV_X2 U11267 ( .A(n17119), .ZN(n17301) );
  OAI21_X2 U11268 ( .B1(n15686), .B2(n15684), .A(n15682), .ZN(n15492) );
  NAND4_X4 U11269 ( .A1(n11733), .A2(n11732), .A3(n11731), .A4(n11730), .ZN(
        n12089) );
  AND4_X2 U11270 ( .A1(n11729), .A2(n11728), .A3(n11727), .A4(n11726), .ZN(
        n11730) );
  NAND2_X2 U11271 ( .A1(n10353), .A2(n11457), .ZN(n10327) );
  NAND2_X1 U11272 ( .A1(n10447), .A2(n11457), .ZN(n10337) );
  NAND2_X2 U11273 ( .A1(n10292), .A2(n10291), .ZN(n10317) );
  AND2_X2 U11274 ( .A1(n13156), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13146) );
  INV_X4 U11275 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10237) );
  NOR2_X2 U11276 ( .A1(n18756), .A2(n18774), .ZN(n18789) );
  INV_X1 U11277 ( .A(n10293), .ZN(n9750) );
  INV_X1 U11278 ( .A(n10797), .ZN(n9752) );
  INV_X1 U11279 ( .A(n10797), .ZN(n9753) );
  BUF_X4 U11280 ( .A(n11083), .Z(n15847) );
  AND2_X1 U11281 ( .A1(n11101), .A2(n19200), .ZN(n9985) );
  XNOR2_X2 U11282 ( .A(n11240), .B(n11542), .ZN(n16371) );
  NAND2_X2 U11283 ( .A1(n11219), .A2(n19170), .ZN(n11240) );
  NAND2_X2 U11284 ( .A1(n10203), .A2(n9833), .ZN(n15579) );
  AOI21_X1 U11285 ( .B1(n14468), .B2(n10196), .A(n10194), .ZN(n10193) );
  NAND2_X1 U11286 ( .A1(n15274), .A2(n10710), .ZN(n10727) );
  NOR2_X1 U11287 ( .A1(n14938), .A2(n9931), .ZN(n14920) );
  AND2_X1 U11288 ( .A1(n14906), .A2(n15109), .ZN(n12061) );
  NAND2_X1 U11289 ( .A1(n11491), .A2(n11164), .ZN(n11277) );
  INV_X2 U11290 ( .A(n17800), .ZN(n17823) );
  OR2_X1 U11291 ( .A1(n17747), .A2(n17872), .ZN(n12788) );
  OR2_X1 U11292 ( .A1(n11338), .A2(n11317), .ZN(n11328) );
  NOR2_X2 U11293 ( .A1(n18959), .A2(n9796), .ZN(n17953) );
  NOR2_X2 U11294 ( .A1(n11309), .A2(n9760), .ZN(n9759) );
  INV_X4 U11295 ( .A(n18787), .ZN(n18755) );
  OR2_X1 U11296 ( .A1(n9779), .A2(n9755), .ZN(n9778) );
  OR2_X1 U11297 ( .A1(n9893), .A2(n11394), .ZN(n11375) );
  AOI21_X1 U11298 ( .B1(n13438), .B2(n11448), .A(n9755), .ZN(n19270) );
  NOR2_X1 U11300 ( .A1(n13102), .A2(n11805), .ZN(n11794) );
  AND2_X1 U11301 ( .A1(n13006), .A2(n12139), .ZN(n13102) );
  CLKBUF_X1 U11303 ( .A(n13083), .Z(n9772) );
  AOI21_X1 U11304 ( .B1(n13099), .B2(n13411), .A(n11780), .ZN(n11781) );
  NAND2_X2 U11305 ( .A1(n14042), .A2(n13547), .ZN(n14540) );
  CLKBUF_X2 U11306 ( .A(n10870), .Z(n11434) );
  NAND2_X1 U11307 ( .A1(n19442), .A2(n10338), .ZN(n10928) );
  CLKBUF_X2 U11308 ( .A(n11915), .Z(n14042) );
  INV_X2 U11309 ( .A(n10353), .ZN(n10338) );
  INV_X1 U11310 ( .A(n11457), .ZN(n19452) );
  OR2_X1 U11311 ( .A1(n11679), .A2(n11678), .ZN(n13917) );
  CLKBUF_X2 U11312 ( .A(n10572), .Z(n10984) );
  AND4_X1 U11313 ( .A1(n10246), .A2(n10245), .A3(n10244), .A4(n10243), .ZN(
        n10247) );
  AND4_X1 U11314 ( .A1(n10241), .A2(n10240), .A3(n10239), .A4(n10238), .ZN(
        n10242) );
  INV_X2 U11315 ( .A(n9757), .ZN(n9777) );
  INV_X1 U11316 ( .A(n20123), .ZN(n9755) );
  CLKBUF_X2 U11317 ( .A(n11847), .Z(n12627) );
  BUF_X2 U11318 ( .A(n11860), .Z(n12498) );
  CLKBUF_X2 U11319 ( .A(n12708), .Z(n17192) );
  CLKBUF_X2 U11321 ( .A(n11830), .Z(n12447) );
  NOR2_X1 U11322 ( .A1(n15538), .A2(n15537), .ZN(n15753) );
  AOI211_X1 U11323 ( .C1(n14456), .C2(n16378), .A(n14455), .B(n14454), .ZN(
        n14457) );
  OAI21_X1 U11324 ( .B1(n14412), .B2(n19385), .A(n10080), .ZN(n10079) );
  NOR2_X1 U11325 ( .A1(n15513), .A2(n15717), .ZN(n15512) );
  XNOR2_X1 U11326 ( .A(n11532), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14456) );
  OAI21_X1 U11327 ( .B1(n15451), .B2(n15454), .A(n10225), .ZN(n11402) );
  AOI21_X1 U11328 ( .B1(n10201), .B2(n10199), .A(n14390), .ZN(n15535) );
  AOI22_X1 U11329 ( .A1(n16335), .A2(n16379), .B1(n19067), .B2(n19382), .ZN(
        n16336) );
  AOI21_X1 U11330 ( .B1(n15547), .B2(n14431), .A(n14430), .ZN(n14473) );
  NAND2_X1 U11331 ( .A1(n15525), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15513) );
  XNOR2_X1 U11332 ( .A(n14824), .B(n14823), .ZN(n14983) );
  INV_X1 U11333 ( .A(n10138), .ZN(n10143) );
  OR2_X1 U11334 ( .A1(n14478), .A2(n14476), .ZN(n14474) );
  OR2_X1 U11335 ( .A1(n15564), .A2(n15748), .ZN(n15547) );
  NAND2_X1 U11336 ( .A1(n9895), .A2(n9894), .ZN(n14478) );
  OR2_X1 U11337 ( .A1(n14815), .A2(n14730), .ZN(n9956) );
  AOI211_X1 U11338 ( .C1(n16141), .C2(n14849), .A(n14848), .B(n14847), .ZN(
        n14850) );
  AOI21_X1 U11339 ( .B1(n14591), .B2(n14603), .A(n14590), .ZN(n14829) );
  NAND2_X1 U11340 ( .A1(n15784), .A2(n9861), .ZN(n15580) );
  NAND2_X1 U11341 ( .A1(n15600), .A2(n11527), .ZN(n15784) );
  XNOR2_X1 U11342 ( .A(n10727), .B(n10728), .ZN(n15268) );
  OR2_X1 U11343 ( .A1(n14851), .A2(n21064), .ZN(n14861) );
  AND2_X1 U11344 ( .A1(n10076), .A2(n10075), .ZN(n10074) );
  CLKBUF_X1 U11346 ( .A(n14644), .Z(n14696) );
  OR2_X1 U11347 ( .A1(n15246), .A2(n15245), .ZN(n10229) );
  NAND2_X1 U11348 ( .A1(n15615), .A2(n11519), .ZN(n15808) );
  AOI21_X1 U11349 ( .B1(n14491), .B2(n19402), .A(n14490), .ZN(n10011) );
  NAND2_X1 U11350 ( .A1(n15616), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15615) );
  NOR2_X1 U11351 ( .A1(n11382), .A2(n9996), .ZN(n9995) );
  OR2_X1 U11352 ( .A1(n13288), .A2(n13289), .ZN(n15241) );
  OAI21_X1 U11353 ( .B1(n11515), .B2(n10231), .A(n11511), .ZN(n9865) );
  NAND2_X1 U11354 ( .A1(n12052), .A2(n12051), .ZN(n14292) );
  NAND2_X1 U11355 ( .A1(n10147), .A2(n10151), .ZN(n10150) );
  NAND2_X1 U11356 ( .A1(n15262), .A2(n15263), .ZN(n13288) );
  INV_X1 U11357 ( .A(n11527), .ZN(n10185) );
  OR2_X1 U11358 ( .A1(n14224), .A2(n12265), .ZN(n14275) );
  AOI21_X1 U11359 ( .B1(n9991), .B2(n15577), .A(n9800), .ZN(n9989) );
  INV_X1 U11360 ( .A(n11282), .ZN(n11517) );
  AND2_X1 U11361 ( .A1(n9925), .A2(n10112), .ZN(n9924) );
  AND2_X1 U11362 ( .A1(n11377), .A2(n11376), .ZN(n16274) );
  XNOR2_X1 U11363 ( .A(n11525), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15601) );
  OR2_X1 U11364 ( .A1(n11520), .A2(n11322), .ZN(n11525) );
  AND2_X1 U11365 ( .A1(n10223), .A2(n11375), .ZN(n11377) );
  NAND2_X1 U11366 ( .A1(n11520), .A2(n10191), .ZN(n11282) );
  NOR2_X1 U11367 ( .A1(n11365), .A2(n9992), .ZN(n9991) );
  OR2_X1 U11368 ( .A1(n15285), .A2(n15286), .ZN(n10230) );
  NAND2_X1 U11369 ( .A1(n10192), .A2(n11275), .ZN(n11520) );
  AOI21_X1 U11370 ( .B1(n14907), .B2(n12061), .A(n12059), .ZN(n15085) );
  NAND2_X1 U11371 ( .A1(n9900), .A2(n9897), .ZN(n14001) );
  NOR2_X1 U11372 ( .A1(n10115), .A2(n10111), .ZN(n10110) );
  AND2_X1 U11373 ( .A1(n11607), .A2(n10081), .ZN(n15301) );
  NOR2_X2 U11374 ( .A1(n16294), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n16293) );
  AND2_X1 U11375 ( .A1(n15519), .A2(n15521), .ZN(n14516) );
  AND3_X1 U11376 ( .A1(n17667), .A2(n17658), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17654) );
  NAND2_X1 U11377 ( .A1(n13772), .A2(n13771), .ZN(n13823) );
  NAND2_X1 U11378 ( .A1(n11367), .A2(n9890), .ZN(n16294) );
  NAND2_X1 U11379 ( .A1(n13785), .A2(n11961), .ZN(n11980) );
  NAND2_X1 U11380 ( .A1(n12191), .A2(n12190), .ZN(n13817) );
  INV_X1 U11381 ( .A(n13244), .ZN(n11050) );
  NAND2_X1 U11382 ( .A1(n11368), .A2(n11375), .ZN(n11367) );
  AND2_X1 U11383 ( .A1(n14155), .A2(n14156), .ZN(n14462) );
  AND2_X1 U11384 ( .A1(n13944), .A2(n9816), .ZN(n14155) );
  AND2_X1 U11385 ( .A1(n19047), .A2(n11396), .ZN(n11333) );
  XNOR2_X1 U11386 ( .A(n12036), .B(n12035), .ZN(n12240) );
  AND2_X1 U11387 ( .A1(n12183), .A2(n12182), .ZN(n13824) );
  OR2_X1 U11388 ( .A1(n12184), .A2(n12338), .ZN(n12191) );
  OAI21_X1 U11389 ( .B1(n20820), .B2(n12338), .A(n12175), .ZN(n13771) );
  AND2_X1 U11390 ( .A1(n13779), .A2(n13942), .ZN(n13944) );
  AND2_X1 U11391 ( .A1(n19070), .A2(n11396), .ZN(n11359) );
  NOR2_X1 U11392 ( .A1(n11171), .A2(n11121), .ZN(n11125) );
  NAND2_X1 U11393 ( .A1(n10016), .A2(n12022), .ZN(n12036) );
  NAND2_X1 U11394 ( .A1(n11999), .A2(n11956), .ZN(n20820) );
  OR2_X1 U11395 ( .A1(n11348), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11337) );
  INV_X1 U11396 ( .A(n14437), .ZN(n11040) );
  INV_X1 U11397 ( .A(n12024), .ZN(n10016) );
  NOR2_X1 U11398 ( .A1(n19790), .A2(n11148), .ZN(n11149) );
  NOR2_X1 U11399 ( .A1(n19790), .A2(n11123), .ZN(n11124) );
  AND2_X1 U11400 ( .A1(n10446), .A2(n13883), .ZN(n13568) );
  OR2_X1 U11401 ( .A1(n19699), .A2(n11103), .ZN(n11104) );
  OR2_X1 U11402 ( .A1(n11110), .A2(n11113), .ZN(n11184) );
  INV_X2 U11403 ( .A(n13793), .ZN(n20281) );
  OR2_X1 U11404 ( .A1(n16396), .A2(n9844), .ZN(n14437) );
  NAND2_X1 U11405 ( .A1(n11954), .A2(n9941), .ZN(n12024) );
  OAI21_X1 U11406 ( .B1(n13731), .B2(n12338), .A(n12145), .ZN(n12146) );
  NAND2_X1 U11407 ( .A1(n13584), .A2(n10421), .ZN(n13569) );
  NAND2_X1 U11408 ( .A1(n11954), .A2(n11953), .ZN(n11999) );
  NAND2_X1 U11409 ( .A1(n9985), .A2(n9984), .ZN(n11177) );
  NAND3_X1 U11410 ( .A1(n9985), .A2(n13588), .A3(n11087), .ZN(n19731) );
  AOI21_X1 U11411 ( .B1(n17802), .B2(n12783), .A(n17804), .ZN(n17759) );
  INV_X1 U11412 ( .A(n9759), .ZN(n11351) );
  AND2_X1 U11413 ( .A1(n13598), .A2(n10417), .ZN(n13585) );
  AND2_X1 U11414 ( .A1(n11953), .A2(n11994), .ZN(n9941) );
  NAND2_X1 U11415 ( .A1(n12152), .A2(n12151), .ZN(n15166) );
  NAND2_X1 U11416 ( .A1(n10403), .A2(n10402), .ZN(n10420) );
  NAND2_X1 U11417 ( .A1(n13646), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13647) );
  INV_X1 U11418 ( .A(n13965), .ZN(n11953) );
  NOR2_X1 U11419 ( .A1(n15344), .A2(n19452), .ZN(n15341) );
  NOR2_X1 U11420 ( .A1(n12782), .A2(n12781), .ZN(n17770) );
  AND2_X1 U11421 ( .A1(n11952), .A2(n11951), .ZN(n13965) );
  XNOR2_X1 U11422 ( .A(n11844), .B(n11843), .ZN(n11909) );
  OR2_X1 U11423 ( .A1(n18270), .A2(n18287), .ZN(n18196) );
  NOR2_X2 U11424 ( .A1(n19453), .A2(n19435), .ZN(n19934) );
  NAND2_X1 U11425 ( .A1(n13613), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11926) );
  NAND2_X1 U11426 ( .A1(n9932), .A2(n9832), .ZN(n11844) );
  AND2_X1 U11427 ( .A1(n15826), .A2(n15825), .ZN(n15828) );
  NOR2_X1 U11428 ( .A1(n11300), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11301) );
  NAND2_X1 U11429 ( .A1(n10414), .A2(n10413), .ZN(n19200) );
  AOI21_X1 U11431 ( .B1(n11921), .B2(n11920), .A(n12044), .ZN(n12148) );
  NAND2_X1 U11432 ( .A1(n11829), .A2(n11828), .ZN(n11931) );
  OR2_X1 U11433 ( .A1(n11829), .A2(n11828), .ZN(n9933) );
  NAND2_X1 U11434 ( .A1(n11846), .A2(n11820), .ZN(n11829) );
  XNOR2_X1 U11435 ( .A(n10424), .B(n10425), .ZN(n10398) );
  NOR2_X1 U11436 ( .A1(n19054), .A2(n10058), .ZN(n19035) );
  XNOR2_X1 U11438 ( .A(n11534), .B(n11536), .ZN(n11533) );
  NAND2_X1 U11439 ( .A1(n10409), .A2(n10410), .ZN(n10414) );
  INV_X1 U11440 ( .A(n10422), .ZN(n10425) );
  NAND3_X1 U11441 ( .A1(n10368), .A2(n10367), .A3(n10366), .ZN(n10409) );
  AND2_X1 U11442 ( .A1(n10436), .A2(n10435), .ZN(n11536) );
  AND2_X1 U11443 ( .A1(n19050), .A2(n19051), .ZN(n19054) );
  CLKBUF_X3 U11444 ( .A(n13180), .Z(n19173) );
  NAND2_X1 U11445 ( .A1(n10397), .A2(n10396), .ZN(n10422) );
  NAND2_X1 U11446 ( .A1(n10390), .A2(n10389), .ZN(n10424) );
  NAND2_X1 U11447 ( .A1(n9886), .A2(n9885), .ZN(n11280) );
  OR2_X1 U11448 ( .A1(n16814), .A2(n9835), .ZN(n10032) );
  NAND2_X1 U11449 ( .A1(n10133), .A2(n10132), .ZN(n10388) );
  OR2_X1 U11450 ( .A1(n10357), .A2(n20119), .ZN(n10367) );
  NAND2_X1 U11451 ( .A1(n16668), .A2(n18972), .ZN(n16682) );
  OR2_X2 U11452 ( .A1(n17538), .A2(n18809), .ZN(n17603) );
  NAND2_X2 U11453 ( .A1(n13206), .A2(n13211), .ZN(n12993) );
  NAND2_X2 U11454 ( .A1(n9762), .A2(n9763), .ZN(n10381) );
  OR2_X1 U11455 ( .A1(n11451), .A2(n10136), .ZN(n10132) );
  AND2_X1 U11456 ( .A1(n10316), .A2(n10850), .ZN(n10859) );
  NAND2_X1 U11457 ( .A1(n9929), .A2(n11786), .ZN(n12986) );
  OR3_X1 U11458 ( .A1(n12895), .A2(n12894), .A3(n15928), .ZN(n18766) );
  NAND2_X1 U11459 ( .A1(n11782), .A2(n11781), .ZN(n11804) );
  AND2_X1 U11460 ( .A1(n11454), .A2(n10825), .ZN(n10370) );
  NAND2_X1 U11461 ( .A1(n10349), .A2(n20109), .ZN(n10850) );
  INV_X1 U11462 ( .A(n11216), .ZN(n9885) );
  AND2_X1 U11463 ( .A1(n13103), .A2(n11785), .ZN(n13110) );
  AND2_X1 U11464 ( .A1(n17687), .A2(n10044), .ZN(n17610) );
  INV_X2 U11465 ( .A(n13091), .ZN(n13064) );
  NOR2_X1 U11466 ( .A1(n11901), .A2(n9918), .ZN(n12044) );
  INV_X1 U11467 ( .A(n12757), .ZN(n17491) );
  INV_X1 U11468 ( .A(n10015), .ZN(n13923) );
  INV_X2 U11469 ( .A(n16573), .ZN(n16623) );
  AND3_X1 U11470 ( .A1(n11799), .A2(n12981), .A3(n12089), .ZN(n11780) );
  OR2_X1 U11471 ( .A1(n11873), .A2(n11872), .ZN(n12047) );
  OR2_X1 U11472 ( .A1(n13917), .A2(n13411), .ZN(n13094) );
  INV_X2 U11473 ( .A(U212), .ZN(n16620) );
  INV_X1 U11474 ( .A(n10317), .ZN(n11446) );
  INV_X1 U11475 ( .A(n11811), .ZN(n11799) );
  INV_X1 U11476 ( .A(n19435), .ZN(n10346) );
  OR2_X1 U11477 ( .A1(n11894), .A2(n11893), .ZN(n11923) );
  OR2_X2 U11478 ( .A1(n11689), .A2(n11688), .ZN(n14360) );
  AND3_X2 U11479 ( .A1(n11701), .A2(n10234), .A3(n11700), .ZN(n11811) );
  NAND2_X4 U11480 ( .A1(n9997), .A2(n10014), .ZN(n10353) );
  AND4_X1 U11481 ( .A1(n11764), .A2(n11763), .A3(n11762), .A4(n11761), .ZN(
        n11775) );
  AND4_X1 U11482 ( .A1(n11750), .A2(n11749), .A3(n11748), .A4(n11747), .ZN(
        n11751) );
  INV_X2 U11483 ( .A(U214), .ZN(n16621) );
  NAND2_X1 U11484 ( .A1(n10242), .A2(n10456), .ZN(n9997) );
  NAND2_X1 U11485 ( .A1(n10247), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10014) );
  NAND2_X1 U11486 ( .A1(n10279), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10280) );
  NAND2_X1 U11487 ( .A1(n9909), .A2(n9910), .ZN(n9908) );
  AND4_X1 U11488 ( .A1(n11760), .A2(n11759), .A3(n11758), .A4(n11757), .ZN(
        n11776) );
  AND4_X1 U11489 ( .A1(n11738), .A2(n11737), .A3(n11736), .A4(n11735), .ZN(
        n11755) );
  INV_X1 U11490 ( .A(n17233), .ZN(n15901) );
  AND4_X1 U11491 ( .A1(n11724), .A2(n11723), .A3(n11722), .A4(n11721), .ZN(
        n11731) );
  AND4_X1 U11492 ( .A1(n11720), .A2(n11719), .A3(n11718), .A4(n11717), .ZN(
        n11732) );
  AND4_X1 U11493 ( .A1(n11746), .A2(n11745), .A3(n11744), .A4(n11743), .ZN(
        n11752) );
  AND4_X1 U11494 ( .A1(n11742), .A2(n11741), .A3(n11740), .A4(n11739), .ZN(
        n11754) );
  AND3_X1 U11495 ( .A1(n10320), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10321), .ZN(n9909) );
  NOR2_X1 U11496 ( .A1(n9799), .A2(n10065), .ZN(n10064) );
  AND4_X1 U11497 ( .A1(n10273), .A2(n10272), .A3(n10271), .A4(n10270), .ZN(
        n10274) );
  NAND2_X2 U11498 ( .A1(n18950), .A2(n21159), .ZN(n18896) );
  AND4_X1 U11499 ( .A1(n10278), .A2(n10277), .A3(n10276), .A4(n10275), .ZN(
        n10279) );
  NAND2_X2 U11500 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20129), .ZN(n20046) );
  INV_X2 U11501 ( .A(n16654), .ZN(U215) );
  CLKBUF_X3 U11502 ( .A(n12688), .Z(n17295) );
  CLKBUF_X3 U11503 ( .A(n12833), .Z(n17277) );
  INV_X2 U11504 ( .A(n16658), .ZN(n16660) );
  NOR2_X1 U11505 ( .A1(n18773), .A2(n12665), .ZN(n13526) );
  OR2_X1 U11506 ( .A1(n18758), .A2(n12665), .ZN(n10227) );
  NOR2_X1 U11507 ( .A1(n12667), .A2(n12668), .ZN(n12833) );
  AND2_X1 U11508 ( .A1(n11663), .A2(n11662), .ZN(n11860) );
  AND2_X2 U11509 ( .A1(n11664), .A2(n11665), .ZN(n11831) );
  AND2_X2 U11510 ( .A1(n11665), .A2(n13681), .ZN(n11852) );
  INV_X2 U11511 ( .A(n19287), .ZN(n19350) );
  AND2_X2 U11512 ( .A1(n11661), .A2(n11665), .ZN(n11940) );
  INV_X2 U11513 ( .A(n18969), .ZN(n18950) );
  NAND2_X1 U11514 ( .A1(n18933), .A2(n21189), .ZN(n12667) );
  NAND2_X1 U11515 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18920), .ZN(
        n12662) );
  AND2_X1 U11516 ( .A1(n11655), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11665) );
  NAND2_X1 U11517 ( .A1(n21189), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n18773) );
  AND2_X2 U11518 ( .A1(n15837), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9771) );
  AND2_X1 U11519 ( .A1(n11802), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11663) );
  NAND2_X1 U11520 ( .A1(n18940), .A2(n18920), .ZN(n12665) );
  INV_X4 U11521 ( .A(n12705), .ZN(n9758) );
  AND2_X2 U11522 ( .A1(n15837), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10804) );
  NAND3_X2 U11523 ( .A1(n21185), .A2(n18971), .A3(n18962), .ZN(n16866) );
  NOR2_X2 U11524 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15837) );
  INV_X1 U11525 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18920) );
  INV_X2 U11526 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n9918) );
  AND2_X2 U11527 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13681) );
  NOR2_X1 U11528 ( .A1(n18334), .A2(n17349), .ZN(n18788) );
  CLKBUF_X1 U11529 ( .A(n10358), .Z(n16502) );
  NAND2_X1 U11530 ( .A1(n10123), .A2(n10122), .ZN(n14852) );
  AND2_X1 U11531 ( .A1(n11394), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n9760) );
  OAI21_X2 U11532 ( .B1(n14882), .B2(n10129), .A(n10128), .ZN(n10127) );
  NOR2_X2 U11533 ( .A1(n11707), .A2(n11706), .ZN(n11712) );
  INV_X1 U11535 ( .A(n11217), .ZN(n9886) );
  AOI21_X1 U11536 ( .B1(n9987), .B2(n11370), .A(n9810), .ZN(n9986) );
  AND2_X2 U11537 ( .A1(n15784), .A2(n9761), .ZN(n14425) );
  AND2_X1 U11538 ( .A1(n9861), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9761) );
  NAND2_X1 U11539 ( .A1(n10349), .A2(n20109), .ZN(n9762) );
  NOR2_X2 U11540 ( .A1(n11778), .A2(n12089), .ZN(n13364) );
  AND2_X1 U11541 ( .A1(n13833), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9764) );
  AND2_X2 U11542 ( .A1(n11403), .A2(n13745), .ZN(n9765) );
  AND2_X2 U11543 ( .A1(n11403), .A2(n13745), .ZN(n10457) );
  AND2_X1 U11544 ( .A1(n10317), .A2(n10345), .ZN(n11454) );
  XNOR2_X2 U11545 ( .A(n11881), .B(n11880), .ZN(n12159) );
  AND2_X2 U11546 ( .A1(n13834), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9766) );
  NOR2_X1 U11547 ( .A1(n14468), .A2(n14467), .ZN(n14466) );
  AND2_X1 U11548 ( .A1(n11663), .A2(n11662), .ZN(n9767) );
  OR2_X2 U11549 ( .A1(n13887), .A2(n10451), .ZN(n10145) );
  NAND2_X1 U11550 ( .A1(n11755), .A2(n9797), .ZN(n9768) );
  NAND2_X1 U11551 ( .A1(n11755), .A2(n9797), .ZN(n9769) );
  NAND2_X2 U11552 ( .A1(n15809), .A2(n11524), .ZN(n15602) );
  NAND2_X2 U11553 ( .A1(n15808), .A2(n15807), .ZN(n15809) );
  NAND2_X2 U11554 ( .A1(n9977), .A2(n11284), .ZN(n15604) );
  NAND2_X2 U11555 ( .A1(n10477), .A2(n10476), .ZN(n13938) );
  AND2_X4 U11556 ( .A1(n13931), .A2(n10511), .ZN(n14023) );
  NOR2_X4 U11557 ( .A1(n13938), .A2(n11016), .ZN(n13931) );
  NAND2_X2 U11558 ( .A1(n13767), .A2(n13766), .ZN(n13765) );
  NAND4_X1 U11559 ( .A1(n11794), .A2(n11800), .A3(n11793), .A4(n11792), .ZN(
        n11795) );
  AND2_X1 U11560 ( .A1(n11403), .A2(n13745), .ZN(n9770) );
  OR2_X1 U11561 ( .A1(n10330), .A2(n11461), .ZN(n10335) );
  NAND2_X1 U11562 ( .A1(n11784), .A2(n9768), .ZN(n13083) );
  NAND2_X1 U11563 ( .A1(n9981), .A2(n9979), .ZN(n11461) );
  INV_X2 U11564 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13745) );
  AND2_X4 U11565 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13834) );
  NAND2_X2 U11566 ( .A1(n10123), .A2(n14873), .ZN(n14816) );
  XNOR2_X1 U11567 ( .A(n11980), .B(n11962), .ZN(n20288) );
  XNOR2_X2 U11568 ( .A(n11506), .B(n11505), .ZN(n14002) );
  INV_X2 U11569 ( .A(n10142), .ZN(n15253) );
  AND2_X4 U11570 ( .A1(n14340), .A2(n14671), .ZN(n14672) );
  NOR2_X4 U11571 ( .A1(n14332), .A2(n14342), .ZN(n14340) );
  OAI21_X2 U11572 ( .B1(n16158), .B2(n9927), .A(n9924), .ZN(n14263) );
  INV_X2 U11573 ( .A(n11915), .ZN(n14138) );
  NAND4_X1 U11574 ( .A1(n11776), .A2(n11775), .A3(n11774), .A4(n11773), .ZN(
        n11915) );
  AOI21_X2 U11575 ( .B1(n11801), .B2(n10235), .A(n9918), .ZN(n11819) );
  NAND2_X2 U11576 ( .A1(n15248), .A2(n15247), .ZN(n15249) );
  NAND2_X1 U11577 ( .A1(n13083), .A2(n13061), .ZN(n13006) );
  NAND2_X2 U11578 ( .A1(n12072), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14832) );
  INV_X1 U11579 ( .A(n10293), .ZN(n9774) );
  OAI222_X1 U11580 ( .A1(n14730), .A2(n14846), .B1(n14694), .B2(n20227), .C1(
        n14995), .C2(n14725), .ZN(P1_U2846) );
  OAI21_X2 U11581 ( .B1(n14614), .B2(n14615), .A(n14602), .ZN(n14846) );
  OR2_X1 U11582 ( .A1(n11101), .A2(n15847), .ZN(n11115) );
  NAND2_X2 U11583 ( .A1(n14883), .A2(n14901), .ZN(n14882) );
  XNOR2_X2 U11584 ( .A(n11927), .B(n11926), .ZN(n13646) );
  NOR2_X2 U11585 ( .A1(n14417), .A2(n14419), .ZN(n14418) );
  NAND2_X2 U11587 ( .A1(n11898), .A2(n11897), .ZN(n11921) );
  NAND2_X1 U11588 ( .A1(n11819), .A2(n11818), .ZN(n11820) );
  OAI21_X2 U11589 ( .B1(n11795), .B2(n12993), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11821) );
  BUF_X4 U11590 ( .A(n11547), .Z(n9775) );
  NAND2_X1 U11591 ( .A1(n11466), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11547) );
  XNOR2_X1 U11592 ( .A(n11914), .B(n11903), .ZN(n12147) );
  OAI21_X2 U11593 ( .B1(n13704), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11859), 
        .ZN(n11914) );
  NOR2_X4 U11594 ( .A1(n14644), .A2(n14645), .ZN(n14627) );
  NOR2_X1 U11595 ( .A1(n13436), .A2(n11466), .ZN(n9779) );
  NAND2_X1 U11596 ( .A1(n13382), .A2(n9748), .ZN(n9780) );
  OR2_X1 U11597 ( .A1(n12996), .A2(n9918), .ZN(n11937) );
  OAI21_X1 U11598 ( .B1(n11804), .B2(n11790), .A(n11788), .ZN(n11793) );
  OR2_X1 U11599 ( .A1(n11858), .A2(n11857), .ZN(n11916) );
  AND2_X1 U11600 ( .A1(n13547), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11899) );
  NAND2_X1 U11601 ( .A1(n11788), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11938) );
  NAND2_X1 U11602 ( .A1(n11198), .A2(n11197), .ZN(n11276) );
  OR2_X1 U11603 ( .A1(n14224), .A2(n14299), .ZN(n12306) );
  AND2_X1 U11604 ( .A1(n11928), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10105) );
  NAND2_X1 U11605 ( .A1(n11811), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12338) );
  OR2_X1 U11606 ( .A1(n14360), .A2(n20839), .ZN(n12638) );
  INV_X1 U11607 ( .A(n10127), .ZN(n10123) );
  NAND2_X1 U11608 ( .A1(n10130), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10129) );
  NAND2_X1 U11609 ( .A1(n15089), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10128) );
  NOR2_X1 U11610 ( .A1(n10100), .A2(n15327), .ZN(n10098) );
  NOR2_X1 U11611 ( .A1(n10629), .A2(n10154), .ZN(n10153) );
  INV_X1 U11612 ( .A(n10532), .ZN(n10154) );
  INV_X1 U11613 ( .A(n15762), .ZN(n10003) );
  OR2_X1 U11614 ( .A1(n10094), .A2(n13762), .ZN(n10093) );
  NAND2_X1 U11615 ( .A1(n10095), .A2(n13638), .ZN(n10094) );
  INV_X1 U11616 ( .A(n13620), .ZN(n10095) );
  NAND2_X1 U11617 ( .A1(n11274), .A2(n11273), .ZN(n11512) );
  OR3_X1 U11618 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18920), .A3(
        n18758), .ZN(n12705) );
  NOR2_X1 U11619 ( .A1(n12662), .A2(n18773), .ZN(n12688) );
  NOR2_X1 U11620 ( .A1(n18773), .A2(n12668), .ZN(n12707) );
  OAI21_X1 U11621 ( .B1(n14852), .B2(n14817), .A(n15089), .ZN(n14843) );
  NAND2_X1 U11622 ( .A1(n14649), .A2(n14630), .ZN(n14632) );
  NAND2_X1 U11623 ( .A1(n13120), .A2(n13422), .ZN(n20314) );
  NAND2_X1 U11624 ( .A1(n13120), .A2(n13107), .ZN(n15050) );
  INV_X1 U11625 ( .A(n14102), .ZN(n10082) );
  INV_X1 U11626 ( .A(n13242), .ZN(n10081) );
  AND2_X1 U11627 ( .A1(n9828), .A2(n15592), .ZN(n10206) );
  OAI21_X1 U11628 ( .B1(n14001), .B2(n14000), .A(n11239), .ZN(n16372) );
  NOR3_X1 U11629 ( .A1(n13288), .A2(n13289), .A3(n15242), .ZN(n15246) );
  AND2_X1 U11630 ( .A1(n11430), .A2(n20123), .ZN(n11650) );
  AOI21_X1 U11631 ( .B1(n12916), .B2(n12918), .A(n12915), .ZN(n18748) );
  NOR2_X2 U11632 ( .A1(n15919), .A2(n12901), .ZN(n17540) );
  NOR2_X1 U11633 ( .A1(n9876), .A2(n9875), .ZN(n9874) );
  AOI21_X1 U11634 ( .B1(n12132), .B2(n14042), .A(n12090), .ZN(n12098) );
  INV_X1 U11635 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n9963) );
  NOR2_X1 U11636 ( .A1(n11842), .A2(n11841), .ZN(n11957) );
  NOR2_X1 U11637 ( .A1(n12139), .A2(n13854), .ZN(n11734) );
  NAND2_X1 U11638 ( .A1(n10984), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n9883) );
  NAND2_X1 U11639 ( .A1(n10896), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n9881) );
  NAND2_X1 U11640 ( .A1(n10986), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n9882) );
  NAND2_X1 U11641 ( .A1(n9759), .A2(n9852), .ZN(n11341) );
  INV_X1 U11642 ( .A(n11431), .ZN(n10825) );
  NOR2_X1 U11643 ( .A1(n11276), .A2(n11512), .ZN(n11275) );
  INV_X1 U11644 ( .A(n11277), .ZN(n10192) );
  INV_X1 U11645 ( .A(n10369), .ZN(n10135) );
  AND3_X1 U11646 ( .A1(n10354), .A2(n9747), .A3(n10928), .ZN(n11452) );
  AND2_X1 U11647 ( .A1(n19442), .A2(n10329), .ZN(n10330) );
  AND2_X1 U11648 ( .A1(n10353), .A2(n9747), .ZN(n10329) );
  NAND2_X1 U11649 ( .A1(n10928), .A2(n11461), .ZN(n10334) );
  AND2_X1 U11650 ( .A1(n10346), .A2(n11457), .ZN(n10333) );
  INV_X1 U11651 ( .A(n10297), .ZN(n9983) );
  NAND2_X1 U11652 ( .A1(n17881), .A2(n12777), .ZN(n12952) );
  INV_X1 U11653 ( .A(n12919), .ZN(n12759) );
  NOR2_X1 U11654 ( .A1(n12446), .A2(n10021), .ZN(n10020) );
  INV_X1 U11655 ( .A(n12410), .ZN(n10021) );
  NOR2_X1 U11656 ( .A1(n12307), .A2(n14282), .ZN(n12324) );
  NOR2_X1 U11657 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n9923), .ZN(
        n9922) );
  INV_X1 U11658 ( .A(n12031), .ZN(n10111) );
  INV_X1 U11659 ( .A(n14244), .ZN(n10115) );
  INV_X1 U11660 ( .A(n14243), .ZN(n10113) );
  INV_X1 U11661 ( .A(n12032), .ZN(n10114) );
  NAND2_X1 U11662 ( .A1(n10110), .A2(n9926), .ZN(n9925) );
  INV_X1 U11663 ( .A(n12009), .ZN(n9926) );
  OR2_X1 U11664 ( .A1(n12019), .A2(n12018), .ZN(n12038) );
  OR2_X1 U11665 ( .A1(n14540), .A2(n13064), .ZN(n13090) );
  OAI21_X1 U11666 ( .B1(n11914), .B2(n14138), .A(n11919), .ZN(n11927) );
  OR2_X1 U11667 ( .A1(n13099), .A2(n13547), .ZN(n11783) );
  NAND2_X1 U11668 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11690) );
  NAND3_X1 U11669 ( .A1(n9916), .A2(n11797), .A3(n9915), .ZN(n9919) );
  AND3_X1 U11670 ( .A1(n19435), .A2(n10317), .A3(n11461), .ZN(n10339) );
  OR2_X1 U11671 ( .A1(n16285), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10223) );
  INV_X1 U11672 ( .A(n15399), .ZN(n10008) );
  NOR2_X2 U11673 ( .A1(n11280), .A2(n11279), .ZN(n11288) );
  NAND2_X1 U11674 ( .A1(n11238), .A2(n9887), .ZN(n11217) );
  INV_X1 U11675 ( .A(n11237), .ZN(n9887) );
  NOR2_X1 U11676 ( .A1(n10085), .A2(n10084), .ZN(n10083) );
  INV_X1 U11677 ( .A(n14026), .ZN(n10084) );
  INV_X1 U11678 ( .A(n10086), .ZN(n10085) );
  NOR2_X1 U11679 ( .A1(n14092), .A2(n10087), .ZN(n10086) );
  INV_X1 U11680 ( .A(n13932), .ZN(n10087) );
  INV_X1 U11681 ( .A(n10354), .ZN(n10363) );
  INV_X1 U11682 ( .A(n14438), .ZN(n11039) );
  NAND2_X1 U11683 ( .A1(n10363), .A2(n10345), .ZN(n10862) );
  INV_X1 U11684 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10065) );
  INV_X1 U11685 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10068) );
  AND2_X1 U11686 ( .A1(n11039), .A2(n11043), .ZN(n10013) );
  INV_X1 U11687 ( .A(n15429), .ZN(n11043) );
  INV_X1 U11688 ( .A(n14467), .ZN(n10195) );
  OR2_X1 U11689 ( .A1(n14445), .A2(n15532), .ZN(n10197) );
  NAND2_X1 U11690 ( .A1(n10199), .A2(n14391), .ZN(n10198) );
  AND2_X1 U11691 ( .A1(n10206), .A2(n10205), .ZN(n10204) );
  INV_X1 U11692 ( .A(n16350), .ZN(n10205) );
  NAND2_X1 U11693 ( .A1(n10204), .A2(n11292), .ZN(n10202) );
  NAND2_X1 U11694 ( .A1(n10006), .A2(n16432), .ZN(n10005) );
  INV_X1 U11695 ( .A(n15812), .ZN(n10006) );
  NOR2_X1 U11696 ( .A1(n10992), .A2(n10991), .ZN(n11215) );
  OAI21_X1 U11697 ( .B1(n10430), .B2(n10456), .A(n10429), .ZN(n11534) );
  NOR2_X1 U11698 ( .A1(n13863), .A2(n13873), .ZN(n9905) );
  NAND2_X1 U11699 ( .A1(n13863), .A2(n13873), .ZN(n9904) );
  NAND2_X1 U11700 ( .A1(n13580), .A2(n11396), .ZN(n9899) );
  NOR2_X1 U11701 ( .A1(n9905), .A2(n9902), .ZN(n9901) );
  INV_X1 U11702 ( .A(n13580), .ZN(n9902) );
  NAND2_X1 U11703 ( .A1(n10426), .A2(n10425), .ZN(n10427) );
  AND3_X1 U11704 ( .A1(n10967), .A2(n10966), .A3(n10965), .ZN(n13574) );
  NOR2_X1 U11705 ( .A1(n15847), .A2(n11087), .ZN(n9984) );
  INV_X1 U11706 ( .A(n12663), .ZN(n17233) );
  NOR2_X1 U11707 ( .A1(n18778), .A2(n12665), .ZN(n12708) );
  NAND2_X1 U11708 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12666) );
  OR2_X1 U11709 ( .A1(n15929), .A2(n12906), .ZN(n12901) );
  AND2_X1 U11710 ( .A1(n12782), .A2(n16508), .ZN(n10177) );
  NAND2_X1 U11711 ( .A1(n12896), .A2(n12893), .ZN(n15919) );
  INV_X1 U11712 ( .A(n12890), .ZN(n9949) );
  INV_X1 U11713 ( .A(n12884), .ZN(n9948) );
  NOR2_X1 U11714 ( .A1(n12888), .A2(n9951), .ZN(n9950) );
  AND2_X1 U11715 ( .A1(n12952), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17791) );
  NOR2_X1 U11716 ( .A1(n12952), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12778) );
  NOR2_X1 U11717 ( .A1(n12937), .A2(n17902), .ZN(n12940) );
  NAND2_X1 U11718 ( .A1(n17942), .A2(n12761), .ZN(n12765) );
  OR2_X1 U11719 ( .A1(n18261), .A2(n12760), .ZN(n12761) );
  AND2_X1 U11720 ( .A1(n13418), .A2(n9856), .ZN(n13422) );
  NAND2_X1 U11721 ( .A1(n12324), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12342) );
  OR2_X1 U11722 ( .A1(n14045), .A2(n11788), .ZN(n14057) );
  INV_X1 U11723 ( .A(n14057), .ZN(n14047) );
  OR3_X1 U11724 ( .A1(n20844), .A2(n20299), .A3(n14034), .ZN(n14112) );
  NOR3_X1 U11725 ( .A1(n14632), .A2(n13087), .A3(n14620), .ZN(n14593) );
  INV_X1 U11726 ( .A(n14540), .ZN(n13560) );
  NAND2_X1 U11727 ( .A1(n14138), .A2(n9769), .ZN(n13604) );
  NAND2_X1 U11728 ( .A1(n12466), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12514) );
  NAND2_X1 U11729 ( .A1(n12411), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12464) );
  NAND2_X1 U11730 ( .A1(n12359), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12375) );
  AND2_X1 U11731 ( .A1(n14318), .A2(n14319), .ZN(n14320) );
  NAND2_X1 U11732 ( .A1(n12201), .A2(n12200), .ZN(n14014) );
  NAND2_X1 U11733 ( .A1(n13656), .A2(n12167), .ZN(n13772) );
  INV_X1 U11734 ( .A(n14620), .ZN(n9962) );
  INV_X1 U11735 ( .A(n14569), .ZN(n9960) );
  NOR3_X1 U11736 ( .A1(n14632), .A2(n13087), .A3(n9961), .ZN(n14570) );
  NAND2_X1 U11737 ( .A1(n9962), .A2(n13092), .ZN(n9961) );
  AOI21_X1 U11738 ( .B1(n10118), .B2(n15089), .A(n10117), .ZN(n10122) );
  INV_X1 U11739 ( .A(n10120), .ZN(n10117) );
  AOI21_X1 U11740 ( .B1(n15089), .B2(n10121), .A(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10120) );
  NOR2_X1 U11741 ( .A1(n13074), .A2(n14700), .ZN(n14649) );
  INV_X1 U11742 ( .A(n10119), .ZN(n14873) );
  NAND2_X1 U11743 ( .A1(n14263), .A2(n12050), .ZN(n12052) );
  OR2_X1 U11744 ( .A1(n14264), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12050) );
  AND2_X1 U11745 ( .A1(n12992), .A2(n13564), .ZN(n13120) );
  NAND2_X1 U11746 ( .A1(n20815), .A2(n9918), .ZN(n11952) );
  NOR2_X1 U11747 ( .A1(n20820), .A2(n13947), .ZN(n20812) );
  OR2_X1 U11748 ( .A1(n13731), .A2(n13965), .ZN(n20672) );
  NAND2_X1 U11749 ( .A1(n12138), .A2(n12137), .ZN(n13429) );
  NAND2_X1 U11750 ( .A1(n12136), .A2(n12974), .ZN(n12137) );
  OAI21_X1 U11751 ( .B1(n12136), .B2(n12134), .A(n12133), .ZN(n12138) );
  NAND2_X1 U11752 ( .A1(n12128), .A2(n12127), .ZN(n12136) );
  NAND2_X1 U11753 ( .A1(n16293), .A2(n20930), .ZN(n16285) );
  NAND2_X1 U11754 ( .A1(n19173), .A2(n16307), .ZN(n10061) );
  NAND2_X1 U11756 ( .A1(n19173), .A2(n19001), .ZN(n10057) );
  INV_X1 U11758 ( .A(n14463), .ZN(n10101) );
  AND2_X1 U11759 ( .A1(n14462), .A2(n10098), .ZN(n15329) );
  AND2_X1 U11760 ( .A1(n11582), .A2(n11581), .ZN(n14102) );
  AND2_X2 U11761 ( .A1(n15348), .A2(n15347), .ZN(n15349) );
  OR2_X1 U11762 ( .A1(n10153), .A2(n10680), .ZN(n10152) );
  NAND2_X1 U11763 ( .A1(n14023), .A2(n9826), .ZN(n10149) );
  INV_X1 U11764 ( .A(n10680), .ZN(n10151) );
  INV_X1 U11765 ( .A(n14023), .ZN(n10147) );
  AND3_X1 U11766 ( .A1(n11013), .A2(n11012), .A3(n11011), .ZN(n15794) );
  NAND2_X1 U11767 ( .A1(n16443), .A2(n11005), .ZN(n15826) );
  NAND2_X1 U11768 ( .A1(n10449), .A2(n10448), .ZN(n13887) );
  NOR2_X1 U11769 ( .A1(n10090), .A2(n10089), .ZN(n10088) );
  INV_X1 U11770 ( .A(n15263), .ZN(n10089) );
  OR3_X1 U11771 ( .A1(n13289), .A2(n15242), .A3(n10091), .ZN(n10090) );
  INV_X1 U11772 ( .A(n12656), .ZN(n10091) );
  OR2_X1 U11773 ( .A1(n10189), .A2(n15639), .ZN(n10188) );
  INV_X1 U11774 ( .A(n11370), .ZN(n9988) );
  NAND2_X1 U11775 ( .A1(n15301), .A2(n11617), .ZN(n15285) );
  INV_X1 U11776 ( .A(n10184), .ZN(n10183) );
  OAI21_X1 U11777 ( .B1(n15601), .B2(n10185), .A(n11530), .ZN(n10184) );
  INV_X1 U11778 ( .A(n14460), .ZN(n10002) );
  INV_X1 U11779 ( .A(n15788), .ZN(n10207) );
  OR2_X1 U11780 ( .A1(n10093), .A2(n10096), .ZN(n10092) );
  INV_X1 U11781 ( .A(n13780), .ZN(n10096) );
  AND2_X1 U11782 ( .A1(n15607), .A2(n15804), .ZN(n11291) );
  OR2_X1 U11783 ( .A1(n15604), .A2(n11292), .ZN(n10208) );
  NAND2_X1 U11784 ( .A1(n9978), .A2(n11241), .ZN(n15618) );
  NAND2_X1 U11785 ( .A1(n14006), .A2(n14506), .ZN(n14507) );
  INV_X1 U11786 ( .A(n9906), .ZN(n9903) );
  NAND2_X1 U11787 ( .A1(n11424), .A2(n10849), .ZN(n16478) );
  OR2_X1 U11788 ( .A1(n15893), .A2(n19274), .ZN(n19725) );
  AND2_X1 U11789 ( .A1(n20072), .A2(n20079), .ZN(n20060) );
  NAND2_X1 U11790 ( .A1(n20119), .A2(n15875), .ZN(n19796) );
  NAND2_X1 U11791 ( .A1(n17029), .A2(n10034), .ZN(n10033) );
  INV_X1 U11792 ( .A(n17693), .ZN(n10034) );
  OR2_X1 U11793 ( .A1(n16814), .A2(n17708), .ZN(n10035) );
  BUF_X1 U11794 ( .A(n17192), .Z(n17248) );
  BUF_X1 U11795 ( .A(n12708), .Z(n17303) );
  NAND2_X1 U11796 ( .A1(n17625), .A2(n17872), .ZN(n16551) );
  AND2_X1 U11797 ( .A1(n12792), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17625) );
  NOR2_X1 U11798 ( .A1(n12792), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17624) );
  AND2_X1 U11799 ( .A1(n17870), .A2(n12782), .ZN(n17803) );
  NAND3_X1 U11800 ( .A1(n18328), .A2(n18236), .A3(n13448), .ZN(n18750) );
  INV_X1 U11801 ( .A(n17906), .ZN(n10175) );
  NAND2_X1 U11802 ( .A1(n10172), .A2(n18231), .ZN(n10171) );
  INV_X1 U11803 ( .A(n17907), .ZN(n10172) );
  AND2_X1 U11804 ( .A1(n17893), .A2(n10171), .ZN(n10170) );
  AND2_X1 U11805 ( .A1(n9814), .A2(n10182), .ZN(n17960) );
  NOR2_X1 U11806 ( .A1(n12756), .A2(n12755), .ZN(n10182) );
  AND2_X1 U11807 ( .A1(n15921), .A2(n12897), .ZN(n9955) );
  NAND2_X1 U11808 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18758) );
  INV_X1 U11809 ( .A(n20194), .ZN(n20206) );
  INV_X1 U11810 ( .A(n20162), .ZN(n20216) );
  OR2_X1 U11811 ( .A1(n12648), .A2(n21154), .ZN(n12649) );
  AND2_X1 U11812 ( .A1(n20139), .A2(n12650), .ZN(n20287) );
  OR2_X1 U11813 ( .A1(n13546), .A2(n15985), .ZN(n20139) );
  INV_X1 U11814 ( .A(n20312), .ZN(n16218) );
  AOI21_X1 U11816 ( .B1(n16254), .B2(n16253), .A(n19972), .ZN(n10078) );
  AND2_X1 U11817 ( .A1(n16256), .A2(n9815), .ZN(n10076) );
  INV_X1 U11818 ( .A(n15541), .ZN(n19031) );
  INV_X1 U11819 ( .A(n20079), .ZN(n19407) );
  XOR2_X1 U11820 ( .A(n11432), .B(n15349), .Z(n15627) );
  NAND2_X1 U11821 ( .A1(n15350), .A2(n9830), .ZN(n15359) );
  AND2_X1 U11822 ( .A1(n19270), .A2(n19452), .ZN(n19263) );
  OAI21_X1 U11823 ( .B1(n15309), .B2(n14529), .A(n14528), .ZN(n14530) );
  INV_X1 U11824 ( .A(n16370), .ZN(n19374) );
  NAND2_X1 U11825 ( .A1(n11652), .A2(n19402), .ZN(n11653) );
  XNOR2_X1 U11826 ( .A(n15246), .B(n12656), .ZN(n15630) );
  OAI21_X1 U11827 ( .B1(n14478), .B2(n9995), .A(n11389), .ZN(n15465) );
  OR2_X1 U11828 ( .A1(n15525), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14523) );
  NAND2_X1 U11829 ( .A1(n9809), .A2(n9789), .ZN(n14412) );
  NOR2_X1 U11830 ( .A1(n14514), .A2(n15533), .ZN(n14393) );
  XNOR2_X1 U11831 ( .A(n14447), .B(n14446), .ZN(n15551) );
  AND2_X1 U11832 ( .A1(n11650), .A2(n20101), .ZN(n16451) );
  AND2_X1 U11833 ( .A1(n14426), .A2(n14427), .ZN(n19396) );
  NOR2_X1 U11834 ( .A1(n17029), .A2(n16699), .ZN(n16712) );
  NOR2_X1 U11835 ( .A1(n16725), .A2(n17029), .ZN(n16718) );
  NAND2_X1 U11836 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17068), .ZN(n17053) );
  INV_X1 U11837 ( .A(n17060), .ZN(n17068) );
  NAND2_X1 U11838 ( .A1(n17356), .A2(n9853), .ZN(n9943) );
  NAND2_X1 U11839 ( .A1(n17358), .A2(n17486), .ZN(n17356) );
  NAND2_X1 U11840 ( .A1(n17361), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n17358) );
  NOR2_X1 U11841 ( .A1(n17565), .A2(n17367), .ZN(n17361) );
  NOR2_X1 U11842 ( .A1(n17432), .A2(n17604), .ZN(n17427) );
  INV_X1 U11843 ( .A(n17392), .ZN(n17424) );
  INV_X1 U11844 ( .A(n17960), .ZN(n10181) );
  AOI21_X1 U11845 ( .B1(n16023), .B2(n16022), .A(n18817), .ZN(n17498) );
  NAND3_X1 U11846 ( .A1(n18748), .A2(n18953), .A3(n16683), .ZN(n16023) );
  INV_X1 U11847 ( .A(n17487), .ZN(n17492) );
  AND2_X1 U11848 ( .A1(n17910), .A2(n17468), .ZN(n17801) );
  INV_X1 U11849 ( .A(n17953), .ZN(n17966) );
  INV_X1 U11850 ( .A(n17910), .ZN(n17965) );
  OAI21_X1 U11851 ( .B1(n12799), .B2(n12798), .A(n12797), .ZN(n16547) );
  OAI22_X1 U11852 ( .A1(n19757), .A2(n11098), .B1(n11097), .B2(n11177), .ZN(
        n11099) );
  XNOR2_X1 U11853 ( .A(n10353), .B(n10447), .ZN(n10852) );
  INV_X1 U11854 ( .A(n12066), .ZN(n10130) );
  INV_X1 U11855 ( .A(n12064), .ZN(n9940) );
  NOR2_X1 U11856 ( .A1(n12064), .A2(n10131), .ZN(n9939) );
  NAND2_X1 U11857 ( .A1(n9813), .A2(n12053), .ZN(n10131) );
  AND2_X1 U11858 ( .A1(n12021), .A2(n12020), .ZN(n12023) );
  OR2_X1 U11859 ( .A1(n13604), .A2(n11786), .ZN(n11787) );
  AOI21_X1 U11860 ( .B1(n12582), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n11768), .ZN(n11774) );
  NOR2_X1 U11861 ( .A1(n11655), .A2(n9918), .ZN(n9917) );
  NAND2_X1 U11862 ( .A1(n11795), .A2(n9917), .ZN(n9916) );
  INV_X1 U11863 ( .A(n12124), .ZN(n12120) );
  AND2_X1 U11864 ( .A1(n12103), .A2(n12102), .ZN(n12107) );
  OR2_X1 U11865 ( .A1(n10964), .A2(n10963), .ZN(n11206) );
  AND2_X1 U11866 ( .A1(n10322), .A2(n10319), .ZN(n9910) );
  AND4_X1 U11867 ( .A1(n10874), .A2(n10873), .A3(n10872), .A4(n10871), .ZN(
        n10889) );
  AND4_X1 U11868 ( .A1(n10878), .A2(n10877), .A3(n10876), .A4(n10875), .ZN(
        n10888) );
  OAI21_X1 U11869 ( .B1(n11277), .B2(n11276), .A(n11512), .ZN(n10191) );
  OAI22_X1 U11870 ( .A1(n11139), .A2(n19731), .B1(n11177), .B2(n11138), .ZN(
        n11140) );
  NAND2_X1 U11871 ( .A1(n10137), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10136) );
  NOR2_X1 U11872 ( .A1(n10327), .A2(n13592), .ZN(n11023) );
  NAND2_X1 U11873 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18940), .ZN(
        n12668) );
  NAND2_X1 U11874 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n9952) );
  OAI22_X1 U11875 ( .A1(n12913), .A2(n12800), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18793), .ZN(n12806) );
  NOR2_X1 U11876 ( .A1(n12762), .A2(n12763), .ZN(n12768) );
  NAND2_X1 U11877 ( .A1(n17491), .A2(n10181), .ZN(n12924) );
  NAND2_X1 U11878 ( .A1(n13560), .A2(n9802), .ZN(n13001) );
  NOR2_X1 U11879 ( .A1(n10030), .A2(n14604), .ZN(n10028) );
  NOR2_X1 U11880 ( .A1(n12305), .A2(n10026), .ZN(n10025) );
  INV_X1 U11881 ( .A(n14251), .ZN(n10026) );
  NAND2_X1 U11882 ( .A1(n14223), .A2(n14225), .ZN(n14224) );
  AND2_X1 U11883 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n12193), .ZN(
        n12202) );
  INV_X1 U11884 ( .A(n12194), .ZN(n12193) );
  INV_X1 U11885 ( .A(n12338), .ZN(n12317) );
  INV_X1 U11886 ( .A(n12070), .ZN(n10121) );
  NAND2_X1 U11887 ( .A1(n14920), .A2(n12056), .ZN(n14907) );
  AND2_X1 U11888 ( .A1(n14918), .A2(n12057), .ZN(n14906) );
  NAND2_X1 U11889 ( .A1(n16209), .A2(n9831), .ZN(n9968) );
  INV_X1 U11890 ( .A(n14232), .ZN(n9964) );
  NOR2_X1 U11891 ( .A1(n14113), .A2(n9966), .ZN(n9965) );
  INV_X1 U11892 ( .A(n14019), .ZN(n9966) );
  INV_X1 U11893 ( .A(n13090), .ZN(n13056) );
  XNOR2_X1 U11894 ( .A(n11999), .B(n11995), .ZN(n12176) );
  NAND2_X1 U11895 ( .A1(n13560), .A2(n13064), .ZN(n13080) );
  OR2_X1 U11896 ( .A1(n13099), .A2(n13061), .ZN(n13103) );
  NAND2_X1 U11897 ( .A1(n11702), .A2(n10022), .ZN(n11707) );
  NAND2_X1 U11898 ( .A1(n12621), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10022) );
  AND3_X1 U11899 ( .A1(n11878), .A2(n11882), .A3(n11877), .ZN(n11903) );
  OAI211_X1 U11900 ( .C1(n11821), .C2(n9930), .A(n11827), .B(n11826), .ZN(
        n11828) );
  OR2_X1 U11901 ( .A1(n11950), .A2(n11949), .ZN(n11975) );
  NAND2_X1 U11902 ( .A1(n11938), .A2(n11937), .ZN(n12132) );
  OAI21_X1 U11903 ( .B1(n16229), .B2(n16233), .A(n14500), .ZN(n13849) );
  AOI22_X1 U11904 ( .A1(n12126), .A2(n12125), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n9918), .ZN(n12127) );
  AND2_X1 U11905 ( .A1(n12132), .A2(n12135), .ZN(n12134) );
  OR2_X1 U11906 ( .A1(n10331), .A2(n15876), .ZN(n10332) );
  AND2_X1 U11907 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20076), .ZN(
        n10832) );
  OR3_X1 U11908 ( .A1(n10943), .A2(n9878), .A3(n9880), .ZN(n11202) );
  NAND3_X1 U11909 ( .A1(n10941), .A2(n9882), .A3(n9881), .ZN(n9880) );
  NAND2_X1 U11910 ( .A1(n11367), .A2(n11366), .ZN(n11373) );
  NAND2_X1 U11911 ( .A1(n11294), .A2(n11564), .ZN(n11300) );
  NOR2_X1 U11912 ( .A1(n11004), .A2(n11003), .ZN(n11278) );
  INV_X1 U11913 ( .A(n10067), .ZN(n10066) );
  NAND2_X1 U11914 ( .A1(n10387), .A2(n9864), .ZN(n9912) );
  NAND2_X1 U11915 ( .A1(n10414), .A2(n10404), .ZN(n9864) );
  OR2_X1 U11916 ( .A1(n10190), .A2(n14494), .ZN(n10189) );
  NAND2_X1 U11917 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10190) );
  INV_X1 U11918 ( .A(n9989), .ZN(n9987) );
  OR2_X1 U11919 ( .A1(n15955), .A2(n11322), .ZN(n11371) );
  AND2_X1 U11920 ( .A1(n10073), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9999) );
  OR2_X1 U11921 ( .A1(n19094), .A2(n11322), .ZN(n11312) );
  NOR2_X1 U11922 ( .A1(n16423), .A2(n15786), .ZN(n10073) );
  OAI21_X1 U11923 ( .B1(n11282), .B2(n11396), .A(n19156), .ZN(n11283) );
  OR2_X1 U11924 ( .A1(n11451), .A2(n11431), .ZN(n10134) );
  OR2_X1 U11925 ( .A1(n10903), .A2(n10902), .ZN(n11492) );
  INV_X1 U11926 ( .A(n10332), .ZN(n10863) );
  OR2_X1 U11927 ( .A1(n11087), .A2(n19381), .ZN(n11109) );
  NAND3_X1 U11928 ( .A1(n20064), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19883), 
        .ZN(n15879) );
  OAI21_X1 U11929 ( .B1(n9983), .B2(n9982), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9981) );
  NAND2_X1 U11930 ( .A1(n9980), .A2(n10456), .ZN(n9979) );
  AND2_X1 U11931 ( .A1(n10049), .A2(n17854), .ZN(n17723) );
  AND2_X1 U11932 ( .A1(n9786), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10049) );
  AND2_X1 U11933 ( .A1(n10222), .A2(n10051), .ZN(n10050) );
  NOR2_X1 U11934 ( .A1(n17810), .A2(n17785), .ZN(n10051) );
  AND2_X1 U11935 ( .A1(n17624), .A2(n10167), .ZN(n12793) );
  AND2_X1 U11936 ( .A1(n17606), .A2(n16536), .ZN(n10167) );
  AND2_X1 U11937 ( .A1(n17625), .A2(n10166), .ZN(n12794) );
  AND2_X1 U11938 ( .A1(n17872), .A2(n16539), .ZN(n10166) );
  AND2_X1 U11939 ( .A1(n12788), .A2(n10165), .ZN(n17701) );
  INV_X1 U11940 ( .A(n17700), .ZN(n10165) );
  AOI22_X1 U11941 ( .A1(n18793), .A2(n21189), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12914) );
  OAI211_X1 U11942 ( .C1(n12910), .C2(n18323), .A(n9954), .B(n9953), .ZN(
        n12912) );
  NAND2_X1 U11943 ( .A1(n12909), .A2(n18323), .ZN(n9953) );
  INV_X1 U11944 ( .A(n12908), .ZN(n9954) );
  AOI21_X1 U11945 ( .B1(n17468), .B2(n12773), .A(n17872), .ZN(n12776) );
  NAND2_X1 U11946 ( .A1(n10169), .A2(n10168), .ZN(n12775) );
  AOI21_X1 U11947 ( .B1(n10170), .B2(n10176), .A(n9807), .ZN(n10169) );
  XNOR2_X1 U11948 ( .A(n12759), .B(n17491), .ZN(n12760) );
  NOR2_X1 U11949 ( .A1(n12912), .A2(n18766), .ZN(n18756) );
  INV_X1 U11950 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14067) );
  OR2_X1 U11951 ( .A1(n14856), .A2(n12636), .ZN(n12536) );
  OR2_X1 U11952 ( .A1(n14789), .A2(n13217), .ZN(n13228) );
  INV_X1 U11953 ( .A(n14327), .ZN(n13927) );
  AND2_X1 U11954 ( .A1(n13421), .A2(n13208), .ZN(n13404) );
  AND2_X1 U11955 ( .A1(n20839), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12644) );
  NOR2_X1 U11956 ( .A1(n12596), .A2(n14827), .ZN(n12597) );
  OR2_X1 U11957 ( .A1(n12555), .A2(n14845), .ZN(n12557) );
  OR2_X1 U11958 ( .A1(n12557), .A2(n12556), .ZN(n12596) );
  AND2_X1 U11959 ( .A1(n12465), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12466) );
  INV_X1 U11960 ( .A(n12464), .ZN(n12465) );
  AND2_X1 U11961 ( .A1(n12495), .A2(n12494), .ZN(n14697) );
  OR2_X1 U11962 ( .A1(n16051), .A2(n12636), .ZN(n12429) );
  NAND2_X1 U11963 ( .A1(n12376), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12430) );
  NOR2_X1 U11964 ( .A1(n12342), .A2(n12341), .ZN(n12359) );
  CLKBUF_X1 U11965 ( .A(n14332), .Z(n14341) );
  OR2_X1 U11966 ( .A1(n12301), .A2(n16095), .ZN(n12307) );
  INV_X1 U11967 ( .A(n12305), .ZN(n10024) );
  AND2_X1 U11968 ( .A1(n12262), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12263) );
  CLKBUF_X1 U11969 ( .A(n14224), .Z(n14272) );
  AND2_X1 U11970 ( .A1(n12202), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12232) );
  INV_X1 U11971 ( .A(n12185), .ZN(n12186) );
  NAND2_X1 U11972 ( .A1(n12186), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12194) );
  NAND2_X1 U11973 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12168) );
  NOR2_X1 U11974 ( .A1(n12168), .A2(n14067), .ZN(n12177) );
  NAND2_X1 U11975 ( .A1(n10107), .A2(n20320), .ZN(n10106) );
  NAND2_X1 U11976 ( .A1(n10108), .A2(n11913), .ZN(n13710) );
  NAND2_X1 U11977 ( .A1(n13710), .A2(n13708), .ZN(n13709) );
  INV_X1 U11978 ( .A(n13654), .ZN(n12166) );
  INV_X1 U11979 ( .A(n10109), .ZN(n14808) );
  AND2_X1 U11980 ( .A1(n14816), .A2(n9934), .ZN(n14820) );
  AOI21_X1 U11981 ( .B1(n14882), .B2(n15138), .A(n10125), .ZN(n10124) );
  NAND2_X1 U11982 ( .A1(n10126), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10125) );
  NAND2_X1 U11983 ( .A1(n15138), .A2(n12066), .ZN(n10126) );
  INV_X1 U11984 ( .A(n14993), .ZN(n9937) );
  NAND2_X1 U11985 ( .A1(n9974), .A2(n9973), .ZN(n9972) );
  INV_X1 U11986 ( .A(n14713), .ZN(n9973) );
  NOR2_X1 U11987 ( .A1(n14663), .A2(n9975), .ZN(n9974) );
  OR2_X1 U11988 ( .A1(n9785), .A2(n14722), .ZN(n14724) );
  OR3_X1 U11989 ( .A1(n9820), .A2(n13043), .A3(n9971), .ZN(n9970) );
  INV_X1 U11990 ( .A(n14677), .ZN(n9971) );
  NAND2_X1 U11991 ( .A1(n12061), .A2(n14917), .ZN(n15086) );
  NOR3_X1 U11992 ( .A1(n14279), .A2(n9820), .A3(n13043), .ZN(n14678) );
  NOR2_X1 U11993 ( .A1(n14279), .A2(n13043), .ZN(n14348) );
  OR2_X1 U11994 ( .A1(n14324), .A2(n14325), .ZN(n14279) );
  NOR2_X1 U11995 ( .A1(n9968), .A2(n9967), .ZN(n14303) );
  INV_X1 U11996 ( .A(n14221), .ZN(n9967) );
  NAND2_X1 U11997 ( .A1(n14303), .A2(n14302), .ZN(n14324) );
  NAND2_X1 U11998 ( .A1(n15138), .A2(n12049), .ZN(n14264) );
  INV_X1 U11999 ( .A(n10110), .ZN(n9927) );
  AOI21_X1 U12000 ( .B1(n14244), .B2(n10114), .A(n10113), .ZN(n10112) );
  NAND2_X1 U12001 ( .A1(n16209), .A2(n9965), .ZN(n14233) );
  NAND2_X1 U12002 ( .A1(n16209), .A2(n14019), .ZN(n14114) );
  NOR2_X1 U12003 ( .A1(n16207), .A2(n16206), .ZN(n16209) );
  NOR2_X1 U12004 ( .A1(n13109), .A2(n14238), .ZN(n15123) );
  OR2_X1 U12005 ( .A1(n13825), .A2(n13819), .ZN(n16207) );
  OR2_X1 U12006 ( .A1(n13827), .A2(n13828), .ZN(n13825) );
  AND2_X1 U12007 ( .A1(n13651), .A2(n13650), .ZN(n13775) );
  NAND2_X1 U12008 ( .A1(n13775), .A2(n13774), .ZN(n13827) );
  NAND2_X1 U12009 ( .A1(n12147), .A2(n12148), .ZN(n12152) );
  NAND2_X1 U12010 ( .A1(n11846), .A2(n13843), .ZN(n13704) );
  NOR2_X1 U12011 ( .A1(n11804), .A2(n11783), .ZN(n12984) );
  NOR2_X1 U12012 ( .A1(n11783), .A2(n14042), .ZN(n10103) );
  INV_X1 U12013 ( .A(n20667), .ZN(n20809) );
  INV_X1 U12014 ( .A(n20642), .ZN(n15236) );
  NOR2_X1 U12015 ( .A1(n20672), .A2(n15166), .ZN(n20811) );
  NOR2_X1 U12016 ( .A1(n11694), .A2(n11693), .ZN(n11701) );
  AND2_X1 U12017 ( .A1(n15166), .A2(n15167), .ZN(n14162) );
  NAND3_X1 U12018 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n9918), .A3(n13849), 
        .ZN(n15178) );
  AOI21_X1 U12019 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20547), .A(n15174), 
        .ZN(n20673) );
  AND2_X1 U12020 ( .A1(n11213), .A2(n11207), .ZN(n11415) );
  NAND2_X1 U12021 ( .A1(n9877), .A2(n9879), .ZN(n11410) );
  NAND2_X1 U12022 ( .A1(n11431), .A2(n11201), .ZN(n9879) );
  NAND2_X1 U12023 ( .A1(n11202), .A2(n10137), .ZN(n9877) );
  OR2_X1 U12024 ( .A1(n11421), .A2(n10858), .ZN(n16477) );
  NAND2_X1 U12025 ( .A1(n11378), .A2(n11379), .ZN(n11384) );
  AND2_X1 U12027 ( .A1(n10061), .A2(n16327), .ZN(n10059) );
  NOR2_X1 U12028 ( .A1(n9891), .A2(n9892), .ZN(n9890) );
  INV_X1 U12029 ( .A(n11366), .ZN(n9891) );
  NAND2_X1 U12030 ( .A1(n11329), .A2(n11315), .ZN(n11338) );
  OR2_X1 U12031 ( .A1(n19035), .A2(n19036), .ZN(n10072) );
  AND2_X1 U12032 ( .A1(n11344), .A2(n11347), .ZN(n19070) );
  INV_X1 U12033 ( .A(n11575), .ZN(n14092) );
  NOR2_X1 U12034 ( .A1(n19175), .A2(n19172), .ZN(n19159) );
  NAND2_X1 U12035 ( .A1(n11212), .A2(n9888), .ZN(n11237) );
  INV_X1 U12036 ( .A(n9889), .ZN(n9888) );
  OAI21_X1 U12037 ( .B1(n11214), .B2(n11213), .A(n11211), .ZN(n9889) );
  NAND2_X1 U12038 ( .A1(n11224), .A2(n11225), .ZN(n11223) );
  INV_X1 U12039 ( .A(n15260), .ZN(n10140) );
  NOR2_X1 U12040 ( .A1(n10792), .A2(n10814), .ZN(n10161) );
  INV_X1 U12041 ( .A(n10814), .ZN(n10162) );
  NOR2_X1 U12042 ( .A1(n15373), .A2(n15364), .ZN(n15366) );
  OR2_X1 U12043 ( .A1(n15383), .A2(n15371), .ZN(n15373) );
  AND2_X1 U12044 ( .A1(n10152), .A2(n10148), .ZN(n10146) );
  INV_X1 U12045 ( .A(n15293), .ZN(n10148) );
  NAND2_X1 U12046 ( .A1(n11050), .A2(n11049), .ZN(n15400) );
  AND2_X1 U12047 ( .A1(n15322), .A2(n15306), .ZN(n15313) );
  NAND2_X1 U12048 ( .A1(n11040), .A2(n11039), .ZN(n15430) );
  NAND2_X1 U12049 ( .A1(n11040), .A2(n10013), .ZN(n15432) );
  NOR2_X1 U12050 ( .A1(n15339), .A2(n15340), .ZN(n15338) );
  OR2_X1 U12051 ( .A1(n16396), .A2(n9822), .ZN(n16384) );
  INV_X1 U12052 ( .A(n13340), .ZN(n15880) );
  INV_X1 U12053 ( .A(n15640), .ZN(n9996) );
  AND2_X1 U12054 ( .A1(n15482), .A2(n15489), .ZN(n9895) );
  AND2_X1 U12055 ( .A1(n9851), .A2(n15390), .ZN(n10007) );
  AND2_X1 U12056 ( .A1(n11040), .A2(n9839), .ZN(n15415) );
  INV_X1 U12057 ( .A(n14396), .ZN(n10012) );
  OR2_X1 U12058 ( .A1(n19017), .A2(n11360), .ZN(n14513) );
  INV_X1 U12059 ( .A(n10193), .ZN(n14514) );
  INV_X1 U12060 ( .A(n10198), .ZN(n10196) );
  OAI21_X1 U12061 ( .B1(n10198), .B2(n10195), .A(n10197), .ZN(n10194) );
  INV_X1 U12062 ( .A(n14466), .ZN(n10201) );
  NOR2_X1 U12063 ( .A1(n14389), .A2(n10200), .ZN(n10199) );
  INV_X1 U12064 ( .A(n14444), .ZN(n10200) );
  OR3_X1 U12065 ( .A1(n19060), .A2(n11322), .A3(n16329), .ZN(n16330) );
  INV_X1 U12066 ( .A(n15555), .ZN(n16328) );
  NAND2_X1 U12067 ( .A1(n15604), .A2(n10204), .ZN(n10203) );
  OR2_X1 U12068 ( .A1(n10005), .A2(n15794), .ZN(n10004) );
  NAND2_X1 U12069 ( .A1(n15602), .A2(n15601), .ZN(n15600) );
  AND2_X1 U12070 ( .A1(n11561), .A2(n11560), .ZN(n13762) );
  XNOR2_X1 U12071 ( .A(n11522), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15807) );
  OR2_X1 U12072 ( .A1(n14507), .A2(n10094), .ZN(n13761) );
  AND2_X1 U12073 ( .A1(n11552), .A2(n11551), .ZN(n13620) );
  NOR2_X1 U12074 ( .A1(n14507), .A2(n13620), .ZN(n13637) );
  NAND2_X1 U12075 ( .A1(n9865), .A2(n11514), .ZN(n15616) );
  AND2_X1 U12076 ( .A1(n13892), .A2(n16442), .ZN(n10009) );
  NAND2_X1 U12077 ( .A1(n10102), .A2(n11537), .ZN(n14008) );
  NAND2_X1 U12078 ( .A1(n11536), .A2(n11535), .ZN(n11537) );
  INV_X1 U12079 ( .A(n9898), .ZN(n9897) );
  OAI21_X1 U12080 ( .B1(n9905), .B2(n9899), .A(n9904), .ZN(n9898) );
  NAND2_X1 U12081 ( .A1(n13891), .A2(n13892), .ZN(n16445) );
  INV_X1 U12082 ( .A(n13592), .ZN(n10932) );
  INV_X1 U12083 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13837) );
  XNOR2_X1 U12084 ( .A(n10420), .B(n10418), .ZN(n13586) );
  AND2_X1 U12085 ( .A1(n20072), .A2(n19407), .ZN(n19695) );
  AND2_X1 U12086 ( .A1(n15893), .A2(n20086), .ZN(n19549) );
  INV_X1 U12087 ( .A(n19695), .ZN(n19692) );
  OR2_X1 U12088 ( .A1(n15893), .A2(n20086), .ZN(n19841) );
  INV_X1 U12089 ( .A(n19725), .ZN(n19789) );
  NOR2_X1 U12090 ( .A1(n15880), .A2(n15879), .ZN(n19450) );
  NOR2_X1 U12091 ( .A1(n15878), .A2(n15879), .ZN(n19451) );
  OR2_X1 U12092 ( .A1(n19841), .A2(n19840), .ZN(n19869) );
  NAND2_X1 U12093 ( .A1(n10274), .A2(n10456), .ZN(n10281) );
  INV_X1 U12094 ( .A(n10447), .ZN(n19442) );
  INV_X1 U12095 ( .A(n19450), .ZN(n19448) );
  INV_X1 U12096 ( .A(n19451), .ZN(n19446) );
  OR2_X1 U12097 ( .A1(n19841), .A2(n15894), .ZN(n19409) );
  OR2_X1 U12098 ( .A1(n19725), .A2(n15894), .ZN(n19870) );
  NAND2_X1 U12099 ( .A1(n16506), .A2(n15875), .ZN(n19453) );
  INV_X1 U12100 ( .A(n15894), .ZN(n15885) );
  NOR2_X1 U12101 ( .A1(n16684), .A2(n16683), .ZN(n18747) );
  AND2_X1 U12102 ( .A1(n10032), .A2(n9829), .ZN(n16790) );
  INV_X1 U12103 ( .A(n12848), .ZN(n9876) );
  NAND2_X1 U12104 ( .A1(n15921), .A2(n18772), .ZN(n16683) );
  OR2_X1 U12105 ( .A1(n12832), .A2(n12831), .ZN(n17500) );
  INV_X1 U12106 ( .A(n17537), .ZN(n17501) );
  NOR3_X1 U12107 ( .A1(n17609), .A2(n16728), .A3(n10048), .ZN(n16524) );
  NOR2_X1 U12108 ( .A1(n17609), .A2(n16749), .ZN(n17608) );
  NOR3_X1 U12109 ( .A1(n17609), .A2(n16749), .A3(n17954), .ZN(n16688) );
  NOR2_X1 U12110 ( .A1(n10047), .A2(n10046), .ZN(n10045) );
  NOR2_X1 U12111 ( .A1(n16695), .A2(n17688), .ZN(n17687) );
  NAND3_X1 U12112 ( .A1(n17723), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16695) );
  AND2_X1 U12113 ( .A1(n17854), .A2(n10050), .ZN(n17775) );
  NAND2_X1 U12114 ( .A1(n17854), .A2(n10222), .ZN(n17808) );
  NOR2_X1 U12115 ( .A1(n17878), .A2(n17879), .ZN(n17854) );
  AND2_X1 U12116 ( .A1(n17901), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17890) );
  NAND2_X1 U12117 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17011) );
  INV_X1 U12118 ( .A(n17011), .ZN(n17923) );
  NOR3_X1 U12119 ( .A1(n16538), .A2(n12795), .A3(n12794), .ZN(n12796) );
  AOI21_X1 U12120 ( .B1(n12793), .B2(n17802), .A(n12794), .ZN(n16009) );
  AND2_X1 U12121 ( .A1(n12788), .A2(n12787), .ZN(n17659) );
  NOR2_X1 U12122 ( .A1(n17701), .A2(n10163), .ZN(n17667) );
  NAND2_X1 U12123 ( .A1(n10164), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10163) );
  INV_X1 U12124 ( .A(n17984), .ZN(n10164) );
  INV_X1 U12125 ( .A(n12788), .ZN(n17712) );
  NOR2_X1 U12126 ( .A1(n9949), .A2(n9948), .ZN(n9947) );
  NAND2_X1 U12127 ( .A1(n17352), .A2(n17349), .ZN(n15928) );
  INV_X1 U12128 ( .A(n18162), .ZN(n18140) );
  INV_X1 U12129 ( .A(n18767), .ZN(n18774) );
  NOR2_X1 U12130 ( .A1(n17828), .A2(n18199), .ZN(n18163) );
  NOR2_X1 U12131 ( .A1(n17869), .A2(n18199), .ZN(n17868) );
  NAND2_X1 U12132 ( .A1(n10178), .A2(n10179), .ZN(n17870) );
  NOR2_X1 U12133 ( .A1(n12778), .A2(n17802), .ZN(n10178) );
  NOR2_X1 U12134 ( .A1(n17791), .A2(n12778), .ZN(n17871) );
  XNOR2_X1 U12135 ( .A(n12775), .B(n12774), .ZN(n17882) );
  INV_X1 U12136 ( .A(n12776), .ZN(n12774) );
  NAND2_X1 U12137 ( .A1(n17882), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17881) );
  NOR2_X1 U12138 ( .A1(n12935), .A2(n17920), .ZN(n17904) );
  NOR2_X1 U12139 ( .A1(n17904), .A2(n17903), .ZN(n17902) );
  NOR2_X1 U12140 ( .A1(n18243), .A2(n17921), .ZN(n17920) );
  XNOR2_X1 U12141 ( .A(n12765), .B(n12764), .ZN(n17928) );
  NAND2_X1 U12142 ( .A1(n17928), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17927) );
  XOR2_X1 U12143 ( .A(n12757), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n17951) );
  AND2_X1 U12144 ( .A1(n9873), .A2(n9872), .ZN(n21180) );
  NAND2_X1 U12145 ( .A1(n21189), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9872) );
  NAND2_X1 U12146 ( .A1(n18940), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9873) );
  OAI21_X1 U12147 ( .B1(n18790), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n9871), .ZN(n21186) );
  OR2_X1 U12148 ( .A1(n18791), .A2(n21180), .ZN(n9871) );
  NOR2_X1 U12149 ( .A1(n18972), .A2(n15923), .ZN(n18785) );
  INV_X1 U12150 ( .A(n18785), .ZN(n18757) );
  NAND2_X1 U12151 ( .A1(n18767), .A2(n18756), .ZN(n18772) );
  INV_X1 U12152 ( .A(n17500), .ZN(n18308) );
  NOR2_X2 U12153 ( .A1(n12822), .A2(n12821), .ZN(n18313) );
  INV_X1 U12154 ( .A(n15929), .ZN(n18318) );
  NOR2_X1 U12155 ( .A1(n12882), .A2(n12881), .ZN(n18328) );
  NOR2_X1 U12156 ( .A1(n12862), .A2(n12861), .ZN(n18334) );
  AOI22_X1 U12157 ( .A1(n18745), .A2(n18744), .B1(n18749), .B2(n16553), .ZN(
        n18753) );
  NAND2_X1 U12158 ( .A1(n14567), .A2(n14565), .ZN(n20844) );
  OR2_X1 U12159 ( .A1(n20203), .A2(n14123), .ZN(n20196) );
  NOR2_X2 U12160 ( .A1(n14037), .A2(n14036), .ZN(n20185) );
  NAND2_X1 U12161 ( .A1(n14047), .A2(n14043), .ZN(n20194) );
  AND2_X1 U12162 ( .A1(n14112), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20193) );
  AND2_X1 U12163 ( .A1(n14037), .A2(n14035), .ZN(n20162) );
  OR2_X1 U12164 ( .A1(n14570), .A2(n13093), .ZN(n14690) );
  INV_X1 U12165 ( .A(n14701), .ZN(n20223) );
  INV_X1 U12166 ( .A(n20227), .ZN(n14716) );
  AND2_X1 U12167 ( .A1(n20227), .A2(n13854), .ZN(n20222) );
  INV_X1 U12168 ( .A(n20222), .ZN(n14725) );
  INV_X1 U12169 ( .A(n14829), .ZN(n14743) );
  INV_X1 U12170 ( .A(n14793), .ZN(n14801) );
  INV_X1 U12171 ( .A(n20250), .ZN(n20228) );
  NOR2_X1 U12172 ( .A1(n20228), .A2(n20847), .ZN(n20239) );
  XNOR2_X1 U12174 ( .A(n14418), .B(n14568), .ZN(n14815) );
  AOI21_X1 U12175 ( .B1(n14419), .B2(n14417), .A(n14418), .ZN(n14689) );
  AOI21_X1 U12176 ( .B1(n14322), .B2(n14321), .A(n14320), .ZN(n16139) );
  AND2_X1 U12177 ( .A1(n14013), .A2(n14015), .ZN(n20224) );
  INV_X1 U12178 ( .A(n14954), .ZN(n20293) );
  INV_X1 U12179 ( .A(n20298), .ZN(n16141) );
  OR2_X1 U12180 ( .A1(n16231), .A2(n13730), .ZN(n14954) );
  INV_X1 U12181 ( .A(n20139), .ZN(n20294) );
  OAI22_X1 U12182 ( .A1(n14570), .A2(n13064), .B1(n14632), .B2(n9958), .ZN(
        n14572) );
  OR2_X1 U12183 ( .A1(n13087), .A2(n9959), .ZN(n9958) );
  NAND2_X1 U12184 ( .A1(n9962), .A2(n9960), .ZN(n9959) );
  NAND2_X1 U12185 ( .A1(n9936), .A2(n15138), .ZN(n14842) );
  NOR2_X1 U12186 ( .A1(n15015), .A2(n13130), .ZN(n15004) );
  NAND2_X1 U12187 ( .A1(n9935), .A2(n14861), .ZN(n14860) );
  OAI21_X1 U12188 ( .B1(n14882), .B2(n12066), .A(n15138), .ZN(n14874) );
  AND2_X1 U12189 ( .A1(n15067), .A2(n10221), .ZN(n15046) );
  NAND2_X1 U12190 ( .A1(n16153), .A2(n12031), .ZN(n10116) );
  AND2_X1 U12191 ( .A1(n15124), .A2(n20314), .ZN(n15100) );
  AND2_X1 U12192 ( .A1(n13120), .A2(n12998), .ZN(n20312) );
  INV_X1 U12193 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20547) );
  NAND2_X1 U12194 ( .A1(n9933), .A2(n11931), .ZN(n13415) );
  OAI22_X1 U12195 ( .A1(n20336), .A2(n20335), .B1(n20520), .B2(n20433), .ZN(
        n20352) );
  NAND2_X1 U12196 ( .A1(n20391), .A2(n13948), .ZN(n20385) );
  INV_X1 U12197 ( .A(n20508), .ZN(n20511) );
  OAI211_X1 U12198 ( .C1(n20541), .C2(n20526), .A(n20525), .B(n20524), .ZN(
        n20544) );
  INV_X1 U12199 ( .A(n20515), .ZN(n20543) );
  INV_X1 U12200 ( .A(n20636), .ZN(n20623) );
  NAND2_X1 U12201 ( .A1(n20812), .A2(n20493), .ZN(n20636) );
  INV_X1 U12202 ( .A(n20410), .ZN(n20692) );
  NOR2_X2 U12203 ( .A1(n20672), .A2(n20327), .ZN(n20721) );
  NOR2_X1 U12204 ( .A1(n13429), .A2(n20526), .ZN(n20803) );
  INV_X1 U12205 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20727) );
  NOR2_X1 U12206 ( .A1(n15952), .A2(n10058), .ZN(n16306) );
  AND2_X1 U12207 ( .A1(n10057), .A2(n10055), .ZN(n10054) );
  INV_X1 U12208 ( .A(n14524), .ZN(n10055) );
  NOR2_X1 U12209 ( .A1(n19010), .A2(n10058), .ZN(n19000) );
  NAND2_X1 U12210 ( .A1(n10071), .A2(n10070), .ZN(n19024) );
  NAND2_X1 U12211 ( .A1(n10058), .A2(n15544), .ZN(n10070) );
  AND2_X1 U12212 ( .A1(n10072), .A2(n19173), .ZN(n19023) );
  CLKBUF_X1 U12213 ( .A(n19211), .Z(n19166) );
  INV_X1 U12214 ( .A(n19187), .ZN(n19199) );
  INV_X1 U12215 ( .A(n19154), .ZN(n19204) );
  CLKBUF_X1 U12216 ( .A(n11101), .Z(n15861) );
  OR2_X1 U12217 ( .A1(n13193), .A2(n13192), .ZN(n19169) );
  NOR2_X1 U12218 ( .A1(n13596), .A2(n13595), .ZN(n19274) );
  NAND2_X1 U12219 ( .A1(n10142), .A2(n10139), .ZN(n15259) );
  NOR2_X1 U12220 ( .A1(n15253), .A2(n10143), .ZN(n15261) );
  NOR2_X1 U12221 ( .A1(n10143), .A2(n10140), .ZN(n10139) );
  INV_X1 U12222 ( .A(n15309), .ZN(n15727) );
  NAND2_X1 U12223 ( .A1(n14462), .A2(n10099), .ZN(n15328) );
  AND2_X1 U12224 ( .A1(n14104), .A2(n14103), .ZN(n19078) );
  AND2_X1 U12225 ( .A1(n9791), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10144) );
  NAND2_X1 U12226 ( .A1(n10145), .A2(n13884), .ZN(n14505) );
  INV_X1 U12227 ( .A(n15341), .ZN(n15337) );
  AND2_X1 U12228 ( .A1(n19270), .A2(n11076), .ZN(n16315) );
  AND2_X1 U12229 ( .A1(n13896), .A2(n15878), .ZN(n19215) );
  AND2_X1 U12230 ( .A1(n13896), .A2(n15880), .ZN(n19217) );
  INV_X1 U12231 ( .A(n19263), .ZN(n19272) );
  AND2_X1 U12232 ( .A1(n13301), .A2(n13187), .ZN(n19357) );
  XNOR2_X1 U12233 ( .A(n9801), .B(n11649), .ZN(n14450) );
  INV_X1 U12234 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19145) );
  NAND2_X1 U12235 ( .A1(n14003), .A2(n11508), .ZN(n16377) );
  INV_X1 U12236 ( .A(n11087), .ZN(n13602) );
  XOR2_X1 U12237 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n15457), .Z(
        n15632) );
  INV_X1 U12238 ( .A(n10010), .ZN(n14492) );
  OAI21_X1 U12239 ( .B1(n15359), .B2(n16433), .A(n10011), .ZN(n10010) );
  AND2_X1 U12240 ( .A1(n10230), .A2(n15287), .ZN(n16324) );
  NOR2_X1 U12241 ( .A1(n16396), .A2(n9787), .ZN(n14459) );
  AND2_X1 U12242 ( .A1(n10208), .A2(n9828), .ZN(n15590) );
  NAND2_X1 U12243 ( .A1(n10208), .A2(n11291), .ZN(n15791) );
  INV_X1 U12244 ( .A(n16433), .ZN(n19391) );
  NOR3_X1 U12245 ( .A1(n19396), .A2(n13875), .A3(n13873), .ZN(n16454) );
  INV_X1 U12246 ( .A(n13196), .ZN(n19185) );
  NAND2_X1 U12247 ( .A1(n9906), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13861) );
  NAND2_X1 U12248 ( .A1(n9903), .A2(n13873), .ZN(n13862) );
  INV_X1 U12249 ( .A(n19274), .ZN(n20086) );
  INV_X1 U12250 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20076) );
  NAND2_X1 U12251 ( .A1(n13598), .A2(n13601), .ZN(n20079) );
  INV_X1 U12252 ( .A(n16478), .ZN(n13749) );
  NAND2_X1 U12253 ( .A1(n13584), .A2(n13587), .ZN(n20072) );
  OR2_X1 U12254 ( .A1(n13586), .A2(n13585), .ZN(n13587) );
  INV_X1 U12255 ( .A(n15835), .ZN(n16494) );
  XNOR2_X1 U12256 ( .A(n13568), .B(n13569), .ZN(n15893) );
  INV_X1 U12257 ( .A(n19496), .ZN(n19514) );
  INV_X1 U12258 ( .A(n19490), .ZN(n19513) );
  OAI21_X1 U12259 ( .B1(n19635), .B2(n19879), .A(n19619), .ZN(n19638) );
  OR2_X1 U12260 ( .A1(n15869), .A2(n15868), .ZN(n19659) );
  OAI21_X1 U12261 ( .B1(n19686), .B2(n19665), .A(n19883), .ZN(n19688) );
  OAI21_X1 U12262 ( .B1(n19734), .B2(n19749), .A(n19883), .ZN(n19752) );
  INV_X1 U12263 ( .A(n19724), .ZN(n19751) );
  INV_X1 U12264 ( .A(n19918), .ZN(n19806) );
  INV_X1 U12265 ( .A(n19937), .ZN(n19815) );
  INV_X1 U12266 ( .A(n19408), .ZN(n19876) );
  INV_X1 U12267 ( .A(n19869), .ZN(n19909) );
  INV_X1 U12268 ( .A(n19847), .ZN(n19917) );
  OAI22_X1 U12269 ( .A1(n19426), .A2(n19446), .B1(n20927), .B2(n19448), .ZN(
        n19924) );
  INV_X1 U12270 ( .A(n19850), .ZN(n19923) );
  OAI22_X1 U12271 ( .A1(n21048), .A2(n19446), .B1(n20915), .B2(n19448), .ZN(
        n19937) );
  INV_X1 U12272 ( .A(n19856), .ZN(n19936) );
  INV_X1 U12273 ( .A(n19901), .ZN(n19935) );
  INV_X1 U12274 ( .A(n19859), .ZN(n19944) );
  INV_X1 U12275 ( .A(n19868), .ZN(n19957) );
  INV_X1 U12276 ( .A(n19409), .ZN(n19960) );
  INV_X1 U12277 ( .A(n19870), .ZN(n19958) );
  XOR2_X1 U12278 ( .A(n18313), .B(n18308), .Z(n18972) );
  NOR2_X1 U12279 ( .A1(n18747), .A2(n17538), .ZN(n18973) );
  INV_X1 U12280 ( .A(n16719), .ZN(n10043) );
  INV_X1 U12281 ( .A(n16724), .ZN(n10040) );
  NAND2_X1 U12282 ( .A1(n10039), .A2(n10038), .ZN(n10037) );
  NOR2_X1 U12283 ( .A1(n16722), .A2(n16721), .ZN(n10038) );
  OR2_X1 U12284 ( .A1(n16732), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n10039) );
  NOR2_X1 U12285 ( .A1(n16768), .A2(n17029), .ZN(n16761) );
  NOR2_X1 U12286 ( .A1(n16761), .A2(n16762), .ZN(n16760) );
  INV_X1 U12287 ( .A(n17050), .ZN(n17057) );
  AND2_X1 U12288 ( .A1(n10035), .A2(n10031), .ZN(n16808) );
  INV_X1 U12289 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17024) );
  NOR2_X1 U12290 ( .A1(n18810), .A2(n16686), .ZN(n17050) );
  INV_X1 U12291 ( .A(n17053), .ZN(n17054) );
  INV_X1 U12292 ( .A(n17371), .ZN(n17368) );
  NAND2_X1 U12293 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17368), .ZN(n17367) );
  NAND2_X1 U12294 ( .A1(n17381), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n17371) );
  NOR2_X1 U12295 ( .A1(n17382), .A2(n17559), .ZN(n17381) );
  NOR2_X1 U12296 ( .A1(n17388), .A2(n17431), .ZN(n17383) );
  NAND2_X1 U12297 ( .A1(n17383), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n17382) );
  NOR4_X1 U12298 ( .A1(n17553), .A2(n17544), .A3(n17426), .A4(n17398), .ZN(
        n17389) );
  NAND2_X1 U12299 ( .A1(n17427), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17426) );
  NAND2_X1 U12300 ( .A1(n9946), .A2(n9944), .ZN(n17432) );
  NOR2_X1 U12301 ( .A1(n17348), .A2(n9945), .ZN(n9944) );
  INV_X1 U12302 ( .A(n17464), .ZN(n9946) );
  INV_X1 U12303 ( .A(n18348), .ZN(n17431) );
  NOR2_X1 U12304 ( .A1(n12743), .A2(n12742), .ZN(n17472) );
  INV_X1 U12305 ( .A(n12921), .ZN(n17475) );
  INV_X1 U12306 ( .A(n12920), .ZN(n12762) );
  CLKBUF_X1 U12307 ( .A(n17514), .Z(n17534) );
  CLKBUF_X1 U12308 ( .A(n18954), .Z(n17535) );
  NOR2_X1 U12309 ( .A1(n18313), .A2(n17600), .ZN(n17593) );
  BUF_X1 U12310 ( .A(n17597), .Z(n17600) );
  CLKBUF_X1 U12311 ( .A(n17593), .Z(n17601) );
  NAND2_X1 U12312 ( .A1(n17687), .A2(n9783), .ZN(n17638) );
  NAND2_X1 U12313 ( .A1(n17687), .A2(n10226), .ZN(n17673) );
  AOI21_X1 U12314 ( .B1(n17732), .B2(n9870), .A(n9868), .ZN(n17722) );
  INV_X1 U12315 ( .A(n18063), .ZN(n9870) );
  OAI21_X1 U12316 ( .B1(n17735), .B2(n20926), .A(n9869), .ZN(n9868) );
  NAND2_X1 U12317 ( .A1(n17873), .A2(n18057), .ZN(n9869) );
  NOR2_X1 U12318 ( .A1(n17769), .A2(n18029), .ZN(n17732) );
  NAND2_X1 U12319 ( .A1(n17854), .A2(n9786), .ZN(n17751) );
  NOR2_X1 U12320 ( .A1(n18159), .A2(n12953), .ZN(n18102) );
  INV_X1 U12321 ( .A(n17862), .ZN(n17834) );
  NAND2_X1 U12322 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17890), .ZN(
        n17878) );
  NOR2_X1 U12323 ( .A1(n9796), .A2(n18313), .ZN(n17910) );
  NOR2_X1 U12324 ( .A1(n17011), .A2(n17024), .ZN(n17901) );
  INV_X1 U12325 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17932) );
  BUF_X1 U12326 ( .A(n18340), .Z(n18349) );
  INV_X1 U12327 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17949) );
  NAND2_X1 U12328 ( .A1(n17624), .A2(n17606), .ZN(n15943) );
  INV_X1 U12329 ( .A(n18196), .ZN(n18125) );
  NAND2_X1 U12330 ( .A1(n18755), .A2(n18757), .ZN(n18270) );
  INV_X1 U12331 ( .A(n18254), .ZN(n18236) );
  NAND2_X1 U12332 ( .A1(n10173), .A2(n10170), .ZN(n17892) );
  NAND2_X1 U12333 ( .A1(n10175), .A2(n10174), .ZN(n10173) );
  NOR2_X1 U12334 ( .A1(n17906), .A2(n17907), .ZN(n17905) );
  INV_X1 U12335 ( .A(n18216), .ZN(n18282) );
  INV_X1 U12336 ( .A(n18789), .ZN(n18287) );
  INV_X1 U12337 ( .A(n18271), .ZN(n18286) );
  INV_X1 U12338 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18935) );
  CLKBUF_X1 U12339 ( .A(n18900), .Z(n18893) );
  AND2_X1 U12340 ( .A1(n13227), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14327)
         );
  INV_X1 U12342 ( .A(n12654), .ZN(n10017) );
  OAI21_X1 U12343 ( .B1(n16252), .B2(n10077), .A(n10074), .ZN(P2_U2826) );
  INV_X1 U12344 ( .A(n10078), .ZN(n10077) );
  NAND2_X1 U12345 ( .A1(n16255), .A2(n19203), .ZN(n10075) );
  OAI21_X1 U12346 ( .B1(n15630), .B2(n15344), .A(n12657), .ZN(n12658) );
  NAND2_X1 U12347 ( .A1(n10867), .A2(n10158), .ZN(n10157) );
  OAI21_X1 U12348 ( .B1(n15722), .B2(n19385), .A(n14531), .ZN(n14532) );
  INV_X1 U12349 ( .A(n14530), .ZN(n14531) );
  INV_X1 U12350 ( .A(n10079), .ZN(n14415) );
  AOI21_X1 U12351 ( .B1(n14414), .B2(n19382), .A(n14413), .ZN(n10080) );
  AOI21_X1 U12352 ( .B1(n15553), .B2(n19382), .A(n15552), .ZN(n9913) );
  NAND2_X1 U12353 ( .A1(n9746), .A2(n16378), .ZN(n9914) );
  NAND2_X1 U12354 ( .A1(n14456), .A2(n16450), .ZN(n10187) );
  AOI211_X1 U12355 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15643), .A(
        n15642), .B(n15641), .ZN(n15646) );
  OAI211_X1 U12356 ( .C1(n19406), .C2(n14412), .A(n9834), .B(n10000), .ZN(
        P2_U3027) );
  AND2_X1 U12357 ( .A1(n15752), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10001) );
  INV_X1 U12358 ( .A(n16668), .ZN(n16663) );
  AOI21_X1 U12359 ( .B1(n16713), .B2(n16712), .A(n16711), .ZN(n16714) );
  NAND2_X1 U12360 ( .A1(n10041), .A2(n10036), .ZN(P3_U2641) );
  NAND2_X1 U12361 ( .A1(n10042), .A2(n17056), .ZN(n10041) );
  NOR2_X1 U12362 ( .A1(n10040), .A2(n10037), .ZN(n10036) );
  XNOR2_X1 U12363 ( .A(n16718), .B(n10043), .ZN(n10042) );
  AOI21_X1 U12364 ( .B1(n9943), .B2(P3_EAX_REG_31__SCAN_IN), .A(n9942), .ZN(
        n17350) );
  AND2_X1 U12365 ( .A1(n17424), .A2(BUF2_REG_31__SCAN_IN), .ZN(n9942) );
  AOI21_X1 U12366 ( .B1(n17493), .B2(BUF2_REG_0__SCAN_IN), .A(n10180), .ZN(
        n16025) );
  AND2_X1 U12367 ( .A1(n17492), .A2(n10181), .ZN(n10180) );
  OAI211_X1 U12368 ( .C1(n16550), .C2(n17966), .A(n12963), .B(n12962), .ZN(
        n12964) );
  AND2_X1 U12369 ( .A1(n11050), .A2(n9849), .ZN(n9781) );
  AND2_X1 U12370 ( .A1(n11050), .A2(n9851), .ZN(n9782) );
  AND2_X1 U12371 ( .A1(n9790), .A2(n10045), .ZN(n9783) );
  OR2_X1 U12372 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n9784) );
  OR2_X1 U12373 ( .A1(n15076), .A2(n15075), .ZN(n9785) );
  NAND2_X1 U12374 ( .A1(n10063), .A2(n10067), .ZN(n13169) );
  NAND2_X1 U12375 ( .A1(n17870), .A2(n10177), .ZN(n12784) );
  OR2_X1 U12376 ( .A1(n14292), .A2(n9813), .ZN(n14945) );
  AND2_X1 U12377 ( .A1(n10050), .A2(n10217), .ZN(n9786) );
  INV_X1 U12378 ( .A(n11431), .ZN(n10137) );
  INV_X1 U12379 ( .A(n15876), .ZN(n20109) );
  OR2_X1 U12380 ( .A1(n9822), .A2(n16385), .ZN(n9787) );
  AND2_X1 U12381 ( .A1(n11396), .A2(n10904), .ZN(n9788) );
  NAND2_X1 U12382 ( .A1(n14833), .A2(n12073), .ZN(n12967) );
  INV_X1 U12383 ( .A(n10176), .ZN(n10174) );
  AND2_X1 U12384 ( .A1(n17907), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10176) );
  NAND2_X1 U12385 ( .A1(n16328), .A2(n14522), .ZN(n9789) );
  NAND2_X1 U12386 ( .A1(n11915), .A2(n13917), .ZN(n13061) );
  AND2_X1 U12387 ( .A1(n15784), .A2(n9999), .ZN(n15581) );
  AND2_X1 U12388 ( .A1(n14672), .A2(n9824), .ZN(n14660) );
  AND2_X1 U12389 ( .A1(n15366), .A2(n13291), .ZN(n15348) );
  OR2_X1 U12390 ( .A1(n15813), .A2(n10005), .ZN(n15792) );
  NAND2_X1 U12391 ( .A1(n13944), .A2(n13932), .ZN(n13933) );
  NAND2_X1 U12392 ( .A1(n13944), .A2(n10083), .ZN(n14025) );
  AND2_X1 U12393 ( .A1(n10226), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9790) );
  AND2_X1 U12394 ( .A1(n13884), .A2(n9854), .ZN(n9791) );
  AND2_X1 U12395 ( .A1(n12073), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9792) );
  OR2_X1 U12396 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13298), .ZN(n9793) );
  OR2_X1 U12397 ( .A1(n10160), .A2(n10161), .ZN(n9794) );
  AND2_X1 U12398 ( .A1(n15260), .A2(n15254), .ZN(n9795) );
  INV_X2 U12399 ( .A(n13504), .ZN(n17267) );
  CLKBUF_X3 U12400 ( .A(n13526), .Z(n17278) );
  OR2_X1 U12401 ( .A1(n18753), .A2(n18817), .ZN(n9796) );
  AND2_X1 U12402 ( .A1(n10794), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10572) );
  AND2_X1 U12403 ( .A1(n11754), .A2(n11753), .ZN(n9797) );
  NAND2_X1 U12404 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13177) );
  NAND2_X1 U12405 ( .A1(n14672), .A2(n12410), .ZN(n14703) );
  NAND2_X1 U12406 ( .A1(n14023), .A2(n10532), .ZN(n14099) );
  INV_X2 U12407 ( .A(n12996), .ZN(n11786) );
  NAND2_X1 U12408 ( .A1(n14945), .A2(n12053), .ZN(n14905) );
  NAND2_X1 U12409 ( .A1(n15784), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15586) );
  AND2_X1 U12410 ( .A1(n14627), .A2(n10028), .ZN(n14588) );
  INV_X2 U12411 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10456) );
  NOR2_X1 U12412 ( .A1(n13173), .A2(n19145), .ZN(n13174) );
  INV_X1 U12414 ( .A(n12690), .ZN(n17218) );
  NOR2_X1 U12415 ( .A1(n9930), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11661) );
  NOR2_X1 U12416 ( .A1(n15493), .A2(n15662), .ZN(n9798) );
  OR2_X1 U12417 ( .A1(n10066), .A2(n16358), .ZN(n9799) );
  NAND2_X1 U12418 ( .A1(n11364), .A2(n15522), .ZN(n9800) );
  OAI21_X1 U12419 ( .B1(n15579), .B2(n15577), .A(n15576), .ZN(n16343) );
  INV_X1 U12420 ( .A(n12089), .ZN(n12083) );
  NAND2_X1 U12421 ( .A1(n15262), .A2(n10088), .ZN(n9801) );
  INV_X1 U12422 ( .A(n15492), .ZN(n9894) );
  AND2_X1 U12423 ( .A1(n16257), .A2(n19173), .ZN(n13283) );
  AND3_X1 U12424 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13175) );
  AND2_X1 U12425 ( .A1(n13064), .A2(n9963), .ZN(n9802) );
  INV_X1 U12426 ( .A(n9893), .ZN(n11295) );
  NAND2_X1 U12427 ( .A1(n11288), .A2(n11286), .ZN(n9893) );
  AND3_X1 U12428 ( .A1(n10014), .A2(n9997), .A3(n19879), .ZN(n9803) );
  INV_X1 U12429 ( .A(n10910), .ZN(n10331) );
  AND2_X1 U12430 ( .A1(n10208), .A2(n10206), .ZN(n9804) );
  NAND2_X1 U12431 ( .A1(n9990), .A2(n9989), .ZN(n15502) );
  INV_X1 U12432 ( .A(n9957), .ZN(n14622) );
  NOR2_X1 U12433 ( .A1(n14632), .A2(n14620), .ZN(n9957) );
  AND4_X1 U12434 ( .A1(n12852), .A2(n12851), .A3(n12850), .A4(n12849), .ZN(
        n9805) );
  OR2_X1 U12435 ( .A1(n14833), .A2(n12074), .ZN(n9806) );
  AND2_X1 U12436 ( .A1(n15269), .A2(n15270), .ZN(n15262) );
  AND2_X1 U12437 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12772), .ZN(
        n9807) );
  AND2_X1 U12438 ( .A1(n10135), .A2(n10134), .ZN(n9808) );
  OR2_X1 U12439 ( .A1(n15537), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9809) );
  NAND2_X1 U12440 ( .A1(n15510), .A2(n10216), .ZN(n9810) );
  NAND2_X1 U12441 ( .A1(n15784), .A2(n10073), .ZN(n15587) );
  AND2_X1 U12442 ( .A1(n14023), .A2(n10153), .ZN(n9811) );
  NAND2_X1 U12443 ( .A1(n14672), .A2(n10020), .ZN(n9812) );
  NOR2_X1 U12444 ( .A1(n15138), .A2(n16189), .ZN(n9813) );
  AND3_X1 U12445 ( .A1(n12747), .A2(n12746), .A3(n12745), .ZN(n9814) );
  AND2_X1 U12446 ( .A1(n14627), .A2(n12537), .ZN(n14614) );
  OR2_X1 U12447 ( .A1(n10229), .A2(n19199), .ZN(n9815) );
  AND2_X1 U12448 ( .A1(n10083), .A2(n10082), .ZN(n9816) );
  OR2_X1 U12449 ( .A1(n15086), .A2(n12063), .ZN(n9817) );
  OR2_X1 U12450 ( .A1(n16262), .A2(n11322), .ZN(n14476) );
  AND2_X1 U12451 ( .A1(n11454), .A2(n10333), .ZN(n9818) );
  AND2_X1 U12452 ( .A1(n10213), .A2(n11653), .ZN(n9819) );
  NAND2_X1 U12453 ( .A1(n9803), .A2(n9747), .ZN(n11030) );
  OR2_X1 U12454 ( .A1(n14344), .A2(n14345), .ZN(n9820) );
  NAND2_X1 U12455 ( .A1(n12306), .A2(n14275), .ZN(n10027) );
  INV_X1 U12456 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11655) );
  NAND2_X1 U12457 ( .A1(n15400), .A2(n13246), .ZN(n9821) );
  NAND2_X1 U12458 ( .A1(n13815), .A2(n14014), .ZN(n14013) );
  NAND2_X1 U12459 ( .A1(n14462), .A2(n14463), .ZN(n14434) );
  NAND2_X1 U12461 ( .A1(n10027), .A2(n10025), .ZN(n14250) );
  NOR2_X1 U12465 ( .A1(n13171), .A2(n19123), .ZN(n13172) );
  NOR2_X1 U12466 ( .A1(n13171), .A2(n9799), .ZN(n13170) );
  NAND2_X1 U12467 ( .A1(n11050), .A2(n10007), .ZN(n15380) );
  OAI22_X1 U12468 ( .A1(n14451), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n20119), 
        .B2(n13141), .ZN(n13180) );
  NOR2_X1 U12469 ( .A1(n10230), .A2(n15277), .ZN(n15269) );
  NOR2_X1 U12470 ( .A1(n14013), .A2(n12243), .ZN(n14223) );
  NOR2_X1 U12471 ( .A1(n16396), .A2(n16397), .ZN(n15761) );
  OR2_X1 U12472 ( .A1(n16397), .A2(n10003), .ZN(n9822) );
  NAND2_X1 U12473 ( .A1(n16158), .A2(n12009), .ZN(n16153) );
  AND2_X1 U12474 ( .A1(n13138), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9823) );
  NAND2_X1 U12475 ( .A1(n10116), .A2(n12032), .ZN(n14242) );
  AND2_X1 U12476 ( .A1(n10020), .A2(n12463), .ZN(n9824) );
  AND2_X1 U12477 ( .A1(n13816), .A2(n13817), .ZN(n13815) );
  AND2_X1 U12478 ( .A1(n9823), .A2(n13139), .ZN(n9825) );
  NOR2_X1 U12479 ( .A1(n14724), .A2(n9972), .ZN(n9976) );
  NOR2_X1 U12480 ( .A1(n13823), .A2(n13824), .ZN(n13816) );
  AND2_X1 U12481 ( .A1(n10153), .A2(n10680), .ZN(n9826) );
  OR3_X1 U12482 ( .A1(n14724), .A2(n14713), .A3(n9975), .ZN(n9827) );
  AND2_X1 U12483 ( .A1(n10207), .A2(n11291), .ZN(n9828) );
  AND2_X1 U12484 ( .A1(n10033), .A2(n10031), .ZN(n9829) );
  OR2_X1 U12485 ( .A1(n15366), .A2(n13291), .ZN(n9830) );
  AND2_X1 U12486 ( .A1(n9965), .A2(n9964), .ZN(n9831) );
  OR2_X1 U12487 ( .A1(n11957), .A2(n11937), .ZN(n9832) );
  AND2_X1 U12488 ( .A1(n10202), .A2(n11308), .ZN(n9833) );
  NAND2_X1 U12489 ( .A1(n13586), .A2(n13585), .ZN(n13584) );
  INV_X1 U12490 ( .A(n10023), .ZN(n14276) );
  NAND2_X1 U12491 ( .A1(n10027), .A2(n10024), .ZN(n10023) );
  NOR2_X1 U12492 ( .A1(n14408), .A2(n10001), .ZN(n9834) );
  INV_X1 U12493 ( .A(n11607), .ZN(n15315) );
  NOR2_X1 U12494 ( .A1(n14398), .A2(n15316), .ZN(n11607) );
  INV_X1 U12495 ( .A(n10030), .ZN(n10029) );
  NAND2_X1 U12496 ( .A1(n12537), .A2(n14615), .ZN(n10030) );
  INV_X1 U12497 ( .A(n10100), .ZN(n10099) );
  OR2_X1 U12498 ( .A1(n14433), .A2(n10101), .ZN(n10100) );
  OR2_X1 U12499 ( .A1(n17693), .A2(n17708), .ZN(n9835) );
  OR2_X1 U12500 ( .A1(n19025), .A2(n19036), .ZN(n9836) );
  AND2_X1 U12501 ( .A1(n14042), .A2(n12089), .ZN(n12080) );
  AND2_X1 U12502 ( .A1(n10098), .A2(n14399), .ZN(n9837) );
  NOR2_X1 U12503 ( .A1(n16306), .A2(n16307), .ZN(n9838) );
  AND2_X1 U12504 ( .A1(n10013), .A2(n10012), .ZN(n9839) );
  AND2_X1 U12505 ( .A1(n12595), .A2(n10028), .ZN(n9840) );
  OR2_X1 U12506 ( .A1(n12074), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9841) );
  AND2_X1 U12507 ( .A1(n9824), .A2(n14697), .ZN(n9842) );
  AND2_X1 U12508 ( .A1(n9825), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9843) );
  OR2_X1 U12509 ( .A1(n9787), .A2(n10002), .ZN(n9844) );
  AND2_X1 U12510 ( .A1(n11130), .A2(n11162), .ZN(n9845) );
  INV_X1 U12511 ( .A(n13802), .ZN(n20257) );
  XOR2_X1 U12512 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n12956), .Z(
        n16696) );
  INV_X1 U12513 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9930) );
  INV_X1 U12514 ( .A(n12643), .ZN(n12636) );
  NOR2_X1 U12515 ( .A1(n13944), .A2(n13943), .ZN(n9846) );
  NOR2_X1 U12516 ( .A1(n20815), .A2(n14046), .ZN(n9847) );
  NOR2_X1 U12517 ( .A1(n15828), .A2(n15827), .ZN(n9848) );
  NAND2_X1 U12518 ( .A1(n10104), .A2(n10103), .ZN(n13211) );
  NAND2_X1 U12519 ( .A1(n10145), .A2(n9791), .ZN(n13623) );
  NOR2_X1 U12520 ( .A1(n16408), .A2(n16409), .ZN(n15774) );
  INV_X1 U12521 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11656) );
  NOR2_X1 U12522 ( .A1(n15813), .A2(n10004), .ZN(n15793) );
  AND2_X1 U12523 ( .A1(n13944), .A2(n10086), .ZN(n14024) );
  NOR2_X1 U12524 ( .A1(n15813), .A2(n15812), .ZN(n15811) );
  AND2_X1 U12525 ( .A1(n13146), .A2(n13138), .ZN(n13148) );
  NOR2_X1 U12526 ( .A1(n14507), .A2(n10092), .ZN(n13779) );
  AND2_X1 U12527 ( .A1(n11049), .A2(n10008), .ZN(n9849) );
  NOR2_X1 U12528 ( .A1(n14008), .A2(n14007), .ZN(n14006) );
  AND2_X1 U12529 ( .A1(n13146), .A2(n9823), .ZN(n13144) );
  AND2_X1 U12530 ( .A1(n11394), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n9850) );
  AND2_X1 U12531 ( .A1(n9849), .A2(n15698), .ZN(n9851) );
  INV_X1 U12532 ( .A(n13411), .ZN(n12981) );
  NAND2_X1 U12533 ( .A1(n11394), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n9852) );
  INV_X1 U12534 ( .A(n15576), .ZN(n9992) );
  XNOR2_X1 U12535 ( .A(n11819), .B(n9919), .ZN(n20392) );
  AND2_X1 U12536 ( .A1(n10173), .A2(n10171), .ZN(n17891) );
  OR2_X1 U12537 ( .A1(n17484), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n9853) );
  INV_X1 U12538 ( .A(n9969), .ZN(n15075) );
  NOR2_X1 U12539 ( .A1(n14279), .A2(n9970), .ZN(n9969) );
  INV_X1 U12540 ( .A(n10160), .ZN(n10159) );
  NOR2_X1 U12541 ( .A1(n10793), .A2(n10162), .ZN(n10160) );
  AND2_X1 U12542 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9854) );
  INV_X1 U12543 ( .A(n9896), .ZN(n13743) );
  AND2_X1 U12544 ( .A1(n10867), .A2(n9794), .ZN(n9855) );
  AND2_X1 U12545 ( .A1(n9929), .A2(n13113), .ZN(n9856) );
  OR2_X1 U12546 ( .A1(n14507), .A2(n10093), .ZN(n10097) );
  NOR2_X1 U12547 ( .A1(n19000), .A2(n19001), .ZN(n9857) );
  AND2_X1 U12548 ( .A1(n12340), .A2(n10025), .ZN(n9858) );
  INV_X1 U12549 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10046) );
  INV_X1 U12550 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n9923) );
  AND2_X1 U12551 ( .A1(n17687), .A2(n9790), .ZN(n9859) );
  AND2_X1 U12552 ( .A1(n13146), .A2(n9825), .ZN(n13143) );
  OR2_X1 U12553 ( .A1(n17609), .A2(n10048), .ZN(n9860) );
  XNOR2_X1 U12555 ( .A(n13140), .B(n21126), .ZN(n14451) );
  AND2_X1 U12556 ( .A1(n9999), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9861) );
  NAND2_X1 U12557 ( .A1(n14522), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9862) );
  INV_X1 U12558 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10047) );
  CLKBUF_X1 U12559 ( .A(n18202), .Z(n9863) );
  NOR3_X1 U12560 ( .A1(n17468), .A2(n18750), .A3(n18286), .ZN(n18202) );
  OR2_X1 U12561 ( .A1(n14458), .A2(n19395), .ZN(n10186) );
  OR2_X1 U12562 ( .A1(n14416), .A2(n19395), .ZN(n10000) );
  OAI211_X1 U12563 ( .C1(n15551), .C2(n9780), .A(n9914), .B(n9913), .ZN(
        P2_U2997) );
  AOI22_X2 U12564 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n15176), .B1(DATAI_18_), 
        .B2(n15177), .ZN(n20654) );
  NOR2_X2 U12565 ( .A1(n9784), .A2(n9793), .ZN(n19198) );
  NOR3_X2 U12566 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18819), .A3(
        n18541), .ZN(n18511) );
  NOR3_X2 U12567 ( .A1(n18819), .A2(n18793), .A3(n18446), .ZN(n18420) );
  NOR2_X2 U12568 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18935), .ZN(n18819) );
  INV_X2 U12569 ( .A(n16866), .ZN(n18285) );
  OR2_X2 U12570 ( .A1(n12652), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20207) );
  NAND2_X1 U12571 ( .A1(n9912), .A2(n10423), .ZN(n10428) );
  XNOR2_X2 U12572 ( .A(n10384), .B(n10385), .ZN(n10404) );
  AND3_X2 U12573 ( .A1(n9998), .A2(n14003), .A3(n11508), .ZN(n11515) );
  NAND2_X2 U12574 ( .A1(n14002), .A2(n20857), .ZN(n14003) );
  NOR2_X2 U12575 ( .A1(n15555), .A2(n9862), .ZN(n15525) );
  NAND2_X1 U12576 ( .A1(n9867), .A2(n9901), .ZN(n9900) );
  OAI21_X2 U12577 ( .B1(n9867), .B2(n13865), .A(n11504), .ZN(n11505) );
  OAI21_X1 U12578 ( .B1(n9867), .B2(n11396), .A(n13580), .ZN(n9906) );
  XNOR2_X1 U12579 ( .A(n9867), .B(n9866), .ZN(n13880) );
  INV_X1 U12580 ( .A(n13865), .ZN(n9866) );
  XNOR2_X2 U12581 ( .A(n10052), .B(n10053), .ZN(n9867) );
  NAND2_X2 U12582 ( .A1(n18933), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n18778) );
  NAND2_X1 U12583 ( .A1(n12902), .A2(n18323), .ZN(n12894) );
  NOR2_X2 U12584 ( .A1(n17500), .A2(n18348), .ZN(n12902) );
  AND2_X2 U12585 ( .A1(n9805), .A2(n9874), .ZN(n18348) );
  NAND3_X1 U12586 ( .A1(n12846), .A2(n12847), .A3(n12845), .ZN(n9875) );
  AND2_X2 U12587 ( .A1(n16682), .A2(n9955), .ZN(n18767) );
  OR2_X2 U12588 ( .A1(n15915), .A2(n17540), .ZN(n16668) );
  NOR2_X2 U12589 ( .A1(n18196), .A2(n18959), .ZN(n18744) );
  AND2_X4 U12590 ( .A1(n13834), .A2(n10237), .ZN(n10801) );
  NAND3_X1 U12591 ( .A1(n9883), .A2(n9884), .A3(n10942), .ZN(n9878) );
  NAND2_X1 U12592 ( .A1(n10469), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n9884) );
  NOR2_X2 U12593 ( .A1(n11223), .A2(n11220), .ZN(n11238) );
  INV_X1 U12594 ( .A(n11374), .ZN(n9892) );
  NOR2_X2 U12596 ( .A1(n11341), .A2(n11314), .ZN(n11329) );
  NAND4_X1 U12597 ( .A1(n10335), .A2(n11445), .A3(n10334), .A4(n10333), .ZN(
        n9896) );
  NAND4_X1 U12598 ( .A1(n10335), .A2(n11445), .A3(n10334), .A4(n9818), .ZN(
        n15840) );
  NAND4_X1 U12599 ( .A1(n9911), .A2(n10323), .A3(n10325), .A4(n10324), .ZN(
        n9907) );
  AND2_X1 U12600 ( .A1(n10326), .A2(n10456), .ZN(n9911) );
  XNOR2_X1 U12601 ( .A(n9912), .B(n10398), .ZN(n11083) );
  AOI21_X2 U12602 ( .B1(n16343), .B2(n16341), .A(n14386), .ZN(n15568) );
  NAND2_X1 U12603 ( .A1(n12993), .A2(n9917), .ZN(n9915) );
  OR2_X2 U12604 ( .A1(n20392), .A2(n11845), .ZN(n11846) );
  NAND3_X1 U12605 ( .A1(n9920), .A2(n10106), .A3(n9921), .ZN(n13708) );
  NAND2_X1 U12606 ( .A1(n13647), .A2(n10105), .ZN(n9920) );
  NAND2_X1 U12607 ( .A1(n13646), .A2(n9922), .ZN(n9921) );
  OAI21_X2 U12608 ( .B1(n14832), .B2(n14851), .A(n14843), .ZN(n14833) );
  OR2_X2 U12609 ( .A1(n14833), .A2(n9841), .ZN(n14807) );
  NAND3_X1 U12610 ( .A1(n14292), .A2(n12053), .A3(n9940), .ZN(n9928) );
  NAND2_X1 U12611 ( .A1(n9929), .A2(n13094), .ZN(n13095) );
  NAND2_X1 U12612 ( .A1(n12140), .A2(n9929), .ZN(n12994) );
  NAND2_X1 U12613 ( .A1(n14934), .A2(n14936), .ZN(n9931) );
  NAND2_X1 U12614 ( .A1(n12054), .A2(n14918), .ZN(n14938) );
  NAND3_X1 U12615 ( .A1(n9933), .A2(n11931), .A3(n9918), .ZN(n9932) );
  NAND2_X1 U12616 ( .A1(n15138), .A2(n14993), .ZN(n9934) );
  INV_X1 U12617 ( .A(n14816), .ZN(n9935) );
  NAND2_X1 U12618 ( .A1(n14816), .A2(n9937), .ZN(n9936) );
  NOR2_X1 U12619 ( .A1(n9939), .A2(n9817), .ZN(n9938) );
  NAND3_X1 U12620 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(P3_EAX_REG_14__SCAN_IN), .ZN(n9945) );
  NAND4_X1 U12621 ( .A1(n12887), .A2(n12886), .A3(n9950), .A4(n9947), .ZN(
        n17349) );
  NAND3_X1 U12622 ( .A1(n12885), .A2(n12889), .A3(n9952), .ZN(n9951) );
  INV_X2 U12623 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21189) );
  AND2_X4 U12624 ( .A1(n13700), .A2(n11662), .ZN(n11725) );
  NOR2_X4 U12625 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11662) );
  NOR2_X4 U12626 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13700) );
  NAND2_X1 U12627 ( .A1(n14688), .A2(n9956), .ZN(P1_U2842) );
  INV_X1 U12628 ( .A(n9968), .ZN(n14234) );
  NOR2_X1 U12629 ( .A1(n14724), .A2(n14713), .ZN(n14715) );
  INV_X1 U12630 ( .A(n14706), .ZN(n9975) );
  INV_X1 U12631 ( .A(n9976), .ZN(n14700) );
  NAND2_X1 U12632 ( .A1(n15618), .A2(n15617), .ZN(n9977) );
  NAND2_X1 U12633 ( .A1(n16371), .A2(n16372), .ZN(n9978) );
  NAND4_X1 U12634 ( .A1(n10301), .A2(n10298), .A3(n10299), .A4(n10300), .ZN(
        n9980) );
  NAND3_X1 U12635 ( .A1(n10295), .A2(n10294), .A3(n10296), .ZN(n9982) );
  NAND2_X1 U12636 ( .A1(n15579), .A2(n9991), .ZN(n9990) );
  OAI21_X2 U12637 ( .B1(n9990), .B2(n9988), .A(n9986), .ZN(n15686) );
  NAND3_X1 U12638 ( .A1(n9994), .A2(n15464), .A3(n9993), .ZN(n15451) );
  NAND2_X1 U12639 ( .A1(n11389), .A2(n9995), .ZN(n9993) );
  NAND2_X1 U12640 ( .A1(n14478), .A2(n11389), .ZN(n9994) );
  INV_X1 U12641 ( .A(n16374), .ZN(n9998) );
  NOR2_X1 U12642 ( .A1(n15828), .A2(n9788), .ZN(n15813) );
  NAND2_X1 U12643 ( .A1(n13891), .A2(n10009), .ZN(n16443) );
  NAND2_X1 U12644 ( .A1(n9747), .A2(n19879), .ZN(n13592) );
  NAND2_X2 U12645 ( .A1(n11777), .A2(n10015), .ZN(n15153) );
  NAND2_X1 U12646 ( .A1(n11786), .A2(n10015), .ZN(n11791) );
  OAI211_X1 U12647 ( .C1(n14965), .C2(n20139), .A(n10018), .B(n10017), .ZN(
        P1_U2968) );
  NAND2_X1 U12648 ( .A1(n14545), .A2(n20293), .ZN(n10018) );
  XNOR2_X2 U12649 ( .A(n10019), .B(n12647), .ZN(n14545) );
  NAND2_X1 U12650 ( .A1(n14418), .A2(n14568), .ZN(n10019) );
  NAND2_X1 U12651 ( .A1(n14672), .A2(n9842), .ZN(n14644) );
  AND4_X4 U12652 ( .A1(n11656), .A2(n11802), .A3(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12621) );
  NAND2_X1 U12653 ( .A1(n10027), .A2(n9858), .ZN(n14332) );
  NAND2_X1 U12654 ( .A1(n14627), .A2(n9840), .ZN(n14417) );
  NAND2_X1 U12655 ( .A1(n14627), .A2(n10029), .ZN(n14602) );
  NAND2_X1 U12656 ( .A1(n10032), .A2(n10033), .ZN(n16807) );
  INV_X1 U12657 ( .A(n10035), .ZN(n16813) );
  AND2_X1 U12658 ( .A1(n9783), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10044) );
  NAND3_X1 U12659 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10048) );
  NAND2_X1 U12660 ( .A1(n11163), .A2(n11162), .ZN(n10052) );
  NAND2_X1 U12661 ( .A1(n11131), .A2(n11130), .ZN(n10053) );
  AND3_X1 U12662 ( .A1(n11131), .A2(n11163), .A3(n9845), .ZN(n11491) );
  XNOR2_X1 U12663 ( .A(n11491), .B(n11164), .ZN(n11506) );
  NAND2_X1 U12665 ( .A1(n10056), .A2(n10057), .ZN(n13239) );
  NAND2_X1 U12666 ( .A1(n10060), .A2(n10061), .ZN(n16298) );
  INV_X1 U12669 ( .A(n13171), .ZN(n10063) );
  NAND2_X1 U12670 ( .A1(n10064), .A2(n10063), .ZN(n13167) );
  NOR2_X1 U12671 ( .A1(n19123), .A2(n10068), .ZN(n10067) );
  NAND2_X1 U12672 ( .A1(n10069), .A2(n11533), .ZN(n10102) );
  XNOR2_X2 U12673 ( .A(n10069), .B(n11533), .ZN(n11101) );
  NAND2_X2 U12674 ( .A1(n10428), .A2(n10427), .ZN(n10069) );
  INV_X1 U12675 ( .A(n10072), .ZN(n19034) );
  NAND2_X1 U12676 ( .A1(n13146), .A2(n9843), .ZN(n13140) );
  INV_X1 U12677 ( .A(n10097), .ZN(n13763) );
  NAND2_X1 U12678 ( .A1(n14462), .A2(n9837), .ZN(n14398) );
  INV_X1 U12679 ( .A(n11804), .ZN(n10104) );
  NAND2_X1 U12680 ( .A1(n11910), .A2(n11955), .ZN(n13731) );
  NAND2_X1 U12681 ( .A1(n13647), .A2(n11928), .ZN(n11929) );
  INV_X1 U12682 ( .A(n11928), .ZN(n10107) );
  NAND3_X1 U12683 ( .A1(n11910), .A2(n11955), .A3(n12080), .ZN(n10108) );
  AND2_X2 U12684 ( .A1(n14807), .A2(n10109), .ZN(n14809) );
  NAND2_X1 U12685 ( .A1(n14833), .A2(n9792), .ZN(n10109) );
  INV_X1 U12686 ( .A(n12071), .ZN(n10118) );
  INV_X1 U12687 ( .A(n10124), .ZN(n14831) );
  NAND2_X1 U12688 ( .A1(n10388), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10383) );
  NAND2_X1 U12689 ( .A1(n10369), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10133) );
  NAND2_X1 U12690 ( .A1(n10138), .A2(n9795), .ZN(n10141) );
  OR2_X2 U12691 ( .A1(n10756), .A2(n10755), .ZN(n10138) );
  OAI22_X2 U12692 ( .A1(n10141), .A2(n15253), .B1(n10142), .B2(n10788), .ZN(
        n15248) );
  AND2_X2 U12693 ( .A1(n10145), .A2(n10144), .ZN(n13767) );
  AND3_X2 U12694 ( .A1(n10150), .A2(n10146), .A3(n10149), .ZN(n15292) );
  NAND3_X1 U12695 ( .A1(n10150), .A2(n10152), .A3(n10149), .ZN(n15294) );
  NAND2_X1 U12696 ( .A1(n15249), .A2(n10161), .ZN(n10155) );
  OAI211_X1 U12697 ( .C1(n15249), .C2(n10162), .A(n10155), .B(n10159), .ZN(
        n12655) );
  OAI211_X1 U12698 ( .C1(n15249), .C2(n10157), .A(n10156), .B(n11082), .ZN(
        P2_U2889) );
  NAND2_X1 U12699 ( .A1(n15249), .A2(n9855), .ZN(n10156) );
  NAND2_X1 U12700 ( .A1(n10159), .A2(n10162), .ZN(n10158) );
  NAND2_X1 U12701 ( .A1(n17906), .A2(n10170), .ZN(n10168) );
  INV_X1 U12702 ( .A(n17791), .ZN(n10179) );
  INV_X2 U12703 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18933) );
  NAND4_X1 U12704 ( .A1(n9998), .A2(n14003), .A3(n11508), .A4(n11517), .ZN(
        n11511) );
  INV_X1 U12705 ( .A(n15693), .ZN(n11531) );
  OAI21_X2 U12706 ( .B1(n15602), .B2(n10185), .A(n10183), .ZN(n15693) );
  NAND3_X1 U12707 ( .A1(n9819), .A2(n10187), .A3(n10186), .ZN(P2_U3015) );
  OR2_X1 U12708 ( .A1(n15493), .A2(n10189), .ZN(n15467) );
  NOR2_X1 U12709 ( .A1(n15493), .A2(n10188), .ZN(n15457) );
  NOR2_X1 U12710 ( .A1(n15493), .A2(n10190), .ZN(n15473) );
  NOR2_X1 U12711 ( .A1(n14466), .A2(n14389), .ZN(n14447) );
  AND2_X4 U12712 ( .A1(n11664), .A2(n13424), .ZN(n11756) );
  NOR2_X4 U12713 ( .A1(n18778), .A2(n12666), .ZN(n15900) );
  CLKBUF_X1 U12714 ( .A(n13704), .Z(n20518) );
  NAND2_X1 U12715 ( .A1(n15268), .A2(n15267), .ZN(n15266) );
  INV_X1 U12716 ( .A(n11909), .ZN(n11907) );
  AND2_X1 U12717 ( .A1(n9811), .A2(n10680), .ZN(n10662) );
  NAND2_X1 U12718 ( .A1(n11452), .A2(n20109), .ZN(n10343) );
  OR2_X1 U12719 ( .A1(n10391), .A2(n11497), .ZN(n10397) );
  AND2_X1 U12720 ( .A1(n12996), .A2(n11899), .ZN(n12124) );
  AND2_X1 U12721 ( .A1(n14360), .A2(n12996), .ZN(n11777) );
  NAND2_X1 U12722 ( .A1(n11651), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10391) );
  NAND2_X1 U12723 ( .A1(n10336), .A2(n15840), .ZN(n11651) );
  AND2_X4 U12724 ( .A1(n11662), .A2(n13424), .ZN(n11861) );
  OR2_X1 U12725 ( .A1(n10708), .A2(n10709), .ZN(n10710) );
  NAND2_X1 U12726 ( .A1(n11531), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15695) );
  INV_X1 U12727 ( .A(n10388), .ZN(n10430) );
  NAND2_X1 U12728 ( .A1(n10388), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10390) );
  AND2_X1 U12729 ( .A1(n14831), .A2(n15138), .ZN(n14851) );
  OR2_X1 U12730 ( .A1(n10386), .A2(n10385), .ZN(n10387) );
  NAND2_X1 U12731 ( .A1(n10431), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10436) );
  INV_X1 U12732 ( .A(n10431), .ZN(n11647) );
  AND2_X1 U12733 ( .A1(n12621), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11694) );
  AOI22_X1 U12734 ( .A1(n12621), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9767), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11672) );
  INV_X1 U12735 ( .A(n14450), .ZN(n11652) );
  INV_X1 U12736 ( .A(n12700), .ZN(n17019) );
  INV_X1 U12737 ( .A(n12707), .ZN(n13525) );
  AND3_X1 U12738 ( .A1(n15624), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16405), .ZN(n10209) );
  INV_X1 U12739 ( .A(n19275), .ZN(n10867) );
  NOR2_X1 U12740 ( .A1(n15280), .A2(n10682), .ZN(n10708) );
  AND2_X1 U12741 ( .A1(n13134), .A2(n10218), .ZN(n10210) );
  AND4_X1 U12742 ( .A1(n10886), .A2(n10885), .A3(n10884), .A4(n10883), .ZN(
        n10211) );
  NOR2_X1 U12743 ( .A1(n11488), .A2(n10209), .ZN(n10212) );
  AND2_X1 U12744 ( .A1(n11489), .A2(n10212), .ZN(n10213) );
  INV_X1 U12745 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20085) );
  AND3_X1 U12746 ( .A1(n12703), .A2(n12702), .A3(n12701), .ZN(n10214) );
  AND4_X1 U12747 ( .A1(n12712), .A2(n12711), .A3(n12710), .A4(n12709), .ZN(
        n10215) );
  OR2_X1 U12748 ( .A1(n11372), .A2(n15704), .ZN(n10216) );
  AND2_X1 U12749 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10217) );
  OR2_X1 U12750 ( .A1(n14961), .A2(n13133), .ZN(n10218) );
  AND2_X1 U12751 ( .A1(n15059), .A2(n15045), .ZN(n10219) );
  INV_X1 U12752 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12075) );
  AND4_X1 U12753 ( .A1(n14388), .A2(n14444), .A3(n16330), .A4(n16341), .ZN(
        n10220) );
  AND2_X1 U12754 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10221) );
  INV_X1 U12755 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20517) );
  INV_X1 U12756 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12780) );
  AND2_X2 U12757 ( .A1(n13215), .A2(n13564), .ZN(n14762) );
  INV_X1 U12758 ( .A(n15174), .ZN(n13970) );
  NAND2_X1 U12759 ( .A1(n9918), .A2(n13849), .ZN(n15174) );
  AND3_X1 U12760 ( .A1(n16903), .A2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10222) );
  AND2_X1 U12761 ( .A1(n10287), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10224) );
  AND2_X1 U12762 ( .A1(n15452), .A2(n15463), .ZN(n10225) );
  AND2_X1 U12763 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10226) );
  INV_X2 U12764 ( .A(n12661), .ZN(n17296) );
  INV_X1 U12765 ( .A(n12750), .ZN(n12661) );
  INV_X1 U12766 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20069) );
  OR2_X1 U12767 ( .A1(n10977), .A2(n10976), .ZN(n11164) );
  AND2_X1 U12768 ( .A1(n12621), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10228) );
  INV_X1 U12769 ( .A(n17486), .ZN(n17375) );
  AND2_X1 U12770 ( .A1(n16382), .A2(n20078), .ZN(n19382) );
  INV_X1 U12771 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n13298) );
  AND2_X1 U12772 ( .A1(n16373), .A2(n11517), .ZN(n10231) );
  AND3_X1 U12773 ( .A1(n11668), .A2(n11667), .A3(n11666), .ZN(n10232) );
  AND4_X1 U12774 ( .A1(n11711), .A2(n11710), .A3(n11709), .A4(n11708), .ZN(
        n10233) );
  BUF_X1 U12775 ( .A(n11831), .Z(n12525) );
  AND4_X1 U12776 ( .A1(n11699), .A2(n11698), .A3(n11697), .A4(n11696), .ZN(
        n10234) );
  AND2_X1 U12777 ( .A1(n11800), .A2(n12997), .ZN(n10235) );
  AND4_X1 U12778 ( .A1(n11660), .A2(n11659), .A3(n11658), .A4(n11657), .ZN(
        n10236) );
  OR2_X1 U12779 ( .A1(n11991), .A2(n11990), .ZN(n12026) );
  AND2_X1 U12780 ( .A1(n11995), .A2(n11996), .ZN(n11994) );
  OR2_X1 U12781 ( .A1(n11914), .A2(n11904), .ZN(n11905) );
  INV_X1 U12782 ( .A(n12023), .ZN(n12022) );
  OR2_X1 U12783 ( .A1(n11972), .A2(n11971), .ZN(n12002) );
  NAND2_X1 U12784 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11702) );
  AND2_X1 U12785 ( .A1(n12124), .A2(n12972), .ZN(n12125) );
  INV_X1 U12786 ( .A(n11276), .ZN(n11199) );
  NAND2_X1 U12787 ( .A1(n12152), .A2(n11905), .ZN(n11908) );
  AND2_X1 U12788 ( .A1(n12068), .A2(n12067), .ZN(n12069) );
  INV_X1 U12789 ( .A(n10728), .ZN(n10729) );
  AND4_X1 U12790 ( .A1(n10882), .A2(n10881), .A3(n10880), .A4(n10879), .ZN(
        n10887) );
  AND2_X1 U12791 ( .A1(n10282), .A2(n10456), .ZN(n10286) );
  INV_X1 U12792 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12779) );
  NAND2_X1 U12793 ( .A1(n12663), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12701) );
  AND2_X1 U12794 ( .A1(n11752), .A2(n11751), .ZN(n11753) );
  INV_X1 U12795 ( .A(n14591), .ZN(n12595) );
  OR2_X1 U12796 ( .A1(n14704), .A2(n14711), .ZN(n12446) );
  NAND2_X1 U12797 ( .A1(n12981), .A2(n13917), .ZN(n12139) );
  AND2_X1 U12798 ( .A1(n13016), .A2(n13015), .ZN(n13819) );
  NAND2_X1 U12799 ( .A1(n12124), .A2(n12080), .ZN(n12133) );
  INV_X1 U12800 ( .A(n11955), .ZN(n11954) );
  AND2_X1 U12801 ( .A1(n10835), .A2(n10834), .ZN(n10842) );
  NAND2_X1 U12802 ( .A1(n10727), .A2(n10729), .ZN(n10730) );
  INV_X1 U12803 ( .A(n11164), .ZN(n11490) );
  AND2_X1 U12804 ( .A1(n10365), .A2(n10364), .ZN(n10366) );
  AND2_X1 U12805 ( .A1(n10947), .A2(n10946), .ZN(n13269) );
  INV_X1 U12806 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n20935) );
  INV_X1 U12807 ( .A(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n20962) );
  NOR2_X1 U12808 ( .A1(n18773), .A2(n12666), .ZN(n12690) );
  NOR2_X1 U12809 ( .A1(n12394), .A2(n16076), .ZN(n12376) );
  INV_X1 U12810 ( .A(n14628), .ZN(n12537) );
  AND4_X1 U12811 ( .A1(n11772), .A2(n11771), .A3(n11770), .A4(n11769), .ZN(
        n11773) );
  OR2_X1 U12812 ( .A1(n14582), .A2(n12636), .ZN(n12617) );
  INV_X1 U12813 ( .A(n14661), .ZN(n12463) );
  INV_X1 U12814 ( .A(n12638), .ZN(n12645) );
  OR2_X1 U12815 ( .A1(n12043), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14244) );
  INV_X1 U12816 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12111) );
  AND2_X1 U12817 ( .A1(n11332), .A2(n11337), .ZN(n19047) );
  AND3_X1 U12818 ( .A1(n11210), .A2(n11209), .A3(n11208), .ZN(n11220) );
  NAND2_X1 U12819 ( .A1(n10844), .A2(n10843), .ZN(n20098) );
  AND2_X1 U12820 ( .A1(n10681), .A2(n10680), .ZN(n10682) );
  AND2_X1 U12821 ( .A1(n11303), .A2(n15786), .ZN(n15788) );
  INV_X1 U12822 ( .A(n10404), .ZN(n10406) );
  OAI21_X1 U12823 ( .B1(n15864), .B2(n20089), .A(n16494), .ZN(n15875) );
  NAND2_X1 U12824 ( .A1(n12690), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12745) );
  NOR2_X1 U12825 ( .A1(n17744), .A2(n12784), .ZN(n17700) );
  NAND2_X1 U12826 ( .A1(n17540), .A2(n18959), .ZN(n15921) );
  NOR2_X1 U12827 ( .A1(n17475), .A2(n12744), .ZN(n12771) );
  NAND2_X1 U12828 ( .A1(n18755), .A2(n18789), .ZN(n18254) );
  AND2_X1 U12829 ( .A1(n12515), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12516) );
  NOR2_X1 U12830 ( .A1(n12430), .A2(n14893), .ZN(n12411) );
  OR2_X1 U12831 ( .A1(n12375), .A2(n12370), .ZN(n12394) );
  INV_X1 U12832 ( .A(n20193), .ZN(n20210) );
  INV_X1 U12833 ( .A(n20189), .ZN(n16031) );
  NAND2_X1 U12834 ( .A1(n11936), .A2(n11935), .ZN(n13901) );
  NAND2_X1 U12835 ( .A1(n14047), .A2(n15993), .ZN(n20203) );
  AND2_X1 U12836 ( .A1(n13008), .A2(n13007), .ZN(n13650) );
  OR2_X1 U12837 ( .A1(n13228), .A2(n13927), .ZN(n14793) );
  XNOR2_X1 U12838 ( .A(n12649), .B(n14559), .ZN(n14037) );
  INV_X1 U12839 ( .A(n14588), .ZN(n14603) );
  OR2_X1 U12840 ( .A1(n16026), .A2(n12636), .ZN(n12495) );
  NOR2_X1 U12841 ( .A1(n12245), .A2(n12244), .ZN(n12262) );
  NAND2_X1 U12842 ( .A1(n12232), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12245) );
  INV_X1 U12843 ( .A(n20287), .ZN(n14950) );
  AND2_X1 U12844 ( .A1(n14935), .A2(n14932), .ZN(n14917) );
  AND2_X1 U12845 ( .A1(n15050), .A2(n16175), .ZN(n15124) );
  OR2_X1 U12846 ( .A1(n15050), .A2(n13642), .ZN(n13108) );
  NAND2_X1 U12847 ( .A1(n13416), .A2(n12141), .ZN(n12997) );
  INV_X1 U12848 ( .A(n20803), .ZN(n14500) );
  AND2_X1 U12849 ( .A1(n20727), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16001) );
  OR2_X1 U12850 ( .A1(n13731), .A2(n11953), .ZN(n14161) );
  AND2_X1 U12851 ( .A1(n20432), .A2(n13970), .ZN(n20525) );
  INV_X1 U12852 ( .A(n15167), .ZN(n15165) );
  INV_X1 U12853 ( .A(n15171), .ZN(n20438) );
  INV_X1 U12854 ( .A(n14360), .ZN(n13854) );
  NOR2_X1 U12855 ( .A1(n15244), .A2(n15243), .ZN(n15245) );
  AND2_X1 U12856 ( .A1(n10724), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13884) );
  INV_X1 U12857 ( .A(n10709), .ZN(n10705) );
  OR2_X1 U12858 ( .A1(n14099), .A2(n15297), .ZN(n15339) );
  AND2_X1 U12859 ( .A1(n11388), .A2(n14477), .ZN(n11389) );
  OR2_X1 U12860 ( .A1(n15677), .A2(n11484), .ZN(n15637) );
  OR2_X1 U12861 ( .A1(n15688), .A2(n15692), .ZN(n15677) );
  OR2_X1 U12862 ( .A1(n11371), .A2(n15717), .ZN(n15510) );
  OR2_X1 U12863 ( .A1(n19041), .A2(n11356), .ZN(n14444) );
  AND2_X1 U12864 ( .A1(n14428), .A2(n16329), .ZN(n14429) );
  INV_X1 U12865 ( .A(n15581), .ZN(n16353) );
  OR2_X1 U12866 ( .A1(n16373), .A2(n11513), .ZN(n11514) );
  INV_X1 U12867 ( .A(n16477), .ZN(n11443) );
  OR2_X1 U12868 ( .A1(n20072), .A2(n19407), .ZN(n15894) );
  OR2_X1 U12869 ( .A1(n20072), .A2(n20079), .ZN(n19840) );
  NOR2_X1 U12870 ( .A1(n18766), .A2(n18318), .ZN(n15915) );
  NAND2_X1 U12871 ( .A1(n18973), .A2(n17500), .ZN(n16686) );
  NOR2_X1 U12872 ( .A1(n18106), .A2(n18118), .ZN(n18105) );
  INV_X1 U12873 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17841) );
  NAND2_X1 U12874 ( .A1(n17797), .A2(n17961), .ZN(n17749) );
  NOR2_X1 U12875 ( .A1(n17872), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12789) );
  NOR2_X1 U12876 ( .A1(n12950), .A2(n17868), .ZN(n18159) );
  NOR2_X1 U12877 ( .A1(n12911), .A2(n12912), .ZN(n18762) );
  NOR2_X1 U12878 ( .A1(n18219), .A2(n17897), .ZN(n17896) );
  INV_X1 U12879 ( .A(n18612), .ZN(n18518) );
  NOR2_X1 U12880 ( .A1(n12844), .A2(n12843), .ZN(n18323) );
  OR2_X1 U12881 ( .A1(n13391), .A2(n20133), .ZN(n14565) );
  NAND2_X1 U12882 ( .A1(n12516), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12555) );
  NOR2_X1 U12883 ( .A1(n14548), .A2(n20196), .ZN(n20158) );
  INV_X1 U12884 ( .A(n13229), .ZN(n13230) );
  INV_X1 U12885 ( .A(n14627), .ZN(n14647) );
  INV_X1 U12886 ( .A(n14762), .ZN(n14789) );
  NAND2_X1 U12887 ( .A1(n12263), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12301) );
  OR2_X1 U12888 ( .A1(n14109), .A2(n14108), .ZN(n14230) );
  NAND2_X1 U12889 ( .A1(n12177), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12185) );
  OR2_X1 U12890 ( .A1(n13429), .A2(n20133), .ZN(n13546) );
  AND2_X1 U12891 ( .A1(n15025), .A2(n13114), .ZN(n14990) );
  OR2_X1 U12892 ( .A1(n15029), .A2(n13127), .ZN(n15015) );
  AND2_X1 U12893 ( .A1(n15046), .A2(n15020), .ZN(n15025) );
  AND2_X1 U12894 ( .A1(n15093), .A2(n13119), .ZN(n15067) );
  NOR2_X1 U12895 ( .A1(n16204), .A2(n13118), .ZN(n15093) );
  NOR2_X1 U12896 ( .A1(n15123), .A2(n15051), .ZN(n16204) );
  INV_X1 U12897 ( .A(n15137), .ZN(n20318) );
  NOR2_X1 U12898 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20804) );
  INV_X1 U12899 ( .A(n20385), .ZN(n20368) );
  AND2_X1 U12900 ( .A1(n20820), .A2(n13731), .ZN(n20391) );
  AND2_X1 U12901 ( .A1(n20391), .A2(n20493), .ZN(n20452) );
  NOR2_X1 U12902 ( .A1(n14161), .A2(n13904), .ZN(n20457) );
  NOR2_X1 U12903 ( .A1(n14161), .A2(n13905), .ZN(n20481) );
  INV_X1 U12904 ( .A(n14161), .ZN(n20817) );
  NOR2_X1 U12905 ( .A1(n15166), .A2(n15165), .ZN(n20516) );
  AND2_X1 U12906 ( .A1(n20812), .A2(n13948), .ZN(n20588) );
  INV_X1 U12907 ( .A(n20627), .ZN(n20618) );
  AND2_X1 U12908 ( .A1(n15166), .A2(n15165), .ZN(n20493) );
  AND2_X1 U12909 ( .A1(n20811), .A2(n15167), .ZN(n20639) );
  AND2_X1 U12910 ( .A1(n20811), .A2(n15165), .ZN(n20658) );
  OAI211_X1 U12911 ( .C1(n13972), .C2(n20655), .A(n13971), .B(n20438), .ZN(
        n20659) );
  AND2_X1 U12912 ( .A1(n19362), .A2(n16501), .ZN(n19203) );
  AND2_X1 U12913 ( .A1(n19357), .A2(n20107), .ZN(n19187) );
  AOI21_X1 U12914 ( .B1(n15351), .B2(n15350), .A(n15349), .ZN(n16255) );
  AND2_X1 U12915 ( .A1(n15338), .A2(n15334), .ZN(n15332) );
  INV_X1 U12916 ( .A(n19270), .ZN(n19262) );
  NOR2_X1 U12918 ( .A1(n15303), .A2(n15302), .ZN(n15962) );
  INV_X2 U12919 ( .A(n10331), .ZN(n19422) );
  INV_X1 U12920 ( .A(n19385), .ZN(n16378) );
  AND2_X1 U12921 ( .A1(n16382), .A2(n19375), .ZN(n16370) );
  AOI21_X1 U12922 ( .B1(n15520), .B2(n14516), .A(n14515), .ZN(n14521) );
  INV_X1 U12923 ( .A(n19406), .ZN(n16450) );
  AND2_X1 U12924 ( .A1(n20064), .A2(n11441), .ZN(n19365) );
  INV_X1 U12925 ( .A(n19402), .ZN(n16411) );
  NOR2_X1 U12926 ( .A1(n13749), .A2(n19879), .ZN(n15835) );
  AND2_X1 U12927 ( .A1(n15893), .A2(n19274), .ZN(n19580) );
  AND2_X1 U12928 ( .A1(n19580), .A2(n20060), .ZN(n19576) );
  AND2_X1 U12929 ( .A1(n19580), .A2(n19834), .ZN(n19637) );
  INV_X1 U12930 ( .A(n19645), .ZN(n19658) );
  AND2_X1 U12931 ( .A1(n19580), .A2(n15885), .ZN(n19683) );
  INV_X1 U12932 ( .A(n19718), .ZN(n19719) );
  INV_X1 U12933 ( .A(n19788), .ZN(n19780) );
  INV_X1 U12934 ( .A(n19794), .ZN(n19824) );
  INV_X1 U12935 ( .A(n19840), .ZN(n19834) );
  INV_X1 U12936 ( .A(n19796), .ZN(n19883) );
  INV_X1 U12937 ( .A(n19889), .ZN(n19833) );
  INV_X1 U12938 ( .A(n19862), .ZN(n19950) );
  INV_X1 U12939 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18926) );
  NAND2_X1 U12940 ( .A1(n16710), .A2(n16709), .ZN(n16711) );
  INV_X1 U12941 ( .A(n16686), .ZN(n16702) );
  INV_X1 U12942 ( .A(n17064), .ZN(n17035) );
  INV_X1 U12943 ( .A(n17065), .ZN(n17048) );
  NOR3_X1 U12944 ( .A1(n17431), .A2(n17544), .A3(n17426), .ZN(n17415) );
  INV_X1 U12945 ( .A(n17769), .ZN(n17755) );
  NAND2_X1 U12946 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18102), .ZN(
        n18028) );
  NOR2_X2 U12947 ( .A1(n17468), .A2(n17965), .ZN(n17873) );
  NAND2_X1 U12948 ( .A1(n17749), .A2(n17823), .ZN(n17955) );
  NOR2_X1 U12949 ( .A1(n12954), .A2(n18028), .ZN(n17967) );
  INV_X1 U12950 ( .A(n17872), .ZN(n17802) );
  NAND2_X1 U12951 ( .A1(n18163), .A2(n18095), .ZN(n18106) );
  OAI21_X2 U12952 ( .B1(n18764), .B2(n18774), .A(n18762), .ZN(n18787) );
  INV_X1 U12953 ( .A(n18750), .ZN(n16553) );
  INV_X1 U12954 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18971) );
  INV_X1 U12955 ( .A(n15880), .ZN(n15878) );
  OR2_X1 U12956 ( .A1(n13546), .A2(n13390), .ZN(n14567) );
  INV_X1 U12957 ( .A(n20205), .ZN(n20191) );
  INV_X1 U12958 ( .A(n20185), .ZN(n16117) );
  INV_X1 U12959 ( .A(n20223), .ZN(n14730) );
  INV_X1 U12960 ( .A(n16135), .ZN(n14339) );
  OR2_X1 U12961 ( .A1(n14789), .A2(n13924), .ZN(n14337) );
  OR3_X1 U12962 ( .A1(n13546), .A2(n13545), .A3(n16017), .ZN(n20250) );
  NOR2_X1 U12963 ( .A1(n14567), .A2(n13605), .ZN(n13802) );
  OAI21_X1 U12964 ( .B1(n14320), .B2(n14277), .A(n10023), .ZN(n14944) );
  OR2_X1 U12965 ( .A1(n20287), .A2(n13617), .ZN(n20298) );
  NAND2_X1 U12966 ( .A1(n13120), .A2(n12995), .ZN(n15137) );
  NAND2_X1 U12967 ( .A1(n20391), .A2(n20516), .ZN(n20372) );
  NAND2_X1 U12968 ( .A1(n20391), .A2(n14162), .ZN(n20425) );
  INV_X1 U12969 ( .A(n20452), .ZN(n20461) );
  INV_X1 U12970 ( .A(n20457), .ZN(n20473) );
  NAND2_X1 U12971 ( .A1(n20817), .A2(n14162), .ZN(n20508) );
  NAND2_X1 U12972 ( .A1(n20812), .A2(n20516), .ZN(n20573) );
  NAND2_X1 U12973 ( .A1(n20812), .A2(n14162), .ZN(n20627) );
  NAND2_X1 U12974 ( .A1(n13966), .A2(n14162), .ZN(n20725) );
  INV_X1 U12975 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20526) );
  AOI21_X1 U12976 ( .B1(n19203), .B2(n15627), .A(n13203), .ZN(n13204) );
  INV_X1 U12977 ( .A(n19203), .ZN(n19182) );
  INV_X1 U12978 ( .A(n12658), .ZN(n12659) );
  INV_X1 U12979 ( .A(n9778), .ZN(n15319) );
  AND2_X1 U12980 ( .A1(n19272), .A2(n19275), .ZN(n19238) );
  INV_X1 U12981 ( .A(n19280), .ZN(n19269) );
  INV_X1 U12982 ( .A(n19293), .ZN(n19319) );
  NAND2_X1 U12983 ( .A1(n19286), .A2(n19980), .ZN(n19352) );
  INV_X1 U12984 ( .A(n19362), .ZN(n19283) );
  NAND2_X1 U12985 ( .A1(n13380), .A2(n13377), .ZN(n16382) );
  INV_X1 U12986 ( .A(n16451), .ZN(n19395) );
  INV_X1 U12987 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20092) );
  NAND2_X1 U12988 ( .A1(n19695), .A2(n19549), .ZN(n19485) );
  NAND2_X1 U12989 ( .A1(n19549), .A2(n20060), .ZN(n19540) );
  INV_X1 U12990 ( .A(n19576), .ZN(n19554) );
  NAND2_X1 U12991 ( .A1(n19549), .A2(n19834), .ZN(n19610) );
  INV_X1 U12992 ( .A(n19637), .ZN(n19634) );
  INV_X1 U12993 ( .A(n19659), .ZN(n19656) );
  INV_X1 U12994 ( .A(n19683), .ZN(n19691) );
  OR2_X1 U12995 ( .A1(n19725), .A2(n19692), .ZN(n19718) );
  OR2_X1 U12996 ( .A1(n19841), .A2(n19692), .ZN(n19724) );
  NAND2_X1 U12997 ( .A1(n19789), .A2(n20060), .ZN(n19788) );
  INV_X1 U12998 ( .A(n19924), .ZN(n19809) );
  INV_X1 U12999 ( .A(n19959), .ZN(n19828) );
  NAND2_X1 U13000 ( .A1(n19789), .A2(n19834), .ZN(n19867) );
  AOI21_X1 U13001 ( .B1(n19878), .B2(n19884), .A(n19875), .ZN(n19914) );
  AOI21_X1 U13002 ( .B1(n15890), .B2(n19873), .A(n15889), .ZN(n19964) );
  AND2_X1 U13003 ( .A1(n17346), .A2(n17431), .ZN(n17343) );
  INV_X1 U13004 ( .A(n14375), .ZN(n17346) );
  INV_X1 U13005 ( .A(n16552), .ZN(n17468) );
  NOR2_X1 U13006 ( .A1(n12733), .A2(n12732), .ZN(n17479) );
  NOR2_X1 U13007 ( .A1(n18954), .A2(n17501), .ZN(n17514) );
  NAND2_X1 U13008 ( .A1(n17539), .A2(n17499), .ZN(n17537) );
  NAND2_X1 U13009 ( .A1(n17834), .A2(n16508), .ZN(n17769) );
  INV_X1 U13010 ( .A(n17873), .ZN(n17837) );
  INV_X1 U13011 ( .A(n17801), .ZN(n17876) );
  INV_X1 U13012 ( .A(n17955), .ZN(n17946) );
  INV_X1 U13013 ( .A(n9863), .ZN(n18175) );
  INV_X1 U13014 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18793) );
  INV_X2 U13015 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18940) );
  INV_X1 U13016 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n20932) );
  OAI21_X1 U13017 ( .B1(n14424), .B2(n15137), .A(n10210), .ZN(P1_U3002) );
  NOR2_X4 U13018 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13833) );
  AND2_X4 U13019 ( .A1(n13834), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10636) );
  AOI22_X1 U13020 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10241) );
  AND2_X2 U13021 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11403) );
  AOI22_X1 U13022 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10457), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10240) );
  AND2_X4 U13023 ( .A1(n13833), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10773) );
  AOI22_X1 U13024 ( .A1(n9764), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10804), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10239) );
  AND3_X4 U13025 ( .A1(n13837), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10806) );
  AND3_X4 U13026 ( .A1(n13745), .A2(n10237), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10805) );
  AOI22_X1 U13027 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10238) );
  AOI22_X1 U13028 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10246) );
  AOI22_X1 U13029 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9765), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10245) );
  AOI22_X1 U13030 ( .A1(n9764), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9771), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10244) );
  AOI22_X1 U13031 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10243) );
  AOI22_X1 U13032 ( .A1(n9750), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n9766), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10251) );
  AOI22_X1 U13033 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10801), .B1(
        n9765), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10250) );
  AOI22_X1 U13034 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10804), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10249) );
  AOI22_X1 U13035 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10248) );
  NAND4_X1 U13036 ( .A1(n10251), .A2(n10250), .A3(n10249), .A4(n10248), .ZN(
        n10252) );
  NAND2_X1 U13037 ( .A1(n10252), .A2(n10456), .ZN(n10259) );
  AOI22_X1 U13038 ( .A1(n9751), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10256) );
  AOI22_X1 U13039 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9770), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U13040 ( .A1(n9764), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9771), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10254) );
  AOI22_X1 U13041 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10253) );
  NAND4_X1 U13042 ( .A1(n10256), .A2(n10255), .A3(n10254), .A4(n10253), .ZN(
        n10257) );
  NAND2_X1 U13043 ( .A1(n10257), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10258) );
  AOI22_X1 U13044 ( .A1(n9751), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n9766), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10263) );
  AOI22_X1 U13045 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9765), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10262) );
  AOI22_X1 U13046 ( .A1(n9764), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10804), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10261) );
  AOI22_X1 U13047 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10260) );
  NAND4_X1 U13048 ( .A1(n10263), .A2(n10262), .A3(n10261), .A4(n10260), .ZN(
        n10269) );
  AOI22_X1 U13049 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10267) );
  AOI22_X1 U13050 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10457), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10266) );
  AOI22_X1 U13051 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9771), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10265) );
  AOI22_X1 U13052 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10264) );
  NAND4_X1 U13053 ( .A1(n10267), .A2(n10266), .A3(n10265), .A4(n10264), .ZN(
        n10268) );
  MUX2_X2 U13054 ( .A(n10269), .B(n10268), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10447) );
  NOR2_X1 U13055 ( .A1(n10327), .A2(n10447), .ZN(n10302) );
  AOI22_X1 U13056 ( .A1(n9750), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10273) );
  AOI22_X1 U13057 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9765), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10272) );
  AOI22_X1 U13058 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10804), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10271) );
  AOI22_X1 U13059 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10270) );
  AOI22_X1 U13060 ( .A1(n9750), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10278) );
  AOI22_X1 U13061 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10804), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10277) );
  AOI22_X1 U13062 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10276) );
  AOI22_X1 U13063 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10457), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10275) );
  NAND2_X2 U13064 ( .A1(n10281), .A2(n10280), .ZN(n19435) );
  AOI22_X1 U13065 ( .A1(n9751), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(n9766), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10282) );
  AOI22_X1 U13066 ( .A1(n9764), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n9771), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10285) );
  AOI22_X1 U13067 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U13068 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9765), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10283) );
  NAND4_X1 U13069 ( .A1(n10286), .A2(n10285), .A3(n10284), .A4(n10283), .ZN(
        n10292) );
  AOI22_X1 U13070 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10804), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10290) );
  AOI22_X1 U13071 ( .A1(n9774), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U13072 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10457), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U13073 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10287) );
  NAND4_X1 U13074 ( .A1(n10290), .A2(n10289), .A3(n10288), .A4(n10224), .ZN(
        n10291) );
  AOI22_X1 U13075 ( .A1(n9750), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U13076 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9770), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10296) );
  AOI22_X1 U13077 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9771), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10295) );
  AOI22_X1 U13078 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10294) );
  AOI22_X1 U13079 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9765), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10300) );
  AOI22_X1 U13080 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10299) );
  AOI22_X1 U13081 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10804), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10298) );
  AOI22_X1 U13082 ( .A1(n10318), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10301) );
  NAND2_X1 U13083 ( .A1(n10302), .A2(n10339), .ZN(n10341) );
  INV_X1 U13084 ( .A(n10341), .ZN(n10358) );
  AOI22_X1 U13085 ( .A1(n9774), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(n9765), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U13086 ( .A1(n10636), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10801), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U13087 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13088 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10804), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10303) );
  NAND4_X1 U13089 ( .A1(n10306), .A2(n10305), .A3(n10304), .A4(n10303), .ZN(
        n10307) );
  NAND2_X1 U13090 ( .A1(n10307), .A2(n10456), .ZN(n10314) );
  AOI22_X1 U13091 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10457), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U13092 ( .A1(n10636), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10801), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10310) );
  AOI22_X1 U13093 ( .A1(n9774), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10804), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10309) );
  AOI22_X1 U13094 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10308) );
  NAND4_X1 U13095 ( .A1(n10311), .A2(n10310), .A3(n10309), .A4(n10308), .ZN(
        n10312) );
  NAND2_X1 U13096 ( .A1(n10312), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10313) );
  NAND2_X2 U13097 ( .A1(n10314), .A2(n10313), .ZN(n15876) );
  NAND2_X1 U13098 ( .A1(n10358), .A2(n15876), .ZN(n10316) );
  NAND4_X1 U13099 ( .A1(n11446), .A2(n19435), .A3(n10338), .A4(n10345), .ZN(
        n10315) );
  NOR2_X2 U13100 ( .A1(n10315), .A2(n10337), .ZN(n10349) );
  AOI22_X1 U13101 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9766), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10322) );
  AOI22_X1 U13102 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10457), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10321) );
  AOI22_X1 U13103 ( .A1(n9751), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(n9771), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U13104 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U13105 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9770), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U13106 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10325) );
  AOI22_X1 U13107 ( .A1(n9774), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U13108 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9771), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10323) );
  INV_X1 U13109 ( .A(n10327), .ZN(n11076) );
  NAND4_X1 U13110 ( .A1(n11454), .A2(n10863), .A3(n11076), .A4(n10447), .ZN(
        n10328) );
  NAND2_X1 U13111 ( .A1(n10381), .A2(n19422), .ZN(n10336) );
  NAND2_X1 U13112 ( .A1(n10332), .A2(n11431), .ZN(n11445) );
  INV_X2 U13113 ( .A(n10391), .ZN(n10431) );
  NAND2_X1 U13114 ( .A1(n10431), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10368) );
  INV_X1 U13115 ( .A(n10337), .ZN(n11066) );
  NAND3_X1 U13116 ( .A1(n10339), .A2(n11066), .A3(n10338), .ZN(n11408) );
  NOR2_X1 U13117 ( .A1(n9747), .A2(n11446), .ZN(n10340) );
  NAND2_X1 U13118 ( .A1(n11408), .A2(n10340), .ZN(n10342) );
  NAND2_X1 U13119 ( .A1(n10342), .A2(n10341), .ZN(n11439) );
  NAND2_X1 U13120 ( .A1(n11439), .A2(n15876), .ZN(n10344) );
  NAND4_X1 U13121 ( .A1(n19452), .A2(n10353), .A3(n19435), .A4(n10447), .ZN(
        n10354) );
  NAND2_X1 U13122 ( .A1(n10344), .A2(n10343), .ZN(n10352) );
  INV_X1 U13123 ( .A(n10928), .ZN(n10906) );
  MUX2_X1 U13124 ( .A(n10447), .B(n11457), .S(n10346), .Z(n10348) );
  AOI21_X1 U13125 ( .B1(n10447), .B2(n10338), .A(n11446), .ZN(n10347) );
  OAI211_X1 U13126 ( .C1(n10345), .C2(n10906), .A(n10348), .B(n10347), .ZN(
        n10351) );
  NOR2_X1 U13127 ( .A1(n10349), .A2(n15876), .ZN(n10350) );
  NAND2_X1 U13128 ( .A1(n10351), .A2(n10350), .ZN(n11450) );
  NAND2_X1 U13129 ( .A1(n10352), .A2(n11450), .ZN(n10369) );
  NAND2_X1 U13130 ( .A1(n10852), .A2(n19435), .ZN(n11458) );
  NAND2_X1 U13131 ( .A1(n10928), .A2(n10346), .ZN(n11456) );
  AND2_X1 U13132 ( .A1(n11461), .A2(n11457), .ZN(n10853) );
  NAND3_X1 U13133 ( .A1(n11458), .A2(n11456), .A3(n10853), .ZN(n10355) );
  NAND2_X1 U13134 ( .A1(n10355), .A2(n10862), .ZN(n11451) );
  NOR2_X1 U13135 ( .A1(n11451), .A2(n11452), .ZN(n10356) );
  NOR2_X1 U13136 ( .A1(n10369), .A2(n10356), .ZN(n10357) );
  NOR2_X1 U13137 ( .A1(n10447), .A2(n20119), .ZN(n13593) );
  NAND2_X1 U13138 ( .A1(n13593), .A2(n10331), .ZN(n10753) );
  NOR2_X1 U13139 ( .A1(n10753), .A2(n20109), .ZN(n10359) );
  AND2_X2 U13140 ( .A1(n16502), .A2(n10359), .ZN(n11635) );
  NOR2_X1 U13141 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11441) );
  INV_X1 U13142 ( .A(n11441), .ZN(n10361) );
  NAND2_X1 U13143 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10360) );
  NAND2_X1 U13144 ( .A1(n10361), .A2(n10360), .ZN(n10362) );
  AOI21_X1 U13145 ( .B1(n11635), .B2(P2_REIP_REG_0__SCAN_IN), .A(n10362), .ZN(
        n10365) );
  NAND2_X1 U13146 ( .A1(n11538), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10364) );
  INV_X1 U13147 ( .A(n10370), .ZN(n10371) );
  NAND2_X1 U13148 ( .A1(n9808), .A2(n10371), .ZN(n10374) );
  NAND2_X1 U13149 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n10372) );
  NAND2_X1 U13150 ( .A1(n9775), .A2(n10372), .ZN(n10373) );
  NAND2_X1 U13151 ( .A1(n10374), .A2(n10373), .ZN(n10377) );
  INV_X1 U13152 ( .A(n15840), .ZN(n10375) );
  AOI22_X1 U13153 ( .A1(n10375), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n11441), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10376) );
  NAND2_X1 U13154 ( .A1(n10377), .A2(n10376), .ZN(n10410) );
  INV_X1 U13155 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19398) );
  NAND2_X1 U13156 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10379) );
  NAND2_X1 U13157 ( .A1(n11635), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10378) );
  OAI211_X1 U13158 ( .C1(n11547), .C2(n13724), .A(n10379), .B(n10378), .ZN(
        n10380) );
  AOI21_X2 U13159 ( .B1(n10431), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10380), .ZN(n10384) );
  AOI22_X1 U13160 ( .A1(n10381), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n11441), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10382) );
  INV_X1 U13161 ( .A(n10384), .ZN(n10386) );
  AOI21_X1 U13162 ( .B1(n20119), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10389) );
  INV_X1 U13163 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11497) );
  INV_X1 U13164 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10394) );
  NAND2_X1 U13165 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10393) );
  NAND2_X1 U13166 ( .A1(n11635), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10392) );
  OAI211_X1 U13167 ( .C1(n9775), .C2(n10394), .A(n10393), .B(n10392), .ZN(
        n10395) );
  INV_X1 U13168 ( .A(n10395), .ZN(n10396) );
  AND2_X1 U13169 ( .A1(n20119), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n10437) );
  NAND2_X1 U13170 ( .A1(n11083), .A2(n10437), .ZN(n10403) );
  NAND2_X1 U13171 ( .A1(n10447), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10399) );
  INV_X1 U13172 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19879) );
  NAND2_X1 U13173 ( .A1(n10399), .A2(n19879), .ZN(n10442) );
  NOR2_X2 U13174 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20064) );
  NAND2_X1 U13175 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19517) );
  NAND2_X1 U13176 ( .A1(n19517), .A2(n20076), .ZN(n10401) );
  NAND2_X1 U13177 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15886) );
  INV_X1 U13178 ( .A(n15886), .ZN(n10400) );
  NAND2_X1 U13179 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10400), .ZN(
        n10438) );
  AND2_X1 U13180 ( .A1(n10401), .A2(n10438), .ZN(n19551) );
  AOI22_X1 U13181 ( .A1(n10442), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n20064), .B2(n19551), .ZN(n10402) );
  INV_X1 U13182 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10686) );
  OR2_X1 U13183 ( .A1(n10753), .A2(n10686), .ZN(n10418) );
  INV_X1 U13184 ( .A(n10414), .ZN(n10405) );
  XNOR2_X2 U13185 ( .A(n10406), .B(n10405), .ZN(n11087) );
  NAND2_X1 U13186 ( .A1(n10442), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10407) );
  NAND2_X1 U13187 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20085), .ZN(
        n19693) );
  NAND2_X1 U13188 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20092), .ZN(
        n19726) );
  AND2_X1 U13189 ( .A1(n19693), .A2(n19726), .ZN(n19550) );
  INV_X1 U13190 ( .A(n19550), .ZN(n19612) );
  NAND2_X1 U13191 ( .A1(n20064), .A2(n19612), .ZN(n19729) );
  NAND2_X1 U13192 ( .A1(n10407), .A2(n19729), .ZN(n10408) );
  AOI21_X1 U13193 ( .B1(n11087), .B2(n10437), .A(n10408), .ZN(n13599) );
  INV_X1 U13194 ( .A(n10409), .ZN(n10412) );
  INV_X1 U13195 ( .A(n10410), .ZN(n10411) );
  NAND2_X1 U13196 ( .A1(n10412), .A2(n10411), .ZN(n10413) );
  INV_X1 U13197 ( .A(n10437), .ZN(n13379) );
  AOI22_X1 U13198 ( .A1(n10442), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20064), .B2(n20092), .ZN(n10415) );
  OAI21_X2 U13199 ( .B1(n19200), .B2(n13379), .A(n10415), .ZN(n13596) );
  INV_X1 U13200 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11105) );
  OR2_X1 U13201 ( .A1(n10753), .A2(n11105), .ZN(n10416) );
  XNOR2_X1 U13202 ( .A(n13596), .B(n10416), .ZN(n13600) );
  NAND2_X1 U13203 ( .A1(n13599), .A2(n13600), .ZN(n13598) );
  INV_X1 U13204 ( .A(n13596), .ZN(n13750) );
  NAND2_X1 U13205 ( .A1(n13750), .A2(n10416), .ZN(n10417) );
  INV_X1 U13206 ( .A(n10418), .ZN(n10419) );
  NAND2_X1 U13207 ( .A1(n10420), .A2(n10419), .ZN(n10421) );
  NAND2_X1 U13208 ( .A1(n10424), .A2(n10422), .ZN(n10423) );
  INV_X1 U13209 ( .A(n10424), .ZN(n10426) );
  NAND2_X1 U13210 ( .A1(n11441), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10429) );
  INV_X1 U13211 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13590) );
  NAND2_X1 U13212 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10433) );
  NAND2_X1 U13213 ( .A1(n11635), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10432) );
  OAI211_X1 U13214 ( .C1(n9775), .C2(n13590), .A(n10433), .B(n10432), .ZN(
        n10434) );
  INV_X1 U13215 ( .A(n10434), .ZN(n10435) );
  NAND2_X1 U13216 ( .A1(n11101), .A2(n10437), .ZN(n10444) );
  INV_X1 U13217 ( .A(n10438), .ZN(n10439) );
  NAND2_X1 U13218 ( .A1(n10439), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19412) );
  OAI211_X1 U13219 ( .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n10439), .A(
        n19412), .B(n20064), .ZN(n10440) );
  INV_X1 U13220 ( .A(n10440), .ZN(n10441) );
  AOI21_X1 U13221 ( .B1(n10442), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10441), .ZN(n10443) );
  NAND2_X1 U13222 ( .A1(n10444), .A2(n10443), .ZN(n10450) );
  INV_X1 U13223 ( .A(n10753), .ZN(n10724) );
  AND2_X1 U13224 ( .A1(n10724), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10445) );
  OR2_X1 U13225 ( .A1(n10450), .A2(n10445), .ZN(n10446) );
  NAND2_X1 U13226 ( .A1(n10450), .A2(n10445), .ZN(n13883) );
  NAND2_X1 U13227 ( .A1(n13569), .A2(n13568), .ZN(n10449) );
  NAND2_X1 U13228 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n10447), .ZN(
        n10448) );
  AND2_X1 U13229 ( .A1(n10450), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10451) );
  AOI22_X1 U13230 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10897), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10455) );
  AND2_X1 U13231 ( .A1(n10806), .A2(n10456), .ZN(n10537) );
  AND2_X1 U13232 ( .A1(n10805), .A2(n10456), .ZN(n10561) );
  AOI22_X1 U13233 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10454) );
  AND2_X2 U13234 ( .A1(n10806), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10891) );
  AND2_X1 U13235 ( .A1(n9771), .A2(n10456), .ZN(n10500) );
  AOI22_X1 U13236 ( .A1(n10891), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10500), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10453) );
  AND2_X1 U13237 ( .A1(n10805), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10890) );
  AOI22_X1 U13238 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10452) );
  NAND4_X1 U13239 ( .A1(n10455), .A2(n10454), .A3(n10453), .A4(n10452), .ZN(
        n10463) );
  AND2_X2 U13240 ( .A1(n10797), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10560) );
  AND2_X1 U13241 ( .A1(n9751), .A2(n10456), .ZN(n10468) );
  AOI22_X1 U13242 ( .A1(n10560), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10461) );
  BUF_X4 U13243 ( .A(n10801), .Z(n10794) );
  AOI22_X1 U13245 ( .A1(n10469), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10896), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10460) );
  AND2_X1 U13246 ( .A1(n9770), .A2(n10456), .ZN(n10492) );
  AOI22_X1 U13247 ( .A1(n10984), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10492), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10459) );
  AND2_X1 U13248 ( .A1(n9766), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10940) );
  AOI22_X1 U13249 ( .A1(n10940), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10458) );
  NAND4_X1 U13250 ( .A1(n10461), .A2(n10460), .A3(n10459), .A4(n10458), .ZN(
        n10462) );
  OR2_X1 U13251 ( .A1(n10463), .A2(n10462), .ZN(n13766) );
  INV_X1 U13252 ( .A(n13765), .ZN(n10477) );
  AOI22_X1 U13253 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10560), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10467) );
  AOI22_X1 U13254 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10537), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10466) );
  AOI22_X1 U13255 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10500), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10465) );
  AOI22_X1 U13256 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10891), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10464) );
  NAND4_X1 U13257 ( .A1(n10467), .A2(n10466), .A3(n10465), .A4(n10464), .ZN(
        n10475) );
  AOI22_X1 U13258 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10468), .B1(
        n10897), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10473) );
  AOI22_X1 U13259 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10896), .B1(
        n10492), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U13260 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10469), .B1(
        n10984), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10471) );
  AOI22_X1 U13261 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10940), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10470) );
  NAND4_X1 U13262 ( .A1(n10473), .A2(n10472), .A3(n10471), .A4(n10470), .ZN(
        n10474) );
  NOR2_X1 U13263 ( .A1(n10475), .A2(n10474), .ZN(n13778) );
  INV_X1 U13264 ( .A(n13778), .ZN(n10476) );
  AOI22_X1 U13265 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10897), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10481) );
  AOI22_X1 U13266 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10500), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10480) );
  AOI22_X1 U13267 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10537), .B1(
        n10891), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U13268 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10561), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10478) );
  NAND4_X1 U13269 ( .A1(n10481), .A2(n10480), .A3(n10479), .A4(n10478), .ZN(
        n10487) );
  AOI22_X1 U13270 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10468), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13271 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10896), .B1(
        n10469), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U13272 ( .A1(n10572), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10492), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10483) );
  AOI22_X1 U13273 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10940), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10482) );
  NAND4_X1 U13274 ( .A1(n10485), .A2(n10484), .A3(n10483), .A4(n10482), .ZN(
        n10486) );
  OR2_X1 U13275 ( .A1(n10487), .A2(n10486), .ZN(n13940) );
  INV_X1 U13276 ( .A(n13940), .ZN(n11016) );
  AOI22_X1 U13277 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10491) );
  AOI22_X1 U13278 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13279 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U13280 ( .A1(n10891), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10488) );
  NAND4_X1 U13281 ( .A1(n10491), .A2(n10490), .A3(n10489), .A4(n10488), .ZN(
        n10498) );
  AOI22_X1 U13282 ( .A1(n10897), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10496) );
  AOI22_X1 U13283 ( .A1(n10492), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10896), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10495) );
  AOI22_X1 U13284 ( .A1(n10469), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10984), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10494) );
  AOI22_X1 U13285 ( .A1(n10940), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10493) );
  NAND4_X1 U13286 ( .A1(n10496), .A2(n10495), .A3(n10494), .A4(n10493), .ZN(
        n10497) );
  OR2_X1 U13287 ( .A1(n10498), .A2(n10497), .ZN(n14094) );
  AOI22_X1 U13288 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10504) );
  AOI22_X1 U13289 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U13290 ( .A1(n10891), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10502) );
  AOI22_X1 U13291 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10501) );
  NAND4_X1 U13292 ( .A1(n10504), .A2(n10503), .A3(n10502), .A4(n10501), .ZN(
        n10510) );
  AOI22_X1 U13293 ( .A1(n10560), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10897), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U13294 ( .A1(n10469), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10896), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U13295 ( .A1(n10984), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10492), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10506) );
  AOI22_X1 U13296 ( .A1(n10940), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10505) );
  NAND4_X1 U13297 ( .A1(n10508), .A2(n10507), .A3(n10506), .A4(n10505), .ZN(
        n10509) );
  OR2_X1 U13298 ( .A1(n10510), .A2(n10509), .ZN(n14093) );
  AND2_X1 U13299 ( .A1(n14094), .A2(n14093), .ZN(n10511) );
  AOI22_X1 U13300 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U13301 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U13302 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U13303 ( .A1(n10891), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10512) );
  NAND4_X1 U13304 ( .A1(n10515), .A2(n10514), .A3(n10513), .A4(n10512), .ZN(
        n10521) );
  AOI22_X1 U13305 ( .A1(n10897), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10519) );
  INV_X1 U13306 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10538) );
  AOI22_X1 U13307 ( .A1(n10492), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10896), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10518) );
  AOI22_X1 U13308 ( .A1(n10469), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10984), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10517) );
  AOI22_X1 U13309 ( .A1(n10940), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10516) );
  NAND4_X1 U13310 ( .A1(n10519), .A2(n10518), .A3(n10517), .A4(n10516), .ZN(
        n10520) );
  OR2_X1 U13311 ( .A1(n10521), .A2(n10520), .ZN(n14098) );
  AOI22_X1 U13312 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10468), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10525) );
  AOI22_X1 U13313 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10561), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10524) );
  AOI22_X1 U13314 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10891), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10523) );
  AOI22_X1 U13315 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10537), .B1(
        n10500), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10522) );
  NAND4_X1 U13316 ( .A1(n10525), .A2(n10524), .A3(n10523), .A4(n10522), .ZN(
        n10531) );
  AOI22_X1 U13317 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10897), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10529) );
  AOI22_X1 U13318 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10469), .B1(
        n10492), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10528) );
  AOI22_X1 U13319 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10896), .B1(
        n10984), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10527) );
  AOI22_X1 U13320 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10940), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10526) );
  NAND4_X1 U13321 ( .A1(n10529), .A2(n10528), .A3(n10527), .A4(n10526), .ZN(
        n10530) );
  OR2_X1 U13322 ( .A1(n10531), .A2(n10530), .ZN(n14100) );
  AND2_X1 U13323 ( .A1(n14098), .A2(n14100), .ZN(n10532) );
  AOI22_X1 U13324 ( .A1(n10897), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13325 ( .A1(n10492), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10896), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13326 ( .A1(n10469), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10984), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10534) );
  AOI22_X1 U13327 ( .A1(n10940), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10533) );
  NAND4_X1 U13328 ( .A1(n10536), .A2(n10535), .A3(n10534), .A4(n10533), .ZN(
        n10545) );
  AOI22_X1 U13329 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10543) );
  AOI22_X1 U13330 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10542) );
  AOI22_X1 U13331 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10541) );
  INV_X1 U13332 ( .A(n10891), .ZN(n10563) );
  INV_X1 U13333 ( .A(n10890), .ZN(n10562) );
  INV_X1 U13334 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11165) );
  OAI22_X1 U13335 ( .A1(n10538), .A2(n10563), .B1(n10562), .B2(n11165), .ZN(
        n10539) );
  INV_X1 U13336 ( .A(n10539), .ZN(n10540) );
  NAND4_X1 U13337 ( .A1(n10543), .A2(n10542), .A3(n10541), .A4(n10540), .ZN(
        n10544) );
  OR2_X1 U13338 ( .A1(n10545), .A2(n10544), .ZN(n15308) );
  AOI22_X1 U13339 ( .A1(n10897), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10549) );
  AOI22_X1 U13340 ( .A1(n10492), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10896), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10548) );
  AOI22_X1 U13341 ( .A1(n10469), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U13342 ( .A1(n10940), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10546) );
  NAND4_X1 U13343 ( .A1(n10549), .A2(n10548), .A3(n10547), .A4(n10546), .ZN(
        n10555) );
  AOI22_X1 U13344 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U13345 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10552) );
  AOI22_X1 U13346 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10551) );
  AOI22_X1 U13347 ( .A1(n10891), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10550) );
  NAND4_X1 U13348 ( .A1(n10553), .A2(n10552), .A3(n10551), .A4(n10550), .ZN(
        n10554) );
  NOR2_X1 U13349 ( .A1(n10555), .A2(n10554), .ZN(n15314) );
  AOI22_X1 U13350 ( .A1(n10897), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10559) );
  AOI22_X1 U13351 ( .A1(n10492), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10896), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10558) );
  AOI22_X1 U13352 ( .A1(n10469), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10984), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10557) );
  AOI22_X1 U13353 ( .A1(n10940), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10556) );
  NAND4_X1 U13354 ( .A1(n10559), .A2(n10558), .A3(n10557), .A4(n10556), .ZN(
        n10571) );
  AOI22_X1 U13355 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U13356 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U13357 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10567) );
  INV_X1 U13358 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10564) );
  INV_X1 U13359 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11142) );
  OAI22_X1 U13360 ( .A1(n10564), .A2(n10563), .B1(n10562), .B2(n11142), .ZN(
        n10565) );
  INV_X1 U13361 ( .A(n10565), .ZN(n10566) );
  NAND4_X1 U13362 ( .A1(n10569), .A2(n10568), .A3(n10567), .A4(n10566), .ZN(
        n10570) );
  OR2_X1 U13363 ( .A1(n10571), .A2(n10570), .ZN(n15321) );
  INV_X1 U13364 ( .A(n15321), .ZN(n15312) );
  NOR2_X1 U13365 ( .A1(n15314), .A2(n15312), .ZN(n15306) );
  AND2_X1 U13366 ( .A1(n15308), .A2(n15306), .ZN(n10583) );
  AOI22_X1 U13367 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10468), .B1(
        n10897), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10576) );
  AOI22_X1 U13368 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10896), .B1(
        n10492), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10575) );
  AOI22_X1 U13369 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10469), .B1(
        n10984), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10574) );
  AOI22_X1 U13370 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10940), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10573) );
  NAND4_X1 U13371 ( .A1(n10576), .A2(n10575), .A3(n10574), .A4(n10573), .ZN(
        n10582) );
  AOI22_X1 U13372 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n10560), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10580) );
  AOI22_X1 U13373 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10579) );
  AOI22_X1 U13374 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10500), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10578) );
  AOI22_X1 U13375 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10891), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10577) );
  NAND4_X1 U13376 ( .A1(n10580), .A2(n10579), .A3(n10578), .A4(n10577), .ZN(
        n10581) );
  OR2_X1 U13377 ( .A1(n10582), .A2(n10581), .ZN(n15326) );
  AND2_X1 U13378 ( .A1(n10583), .A2(n15326), .ZN(n15298) );
  AOI22_X1 U13379 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10499), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10587) );
  AOI22_X1 U13380 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n10537), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10586) );
  AOI22_X1 U13381 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10500), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10585) );
  AOI22_X1 U13382 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10891), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10584) );
  NAND4_X1 U13383 ( .A1(n10587), .A2(n10586), .A3(n10585), .A4(n10584), .ZN(
        n10593) );
  AOI22_X1 U13384 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10468), .B1(
        n10897), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10591) );
  AOI22_X1 U13385 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10896), .B1(
        n10492), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10590) );
  AOI22_X1 U13386 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10469), .B1(
        n10984), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U13387 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10940), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10588) );
  NAND4_X1 U13388 ( .A1(n10591), .A2(n10590), .A3(n10589), .A4(n10588), .ZN(
        n10592) );
  NOR2_X1 U13389 ( .A1(n10593), .A2(n10592), .ZN(n15299) );
  INV_X1 U13390 ( .A(n15299), .ZN(n10594) );
  AND2_X1 U13391 ( .A1(n15298), .A2(n10594), .ZN(n10605) );
  AOI22_X1 U13392 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10468), .B1(
        n10897), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10598) );
  AOI22_X1 U13393 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10896), .B1(
        n10492), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10597) );
  AOI22_X1 U13394 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10469), .B1(
        n10984), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10596) );
  AOI22_X1 U13395 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10940), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10595) );
  NAND4_X1 U13396 ( .A1(n10598), .A2(n10597), .A3(n10596), .A4(n10595), .ZN(
        n10604) );
  AOI22_X1 U13397 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10560), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10602) );
  AOI22_X1 U13398 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10537), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10601) );
  AOI22_X1 U13399 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10500), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10600) );
  AOI22_X1 U13400 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10891), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10599) );
  NAND4_X1 U13401 ( .A1(n10602), .A2(n10601), .A3(n10600), .A4(n10599), .ZN(
        n10603) );
  OR2_X1 U13402 ( .A1(n10604), .A2(n10603), .ZN(n15334) );
  NAND2_X1 U13403 ( .A1(n10605), .A2(n15334), .ZN(n10616) );
  AOI22_X1 U13404 ( .A1(n10897), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10609) );
  AOI22_X1 U13405 ( .A1(n10492), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10896), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10608) );
  AOI22_X1 U13406 ( .A1(n10469), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10984), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U13407 ( .A1(n10940), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10606) );
  NAND4_X1 U13408 ( .A1(n10609), .A2(n10608), .A3(n10607), .A4(n10606), .ZN(
        n10615) );
  AOI22_X1 U13409 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10613) );
  AOI22_X1 U13410 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10612) );
  AOI22_X1 U13411 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10611) );
  AOI22_X1 U13412 ( .A1(n10891), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10610) );
  NAND4_X1 U13413 ( .A1(n10613), .A2(n10612), .A3(n10611), .A4(n10610), .ZN(
        n10614) );
  NOR2_X1 U13414 ( .A1(n10615), .A2(n10614), .ZN(n15340) );
  OR2_X1 U13415 ( .A1(n10616), .A2(n15340), .ZN(n10628) );
  AOI22_X1 U13416 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n10560), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10621) );
  AOI22_X1 U13417 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10537), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U13418 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10500), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13419 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n10891), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10618) );
  NAND4_X1 U13420 ( .A1(n10621), .A2(n10620), .A3(n10619), .A4(n10618), .ZN(
        n10627) );
  AOI22_X1 U13421 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10468), .B1(
        n10897), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10625) );
  AOI22_X1 U13422 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10896), .B1(
        n10492), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10624) );
  AOI22_X1 U13423 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10469), .B1(
        n10984), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10623) );
  AOI22_X1 U13424 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10940), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10622) );
  NAND4_X1 U13425 ( .A1(n10625), .A2(n10624), .A3(n10623), .A4(n10622), .ZN(
        n10626) );
  OR2_X1 U13426 ( .A1(n10627), .A2(n10626), .ZN(n11034) );
  INV_X1 U13427 ( .A(n11034), .ZN(n15297) );
  OR2_X1 U13428 ( .A1(n10628), .A2(n15297), .ZN(n10629) );
  INV_X1 U13429 ( .A(n10773), .ZN(n10778) );
  INV_X1 U13430 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10631) );
  INV_X1 U13431 ( .A(n10804), .ZN(n10777) );
  INV_X1 U13432 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10630) );
  OAI22_X1 U13433 ( .A1(n10778), .A2(n10631), .B1(n10777), .B2(n10630), .ZN(
        n10635) );
  INV_X1 U13434 ( .A(n10805), .ZN(n10780) );
  INV_X1 U13435 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10633) );
  INV_X1 U13436 ( .A(n10806), .ZN(n10779) );
  INV_X1 U13437 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10632) );
  OAI22_X1 U13438 ( .A1(n10780), .A2(n10633), .B1(n10779), .B2(n10632), .ZN(
        n10634) );
  NOR2_X1 U13439 ( .A1(n10635), .A2(n10634), .ZN(n10639) );
  INV_X1 U13440 ( .A(n10636), .ZN(n15842) );
  AOI22_X1 U13441 ( .A1(n10797), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10638) );
  AOI22_X1 U13442 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10457), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10637) );
  XNOR2_X1 U13443 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10798) );
  NAND4_X1 U13444 ( .A1(n10639), .A2(n10638), .A3(n10637), .A4(n10798), .ZN(
        n10650) );
  INV_X1 U13445 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10641) );
  INV_X1 U13446 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10640) );
  OAI22_X1 U13447 ( .A1(n10778), .A2(n10641), .B1(n10777), .B2(n10640), .ZN(
        n10645) );
  INV_X1 U13448 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10643) );
  INV_X1 U13449 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10642) );
  OAI22_X1 U13450 ( .A1(n10780), .A2(n10643), .B1(n10779), .B2(n10642), .ZN(
        n10644) );
  NOR2_X1 U13451 ( .A1(n10645), .A2(n10644), .ZN(n10648) );
  INV_X1 U13452 ( .A(n10798), .ZN(n10807) );
  AOI22_X1 U13453 ( .A1(n10797), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10647) );
  AOI22_X1 U13454 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9770), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10646) );
  NAND4_X1 U13455 ( .A1(n10648), .A2(n10807), .A3(n10647), .A4(n10646), .ZN(
        n10649) );
  AND2_X1 U13456 ( .A1(n10650), .A2(n10649), .ZN(n10678) );
  NAND2_X1 U13457 ( .A1(n9748), .A2(n10678), .ZN(n10661) );
  AOI22_X1 U13458 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10468), .B1(
        n10897), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10654) );
  AOI22_X1 U13459 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10469), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U13460 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10896), .B1(
        n10492), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U13461 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10940), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10651) );
  NAND4_X1 U13462 ( .A1(n10654), .A2(n10653), .A3(n10652), .A4(n10651), .ZN(
        n10660) );
  AOI22_X1 U13463 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n10560), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U13464 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10891), .B1(
        n10500), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U13465 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10537), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10656) );
  AOI22_X1 U13466 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10617), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10655) );
  NAND4_X1 U13467 ( .A1(n10658), .A2(n10657), .A3(n10656), .A4(n10655), .ZN(
        n10659) );
  OR2_X1 U13468 ( .A1(n10660), .A2(n10659), .ZN(n10675) );
  XNOR2_X1 U13469 ( .A(n10661), .B(n10675), .ZN(n10680) );
  NAND2_X1 U13470 ( .A1(n19422), .A2(n10678), .ZN(n15293) );
  NOR2_X2 U13471 ( .A1(n15292), .A2(n10662), .ZN(n15282) );
  INV_X1 U13472 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11085) );
  OAI22_X1 U13473 ( .A1(n10778), .A2(n11105), .B1(n10777), .B2(n11085), .ZN(
        n10664) );
  INV_X1 U13474 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11089) );
  INV_X1 U13475 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11116) );
  OAI22_X1 U13476 ( .A1(n10780), .A2(n11089), .B1(n10779), .B2(n11116), .ZN(
        n10663) );
  NOR2_X1 U13477 ( .A1(n10664), .A2(n10663), .ZN(n10667) );
  AOI22_X1 U13478 ( .A1(n10797), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10666) );
  AOI22_X1 U13479 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9765), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10665) );
  NAND4_X1 U13480 ( .A1(n10667), .A2(n10666), .A3(n10665), .A4(n10798), .ZN(
        n10674) );
  INV_X1 U13481 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11097) );
  INV_X1 U13482 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11094) );
  OAI22_X1 U13483 ( .A1(n10778), .A2(n11097), .B1(n10777), .B2(n11094), .ZN(
        n10669) );
  INV_X1 U13484 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11121) );
  INV_X1 U13485 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11103) );
  OAI22_X1 U13486 ( .A1(n10780), .A2(n11121), .B1(n10779), .B2(n11103), .ZN(
        n10668) );
  NOR2_X1 U13487 ( .A1(n10669), .A2(n10668), .ZN(n10672) );
  AOI22_X1 U13488 ( .A1(n10797), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U13489 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9765), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10670) );
  NAND4_X1 U13490 ( .A1(n10672), .A2(n10807), .A3(n10671), .A4(n10670), .ZN(
        n10673) );
  NAND2_X1 U13491 ( .A1(n10674), .A2(n10673), .ZN(n10683) );
  NAND2_X1 U13492 ( .A1(n10675), .A2(n10678), .ZN(n10684) );
  XOR2_X1 U13493 ( .A(n10683), .B(n10684), .Z(n10676) );
  NAND2_X1 U13494 ( .A1(n10676), .A2(n10724), .ZN(n15281) );
  NOR2_X1 U13495 ( .A1(n15282), .A2(n15281), .ZN(n15280) );
  INV_X1 U13496 ( .A(n10683), .ZN(n10677) );
  NAND2_X1 U13497 ( .A1(n19422), .A2(n10677), .ZN(n15284) );
  INV_X1 U13498 ( .A(n10678), .ZN(n10679) );
  NOR2_X1 U13499 ( .A1(n15284), .A2(n10679), .ZN(n10681) );
  NOR2_X1 U13500 ( .A1(n10684), .A2(n10683), .ZN(n10704) );
  INV_X1 U13501 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10685) );
  OAI22_X1 U13502 ( .A1(n10778), .A2(n10686), .B1(n10777), .B2(n10685), .ZN(
        n10690) );
  INV_X1 U13503 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10688) );
  INV_X1 U13504 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10687) );
  OAI22_X1 U13505 ( .A1(n10780), .A2(n10688), .B1(n10779), .B2(n10687), .ZN(
        n10689) );
  NOR2_X1 U13506 ( .A1(n10690), .A2(n10689), .ZN(n10693) );
  AOI22_X1 U13507 ( .A1(n10797), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U13508 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9765), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10691) );
  NAND4_X1 U13509 ( .A1(n10693), .A2(n10692), .A3(n10691), .A4(n10798), .ZN(
        n10703) );
  INV_X1 U13510 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10694) );
  INV_X1 U13511 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n21076) );
  OAI22_X1 U13512 ( .A1(n9752), .A2(n10694), .B1(n10777), .B2(n21076), .ZN(
        n10698) );
  INV_X1 U13513 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10696) );
  INV_X1 U13514 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10695) );
  OAI22_X1 U13515 ( .A1(n10780), .A2(n10696), .B1(n10779), .B2(n10695), .ZN(
        n10697) );
  NOR2_X1 U13516 ( .A1(n10698), .A2(n10697), .ZN(n10701) );
  INV_X1 U13517 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n21107) );
  AOI22_X1 U13518 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10700) );
  AOI22_X1 U13519 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10457), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10699) );
  NAND4_X1 U13520 ( .A1(n10701), .A2(n10807), .A3(n10700), .A4(n10699), .ZN(
        n10702) );
  AND2_X1 U13521 ( .A1(n10703), .A2(n10702), .ZN(n10706) );
  NAND2_X1 U13522 ( .A1(n10704), .A2(n10706), .ZN(n10732) );
  OAI211_X1 U13523 ( .C1(n10704), .C2(n10706), .A(n10732), .B(n10724), .ZN(
        n10709) );
  XNOR2_X1 U13524 ( .A(n10708), .B(n10705), .ZN(n15276) );
  INV_X1 U13525 ( .A(n10706), .ZN(n10707) );
  NOR2_X1 U13526 ( .A1(n9748), .A2(n10707), .ZN(n15275) );
  NAND2_X1 U13527 ( .A1(n15276), .A2(n15275), .ZN(n15274) );
  INV_X1 U13528 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11136) );
  OAI22_X1 U13529 ( .A1(n10778), .A2(n10564), .B1(n10777), .B2(n11136), .ZN(
        n10713) );
  INV_X1 U13530 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11137) );
  INV_X1 U13531 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10711) );
  OAI22_X1 U13532 ( .A1(n10780), .A2(n11137), .B1(n10779), .B2(n10711), .ZN(
        n10712) );
  NOR2_X1 U13533 ( .A1(n10713), .A2(n10712), .ZN(n10716) );
  AOI22_X1 U13534 ( .A1(n10797), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10715) );
  AOI22_X1 U13535 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9770), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10714) );
  NAND4_X1 U13536 ( .A1(n10716), .A2(n10715), .A3(n10714), .A4(n10798), .ZN(
        n10723) );
  INV_X1 U13537 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11138) );
  OAI22_X1 U13538 ( .A1(n10778), .A2(n11138), .B1(n10777), .B2(n11142), .ZN(
        n10718) );
  INV_X1 U13539 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11134) );
  INV_X1 U13540 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11143) );
  OAI22_X1 U13541 ( .A1(n10780), .A2(n11134), .B1(n10779), .B2(n11143), .ZN(
        n10717) );
  NOR2_X1 U13542 ( .A1(n10718), .A2(n10717), .ZN(n10721) );
  AOI22_X1 U13543 ( .A1(n10797), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U13544 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10457), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10719) );
  NAND4_X1 U13545 ( .A1(n10721), .A2(n10807), .A3(n10720), .A4(n10719), .ZN(
        n10722) );
  AND2_X1 U13546 ( .A1(n10723), .A2(n10722), .ZN(n10726) );
  XNOR2_X1 U13547 ( .A(n10732), .B(n10726), .ZN(n10725) );
  NAND2_X1 U13548 ( .A1(n10725), .A2(n10724), .ZN(n10728) );
  INV_X1 U13549 ( .A(n10726), .ZN(n10731) );
  NOR2_X1 U13550 ( .A1(n9748), .A2(n10731), .ZN(n15267) );
  OR2_X1 U13551 ( .A1(n10732), .A2(n10731), .ZN(n10754) );
  INV_X1 U13552 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10734) );
  INV_X1 U13553 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10733) );
  OAI22_X1 U13554 ( .A1(n10778), .A2(n10734), .B1(n10777), .B2(n10733), .ZN(
        n10738) );
  INV_X1 U13555 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10736) );
  INV_X1 U13556 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10735) );
  OAI22_X1 U13557 ( .A1(n10780), .A2(n10736), .B1(n10779), .B2(n10735), .ZN(
        n10737) );
  NOR2_X1 U13558 ( .A1(n10738), .A2(n10737), .ZN(n10741) );
  AOI22_X1 U13559 ( .A1(n10797), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10740) );
  AOI22_X1 U13560 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9765), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10739) );
  NAND4_X1 U13561 ( .A1(n10741), .A2(n10740), .A3(n10739), .A4(n10798), .ZN(
        n10752) );
  INV_X1 U13562 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10743) );
  INV_X1 U13563 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10742) );
  OAI22_X1 U13564 ( .A1(n10778), .A2(n10743), .B1(n10777), .B2(n10742), .ZN(
        n10747) );
  INV_X1 U13565 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10745) );
  INV_X1 U13566 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10744) );
  OAI22_X1 U13567 ( .A1(n10780), .A2(n10745), .B1(n10779), .B2(n10744), .ZN(
        n10746) );
  NOR2_X1 U13568 ( .A1(n10747), .A2(n10746), .ZN(n10750) );
  AOI22_X1 U13569 ( .A1(n10797), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U13570 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10457), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10748) );
  NAND4_X1 U13571 ( .A1(n10750), .A2(n10807), .A3(n10749), .A4(n10748), .ZN(
        n10751) );
  NAND2_X1 U13572 ( .A1(n10752), .A2(n10751), .ZN(n10757) );
  NOR2_X1 U13573 ( .A1(n10754), .A2(n10757), .ZN(n15252) );
  AOI211_X1 U13574 ( .C1(n10754), .C2(n10757), .A(n10753), .B(n15252), .ZN(
        n10755) );
  NOR2_X1 U13575 ( .A1(n9748), .A2(n10757), .ZN(n15260) );
  INV_X1 U13576 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11175) );
  OAI22_X1 U13577 ( .A1(n10778), .A2(n10538), .B1(n10777), .B2(n11175), .ZN(
        n10760) );
  INV_X1 U13578 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11186) );
  INV_X1 U13579 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10758) );
  OAI22_X1 U13580 ( .A1(n10780), .A2(n11186), .B1(n10779), .B2(n10758), .ZN(
        n10759) );
  NOR2_X1 U13581 ( .A1(n10760), .A2(n10759), .ZN(n10763) );
  AOI22_X1 U13582 ( .A1(n9774), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U13583 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10457), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10761) );
  NAND4_X1 U13584 ( .A1(n10763), .A2(n10762), .A3(n10761), .A4(n10798), .ZN(
        n10770) );
  INV_X1 U13585 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11178) );
  OAI22_X1 U13586 ( .A1(n10778), .A2(n11178), .B1(n10777), .B2(n11165), .ZN(
        n10765) );
  INV_X1 U13587 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11172) );
  INV_X1 U13588 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11167) );
  OAI22_X1 U13589 ( .A1(n10780), .A2(n11172), .B1(n10779), .B2(n11167), .ZN(
        n10764) );
  NOR2_X1 U13590 ( .A1(n10765), .A2(n10764), .ZN(n10768) );
  AOI22_X1 U13591 ( .A1(n10797), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10767) );
  AOI22_X1 U13592 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9765), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10766) );
  NAND4_X1 U13593 ( .A1(n10768), .A2(n10807), .A3(n10767), .A4(n10766), .ZN(
        n10769) );
  NAND2_X1 U13594 ( .A1(n10770), .A2(n10769), .ZN(n10788) );
  INV_X1 U13595 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11258) );
  INV_X1 U13596 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11251) );
  OAI22_X1 U13597 ( .A1(n9753), .A2(n11258), .B1(n10780), .B2(n11251), .ZN(
        n10772) );
  INV_X1 U13598 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11260) );
  INV_X1 U13599 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11259) );
  OAI22_X1 U13600 ( .A1(n10777), .A2(n11260), .B1(n10779), .B2(n11259), .ZN(
        n10771) );
  NOR2_X1 U13601 ( .A1(n10772), .A2(n10771), .ZN(n10776) );
  AOI22_X1 U13602 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10775) );
  AOI22_X1 U13603 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10457), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10774) );
  NAND4_X1 U13604 ( .A1(n10776), .A2(n10775), .A3(n10774), .A4(n10798), .ZN(
        n10787) );
  INV_X1 U13605 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11253) );
  INV_X1 U13606 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11242) );
  OAI22_X1 U13607 ( .A1(n10778), .A2(n11253), .B1(n10777), .B2(n11242), .ZN(
        n10782) );
  INV_X1 U13608 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11248) );
  INV_X1 U13609 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11244) );
  OAI22_X1 U13610 ( .A1(n10780), .A2(n11248), .B1(n10779), .B2(n11244), .ZN(
        n10781) );
  NOR2_X1 U13611 ( .A1(n10782), .A2(n10781), .ZN(n10785) );
  AOI22_X1 U13612 ( .A1(n9750), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10794), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10784) );
  AOI22_X1 U13613 ( .A1(n10636), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9770), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10783) );
  NAND4_X1 U13614 ( .A1(n10785), .A2(n10807), .A3(n10784), .A4(n10783), .ZN(
        n10786) );
  NAND2_X1 U13615 ( .A1(n10787), .A2(n10786), .ZN(n10791) );
  INV_X1 U13616 ( .A(n10788), .ZN(n15254) );
  AND2_X1 U13617 ( .A1(n9748), .A2(n15254), .ZN(n10789) );
  NAND2_X1 U13618 ( .A1(n15252), .A2(n10789), .ZN(n10790) );
  NOR2_X1 U13619 ( .A1(n10790), .A2(n10791), .ZN(n10792) );
  AOI21_X1 U13620 ( .B1(n10791), .B2(n10790), .A(n10792), .ZN(n15247) );
  INV_X1 U13621 ( .A(n10792), .ZN(n10793) );
  AOI22_X1 U13622 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10796) );
  AOI22_X1 U13623 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10457), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10795) );
  NAND2_X1 U13624 ( .A1(n10796), .A2(n10795), .ZN(n10813) );
  AOI22_X1 U13625 ( .A1(n9774), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(n9771), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10800) );
  AOI22_X1 U13626 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10799) );
  NAND3_X1 U13627 ( .A1(n10800), .A2(n10799), .A3(n10798), .ZN(n10812) );
  AOI22_X1 U13628 ( .A1(n10797), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U13629 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9765), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10802) );
  NAND2_X1 U13630 ( .A1(n10803), .A2(n10802), .ZN(n10811) );
  AOI22_X1 U13631 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9771), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U13632 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10808) );
  NAND3_X1 U13633 ( .A1(n10809), .A2(n10808), .A3(n10807), .ZN(n10810) );
  OAI22_X1 U13634 ( .A1(n10813), .A2(n10812), .B1(n10811), .B2(n10810), .ZN(
        n10814) );
  NAND2_X1 U13635 ( .A1(n15876), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19289) );
  NAND2_X1 U13636 ( .A1(n19289), .A2(n9748), .ZN(n10818) );
  MUX2_X1 U13637 ( .A(n20085), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n10819) );
  NAND2_X1 U13638 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20092), .ZN(
        n10820) );
  INV_X1 U13639 ( .A(n10820), .ZN(n10815) );
  NAND2_X1 U13640 ( .A1(n10819), .A2(n10815), .ZN(n10821) );
  NAND2_X1 U13641 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20085), .ZN(
        n10816) );
  NAND2_X1 U13642 ( .A1(n10821), .A2(n10816), .ZN(n10833) );
  XNOR2_X1 U13643 ( .A(n20076), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10817) );
  XNOR2_X1 U13644 ( .A(n10833), .B(n10817), .ZN(n11201) );
  MUX2_X1 U13645 ( .A(n10818), .B(n11431), .S(n11201), .Z(n10831) );
  OAI21_X1 U13646 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20092), .A(
        n10820), .ZN(n10827) );
  INV_X1 U13647 ( .A(n10827), .ZN(n11411) );
  INV_X1 U13648 ( .A(n10819), .ZN(n10826) );
  NAND2_X1 U13649 ( .A1(n10826), .A2(n10820), .ZN(n11412) );
  AND2_X1 U13650 ( .A1(n11412), .A2(n10821), .ZN(n10860) );
  OAI21_X1 U13651 ( .B1(n9748), .B2(n11411), .A(n10860), .ZN(n10823) );
  NAND2_X1 U13652 ( .A1(n19422), .A2(n11201), .ZN(n10822) );
  NAND2_X1 U13653 ( .A1(n10823), .A2(n10822), .ZN(n10824) );
  NAND2_X1 U13654 ( .A1(n10824), .A2(n20109), .ZN(n10829) );
  OAI21_X1 U13655 ( .B1(n10827), .B2(n10826), .A(n10825), .ZN(n10828) );
  NAND2_X1 U13656 ( .A1(n10829), .A2(n10828), .ZN(n10830) );
  NAND2_X1 U13657 ( .A1(n10831), .A2(n10830), .ZN(n10840) );
  OAI22_X1 U13658 ( .A1(n10833), .A2(n10832), .B1(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20076), .ZN(n10839) );
  MUX2_X1 U13659 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n20069), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10837) );
  OR2_X1 U13660 ( .A1(n10839), .A2(n10837), .ZN(n10835) );
  NAND2_X1 U13661 ( .A1(n20069), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10834) );
  INV_X1 U13662 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16493) );
  NOR2_X1 U13663 ( .A1(n16493), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10836) );
  NAND2_X1 U13664 ( .A1(n10842), .A2(n10836), .ZN(n11213) );
  INV_X1 U13665 ( .A(n10837), .ZN(n10838) );
  XNOR2_X1 U13666 ( .A(n10839), .B(n10838), .ZN(n11207) );
  MUX2_X1 U13667 ( .A(n11431), .B(n10840), .S(n11415), .Z(n10845) );
  NAND2_X1 U13668 ( .A1(n16493), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10841) );
  NAND2_X1 U13669 ( .A1(n10842), .A2(n10841), .ZN(n10844) );
  INV_X1 U13670 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13444) );
  NAND2_X1 U13671 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13444), .ZN(
        n10843) );
  NAND2_X1 U13672 ( .A1(n10845), .A2(n20098), .ZN(n10846) );
  MUX2_X1 U13673 ( .A(n10846), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n20119), .Z(n11424) );
  INV_X1 U13674 ( .A(n20098), .ZN(n10848) );
  INV_X1 U13675 ( .A(n19289), .ZN(n10847) );
  NAND2_X1 U13676 ( .A1(n10848), .A2(n10847), .ZN(n10849) );
  NAND2_X1 U13677 ( .A1(n11456), .A2(n10317), .ZN(n10851) );
  NAND2_X1 U13678 ( .A1(n10850), .A2(n10851), .ZN(n10857) );
  AND2_X1 U13679 ( .A1(n19422), .A2(n15876), .ZN(n20106) );
  OAI21_X1 U13680 ( .B1(n10852), .B2(n19452), .A(n20106), .ZN(n11460) );
  NAND2_X1 U13681 ( .A1(n10346), .A2(n19422), .ZN(n10858) );
  NAND2_X1 U13682 ( .A1(n10858), .A2(n20109), .ZN(n10854) );
  NAND2_X1 U13683 ( .A1(n10854), .A2(n10853), .ZN(n10855) );
  NAND2_X1 U13684 ( .A1(n10855), .A2(n10317), .ZN(n10856) );
  NAND4_X1 U13685 ( .A1(n10857), .A2(n11460), .A3(n11458), .A4(n10856), .ZN(
        n11421) );
  AND2_X1 U13686 ( .A1(n11201), .A2(n11415), .ZN(n11406) );
  NAND2_X1 U13687 ( .A1(n10860), .A2(n11406), .ZN(n10861) );
  NAND2_X1 U13688 ( .A1(n20098), .A2(n10861), .ZN(n16473) );
  NOR2_X1 U13689 ( .A1(n10859), .A2(n16473), .ZN(n13309) );
  NAND2_X1 U13690 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20118) );
  AND2_X1 U13691 ( .A1(n11445), .A2(n20118), .ZN(n13311) );
  AOI22_X1 U13692 ( .A1(n16478), .A2(n11443), .B1(n13309), .B2(n13311), .ZN(
        n13438) );
  INV_X1 U13693 ( .A(n10862), .ZN(n10865) );
  AND2_X1 U13694 ( .A1(n10863), .A2(n10317), .ZN(n10864) );
  NAND2_X1 U13695 ( .A1(n10865), .A2(n10864), .ZN(n11448) );
  NAND2_X1 U13696 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13298), .ZN(n13195) );
  INV_X1 U13697 ( .A(n13195), .ZN(n10866) );
  AND2_X1 U13698 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10866), .ZN(n20123) );
  NAND2_X1 U13699 ( .A1(n19270), .A2(n10906), .ZN(n19275) );
  NAND2_X1 U13700 ( .A1(n11433), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n10869) );
  NOR2_X1 U13701 ( .A1(n9747), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10914) );
  BUF_X1 U13702 ( .A(n10914), .Z(n11063) );
  NOR2_X1 U13703 ( .A1(n11457), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10870) );
  AOI22_X1 U13704 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n10868) );
  NAND2_X1 U13705 ( .A1(n10869), .A2(n10868), .ZN(n11432) );
  AOI222_X1 U13706 ( .A1(n11433), .A2(P2_REIP_REG_7__SCAN_IN), .B1(n11063), 
        .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n11434), .C2(
        P2_EAX_REG_7__SCAN_IN), .ZN(n15812) );
  NAND2_X1 U13707 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10874) );
  NAND2_X1 U13708 ( .A1(n10560), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10873) );
  NAND2_X1 U13709 ( .A1(n10891), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10872) );
  NAND2_X1 U13710 ( .A1(n10890), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10871) );
  NAND2_X1 U13711 ( .A1(n10897), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10878) );
  NAND2_X1 U13712 ( .A1(n10468), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10877) );
  NAND2_X1 U13713 ( .A1(n10492), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10876) );
  NAND2_X1 U13714 ( .A1(n10896), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10875) );
  NAND2_X1 U13715 ( .A1(n10561), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10882) );
  NAND2_X1 U13716 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10881) );
  NAND2_X1 U13717 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10880) );
  NAND2_X1 U13718 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10879) );
  NAND2_X1 U13719 ( .A1(n10469), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10886) );
  NAND2_X1 U13720 ( .A1(n10984), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10885) );
  NAND2_X1 U13721 ( .A1(n10940), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10884) );
  NAND2_X1 U13722 ( .A1(n10986), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10883) );
  NAND4_X1 U13723 ( .A1(n10889), .A2(n10888), .A3(n10887), .A4(n10211), .ZN(
        n11200) );
  INV_X1 U13724 ( .A(n11200), .ZN(n11322) );
  INV_X1 U13725 ( .A(n11030), .ZN(n10904) );
  AOI22_X1 U13726 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U13727 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U13728 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10893) );
  AOI22_X1 U13729 ( .A1(n10891), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10892) );
  NAND4_X1 U13730 ( .A1(n10895), .A2(n10894), .A3(n10893), .A4(n10892), .ZN(
        n10903) );
  AOI22_X1 U13731 ( .A1(n10469), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10901) );
  AOI22_X1 U13732 ( .A1(n10492), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10896), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10900) );
  AOI22_X1 U13733 ( .A1(n10897), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10899) );
  AOI22_X1 U13734 ( .A1(n10940), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10898) );
  NAND4_X1 U13735 ( .A1(n10901), .A2(n10900), .A3(n10899), .A4(n10898), .ZN(
        n10902) );
  NAND2_X1 U13736 ( .A1(n10904), .A2(n11492), .ZN(n10908) );
  AND2_X1 U13737 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10905) );
  NOR2_X1 U13738 ( .A1(n10870), .A2(n10905), .ZN(n10907) );
  NAND2_X1 U13739 ( .A1(n10914), .A2(n10906), .ZN(n10944) );
  NAND3_X1 U13740 ( .A1(n10908), .A2(n10907), .A3(n10944), .ZN(n13254) );
  NAND2_X1 U13741 ( .A1(n11023), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10913) );
  INV_X1 U13742 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19399) );
  NAND2_X1 U13743 ( .A1(n19452), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n10909) );
  OAI211_X1 U13744 ( .C1(n9747), .C2(n19399), .A(n10909), .B(n19879), .ZN(
        n10911) );
  INV_X1 U13745 ( .A(n10911), .ZN(n10912) );
  NAND2_X1 U13746 ( .A1(n10913), .A2(n10912), .ZN(n13255) );
  NAND2_X1 U13747 ( .A1(n13254), .A2(n13255), .ZN(n13258) );
  NAND2_X1 U13748 ( .A1(n11023), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U13749 ( .A1(n10914), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n10870), .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n10915) );
  AND2_X1 U13750 ( .A1(n10916), .A2(n10915), .ZN(n10934) );
  INV_X1 U13751 ( .A(n10934), .ZN(n10917) );
  XNOR2_X1 U13752 ( .A(n13258), .B(n10917), .ZN(n13716) );
  AOI22_X1 U13753 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n10560), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10921) );
  AOI22_X1 U13754 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10537), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10920) );
  AOI22_X1 U13755 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10492), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10919) );
  AOI22_X1 U13756 ( .A1(n10897), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10896), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10918) );
  NAND4_X1 U13757 ( .A1(n10921), .A2(n10920), .A3(n10919), .A4(n10918), .ZN(
        n10927) );
  AOI22_X1 U13758 ( .A1(n10468), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10469), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10925) );
  AOI22_X1 U13759 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n10891), .B1(
        n10500), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U13760 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10572), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U13761 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10940), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10922) );
  NAND4_X1 U13762 ( .A1(n10925), .A2(n10924), .A3(n10923), .A4(n10922), .ZN(
        n10926) );
  NOR2_X1 U13763 ( .A1(n10927), .A2(n10926), .ZN(n11493) );
  INV_X1 U13765 ( .A(n11205), .ZN(n10933) );
  NAND2_X1 U13766 ( .A1(n10928), .A2(n11457), .ZN(n10929) );
  MUX2_X1 U13767 ( .A(n10929), .B(n20085), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10930) );
  INV_X1 U13768 ( .A(n10930), .ZN(n10931) );
  AOI21_X1 U13769 ( .B1(n10933), .B2(n10932), .A(n10931), .ZN(n13717) );
  NAND2_X1 U13770 ( .A1(n13716), .A2(n13717), .ZN(n13721) );
  NAND2_X1 U13771 ( .A1(n10934), .A2(n13258), .ZN(n10935) );
  NAND2_X1 U13772 ( .A1(n13721), .A2(n10935), .ZN(n10949) );
  AOI22_X1 U13773 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10468), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U13774 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n10891), .B1(
        n10500), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U13775 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10537), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U13776 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10561), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10936) );
  NAND4_X1 U13777 ( .A1(n10939), .A2(n10938), .A3(n10937), .A4(n10936), .ZN(
        n10943) );
  AOI22_X1 U13778 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10897), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U13779 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10492), .B1(
        n10940), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10941) );
  INV_X1 U13780 ( .A(n11202), .ZN(n11500) );
  OR2_X1 U13781 ( .A1(n11030), .A2(n11500), .ZN(n10945) );
  OAI211_X1 U13782 ( .C1(n19879), .C2(n20076), .A(n10945), .B(n10944), .ZN(
        n10948) );
  XNOR2_X1 U13783 ( .A(n10949), .B(n10948), .ZN(n13270) );
  NAND2_X1 U13784 ( .A1(n11433), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10947) );
  AOI22_X1 U13785 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n10946) );
  NAND2_X1 U13786 ( .A1(n13270), .A2(n13269), .ZN(n13271) );
  INV_X1 U13787 ( .A(n10948), .ZN(n10950) );
  NAND2_X1 U13788 ( .A1(n10950), .A2(n10949), .ZN(n10951) );
  NAND2_X1 U13789 ( .A1(n13271), .A2(n10951), .ZN(n13573) );
  NAND2_X1 U13790 ( .A1(n11433), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10967) );
  NAND2_X1 U13791 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10954) );
  NOR2_X1 U13792 ( .A1(n20069), .A2(n19879), .ZN(n10952) );
  AOI21_X1 U13793 ( .B1(n11434), .B2(P2_EAX_REG_3__SCAN_IN), .A(n10952), .ZN(
        n10953) );
  AND2_X1 U13794 ( .A1(n10954), .A2(n10953), .ZN(n10966) );
  AOI22_X1 U13795 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10897), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10958) );
  AOI22_X1 U13796 ( .A1(n10891), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10500), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U13797 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10956) );
  AOI22_X1 U13798 ( .A1(n10561), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10955) );
  NAND4_X1 U13799 ( .A1(n10958), .A2(n10957), .A3(n10956), .A4(n10955), .ZN(
        n10964) );
  AOI22_X1 U13800 ( .A1(n10560), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10962) );
  AOI22_X1 U13801 ( .A1(n10469), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10492), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10961) );
  AOI22_X1 U13802 ( .A1(n10984), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10940), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U13803 ( .A1(n10896), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10959) );
  NAND4_X1 U13804 ( .A1(n10962), .A2(n10961), .A3(n10960), .A4(n10959), .ZN(
        n10963) );
  INV_X1 U13805 ( .A(n11206), .ZN(n11161) );
  OR2_X1 U13806 ( .A1(n11030), .A2(n11161), .ZN(n10965) );
  AOI22_X1 U13807 ( .A1(n10560), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10971) );
  AOI22_X1 U13808 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U13809 ( .A1(n10891), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10500), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10969) );
  AOI22_X1 U13810 ( .A1(n10561), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10968) );
  NAND4_X1 U13811 ( .A1(n10971), .A2(n10970), .A3(n10969), .A4(n10968), .ZN(
        n10977) );
  AOI22_X1 U13812 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10897), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10975) );
  AOI22_X1 U13813 ( .A1(n10469), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10984), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10974) );
  AOI22_X1 U13814 ( .A1(n10492), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10896), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10973) );
  AOI22_X1 U13815 ( .A1(n10940), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10972) );
  NAND4_X1 U13816 ( .A1(n10975), .A2(n10974), .A3(n10973), .A4(n10972), .ZN(
        n10976) );
  NAND2_X1 U13817 ( .A1(n11433), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n10979) );
  AOI22_X1 U13818 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n10978) );
  OAI211_X1 U13819 ( .C1(n11030), .C2(n11490), .A(n10979), .B(n10978), .ZN(
        n13892) );
  AOI22_X1 U13820 ( .A1(n10499), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10983) );
  AOI22_X1 U13821 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10982) );
  AOI22_X1 U13822 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10981) );
  AOI22_X1 U13823 ( .A1(n10891), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10980) );
  NAND4_X1 U13824 ( .A1(n10983), .A2(n10982), .A3(n10981), .A4(n10980), .ZN(
        n10992) );
  AOI22_X1 U13825 ( .A1(n10897), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10990) );
  AOI22_X1 U13826 ( .A1(n10492), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10896), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10989) );
  INV_X1 U13827 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n20948) );
  AOI22_X1 U13828 ( .A1(n10469), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10984), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10988) );
  AOI22_X1 U13829 ( .A1(n10940), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10987) );
  NAND4_X1 U13830 ( .A1(n10990), .A2(n10989), .A3(n10988), .A4(n10987), .ZN(
        n10991) );
  NAND2_X1 U13831 ( .A1(n11433), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U13832 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n10993) );
  OAI211_X1 U13833 ( .C1(n11030), .C2(n11215), .A(n10994), .B(n10993), .ZN(
        n16442) );
  AOI22_X1 U13834 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10560), .B1(
        n10499), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U13835 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10537), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10997) );
  AOI22_X1 U13836 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10500), .B1(
        n10617), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10996) );
  AOI22_X1 U13837 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n10891), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10995) );
  NAND4_X1 U13838 ( .A1(n10998), .A2(n10997), .A3(n10996), .A4(n10995), .ZN(
        n11004) );
  AOI22_X1 U13839 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10897), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11002) );
  AOI22_X1 U13840 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10492), .B1(
        n10896), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11001) );
  AOI22_X1 U13841 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10469), .B1(
        n10984), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U13842 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10940), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10999) );
  NAND4_X1 U13843 ( .A1(n11002), .A2(n11001), .A3(n11000), .A4(n10999), .ZN(
        n11003) );
  OR2_X1 U13844 ( .A1(n11030), .A2(n11278), .ZN(n11005) );
  NAND2_X1 U13845 ( .A1(n11433), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11007) );
  AOI22_X1 U13846 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n11006) );
  NAND2_X1 U13847 ( .A1(n11007), .A2(n11006), .ZN(n15825) );
  INV_X1 U13848 ( .A(n13766), .ZN(n11010) );
  NAND2_X1 U13849 ( .A1(n11433), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11009) );
  AOI22_X1 U13850 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n11008) );
  OAI211_X1 U13851 ( .C1(n11030), .C2(n11010), .A(n11009), .B(n11008), .ZN(
        n16432) );
  NAND2_X1 U13852 ( .A1(n11433), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11013) );
  AOI22_X1 U13853 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n11012) );
  OR2_X1 U13854 ( .A1(n11030), .A2(n13778), .ZN(n11011) );
  NAND2_X1 U13855 ( .A1(n11433), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11015) );
  AOI22_X1 U13856 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n11014) );
  OAI211_X1 U13857 ( .C1(n11030), .C2(n11016), .A(n11015), .B(n11014), .ZN(
        n16421) );
  NAND2_X1 U13858 ( .A1(n15793), .A2(n16421), .ZN(n16408) );
  INV_X1 U13859 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n11018) );
  AOI22_X1 U13860 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n11017) );
  OAI21_X1 U13861 ( .B1(n11065), .B2(n11018), .A(n11017), .ZN(n11019) );
  AOI21_X1 U13862 ( .B1(n10904), .B2(n14094), .A(n11019), .ZN(n16409) );
  INV_X1 U13863 ( .A(n14093), .ZN(n11022) );
  NAND2_X1 U13864 ( .A1(n11433), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11021) );
  AOI22_X1 U13865 ( .A1(n10914), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n11020) );
  OAI211_X1 U13866 ( .C1(n11030), .C2(n11022), .A(n11021), .B(n11020), .ZN(
        n15775) );
  NAND2_X1 U13867 ( .A1(n15774), .A2(n15775), .ZN(n16396) );
  INV_X1 U13868 ( .A(n11023), .ZN(n11065) );
  INV_X1 U13869 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n11025) );
  AOI22_X1 U13870 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n11024) );
  OAI21_X1 U13871 ( .B1(n11065), .B2(n11025), .A(n11024), .ZN(n11026) );
  AOI21_X1 U13872 ( .B1(n10904), .B2(n14098), .A(n11026), .ZN(n16397) );
  INV_X1 U13873 ( .A(n14100), .ZN(n11029) );
  NAND2_X1 U13874 ( .A1(n11433), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11028) );
  AOI22_X1 U13875 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n11027) );
  OAI211_X1 U13876 ( .C1(n11030), .C2(n11029), .A(n11028), .B(n11027), .ZN(
        n15762) );
  INV_X1 U13877 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n11032) );
  AOI22_X1 U13878 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n11031) );
  OAI21_X1 U13879 ( .B1(n11065), .B2(n11032), .A(n11031), .ZN(n11033) );
  AOI21_X1 U13880 ( .B1(n10904), .B2(n11034), .A(n11033), .ZN(n16385) );
  NAND2_X1 U13881 ( .A1(n11433), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11036) );
  AOI22_X1 U13882 ( .A1(n10914), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n11035) );
  NAND2_X1 U13883 ( .A1(n11036), .A2(n11035), .ZN(n14460) );
  NAND2_X1 U13884 ( .A1(n11433), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11038) );
  AOI22_X1 U13885 ( .A1(n10914), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n11037) );
  AND2_X1 U13886 ( .A1(n11038), .A2(n11037), .ZN(n14438) );
  NAND2_X1 U13887 ( .A1(n11433), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11042) );
  AOI22_X1 U13888 ( .A1(n10914), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n11041) );
  AND2_X1 U13889 ( .A1(n11042), .A2(n11041), .ZN(n15429) );
  NAND2_X1 U13890 ( .A1(n11433), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11045) );
  AOI22_X1 U13891 ( .A1(n10914), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n11044) );
  AND2_X1 U13892 ( .A1(n11045), .A2(n11044), .ZN(n14396) );
  INV_X1 U13893 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20025) );
  AOI22_X1 U13894 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n11046) );
  OAI21_X1 U13895 ( .B1(n11065), .B2(n20025), .A(n11046), .ZN(n15414) );
  NAND2_X1 U13896 ( .A1(n15415), .A2(n15414), .ZN(n13244) );
  NAND2_X1 U13897 ( .A1(n11433), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11048) );
  AOI22_X1 U13898 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n11047) );
  AND2_X1 U13899 ( .A1(n11048), .A2(n11047), .ZN(n13245) );
  INV_X1 U13900 ( .A(n13245), .ZN(n11049) );
  NAND2_X1 U13901 ( .A1(n11433), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11052) );
  AOI22_X1 U13902 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n11051) );
  AND2_X1 U13903 ( .A1(n11052), .A2(n11051), .ZN(n15399) );
  NAND2_X1 U13904 ( .A1(n11433), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U13905 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n11053) );
  NAND2_X1 U13906 ( .A1(n11054), .A2(n11053), .ZN(n15698) );
  INV_X1 U13907 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20033) );
  AOI22_X1 U13908 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n11055) );
  OAI21_X1 U13909 ( .B1(n11065), .B2(n20033), .A(n11055), .ZN(n15390) );
  NAND2_X1 U13910 ( .A1(n11433), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11057) );
  AOI22_X1 U13911 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n11056) );
  AND2_X1 U13912 ( .A1(n11057), .A2(n11056), .ZN(n15381) );
  NAND2_X1 U13913 ( .A1(n11433), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11059) );
  AOI22_X1 U13914 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n11058) );
  AND2_X1 U13915 ( .A1(n11059), .A2(n11058), .ZN(n15371) );
  NAND2_X1 U13916 ( .A1(n11433), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11061) );
  AOI22_X1 U13917 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n11060) );
  AND2_X1 U13918 ( .A1(n11061), .A2(n11060), .ZN(n15364) );
  INV_X1 U13919 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20041) );
  AOI22_X1 U13920 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n11062) );
  OAI21_X1 U13921 ( .B1(n11065), .B2(n20041), .A(n11062), .ZN(n13291) );
  INV_X1 U13922 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20043) );
  AOI22_X1 U13923 ( .A1(n11063), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n11064) );
  OAI21_X1 U13924 ( .B1(n11065), .B2(n20043), .A(n11064), .ZN(n15347) );
  AND2_X1 U13925 ( .A1(n11066), .A2(n19270), .ZN(n13896) );
  NOR4_X1 U13926 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n11070) );
  NOR4_X1 U13927 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n11069) );
  NOR4_X1 U13928 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n11068) );
  NOR4_X1 U13929 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n11067) );
  NAND4_X1 U13930 ( .A1(n11070), .A2(n11069), .A3(n11068), .A4(n11067), .ZN(
        n11075) );
  NOR4_X1 U13931 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_15__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n11073) );
  NOR4_X1 U13932 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n11072) );
  NOR4_X1 U13933 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n11071) );
  INV_X1 U13934 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19997) );
  NAND4_X1 U13935 ( .A1(n11073), .A2(n11072), .A3(n11071), .A4(n19997), .ZN(
        n11074) );
  OAI21_X1 U13936 ( .B1(n11075), .B2(n11074), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13340) );
  INV_X1 U13937 ( .A(n19215), .ZN(n11080) );
  INV_X1 U13938 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n11079) );
  MUX2_X1 U13939 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n15878), .Z(n19356) );
  AOI22_X1 U13940 ( .A1(n16315), .A2(n19356), .B1(n19262), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n11078) );
  NAND2_X1 U13941 ( .A1(n19217), .A2(BUF1_REG_30__SCAN_IN), .ZN(n11077) );
  OAI211_X1 U13942 ( .C1(n11080), .C2(n11079), .A(n11078), .B(n11077), .ZN(
        n11081) );
  AOI21_X1 U13943 ( .B1(n15627), .B2(n19263), .A(n11081), .ZN(n11082) );
  INV_X1 U13944 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11086) );
  INV_X1 U13945 ( .A(n11101), .ZN(n11084) );
  NAND2_X2 U13946 ( .A1(n11084), .A2(n15847), .ZN(n11110) );
  INV_X1 U13947 ( .A(n19200), .ZN(n19381) );
  AND2_X1 U13948 ( .A1(n10404), .A2(n19381), .ZN(n11092) );
  INV_X1 U13949 ( .A(n11092), .ZN(n11108) );
  OR2_X1 U13950 ( .A1(n10404), .A2(n19200), .ZN(n11114) );
  OAI22_X1 U13951 ( .A1(n11086), .A2(n15866), .B1(n19585), .B2(n11085), .ZN(
        n11091) );
  NAND2_X1 U13952 ( .A1(n11087), .A2(n19200), .ZN(n11113) );
  INV_X1 U13953 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11088) );
  OAI22_X1 U13954 ( .A1(n11089), .A2(n11184), .B1(n19731), .B2(n11088), .ZN(
        n11090) );
  NOR2_X1 U13955 ( .A1(n11091), .A2(n11090), .ZN(n11129) );
  INV_X1 U13956 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11095) );
  NAND2_X1 U13957 ( .A1(n11101), .A2(n11092), .ZN(n11096) );
  INV_X1 U13958 ( .A(n15847), .ZN(n13588) );
  INV_X1 U13959 ( .A(n11114), .ZN(n11093) );
  NAND2_X1 U13960 ( .A1(n11101), .A2(n11093), .ZN(n11102) );
  OAI22_X1 U13961 ( .A1(n11095), .A2(n15888), .B1(n19829), .B2(n11094), .ZN(
        n11100) );
  INV_X1 U13962 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11098) );
  OR2_X1 U13963 ( .A1(n11100), .A2(n11099), .ZN(n11107) );
  NOR2_X2 U13964 ( .A1(n11115), .A2(n11109), .ZN(n19415) );
  INV_X1 U13965 ( .A(n19415), .ZN(n11185) );
  OAI211_X1 U13967 ( .C1(n11185), .C2(n11105), .A(n11104), .B(n9748), .ZN(
        n11106) );
  NOR2_X1 U13968 ( .A1(n11107), .A2(n11106), .ZN(n11128) );
  INV_X1 U13969 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11112) );
  OR2_X2 U13970 ( .A1(n11115), .A2(n11108), .ZN(n19519) );
  INV_X1 U13971 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11111) );
  OAI22_X1 U13972 ( .A1(n11112), .A2(n19519), .B1(n19556), .B2(n11111), .ZN(
        n11119) );
  INV_X1 U13973 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11117) );
  OR2_X2 U13974 ( .A1(n11115), .A2(n11113), .ZN(n19486) );
  NOR2_X2 U13975 ( .A1(n11115), .A2(n11114), .ZN(n19460) );
  INV_X1 U13976 ( .A(n19460), .ZN(n11257) );
  OAI22_X1 U13977 ( .A1(n11117), .A2(n19486), .B1(n11257), .B2(n11116), .ZN(
        n11118) );
  NOR2_X1 U13978 ( .A1(n11119), .A2(n11118), .ZN(n11127) );
  NAND2_X1 U13979 ( .A1(n9985), .A2(n15847), .ZN(n11122) );
  NOR2_X2 U13980 ( .A1(n11122), .A2(n13602), .ZN(n11120) );
  INV_X1 U13981 ( .A(n11120), .ZN(n11171) );
  OR2_X2 U13982 ( .A1(n11122), .A2(n11087), .ZN(n19790) );
  INV_X1 U13983 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11123) );
  NOR2_X1 U13984 ( .A1(n11125), .A2(n11124), .ZN(n11126) );
  NAND4_X1 U13985 ( .A1(n11129), .A2(n11128), .A3(n11127), .A4(n11126), .ZN(
        n11131) );
  NAND2_X1 U13986 ( .A1(n11492), .A2(n19422), .ZN(n13253) );
  OR2_X1 U13987 ( .A1(n11493), .A2(n13253), .ZN(n11498) );
  NAND2_X1 U13988 ( .A1(n11498), .A2(n11500), .ZN(n11130) );
  NAND2_X1 U13989 ( .A1(n19460), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11133) );
  NAND2_X1 U13990 ( .A1(n19415), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11132) );
  OAI211_X1 U13991 ( .C1(n11171), .C2(n11134), .A(n11133), .B(n11132), .ZN(
        n11135) );
  INV_X1 U13992 ( .A(n11135), .ZN(n11160) );
  OAI22_X1 U13993 ( .A1(n11137), .A2(n11184), .B1(n19585), .B2(n11136), .ZN(
        n11141) );
  INV_X1 U13994 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11139) );
  NOR2_X1 U13995 ( .A1(n11141), .A2(n11140), .ZN(n11159) );
  OAI22_X1 U13996 ( .A1(n11143), .A2(n19699), .B1(n19829), .B2(n11142), .ZN(
        n11147) );
  INV_X1 U13997 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11145) );
  INV_X1 U13998 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11144) );
  OAI22_X1 U13999 ( .A1(n11145), .A2(n19757), .B1(n15888), .B2(n11144), .ZN(
        n11146) );
  OR2_X1 U14000 ( .A1(n11147), .A2(n11146), .ZN(n11150) );
  INV_X1 U14001 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11148) );
  NOR2_X1 U14002 ( .A1(n11150), .A2(n11149), .ZN(n11158) );
  INV_X1 U14003 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11152) );
  INV_X1 U14004 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11151) );
  OAI22_X1 U14005 ( .A1(n11152), .A2(n19556), .B1(n15866), .B2(n11151), .ZN(
        n11156) );
  INV_X1 U14006 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11154) );
  INV_X1 U14007 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11153) );
  OAI22_X1 U14008 ( .A1(n11154), .A2(n19519), .B1(n19486), .B2(n11153), .ZN(
        n11155) );
  NOR2_X1 U14009 ( .A1(n11156), .A2(n11155), .ZN(n11157) );
  NAND4_X1 U14010 ( .A1(n11160), .A2(n11159), .A3(n11158), .A4(n11157), .ZN(
        n11163) );
  NAND2_X1 U14011 ( .A1(n11161), .A2(n19422), .ZN(n11162) );
  INV_X1 U14012 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11166) );
  OAI22_X1 U14013 ( .A1(n11166), .A2(n15888), .B1(n19829), .B2(n11165), .ZN(
        n11170) );
  INV_X1 U14014 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11168) );
  OAI22_X1 U14015 ( .A1(n11168), .A2(n19757), .B1(n19699), .B2(n11167), .ZN(
        n11169) );
  OR2_X1 U14016 ( .A1(n11170), .A2(n11169), .ZN(n11174) );
  NOR2_X1 U14017 ( .A1(n11171), .A2(n11172), .ZN(n11173) );
  NOR2_X1 U14018 ( .A1(n11174), .A2(n11173), .ZN(n11196) );
  INV_X1 U14019 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11176) );
  OAI22_X1 U14020 ( .A1(n11176), .A2(n15866), .B1(n19585), .B2(n11175), .ZN(
        n11181) );
  INV_X1 U14021 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11179) );
  OAI22_X1 U14022 ( .A1(n11179), .A2(n19731), .B1(n11177), .B2(n11178), .ZN(
        n11180) );
  NOR2_X1 U14023 ( .A1(n11181), .A2(n11180), .ZN(n11195) );
  INV_X1 U14024 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11183) );
  INV_X1 U14025 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11182) );
  OAI22_X1 U14026 ( .A1(n11183), .A2(n19519), .B1(n19486), .B2(n11182), .ZN(
        n11188) );
  OAI22_X1 U14027 ( .A1(n11186), .A2(n11184), .B1(n11185), .B2(n10538), .ZN(
        n11187) );
  NOR2_X1 U14028 ( .A1(n11188), .A2(n11187), .ZN(n11194) );
  INV_X1 U14029 ( .A(n19556), .ZN(n11189) );
  NAND2_X1 U14030 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11191) );
  NAND2_X1 U14031 ( .A1(n19460), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11190) );
  OAI211_X1 U14032 ( .C1(n19790), .C2(n20948), .A(n11191), .B(n11190), .ZN(
        n11192) );
  INV_X1 U14033 ( .A(n11192), .ZN(n11193) );
  NAND4_X1 U14034 ( .A1(n11196), .A2(n11195), .A3(n11194), .A4(n11193), .ZN(
        n11198) );
  NAND2_X1 U14035 ( .A1(n11215), .A2(n19422), .ZN(n11197) );
  XNOR2_X2 U14036 ( .A(n11277), .B(n11199), .ZN(n11509) );
  NAND2_X1 U14037 ( .A1(n11509), .A2(n11322), .ZN(n11219) );
  INV_X2 U14038 ( .A(n10338), .ZN(n11394) );
  MUX2_X1 U14039 ( .A(n11410), .B(n10394), .S(n11394), .Z(n11224) );
  INV_X1 U14040 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13724) );
  INV_X1 U14041 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n11203) );
  NAND3_X1 U14042 ( .A1(n11394), .A2(n13724), .A3(n11203), .ZN(n11204) );
  NOR2_X1 U14043 ( .A1(n11431), .A2(n11394), .ZN(n11229) );
  NAND2_X1 U14044 ( .A1(n11229), .A2(n11206), .ZN(n11210) );
  AND2_X1 U14045 ( .A1(n10338), .A2(n11431), .ZN(n11230) );
  NAND2_X1 U14046 ( .A1(n11230), .A2(n11207), .ZN(n11209) );
  NAND2_X1 U14047 ( .A1(n11394), .A2(n13590), .ZN(n11208) );
  INV_X1 U14048 ( .A(n11230), .ZN(n11214) );
  NAND2_X1 U14049 ( .A1(n11229), .A2(n11490), .ZN(n11212) );
  NAND2_X1 U14050 ( .A1(n11394), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11211) );
  MUX2_X1 U14051 ( .A(n11215), .B(P2_EBX_REG_5__SCAN_IN), .S(n11394), .Z(
        n11216) );
  NAND2_X1 U14052 ( .A1(n11217), .A2(n11216), .ZN(n11218) );
  NAND2_X1 U14053 ( .A1(n11280), .A2(n11218), .ZN(n19170) );
  INV_X1 U14054 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11542) );
  INV_X1 U14055 ( .A(n11322), .ZN(n11396) );
  INV_X1 U14056 ( .A(n11238), .ZN(n11222) );
  NAND2_X1 U14057 ( .A1(n11223), .A2(n11220), .ZN(n11221) );
  NAND2_X1 U14058 ( .A1(n11222), .A2(n11221), .ZN(n13580) );
  OAI21_X1 U14059 ( .B1(n11225), .B2(n11224), .A(n11223), .ZN(n13633) );
  XNOR2_X1 U14060 ( .A(n13633), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13275) );
  INV_X1 U14061 ( .A(n11225), .ZN(n11228) );
  AND2_X1 U14062 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n11226) );
  NAND2_X1 U14063 ( .A1(n11394), .A2(n11226), .ZN(n11227) );
  NAND2_X1 U14064 ( .A1(n11228), .A2(n11227), .ZN(n13722) );
  NAND2_X1 U14065 ( .A1(n11229), .A2(n11492), .ZN(n11232) );
  NAND2_X1 U14066 ( .A1(n11230), .A2(n11411), .ZN(n11231) );
  OAI211_X1 U14067 ( .C1(n11203), .C2(n10338), .A(n11232), .B(n11231), .ZN(
        n19201) );
  NAND2_X1 U14068 ( .A1(n19201), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13395) );
  OAI21_X1 U14069 ( .B1(n13722), .B2(n19398), .A(n13395), .ZN(n11234) );
  NAND2_X1 U14070 ( .A1(n13722), .A2(n19398), .ZN(n11233) );
  AND2_X1 U14071 ( .A1(n11234), .A2(n11233), .ZN(n13274) );
  NAND2_X1 U14072 ( .A1(n13275), .A2(n13274), .ZN(n13273) );
  INV_X1 U14073 ( .A(n13633), .ZN(n11235) );
  NAND2_X1 U14074 ( .A1(n11235), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11236) );
  AND2_X1 U14075 ( .A1(n13273), .A2(n11236), .ZN(n13863) );
  INV_X1 U14076 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13873) );
  XNOR2_X1 U14077 ( .A(n11238), .B(n11237), .ZN(n19180) );
  XNOR2_X1 U14078 ( .A(n19180), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14000) );
  NAND2_X1 U14079 ( .A1(n19180), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11239) );
  NAND2_X1 U14080 ( .A1(n11240), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11241) );
  INV_X1 U14081 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11243) );
  OAI22_X1 U14082 ( .A1(n11243), .A2(n19757), .B1(n19829), .B2(n11242), .ZN(
        n11247) );
  INV_X1 U14083 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11245) );
  OAI22_X1 U14084 ( .A1(n11245), .A2(n15888), .B1(n19699), .B2(n11244), .ZN(
        n11246) );
  OR2_X1 U14085 ( .A1(n11247), .A2(n11246), .ZN(n11250) );
  NOR2_X1 U14086 ( .A1(n11171), .A2(n11248), .ZN(n11249) );
  NOR2_X1 U14087 ( .A1(n11250), .A2(n11249), .ZN(n11272) );
  INV_X1 U14088 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11252) );
  OAI22_X1 U14089 ( .A1(n11252), .A2(n19519), .B1(n11184), .B2(n11251), .ZN(
        n11256) );
  INV_X1 U14090 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11254) );
  OAI22_X1 U14091 ( .A1(n11254), .A2(n19731), .B1(n11177), .B2(n11253), .ZN(
        n11255) );
  NOR2_X1 U14092 ( .A1(n11256), .A2(n11255), .ZN(n11271) );
  OAI22_X1 U14093 ( .A1(n11259), .A2(n11257), .B1(n19556), .B2(n11258), .ZN(
        n11263) );
  INV_X1 U14094 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11261) );
  OAI22_X1 U14095 ( .A1(n11261), .A2(n19486), .B1(n19585), .B2(n11260), .ZN(
        n11262) );
  NOR2_X1 U14096 ( .A1(n11263), .A2(n11262), .ZN(n11270) );
  INV_X1 U14097 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11267) );
  INV_X1 U14098 ( .A(n15866), .ZN(n11264) );
  NAND2_X1 U14099 ( .A1(n11264), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11266) );
  NAND2_X1 U14100 ( .A1(n19415), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11265) );
  OAI211_X1 U14101 ( .C1(n19790), .C2(n11267), .A(n11266), .B(n11265), .ZN(
        n11268) );
  INV_X1 U14102 ( .A(n11268), .ZN(n11269) );
  NAND4_X1 U14103 ( .A1(n11272), .A2(n11271), .A3(n11270), .A4(n11269), .ZN(
        n11274) );
  NAND2_X1 U14104 ( .A1(n11278), .A2(n19422), .ZN(n11273) );
  MUX2_X1 U14105 ( .A(n11278), .B(P2_EBX_REG_6__SCAN_IN), .S(n11394), .Z(
        n11279) );
  AND2_X1 U14106 ( .A1(n11280), .A2(n11279), .ZN(n11281) );
  OR2_X1 U14107 ( .A1(n11281), .A2(n11288), .ZN(n19156) );
  INV_X1 U14108 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11546) );
  XNOR2_X1 U14109 ( .A(n11283), .B(n11546), .ZN(n15617) );
  NAND2_X1 U14110 ( .A1(n11283), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11284) );
  INV_X1 U14111 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n11555) );
  MUX2_X1 U14112 ( .A(n11200), .B(n11555), .S(n11394), .Z(n11286) );
  XNOR2_X1 U14113 ( .A(n11295), .B(n9850), .ZN(n19132) );
  AND2_X1 U14114 ( .A1(n11396), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11285) );
  NAND2_X1 U14115 ( .A1(n19132), .A2(n11285), .ZN(n15606) );
  INV_X1 U14116 ( .A(n11286), .ZN(n11287) );
  XNOR2_X1 U14117 ( .A(n11288), .B(n11287), .ZN(n19142) );
  NAND2_X1 U14118 ( .A1(n19142), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15805) );
  NAND2_X1 U14119 ( .A1(n15606), .A2(n15805), .ZN(n11292) );
  NAND2_X1 U14120 ( .A1(n19132), .A2(n11396), .ZN(n11289) );
  INV_X1 U14121 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16434) );
  NAND2_X1 U14122 ( .A1(n11289), .A2(n16434), .ZN(n15607) );
  INV_X1 U14123 ( .A(n19142), .ZN(n11290) );
  INV_X1 U14124 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n20950) );
  NAND2_X1 U14125 ( .A1(n11290), .A2(n20950), .ZN(n15804) );
  AND2_X1 U14126 ( .A1(n11394), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11293) );
  XNOR2_X1 U14127 ( .A(n11294), .B(n11293), .ZN(n19121) );
  NAND2_X1 U14128 ( .A1(n19121), .A2(n11396), .ZN(n11303) );
  INV_X1 U14129 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15786) );
  INV_X1 U14130 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11564) );
  OR2_X1 U14131 ( .A1(n11300), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11299) );
  NAND2_X1 U14132 ( .A1(n11300), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11296) );
  OAI21_X1 U14133 ( .B1(n11296), .B2(n10338), .A(n11375), .ZN(n11297) );
  INV_X1 U14134 ( .A(n11297), .ZN(n11298) );
  NAND2_X1 U14135 ( .A1(n11299), .A2(n11298), .ZN(n19112) );
  INV_X1 U14136 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16423) );
  OAI21_X1 U14137 ( .B1(n19112), .B2(n11322), .A(n16423), .ZN(n15592) );
  INV_X1 U14138 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13935) );
  NAND2_X1 U14139 ( .A1(n13935), .A2(n11301), .ZN(n11310) );
  AND2_X2 U14140 ( .A1(n11375), .A2(n11310), .ZN(n11309) );
  NAND3_X1 U14141 ( .A1(n11394), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n11299), 
        .ZN(n11302) );
  AND2_X1 U14142 ( .A1(n11309), .A2(n11302), .ZN(n19100) );
  AOI21_X1 U14143 ( .B1(n19100), .B2(n11396), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16350) );
  OR2_X1 U14144 ( .A1(n11303), .A2(n15786), .ZN(n15589) );
  INV_X1 U14145 ( .A(n19112), .ZN(n11305) );
  AND2_X1 U14146 ( .A1(n11396), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11304) );
  NAND2_X1 U14147 ( .A1(n11305), .A2(n11304), .ZN(n15591) );
  NAND2_X1 U14148 ( .A1(n15589), .A2(n15591), .ZN(n16348) );
  INV_X1 U14149 ( .A(n19100), .ZN(n11307) );
  NAND2_X1 U14150 ( .A1(n11396), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11306) );
  NOR2_X1 U14151 ( .A1(n11307), .A2(n11306), .ZN(n16349) );
  NOR2_X1 U14152 ( .A1(n16348), .A2(n16349), .ZN(n11308) );
  NAND3_X1 U14153 ( .A1(n11394), .A2(P2_EBX_REG_12__SCAN_IN), .A3(n11310), 
        .ZN(n11311) );
  NAND2_X1 U14154 ( .A1(n11351), .A2(n11311), .ZN(n19094) );
  INV_X1 U14155 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n20867) );
  NOR2_X1 U14156 ( .A1(n11312), .A2(n20867), .ZN(n15577) );
  NAND2_X1 U14157 ( .A1(n11312), .A2(n20867), .ZN(n15576) );
  INV_X1 U14158 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n14107) );
  INV_X1 U14159 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11585) );
  NAND2_X1 U14160 ( .A1(n14107), .A2(n11585), .ZN(n11313) );
  AND2_X1 U14161 ( .A1(n11394), .A2(n11313), .ZN(n11314) );
  OAI21_X1 U14162 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(P2_EBX_REG_16__SCAN_IN), 
        .A(n11394), .ZN(n11315) );
  INV_X1 U14163 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n15323) );
  INV_X1 U14164 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n11598) );
  NAND2_X1 U14165 ( .A1(n15323), .A2(n11598), .ZN(n11316) );
  AND2_X1 U14166 ( .A1(n11394), .A2(n11316), .ZN(n11317) );
  NOR2_X2 U14167 ( .A1(n11328), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11319) );
  INV_X1 U14168 ( .A(n11319), .ZN(n11318) );
  AND3_X1 U14169 ( .A1(n11318), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n11394), .ZN(
        n11320) );
  INV_X1 U14170 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n11610) );
  NAND2_X1 U14171 ( .A1(n11319), .A2(n11610), .ZN(n11368) );
  OR2_X1 U14172 ( .A1(n11320), .A2(n11367), .ZN(n13241) );
  INV_X1 U14173 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15730) );
  OAI21_X1 U14174 ( .B1(n13241), .B2(n11322), .A(n15730), .ZN(n14518) );
  OAI211_X1 U14175 ( .C1(n11338), .C2(P2_EBX_REG_18__SCAN_IN), .A(
        P2_EBX_REG_19__SCAN_IN), .B(n11394), .ZN(n11321) );
  NAND2_X1 U14176 ( .A1(n11321), .A2(n11328), .ZN(n19017) );
  OR2_X1 U14177 ( .A1(n19017), .A2(n11322), .ZN(n11323) );
  INV_X1 U14178 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11600) );
  NAND2_X1 U14179 ( .A1(n11323), .A2(n11600), .ZN(n14385) );
  NAND2_X1 U14180 ( .A1(n11394), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11324) );
  XNOR2_X1 U14181 ( .A(n11338), .B(n11324), .ZN(n19026) );
  NAND2_X1 U14182 ( .A1(n19026), .A2(n11396), .ZN(n11326) );
  INV_X1 U14183 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11325) );
  NAND2_X1 U14184 ( .A1(n11326), .A2(n11325), .ZN(n14392) );
  AND2_X1 U14185 ( .A1(n14385), .A2(n14392), .ZN(n15519) );
  NAND2_X1 U14186 ( .A1(n11394), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11327) );
  XNOR2_X1 U14187 ( .A(n11328), .B(n11327), .ZN(n19002) );
  NAND2_X1 U14188 ( .A1(n19002), .A2(n11396), .ZN(n11362) );
  INV_X1 U14189 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15526) );
  NAND2_X1 U14190 ( .A1(n11362), .A2(n15526), .ZN(n15521) );
  INV_X1 U14191 ( .A(n11329), .ZN(n11348) );
  AND2_X1 U14192 ( .A1(n11394), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11331) );
  INV_X1 U14193 ( .A(n11375), .ZN(n11330) );
  AOI21_X1 U14194 ( .B1(n11348), .B2(n11331), .A(n11330), .ZN(n11332) );
  NAND2_X1 U14195 ( .A1(n11333), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14388) );
  INV_X1 U14196 ( .A(n11333), .ZN(n11334) );
  INV_X1 U14197 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15554) );
  NAND2_X1 U14198 ( .A1(n11334), .A2(n15554), .ZN(n11335) );
  NAND2_X1 U14199 ( .A1(n14388), .A2(n11335), .ZN(n14467) );
  AND2_X1 U14200 ( .A1(n11394), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11336) );
  NAND2_X1 U14201 ( .A1(n11337), .A2(n11336), .ZN(n11339) );
  NAND2_X1 U14202 ( .A1(n11339), .A2(n11338), .ZN(n19041) );
  OR2_X1 U14203 ( .A1(n19041), .A2(n11322), .ZN(n11340) );
  INV_X1 U14204 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15749) );
  NAND2_X1 U14205 ( .A1(n11340), .A2(n15749), .ZN(n14445) );
  NAND2_X1 U14206 ( .A1(n11394), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11342) );
  INV_X1 U14207 ( .A(n11341), .ZN(n11343) );
  MUX2_X1 U14208 ( .A(n11342), .B(n11394), .S(n11343), .Z(n11344) );
  NAND2_X1 U14209 ( .A1(n11343), .A2(n14107), .ZN(n11347) );
  INV_X1 U14210 ( .A(n11359), .ZN(n11345) );
  INV_X1 U14211 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15759) );
  NAND2_X1 U14212 ( .A1(n11345), .A2(n15759), .ZN(n15565) );
  AND2_X1 U14213 ( .A1(n11394), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11346) );
  NAND2_X1 U14214 ( .A1(n11347), .A2(n11346), .ZN(n11349) );
  NAND2_X1 U14215 ( .A1(n11349), .A2(n11348), .ZN(n19060) );
  OR2_X1 U14216 ( .A1(n19060), .A2(n11322), .ZN(n11350) );
  INV_X1 U14217 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16329) );
  NAND2_X1 U14218 ( .A1(n11350), .A2(n16329), .ZN(n16331) );
  XNOR2_X1 U14219 ( .A(n11351), .B(n9852), .ZN(n19081) );
  NAND2_X1 U14220 ( .A1(n19081), .A2(n11396), .ZN(n11352) );
  INV_X1 U14221 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16394) );
  NAND2_X1 U14222 ( .A1(n11352), .A2(n16394), .ZN(n16342) );
  NAND4_X1 U14223 ( .A1(n14445), .A2(n15565), .A3(n16331), .A4(n16342), .ZN(
        n11353) );
  NOR2_X1 U14224 ( .A1(n14467), .A2(n11353), .ZN(n11354) );
  NAND3_X1 U14225 ( .A1(n14518), .A2(n14516), .A3(n11354), .ZN(n11365) );
  NAND2_X1 U14226 ( .A1(n11396), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11355) );
  NOR2_X1 U14227 ( .A1(n13241), .A2(n11355), .ZN(n14517) );
  NAND2_X1 U14228 ( .A1(n11396), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11356) );
  AND2_X1 U14229 ( .A1(n11396), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11357) );
  NAND2_X1 U14230 ( .A1(n19081), .A2(n11357), .ZN(n16341) );
  AND2_X1 U14231 ( .A1(n11396), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11358) );
  NAND2_X1 U14232 ( .A1(n19026), .A2(n11358), .ZN(n14391) );
  NAND2_X1 U14233 ( .A1(n11359), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15566) );
  NAND2_X1 U14234 ( .A1(n11396), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11360) );
  NAND4_X1 U14235 ( .A1(n10220), .A2(n14391), .A3(n15566), .A4(n14513), .ZN(
        n11361) );
  NOR2_X1 U14236 ( .A1(n14517), .A2(n11361), .ZN(n11364) );
  INV_X1 U14237 ( .A(n11362), .ZN(n11363) );
  NAND2_X1 U14238 ( .A1(n11363), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15522) );
  NAND2_X1 U14239 ( .A1(n11394), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11366) );
  NAND3_X1 U14240 ( .A1(n11368), .A2(n11394), .A3(P2_EBX_REG_22__SCAN_IN), 
        .ZN(n11369) );
  NAND2_X1 U14241 ( .A1(n11373), .A2(n11369), .ZN(n15955) );
  INV_X1 U14242 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15717) );
  NAND2_X1 U14243 ( .A1(n11371), .A2(n15717), .ZN(n15509) );
  NAND2_X1 U14244 ( .A1(n11394), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11374) );
  XNOR2_X1 U14245 ( .A(n11373), .B(n11374), .ZN(n16308) );
  NAND2_X1 U14246 ( .A1(n16308), .A2(n11396), .ZN(n11372) );
  XNOR2_X1 U14247 ( .A(n11372), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15504) );
  AND2_X1 U14248 ( .A1(n15509), .A2(n15504), .ZN(n11370) );
  INV_X1 U14249 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15704) );
  NAND2_X1 U14250 ( .A1(n11375), .A2(n11396), .ZN(n11399) );
  INV_X1 U14251 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15692) );
  NOR2_X1 U14252 ( .A1(n11399), .A2(n15692), .ZN(n15684) );
  NAND2_X1 U14253 ( .A1(n11399), .A2(n15692), .ZN(n15682) );
  INV_X1 U14254 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n20930) );
  NAND3_X1 U14255 ( .A1(n11394), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n16285), 
        .ZN(n11376) );
  NAND2_X1 U14256 ( .A1(n16274), .A2(n11200), .ZN(n11386) );
  XNOR2_X1 U14257 ( .A(n11386), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15482) );
  INV_X1 U14258 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n20936) );
  NAND2_X1 U14259 ( .A1(n11399), .A2(n20936), .ZN(n15489) );
  INV_X1 U14260 ( .A(n11377), .ZN(n11378) );
  NAND2_X1 U14261 ( .A1(n11394), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11379) );
  INV_X1 U14262 ( .A(n11379), .ZN(n11380) );
  NAND2_X1 U14263 ( .A1(n11380), .A2(n10223), .ZN(n11381) );
  NAND2_X1 U14264 ( .A1(n11384), .A2(n11381), .ZN(n16262) );
  INV_X1 U14265 ( .A(n14476), .ZN(n11382) );
  AND2_X1 U14266 ( .A1(n11394), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11383) );
  OR2_X2 U14267 ( .A1(n11384), .A2(n11383), .ZN(n11393) );
  NAND2_X1 U14268 ( .A1(n11384), .A2(n11383), .ZN(n11385) );
  NAND2_X1 U14269 ( .A1(n11393), .A2(n11385), .ZN(n13287) );
  NOR2_X1 U14270 ( .A1(n13287), .A2(n11322), .ZN(n14480) );
  INV_X1 U14271 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14494) );
  INV_X1 U14272 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15655) );
  NAND2_X1 U14273 ( .A1(n14494), .A2(n15655), .ZN(n14489) );
  NAND2_X1 U14274 ( .A1(n14480), .A2(n14489), .ZN(n11388) );
  INV_X1 U14275 ( .A(n11386), .ZN(n11387) );
  NOR2_X1 U14276 ( .A1(n11399), .A2(n20936), .ZN(n15488) );
  AOI21_X1 U14277 ( .B1(n11387), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15488), .ZN(n14477) );
  NAND2_X1 U14278 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15640) );
  INV_X1 U14279 ( .A(n11393), .ZN(n11391) );
  NAND2_X1 U14280 ( .A1(n11394), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11390) );
  XNOR2_X1 U14281 ( .A(n11391), .B(n11390), .ZN(n11398) );
  INV_X1 U14282 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15639) );
  OAI21_X1 U14283 ( .B1(n11398), .B2(n11322), .A(n15639), .ZN(n15464) );
  AND2_X1 U14284 ( .A1(n11394), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11392) );
  OR2_X2 U14285 ( .A1(n11393), .A2(n11392), .ZN(n16241) );
  NAND2_X1 U14286 ( .A1(n11394), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11395) );
  XNOR2_X1 U14287 ( .A(n16241), .B(n11395), .ZN(n13191) );
  AOI21_X1 U14288 ( .B1(n13191), .B2(n11396), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15454) );
  AND2_X1 U14289 ( .A1(n11396), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11397) );
  NAND2_X1 U14290 ( .A1(n13191), .A2(n11397), .ZN(n15452) );
  INV_X1 U14291 ( .A(n11398), .ZN(n16249) );
  NAND3_X1 U14292 ( .A1(n16249), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11396), .ZN(n15463) );
  INV_X1 U14293 ( .A(n11399), .ZN(n11400) );
  XOR2_X1 U14294 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11400), .Z(
        n11401) );
  XNOR2_X1 U14295 ( .A(n11402), .B(n11401), .ZN(n14458) );
  NAND2_X1 U14296 ( .A1(n11403), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11404) );
  NAND2_X1 U14297 ( .A1(n11404), .A2(n13444), .ZN(n13441) );
  OR2_X1 U14298 ( .A1(n10891), .A2(n13441), .ZN(n11405) );
  INV_X1 U14299 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n21077) );
  NAND2_X1 U14300 ( .A1(n11405), .A2(n21077), .ZN(n20088) );
  AOI21_X1 U14301 ( .B1(n11411), .B2(n11406), .A(n16473), .ZN(n11407) );
  MUX2_X1 U14302 ( .A(n20088), .B(n11407), .S(n13298), .Z(n16020) );
  INV_X1 U14303 ( .A(n11408), .ZN(n11409) );
  NAND3_X1 U14304 ( .A1(n16020), .A2(n11409), .A3(n9748), .ZN(n11419) );
  INV_X1 U14305 ( .A(n11410), .ZN(n11414) );
  NAND2_X1 U14306 ( .A1(n11412), .A2(n11411), .ZN(n11413) );
  NAND2_X1 U14307 ( .A1(n11414), .A2(n11413), .ZN(n11416) );
  NAND2_X1 U14308 ( .A1(n11416), .A2(n11415), .ZN(n20097) );
  INV_X1 U14309 ( .A(n20106), .ZN(n11417) );
  NOR2_X1 U14310 ( .A1(n11408), .A2(n11417), .ZN(n20095) );
  NAND3_X1 U14311 ( .A1(n20097), .A2(n20095), .A3(n20098), .ZN(n11418) );
  NAND2_X1 U14312 ( .A1(n11419), .A2(n11418), .ZN(n13314) );
  INV_X1 U14313 ( .A(n13314), .ZN(n11429) );
  INV_X1 U14314 ( .A(n16473), .ZN(n13186) );
  INV_X1 U14315 ( .A(n20118), .ZN(n20114) );
  INV_X1 U14316 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20958) );
  INV_X1 U14317 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20966) );
  NOR2_X1 U14318 ( .A1(n20958), .A2(n20966), .ZN(n19986) );
  NAND2_X1 U14319 ( .A1(n20958), .A2(n20966), .ZN(n19988) );
  INV_X1 U14320 ( .A(n19988), .ZN(n19975) );
  NOR3_X1 U14321 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19986), .A3(n19975), 
        .ZN(n19980) );
  INV_X1 U14322 ( .A(n19980), .ZN(n20108) );
  NOR2_X1 U14323 ( .A1(n20114), .A2(n20108), .ZN(n13310) );
  AND3_X1 U14324 ( .A1(n13186), .A2(n16502), .A3(n13310), .ZN(n11420) );
  NOR2_X1 U14325 ( .A1(n11421), .A2(n11420), .ZN(n13434) );
  MUX2_X1 U14326 ( .A(n16502), .B(n11446), .S(n19422), .Z(n11422) );
  NAND3_X1 U14327 ( .A1(n11422), .A2(n13186), .A3(n20118), .ZN(n11423) );
  AND2_X1 U14328 ( .A1(n13434), .A2(n11423), .ZN(n11428) );
  NAND2_X1 U14329 ( .A1(n16478), .A2(n9748), .ZN(n19285) );
  AOI21_X1 U14330 ( .B1(n11424), .B2(n20109), .A(n19435), .ZN(n11425) );
  NAND2_X1 U14331 ( .A1(n19285), .A2(n11425), .ZN(n11427) );
  INV_X1 U14332 ( .A(n13310), .ZN(n13433) );
  OR3_X1 U14333 ( .A1(n19285), .A2(n10317), .A3(n13433), .ZN(n11426) );
  NAND4_X1 U14334 ( .A1(n11429), .A2(n11428), .A3(n11427), .A4(n11426), .ZN(
        n11430) );
  NOR2_X1 U14335 ( .A1(n11408), .A2(n11431), .ZN(n20101) );
  NAND2_X1 U14336 ( .A1(n15349), .A2(n11432), .ZN(n11438) );
  NAND2_X1 U14337 ( .A1(n11433), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U14338 ( .A1(n10914), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n11434), .B2(P2_EAX_REG_31__SCAN_IN), .ZN(n11435) );
  NAND2_X1 U14339 ( .A1(n11436), .A2(n11435), .ZN(n11437) );
  XNOR2_X1 U14340 ( .A(n11438), .B(n11437), .ZN(n19216) );
  NAND2_X1 U14341 ( .A1(n13743), .A2(n11439), .ZN(n16472) );
  OAI21_X1 U14342 ( .B1(n10859), .B2(n19422), .A(n16472), .ZN(n11440) );
  NAND2_X1 U14343 ( .A1(n11650), .A2(n11440), .ZN(n16433) );
  NAND2_X1 U14344 ( .A1(n19365), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14453) );
  INV_X1 U14345 ( .A(n14453), .ZN(n11442) );
  AOI21_X1 U14346 ( .B1(n19216), .B2(n19391), .A(n11442), .ZN(n11489) );
  NOR2_X1 U14347 ( .A1(n20950), .A2(n16434), .ZN(n16431) );
  NAND2_X1 U14348 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16453) );
  NOR2_X1 U14349 ( .A1(n11546), .A2(n16453), .ZN(n15814) );
  NAND2_X1 U14350 ( .A1(n11650), .A2(n11443), .ZN(n14426) );
  INV_X1 U14351 ( .A(n11454), .ZN(n11444) );
  NAND2_X1 U14352 ( .A1(n11444), .A2(n19435), .ZN(n11447) );
  INV_X1 U14353 ( .A(n11445), .ZN(n14536) );
  AOI22_X1 U14354 ( .A1(n11447), .A2(n14536), .B1(n15876), .B2(n11446), .ZN(
        n11449) );
  AND3_X1 U14355 ( .A1(n11450), .A2(n11449), .A3(n11448), .ZN(n11465) );
  INV_X1 U14356 ( .A(n11451), .ZN(n11455) );
  INV_X1 U14357 ( .A(n11452), .ZN(n11453) );
  NAND3_X1 U14358 ( .A1(n11455), .A2(n11454), .A3(n11453), .ZN(n11464) );
  NAND3_X1 U14359 ( .A1(n11458), .A2(n11457), .A3(n11456), .ZN(n11459) );
  NAND2_X1 U14360 ( .A1(n11459), .A2(n9748), .ZN(n13744) );
  NAND2_X1 U14361 ( .A1(n13744), .A2(n11460), .ZN(n11462) );
  NAND2_X1 U14362 ( .A1(n11462), .A2(n11461), .ZN(n11463) );
  AND3_X1 U14363 ( .A1(n11465), .A2(n11464), .A3(n11463), .ZN(n13832) );
  INV_X1 U14364 ( .A(n11466), .ZN(n15839) );
  NAND2_X1 U14365 ( .A1(n13832), .A2(n15839), .ZN(n11467) );
  NAND2_X1 U14366 ( .A1(n11650), .A2(n11467), .ZN(n14427) );
  NAND2_X1 U14367 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13266) );
  INV_X1 U14368 ( .A(n13266), .ZN(n19397) );
  INV_X1 U14369 ( .A(n14426), .ZN(n11468) );
  NAND2_X1 U14370 ( .A1(n11497), .A2(n13266), .ZN(n13264) );
  AOI22_X1 U14371 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19397), .B1(
        n11468), .B2(n13264), .ZN(n13875) );
  NAND2_X1 U14372 ( .A1(n15814), .A2(n16454), .ZN(n16430) );
  INV_X1 U14373 ( .A(n16430), .ZN(n11469) );
  NAND2_X1 U14374 ( .A1(n16431), .A2(n11469), .ZN(n15800) );
  AND2_X1 U14375 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15758) );
  AND2_X1 U14376 ( .A1(n15758), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15760) );
  AND2_X1 U14377 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16415) );
  AND2_X1 U14378 ( .A1(n16415), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11470) );
  AND2_X1 U14379 ( .A1(n15760), .A2(n11470), .ZN(n14436) );
  NAND2_X1 U14380 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15748) );
  NAND2_X1 U14381 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14404) );
  NOR2_X1 U14382 ( .A1(n15748), .A2(n14404), .ZN(n11471) );
  NAND2_X1 U14383 ( .A1(n14436), .A2(n11471), .ZN(n14401) );
  NAND2_X1 U14384 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11472) );
  NOR2_X1 U14385 ( .A1(n14401), .A2(n11472), .ZN(n15723) );
  NAND2_X1 U14386 ( .A1(n15723), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11529) );
  NOR2_X1 U14387 ( .A1(n15800), .A2(n11529), .ZN(n15718) );
  NAND2_X1 U14388 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11528) );
  INV_X1 U14389 ( .A(n11528), .ZN(n11480) );
  NAND2_X1 U14390 ( .A1(n15718), .A2(n11480), .ZN(n15688) );
  NAND2_X1 U14391 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11484) );
  INV_X1 U14392 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11641) );
  NOR2_X1 U14393 ( .A1(n15639), .A2(n15640), .ZN(n15638) );
  INV_X1 U14394 ( .A(n15638), .ZN(n15623) );
  NOR4_X1 U14395 ( .A1(n15637), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n11641), .A4(n15623), .ZN(n11488) );
  OR2_X1 U14396 ( .A1(n14427), .A2(n19397), .ZN(n11474) );
  INV_X1 U14397 ( .A(n11650), .ZN(n11473) );
  NAND2_X1 U14398 ( .A1(n11473), .A2(n13196), .ZN(n13251) );
  AND2_X1 U14399 ( .A1(n11474), .A2(n13251), .ZN(n13265) );
  OR2_X1 U14400 ( .A1(n14427), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11475) );
  NAND2_X1 U14401 ( .A1(n13265), .A2(n11475), .ZN(n13871) );
  INV_X1 U14402 ( .A(n13871), .ZN(n11478) );
  INV_X1 U14403 ( .A(n19396), .ZN(n15815) );
  NAND4_X1 U14404 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15814), .A3(
        n16431), .A4(n13264), .ZN(n11476) );
  NAND2_X1 U14405 ( .A1(n15815), .A2(n11476), .ZN(n11477) );
  NAND2_X1 U14406 ( .A1(n11478), .A2(n11477), .ZN(n15798) );
  OR2_X1 U14407 ( .A1(n15798), .A2(n11529), .ZN(n11479) );
  NAND2_X1 U14408 ( .A1(n19396), .A2(n13251), .ZN(n16405) );
  NAND2_X1 U14409 ( .A1(n11479), .A2(n16405), .ZN(n15731) );
  OAI21_X1 U14410 ( .B1(n19396), .B2(n11480), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11481) );
  INV_X1 U14411 ( .A(n11481), .ZN(n11482) );
  AND2_X1 U14412 ( .A1(n15731), .A2(n11482), .ZN(n15687) );
  INV_X1 U14413 ( .A(n15687), .ZN(n11483) );
  NAND2_X1 U14414 ( .A1(n11483), .A2(n16405), .ZN(n15673) );
  NAND2_X1 U14415 ( .A1(n16405), .A2(n11484), .ZN(n11485) );
  NAND2_X1 U14416 ( .A1(n15673), .A2(n11485), .ZN(n15643) );
  NAND2_X1 U14417 ( .A1(n16405), .A2(n15623), .ZN(n11486) );
  NAND2_X1 U14418 ( .A1(n11486), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11487) );
  OR2_X1 U14419 ( .A1(n15643), .A2(n11487), .ZN(n15624) );
  NAND2_X1 U14420 ( .A1(n13253), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13252) );
  INV_X1 U14421 ( .A(n13252), .ZN(n11494) );
  XNOR2_X1 U14422 ( .A(n11493), .B(n11492), .ZN(n11495) );
  NAND2_X1 U14423 ( .A1(n11494), .A2(n11495), .ZN(n11496) );
  XNOR2_X1 U14424 ( .A(n13252), .B(n11495), .ZN(n13397) );
  NAND2_X1 U14425 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13397), .ZN(
        n13398) );
  NAND2_X1 U14426 ( .A1(n11496), .A2(n13398), .ZN(n11501) );
  XNOR2_X1 U14427 ( .A(n11497), .B(n11501), .ZN(n13278) );
  INV_X1 U14428 ( .A(n11498), .ZN(n11499) );
  XOR2_X1 U14429 ( .A(n11500), .B(n11499), .Z(n13277) );
  NAND2_X1 U14430 ( .A1(n13278), .A2(n13277), .ZN(n13276) );
  NAND2_X1 U14431 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11501), .ZN(
        n11502) );
  NAND2_X1 U14432 ( .A1(n13276), .A2(n11502), .ZN(n11503) );
  XNOR2_X1 U14433 ( .A(n11503), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13865) );
  NAND2_X1 U14434 ( .A1(n11503), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11504) );
  INV_X1 U14435 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20857) );
  INV_X1 U14436 ( .A(n11505), .ZN(n11507) );
  NAND2_X1 U14437 ( .A1(n11507), .A2(n11506), .ZN(n11508) );
  INV_X1 U14438 ( .A(n11509), .ZN(n11510) );
  AND2_X1 U14439 ( .A1(n11510), .A2(n11542), .ZN(n16374) );
  NAND2_X1 U14440 ( .A1(n11509), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16373) );
  INV_X1 U14441 ( .A(n11512), .ZN(n11513) );
  INV_X1 U14442 ( .A(n11515), .ZN(n11516) );
  NAND2_X1 U14443 ( .A1(n11516), .A2(n16373), .ZN(n11518) );
  NAND2_X1 U14444 ( .A1(n11518), .A2(n11517), .ZN(n11519) );
  NAND2_X1 U14445 ( .A1(n11520), .A2(n11322), .ZN(n11521) );
  NAND2_X1 U14446 ( .A1(n11525), .A2(n11521), .ZN(n11522) );
  INV_X1 U14447 ( .A(n11522), .ZN(n11523) );
  NAND2_X1 U14448 ( .A1(n11523), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11524) );
  INV_X1 U14449 ( .A(n11525), .ZN(n11526) );
  NAND2_X1 U14450 ( .A1(n11526), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11527) );
  NOR2_X1 U14451 ( .A1(n11529), .A2(n11528), .ZN(n11530) );
  OR2_X2 U14452 ( .A1(n15695), .A2(n20936), .ZN(n15493) );
  INV_X1 U14453 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15662) );
  NAND2_X1 U14454 ( .A1(n15457), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11532) );
  NAND2_X1 U14455 ( .A1(n11650), .A2(n20095), .ZN(n19406) );
  INV_X1 U14456 ( .A(n11534), .ZN(n11535) );
  AOI22_X1 U14457 ( .A1(n11644), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11540) );
  NAND2_X1 U14458 ( .A1(n11538), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11539) );
  OAI211_X1 U14459 ( .C1(n11647), .C2(n20857), .A(n11540), .B(n11539), .ZN(
        n11541) );
  INV_X1 U14460 ( .A(n11541), .ZN(n14007) );
  INV_X1 U14461 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n11545) );
  OR2_X1 U14462 ( .A1(n11647), .A2(n11542), .ZN(n11544) );
  AOI22_X1 U14463 ( .A1(n11644), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11543) );
  OAI211_X1 U14464 ( .C1(n11545), .C2(n9775), .A(n11544), .B(n11543), .ZN(
        n14506) );
  OR2_X1 U14465 ( .A1(n11647), .A2(n11546), .ZN(n11552) );
  INV_X1 U14466 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19155) );
  NAND2_X1 U14467 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11549) );
  NAND2_X1 U14468 ( .A1(n11644), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11548) );
  OAI211_X1 U14469 ( .C1(n9775), .C2(n19155), .A(n11549), .B(n11548), .ZN(
        n11550) );
  INV_X1 U14470 ( .A(n11550), .ZN(n11551) );
  OR2_X1 U14471 ( .A1(n11647), .A2(n20950), .ZN(n11554) );
  AOI22_X1 U14472 ( .A1(n11644), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11553) );
  OAI211_X1 U14473 ( .C1(n9775), .C2(n11555), .A(n11554), .B(n11553), .ZN(
        n13638) );
  OR2_X1 U14474 ( .A1(n11647), .A2(n16434), .ZN(n11561) );
  INV_X1 U14475 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n11558) );
  NAND2_X1 U14476 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11557) );
  NAND2_X1 U14477 ( .A1(n11644), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11556) );
  OAI211_X1 U14478 ( .C1(n9775), .C2(n11558), .A(n11557), .B(n11556), .ZN(
        n11559) );
  INV_X1 U14479 ( .A(n11559), .ZN(n11560) );
  OR2_X1 U14480 ( .A1(n11647), .A2(n15786), .ZN(n11567) );
  NAND2_X1 U14481 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11563) );
  NAND2_X1 U14482 ( .A1(n11644), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11562) );
  OAI211_X1 U14483 ( .C1(n9775), .C2(n11564), .A(n11563), .B(n11562), .ZN(
        n11565) );
  INV_X1 U14484 ( .A(n11565), .ZN(n11566) );
  NAND2_X1 U14485 ( .A1(n11567), .A2(n11566), .ZN(n13780) );
  INV_X1 U14486 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n11570) );
  OR2_X1 U14487 ( .A1(n11647), .A2(n16423), .ZN(n11569) );
  AOI22_X1 U14488 ( .A1(n11644), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11568) );
  OAI211_X1 U14489 ( .C1(n11570), .C2(n9775), .A(n11569), .B(n11568), .ZN(
        n13942) );
  INV_X1 U14490 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16354) );
  OR2_X1 U14491 ( .A1(n11647), .A2(n16354), .ZN(n11572) );
  AOI22_X1 U14492 ( .A1(n11644), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11571) );
  OAI211_X1 U14493 ( .C1(n13935), .C2(n9775), .A(n11572), .B(n11571), .ZN(
        n13932) );
  AOI22_X1 U14494 ( .A1(n11644), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11574) );
  NAND2_X1 U14495 ( .A1(n11538), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11573) );
  OAI211_X1 U14496 ( .C1(n11647), .C2(n20867), .A(n11574), .B(n11573), .ZN(
        n11575) );
  AOI22_X1 U14497 ( .A1(n11644), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11577) );
  NAND2_X1 U14498 ( .A1(n11538), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11576) );
  OAI211_X1 U14499 ( .C1(n11647), .C2(n16394), .A(n11577), .B(n11576), .ZN(
        n14026) );
  OR2_X1 U14500 ( .A1(n11647), .A2(n15759), .ZN(n11582) );
  NAND2_X1 U14501 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11579) );
  NAND2_X1 U14502 ( .A1(n11644), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11578) );
  OAI211_X1 U14503 ( .C1(n9775), .C2(n14107), .A(n11579), .B(n11578), .ZN(
        n11580) );
  INV_X1 U14504 ( .A(n11580), .ZN(n11581) );
  OR2_X1 U14505 ( .A1(n11647), .A2(n16329), .ZN(n11584) );
  AOI22_X1 U14506 ( .A1(n11644), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11583) );
  OAI211_X1 U14507 ( .C1(n11585), .C2(n9775), .A(n11584), .B(n11583), .ZN(
        n14156) );
  OR2_X1 U14508 ( .A1(n11647), .A2(n15554), .ZN(n11591) );
  INV_X1 U14509 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11588) );
  NAND2_X1 U14510 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11587) );
  NAND2_X1 U14511 ( .A1(n11644), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11586) );
  OAI211_X1 U14512 ( .C1(n9775), .C2(n11588), .A(n11587), .B(n11586), .ZN(
        n11589) );
  INV_X1 U14513 ( .A(n11589), .ZN(n11590) );
  NAND2_X1 U14514 ( .A1(n11591), .A2(n11590), .ZN(n14463) );
  INV_X1 U14515 ( .A(n11647), .ZN(n11640) );
  INV_X1 U14516 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n11594) );
  NAND2_X1 U14517 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11593) );
  NAND2_X1 U14518 ( .A1(n11644), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11592) );
  OAI211_X1 U14519 ( .C1(n9775), .C2(n11594), .A(n11593), .B(n11592), .ZN(
        n11595) );
  AOI21_X1 U14520 ( .B1(n11640), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11595), .ZN(n14433) );
  NAND2_X1 U14521 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11597) );
  NAND2_X1 U14522 ( .A1(n11644), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11596) );
  OAI211_X1 U14523 ( .C1(n9775), .C2(n11598), .A(n11597), .B(n11596), .ZN(
        n11599) );
  AOI21_X1 U14524 ( .B1(n11640), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n11599), .ZN(n15327) );
  OR2_X1 U14525 ( .A1(n11647), .A2(n11600), .ZN(n11602) );
  AOI22_X1 U14526 ( .A1(n11644), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11601) );
  OAI211_X1 U14527 ( .C1(n9775), .C2(n15323), .A(n11602), .B(n11601), .ZN(
        n14399) );
  INV_X1 U14528 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n11605) );
  NAND2_X1 U14529 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11604) );
  NAND2_X1 U14530 ( .A1(n11644), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11603) );
  OAI211_X1 U14531 ( .C1(n9775), .C2(n11605), .A(n11604), .B(n11603), .ZN(
        n11606) );
  AOI21_X1 U14532 ( .B1(n11640), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11606), .ZN(n15316) );
  NAND2_X1 U14533 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11609) );
  NAND2_X1 U14534 ( .A1(n11644), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11608) );
  OAI211_X1 U14535 ( .C1(n9775), .C2(n11610), .A(n11609), .B(n11608), .ZN(
        n11611) );
  AOI21_X1 U14536 ( .B1(n11640), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11611), .ZN(n13242) );
  INV_X1 U14537 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11614) );
  OR2_X1 U14538 ( .A1(n11647), .A2(n15704), .ZN(n11613) );
  AOI22_X1 U14539 ( .A1(n11644), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11612) );
  OAI211_X1 U14540 ( .C1(n9775), .C2(n11614), .A(n11613), .B(n11612), .ZN(
        n15290) );
  INV_X1 U14541 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15954) );
  OR2_X1 U14542 ( .A1(n11647), .A2(n15717), .ZN(n11616) );
  AOI22_X1 U14543 ( .A1(n11644), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11615) );
  OAI211_X1 U14544 ( .C1(n9775), .C2(n15954), .A(n11616), .B(n11615), .ZN(
        n15300) );
  AND2_X1 U14545 ( .A1(n15290), .A2(n15300), .ZN(n11617) );
  INV_X1 U14546 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n11620) );
  NAND2_X1 U14547 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11619) );
  NAND2_X1 U14548 ( .A1(n11635), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11618) );
  OAI211_X1 U14549 ( .C1(n9775), .C2(n11620), .A(n11619), .B(n11618), .ZN(
        n11621) );
  AOI21_X1 U14550 ( .B1(n11640), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11621), .ZN(n15286) );
  NAND2_X1 U14551 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11623) );
  NAND2_X1 U14552 ( .A1(n11635), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11622) );
  OAI211_X1 U14553 ( .C1(n9775), .C2(n20930), .A(n11623), .B(n11622), .ZN(
        n11624) );
  AOI21_X1 U14554 ( .B1(n11640), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n11624), .ZN(n15277) );
  INV_X1 U14555 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n11627) );
  OR2_X1 U14556 ( .A1(n11647), .A2(n15662), .ZN(n11626) );
  AOI22_X1 U14557 ( .A1(n11644), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11625) );
  OAI211_X1 U14558 ( .C1(n9775), .C2(n11627), .A(n11626), .B(n11625), .ZN(
        n15270) );
  INV_X1 U14559 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n11630) );
  OR2_X1 U14560 ( .A1(n11647), .A2(n15655), .ZN(n11629) );
  AOI22_X1 U14561 ( .A1(n11644), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11628) );
  OAI211_X1 U14562 ( .C1(n9775), .C2(n11630), .A(n11629), .B(n11628), .ZN(
        n15263) );
  INV_X1 U14563 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11633) );
  NAND2_X1 U14564 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11632) );
  NAND2_X1 U14565 ( .A1(n11635), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11631) );
  OAI211_X1 U14566 ( .C1(n9775), .C2(n11633), .A(n11632), .B(n11631), .ZN(
        n11634) );
  AOI21_X1 U14567 ( .B1(n11640), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11634), .ZN(n13289) );
  INV_X1 U14568 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n11638) );
  NAND2_X1 U14569 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11637) );
  NAND2_X1 U14570 ( .A1(n11635), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11636) );
  OAI211_X1 U14571 ( .C1(n9775), .C2(n11638), .A(n11637), .B(n11636), .ZN(
        n11639) );
  AOI21_X1 U14572 ( .B1(n11640), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11639), .ZN(n15242) );
  INV_X1 U14573 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n16239) );
  OR2_X1 U14574 ( .A1(n11647), .A2(n11641), .ZN(n11643) );
  AOI22_X1 U14575 ( .A1(n11644), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11642) );
  OAI211_X1 U14576 ( .C1(n9775), .C2(n16239), .A(n11643), .B(n11642), .ZN(
        n12656) );
  INV_X1 U14577 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13141) );
  AOI22_X1 U14578 ( .A1(n11644), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11646) );
  NAND2_X1 U14579 ( .A1(n11538), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n11645) );
  OAI211_X1 U14580 ( .C1(n11647), .C2(n13141), .A(n11646), .B(n11645), .ZN(
        n11648) );
  INV_X1 U14581 ( .A(n11648), .ZN(n11649) );
  AND2_X1 U14582 ( .A1(n11651), .A2(n11650), .ZN(n19402) );
  INV_X2 U14583 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11654) );
  NOR2_X4 U14584 ( .A1(n11654), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11664) );
  AND2_X4 U14585 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13424) );
  AOI22_X1 U14586 ( .A1(n11831), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11836), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14587 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11659) );
  AND2_X2 U14588 ( .A1(n11661), .A2(n13700), .ZN(n11695) );
  AND2_X4 U14589 ( .A1(n13700), .A2(n13681), .ZN(n12622) );
  AOI22_X1 U14590 ( .A1(n11695), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11658) );
  AND2_X4 U14591 ( .A1(n13424), .A2(n13681), .ZN(n12582) );
  AOI22_X1 U14592 ( .A1(n11888), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14593 ( .A1(n11830), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11669) );
  AOI22_X1 U14594 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U14595 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11860), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U14596 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11852), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11666) );
  NAND3_X2 U14597 ( .A1(n10236), .A2(n11669), .A3(n10232), .ZN(n13411) );
  AOI22_X1 U14598 ( .A1(n11830), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U14599 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11847), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11671) );
  AOI22_X1 U14600 ( .A1(n11831), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11670) );
  NAND4_X1 U14601 ( .A1(n11673), .A2(n11672), .A3(n11671), .A4(n11670), .ZN(
        n11679) );
  AOI22_X1 U14602 ( .A1(n11888), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11836), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U14603 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14604 ( .A1(n11695), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11675) );
  AOI22_X1 U14605 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11674) );
  NAND4_X1 U14606 ( .A1(n11677), .A2(n11676), .A3(n11675), .A4(n11674), .ZN(
        n11678) );
  AOI22_X1 U14607 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11695), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14608 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U14609 ( .A1(n11830), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11836), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U14610 ( .A1(n11888), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11680) );
  NAND4_X1 U14611 ( .A1(n11683), .A2(n11682), .A3(n11681), .A4(n11680), .ZN(
        n11689) );
  AOI22_X1 U14612 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11852), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14613 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11847), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U14614 ( .A1(n11725), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U14615 ( .A1(n11831), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11684) );
  NAND4_X1 U14616 ( .A1(n11687), .A2(n11686), .A3(n11685), .A4(n11684), .ZN(
        n11688) );
  AOI22_X1 U14617 ( .A1(n11830), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14618 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11691) );
  NAND3_X1 U14619 ( .A1(n11692), .A2(n11691), .A3(n11690), .ZN(n11693) );
  AOI22_X1 U14620 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11831), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U14621 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11695), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14622 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U14623 ( .A1(n11888), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11836), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14624 ( .A1(n11725), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U14625 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11847), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U14626 ( .A1(n11831), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11704) );
  AOI22_X1 U14627 ( .A1(n11830), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11703) );
  NAND3_X1 U14628 ( .A1(n11705), .A2(n11704), .A3(n11703), .ZN(n11706) );
  AOI22_X1 U14629 ( .A1(n11888), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11836), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14630 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U14631 ( .A1(n11695), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14632 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11708) );
  NAND2_X2 U14633 ( .A1(n11712), .A2(n10233), .ZN(n12996) );
  NAND2_X1 U14634 ( .A1(n11811), .A2(n11786), .ZN(n11778) );
  NAND2_X1 U14635 ( .A1(n11830), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11715) );
  NAND2_X1 U14636 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11714) );
  NAND2_X1 U14637 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11713) );
  NAND3_X1 U14638 ( .A1(n11715), .A2(n11714), .A3(n11713), .ZN(n11716) );
  NOR2_X1 U14639 ( .A1(n10228), .A2(n11716), .ZN(n11733) );
  NAND2_X1 U14640 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11720) );
  NAND2_X1 U14641 ( .A1(n11831), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11719) );
  NAND2_X1 U14642 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11718) );
  NAND2_X1 U14643 ( .A1(n11861), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11717) );
  NAND2_X1 U14644 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11724) );
  NAND2_X1 U14645 ( .A1(n11888), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11723) );
  NAND2_X1 U14646 ( .A1(n11836), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11722) );
  NAND2_X1 U14647 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11721) );
  NAND2_X1 U14648 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11729) );
  NAND2_X1 U14649 ( .A1(n11695), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11728) );
  NAND2_X1 U14650 ( .A1(n11725), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11727) );
  NAND2_X1 U14651 ( .A1(n12622), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11726) );
  NAND2_X1 U14652 ( .A1(n11734), .A2(n13364), .ZN(n12977) );
  NAND2_X1 U14653 ( .A1(n11830), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11738) );
  NAND2_X1 U14654 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11737) );
  NAND2_X1 U14655 ( .A1(n12621), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11736) );
  NAND2_X1 U14656 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11735) );
  NAND2_X1 U14657 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11742) );
  NAND2_X1 U14658 ( .A1(n11695), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11741) );
  NAND2_X1 U14659 ( .A1(n11725), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11740) );
  NAND2_X1 U14660 ( .A1(n12622), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11739) );
  NAND2_X1 U14661 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11746) );
  NAND2_X1 U14662 ( .A1(n11888), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11745) );
  NAND2_X1 U14663 ( .A1(n11836), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11744) );
  NAND2_X1 U14664 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11743) );
  NAND2_X1 U14665 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11750) );
  NAND2_X1 U14666 ( .A1(n11831), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11749) );
  NAND2_X1 U14667 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11748) );
  NAND2_X1 U14668 ( .A1(n11861), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11747) );
  NAND2_X4 U14669 ( .A1(n11755), .A2(n9797), .ZN(n13547) );
  NAND2_X1 U14670 ( .A1(n11830), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11760) );
  NAND2_X1 U14671 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11759) );
  NAND2_X1 U14672 ( .A1(n12621), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11758) );
  NAND2_X1 U14673 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11757) );
  NAND2_X1 U14674 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11764) );
  NAND2_X1 U14675 ( .A1(n11831), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11763) );
  NAND2_X1 U14676 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11762) );
  NAND2_X1 U14677 ( .A1(n11861), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11761) );
  NAND2_X1 U14678 ( .A1(n11888), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11767) );
  NAND2_X1 U14679 ( .A1(n11836), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11766) );
  NAND2_X1 U14680 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11765) );
  NAND3_X1 U14681 ( .A1(n11767), .A2(n11766), .A3(n11765), .ZN(n11768) );
  NAND2_X1 U14682 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11772) );
  NAND2_X1 U14683 ( .A1(n11695), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11771) );
  NAND2_X1 U14684 ( .A1(n11725), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11770) );
  NAND2_X1 U14685 ( .A1(n12622), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11769) );
  OR2_X2 U14686 ( .A1(n12977), .A2(n14540), .ZN(n13206) );
  INV_X1 U14687 ( .A(n13917), .ZN(n11784) );
  NAND3_X1 U14688 ( .A1(n11778), .A2(n11784), .A3(n14360), .ZN(n11779) );
  NAND2_X1 U14689 ( .A1(n15153), .A2(n11779), .ZN(n11782) );
  NAND2_X2 U14690 ( .A1(n11786), .A2(n12089), .ZN(n13099) );
  NAND2_X1 U14691 ( .A1(n13411), .A2(n13547), .ZN(n11785) );
  NAND2_X1 U14692 ( .A1(n13110), .A2(n11787), .ZN(n11805) );
  NOR2_X2 U14693 ( .A1(n12977), .A2(n11788), .ZN(n13361) );
  INV_X1 U14694 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n11789) );
  XNOR2_X1 U14695 ( .A(n11789), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n12975) );
  NAND2_X1 U14696 ( .A1(n13361), .A2(n12975), .ZN(n11800) );
  NAND2_X1 U14697 ( .A1(n13094), .A2(n14138), .ZN(n11790) );
  NAND2_X1 U14698 ( .A1(n12083), .A2(n11799), .ZN(n13209) );
  NAND2_X1 U14699 ( .A1(n12986), .A2(n15153), .ZN(n11792) );
  INV_X1 U14700 ( .A(n16001), .ZN(n15994) );
  NAND2_X1 U14701 ( .A1(n15994), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11817) );
  NAND2_X1 U14702 ( .A1(n20804), .A2(n9918), .ZN(n12652) );
  NAND2_X1 U14703 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11823) );
  OAI21_X1 U14704 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n11823), .ZN(n20332) );
  OR2_X1 U14705 ( .A1(n12652), .A2(n20332), .ZN(n11796) );
  AND2_X1 U14706 ( .A1(n11817), .A2(n11796), .ZN(n11797) );
  INV_X1 U14707 ( .A(n12993), .ZN(n11801) );
  NOR2_X1 U14708 ( .A1(n13094), .A2(n12089), .ZN(n11798) );
  NOR2_X1 U14709 ( .A1(n13547), .A2(n14042), .ZN(n11806) );
  AND2_X1 U14710 ( .A1(n11798), .A2(n11806), .ZN(n13416) );
  AND2_X1 U14711 ( .A1(n11799), .A2(n14360), .ZN(n12141) );
  MUX2_X1 U14712 ( .A(n12652), .B(n16001), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11803) );
  OAI21_X2 U14713 ( .B1(n11821), .B2(n11802), .A(n11803), .ZN(n11881) );
  NAND3_X1 U14714 ( .A1(n12986), .A2(n14042), .A3(n15153), .ZN(n11816) );
  NAND2_X1 U14715 ( .A1(n11804), .A2(n11806), .ZN(n13097) );
  INV_X1 U14716 ( .A(n11805), .ZN(n11815) );
  AND2_X1 U14717 ( .A1(n13923), .A2(n13917), .ZN(n11810) );
  INV_X1 U14718 ( .A(n11806), .ZN(n14038) );
  NAND2_X1 U14719 ( .A1(n14038), .A2(n13064), .ZN(n13392) );
  INV_X1 U14720 ( .A(n11807), .ZN(n11808) );
  INV_X1 U14721 ( .A(n13604), .ZN(n20841) );
  NAND2_X1 U14722 ( .A1(n11808), .A2(n20841), .ZN(n11809) );
  OAI21_X1 U14723 ( .B1(n11810), .B2(n13392), .A(n11809), .ZN(n11813) );
  INV_X1 U14724 ( .A(n13094), .ZN(n13687) );
  NAND2_X1 U14725 ( .A1(n13687), .A2(n11811), .ZN(n13105) );
  NAND2_X1 U14726 ( .A1(n11788), .A2(n14042), .ZN(n14044) );
  NAND4_X1 U14727 ( .A1(n13105), .A2(n20804), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .A4(n14044), .ZN(n11812) );
  NOR2_X1 U14728 ( .A1(n11813), .A2(n11812), .ZN(n11814) );
  NAND4_X1 U14729 ( .A1(n11816), .A2(n13097), .A3(n11815), .A4(n11814), .ZN(
        n11879) );
  NAND2_X1 U14730 ( .A1(n11881), .A2(n11879), .ZN(n11845) );
  NAND2_X1 U14731 ( .A1(n11817), .A2(n11655), .ZN(n11818) );
  INV_X1 U14732 ( .A(n11823), .ZN(n11822) );
  NAND2_X1 U14733 ( .A1(n11822), .A2(n12111), .ZN(n20594) );
  NAND2_X1 U14734 ( .A1(n11823), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11824) );
  NAND2_X1 U14735 ( .A1(n20594), .A2(n11824), .ZN(n13953) );
  INV_X1 U14736 ( .A(n12652), .ZN(n11825) );
  NAND2_X1 U14737 ( .A1(n13953), .A2(n11825), .ZN(n11827) );
  NAND2_X1 U14738 ( .A1(n15994), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11826) );
  AOI22_X1 U14739 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11835) );
  AOI22_X1 U14740 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11834) );
  AOI22_X1 U14741 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U14742 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11832) );
  NAND4_X1 U14743 ( .A1(n11835), .A2(n11834), .A3(n11833), .A4(n11832), .ZN(
        n11842) );
  INV_X1 U14744 ( .A(n11836), .ZN(n11866) );
  INV_X2 U14745 ( .A(n11866), .ZN(n12620) );
  AOI22_X1 U14746 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11840) );
  AOI22_X1 U14747 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U14748 ( .A1(n12559), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U14749 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11837) );
  NAND4_X1 U14750 ( .A1(n11840), .A2(n11839), .A3(n11838), .A4(n11837), .ZN(
        n11841) );
  INV_X1 U14751 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20912) );
  OAI22_X1 U14752 ( .A1(n12120), .A2(n20912), .B1(n11938), .B2(n11957), .ZN(
        n11843) );
  NAND2_X1 U14753 ( .A1(n20392), .A2(n11845), .ZN(n13843) );
  INV_X1 U14754 ( .A(n11937), .ZN(n11875) );
  AOI22_X1 U14755 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11851) );
  AOI22_X1 U14756 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U14757 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U14758 ( .A1(n11831), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11848) );
  NAND4_X1 U14759 ( .A1(n11851), .A2(n11850), .A3(n11849), .A4(n11848), .ZN(
        n11858) );
  AOI22_X1 U14760 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12559), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11856) );
  BUF_X1 U14761 ( .A(n11852), .Z(n11887) );
  AOI22_X1 U14762 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11855) );
  AOI22_X1 U14763 ( .A1(n12621), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11854) );
  AOI22_X1 U14764 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11853) );
  NAND4_X1 U14765 ( .A1(n11856), .A2(n11855), .A3(n11854), .A4(n11853), .ZN(
        n11857) );
  NAND2_X1 U14766 ( .A1(n11875), .A2(n11916), .ZN(n11859) );
  NAND2_X1 U14767 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11878) );
  AOI22_X1 U14768 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U14769 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U14770 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11847), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11863) );
  AOI22_X1 U14771 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11862) );
  NAND4_X1 U14772 ( .A1(n11865), .A2(n11864), .A3(n11863), .A4(n11862), .ZN(
        n11873) );
  AOI22_X1 U14773 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11871) );
  BUF_X1 U14774 ( .A(n11940), .Z(n11867) );
  AOI22_X1 U14775 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U14776 ( .A1(n12559), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U14777 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11868) );
  NAND4_X1 U14778 ( .A1(n11871), .A2(n11870), .A3(n11869), .A4(n11868), .ZN(
        n11872) );
  INV_X1 U14779 ( .A(n12047), .ZN(n11874) );
  NAND2_X1 U14780 ( .A1(n11875), .A2(n11874), .ZN(n11882) );
  INV_X1 U14781 ( .A(n11938), .ZN(n11876) );
  NAND2_X1 U14782 ( .A1(n11876), .A2(n11916), .ZN(n11877) );
  INV_X1 U14783 ( .A(n11879), .ZN(n11880) );
  NAND2_X1 U14784 ( .A1(n12159), .A2(n9918), .ZN(n11898) );
  NAND2_X1 U14785 ( .A1(n11786), .A2(n12047), .ZN(n11901) );
  INV_X1 U14786 ( .A(n11882), .ZN(n11895) );
  AOI22_X1 U14787 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U14788 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9767), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11885) );
  AOI22_X1 U14789 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11695), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U14790 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11883) );
  NAND4_X1 U14791 ( .A1(n11886), .A2(n11885), .A3(n11884), .A4(n11883), .ZN(
        n11894) );
  AOI22_X1 U14792 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U14793 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U14794 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U14795 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11889) );
  NAND4_X1 U14796 ( .A1(n11892), .A2(n11891), .A3(n11890), .A4(n11889), .ZN(
        n11893) );
  MUX2_X1 U14797 ( .A(n12044), .B(n11895), .S(n11923), .Z(n11896) );
  INV_X1 U14798 ( .A(n11896), .ZN(n11897) );
  INV_X1 U14799 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11902) );
  INV_X1 U14800 ( .A(n11899), .ZN(n12086) );
  OAI21_X1 U14801 ( .B1(n11923), .B2(n9918), .A(n12086), .ZN(n11900) );
  OAI211_X1 U14802 ( .C1(n12120), .C2(n11902), .A(n11901), .B(n11900), .ZN(
        n11920) );
  INV_X1 U14803 ( .A(n11903), .ZN(n11904) );
  INV_X1 U14804 ( .A(n11908), .ZN(n11906) );
  NAND2_X2 U14805 ( .A1(n11907), .A2(n11906), .ZN(n11955) );
  NAND2_X1 U14806 ( .A1(n11908), .A2(n11909), .ZN(n11910) );
  INV_X1 U14807 ( .A(n12080), .ZN(n12001) );
  NAND2_X1 U14808 ( .A1(n11916), .A2(n11923), .ZN(n11958) );
  XNOR2_X1 U14809 ( .A(n11958), .B(n11957), .ZN(n11912) );
  NAND2_X1 U14810 ( .A1(n11788), .A2(n13917), .ZN(n11922) );
  INV_X1 U14811 ( .A(n11922), .ZN(n11911) );
  AOI21_X1 U14812 ( .B1(n11912), .B2(n20841), .A(n11911), .ZN(n11913) );
  OAI21_X1 U14813 ( .B1(n11923), .B2(n11916), .A(n11958), .ZN(n11917) );
  INV_X1 U14814 ( .A(n12139), .ZN(n13365) );
  OAI211_X1 U14815 ( .C1(n11917), .C2(n13604), .A(n13365), .B(n12089), .ZN(
        n11918) );
  INV_X1 U14816 ( .A(n11918), .ZN(n11919) );
  OAI21_X1 U14817 ( .B1(n13604), .B2(n11923), .A(n11922), .ZN(n11924) );
  INV_X1 U14818 ( .A(n11924), .ZN(n11925) );
  OAI21_X2 U14819 ( .B1(n12157), .B2(n12001), .A(n11925), .ZN(n13613) );
  INV_X1 U14820 ( .A(n11926), .ZN(n13614) );
  NAND2_X1 U14821 ( .A1(n13614), .A2(n11927), .ZN(n11928) );
  INV_X1 U14822 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20320) );
  NAND2_X1 U14823 ( .A1(n11929), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11930) );
  INV_X1 U14824 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13789) );
  INV_X1 U14825 ( .A(n11821), .ZN(n11932) );
  NAND2_X1 U14826 ( .A1(n11932), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11936) );
  INV_X1 U14827 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20825) );
  NOR3_X1 U14828 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12111), .A3(
        n20517), .ZN(n20492) );
  NAND2_X1 U14829 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20492), .ZN(
        n20486) );
  NAND2_X1 U14830 ( .A1(n20825), .A2(n20486), .ZN(n11933) );
  NAND3_X1 U14831 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20666) );
  INV_X1 U14832 ( .A(n20666), .ZN(n20675) );
  NAND2_X1 U14833 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20675), .ZN(
        n20663) );
  NAND2_X1 U14834 ( .A1(n11933), .A2(n20663), .ZN(n20331) );
  OAI22_X1 U14835 ( .A1(n12652), .A2(n20331), .B1(n16001), .B2(n20825), .ZN(
        n11934) );
  INV_X1 U14836 ( .A(n11934), .ZN(n11935) );
  XNOR2_X2 U14837 ( .A(n11931), .B(n13901), .ZN(n20815) );
  AOI22_X1 U14838 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11944) );
  AOI22_X1 U14839 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U14840 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11942) );
  AOI22_X1 U14841 ( .A1(n12559), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11941) );
  NAND4_X1 U14842 ( .A1(n11944), .A2(n11943), .A3(n11942), .A4(n11941), .ZN(
        n11950) );
  AOI22_X1 U14843 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U14844 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11947) );
  AOI22_X1 U14845 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11946) );
  AOI22_X1 U14846 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11945) );
  NAND4_X1 U14847 ( .A1(n11948), .A2(n11947), .A3(n11946), .A4(n11945), .ZN(
        n11949) );
  AOI22_X1 U14848 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12124), .B1(
        n12132), .B2(n11975), .ZN(n11951) );
  NAND2_X1 U14849 ( .A1(n11955), .A2(n13965), .ZN(n11956) );
  NAND2_X1 U14850 ( .A1(n11958), .A2(n11957), .ZN(n11976) );
  XNOR2_X1 U14851 ( .A(n11976), .B(n11975), .ZN(n11959) );
  OAI22_X1 U14852 ( .A1(n20820), .A2(n12001), .B1(n13604), .B2(n11959), .ZN(
        n13786) );
  NAND2_X1 U14853 ( .A1(n13784), .A2(n13786), .ZN(n13785) );
  NAND2_X1 U14854 ( .A1(n11960), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11961) );
  INV_X1 U14855 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11962) );
  NAND2_X1 U14856 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11974) );
  AOI22_X1 U14857 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U14858 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11965) );
  AOI22_X1 U14859 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n9776), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11964) );
  AOI22_X1 U14860 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11963) );
  NAND4_X1 U14861 ( .A1(n11966), .A2(n11965), .A3(n11964), .A4(n11963), .ZN(
        n11972) );
  AOI22_X1 U14862 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n9777), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11970) );
  AOI22_X1 U14863 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11867), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11969) );
  AOI22_X1 U14864 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12559), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11968) );
  AOI22_X1 U14865 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11967) );
  NAND4_X1 U14866 ( .A1(n11970), .A2(n11969), .A3(n11968), .A4(n11967), .ZN(
        n11971) );
  NAND2_X1 U14867 ( .A1(n12132), .A2(n12002), .ZN(n11973) );
  NAND2_X1 U14868 ( .A1(n11974), .A2(n11973), .ZN(n11995) );
  NAND2_X1 U14869 ( .A1(n12176), .A2(n12080), .ZN(n11979) );
  NAND2_X1 U14870 ( .A1(n11976), .A2(n11975), .ZN(n12004) );
  XNOR2_X1 U14871 ( .A(n12004), .B(n12002), .ZN(n11977) );
  NAND2_X1 U14872 ( .A1(n11977), .A2(n20841), .ZN(n11978) );
  NAND2_X1 U14873 ( .A1(n11979), .A2(n11978), .ZN(n20290) );
  NAND2_X1 U14874 ( .A1(n20288), .A2(n20290), .ZN(n20289) );
  NAND2_X1 U14875 ( .A1(n11980), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11981) );
  NAND2_X1 U14876 ( .A1(n20289), .A2(n11981), .ZN(n16160) );
  INV_X1 U14877 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U14878 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11985) );
  AOI22_X1 U14879 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11984) );
  AOI22_X1 U14880 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U14881 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11982) );
  NAND4_X1 U14882 ( .A1(n11985), .A2(n11984), .A3(n11983), .A4(n11982), .ZN(
        n11991) );
  AOI22_X1 U14883 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12559), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U14884 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U14885 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11987) );
  AOI22_X1 U14886 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11986) );
  NAND4_X1 U14887 ( .A1(n11989), .A2(n11988), .A3(n11987), .A4(n11986), .ZN(
        n11990) );
  NAND2_X1 U14888 ( .A1(n12132), .A2(n12026), .ZN(n11992) );
  OAI21_X1 U14889 ( .B1(n12120), .B2(n11993), .A(n11992), .ZN(n11996) );
  INV_X1 U14890 ( .A(n11995), .ZN(n11998) );
  INV_X1 U14891 ( .A(n11996), .ZN(n11997) );
  OAI21_X1 U14892 ( .B1(n11999), .B2(n11998), .A(n11997), .ZN(n12000) );
  NAND2_X1 U14893 ( .A1(n12024), .A2(n12000), .ZN(n12184) );
  OR2_X1 U14894 ( .A1(n12184), .A2(n12001), .ZN(n12007) );
  INV_X1 U14895 ( .A(n12002), .ZN(n12003) );
  OR2_X1 U14896 ( .A1(n12004), .A2(n12003), .ZN(n12025) );
  XNOR2_X1 U14897 ( .A(n12025), .B(n12026), .ZN(n12005) );
  NAND2_X1 U14898 ( .A1(n12005), .A2(n20841), .ZN(n12006) );
  NAND2_X1 U14899 ( .A1(n12007), .A2(n12006), .ZN(n12008) );
  INV_X1 U14900 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13109) );
  XNOR2_X1 U14901 ( .A(n12008), .B(n13109), .ZN(n16159) );
  NAND2_X1 U14902 ( .A1(n16160), .A2(n16159), .ZN(n16158) );
  NAND2_X1 U14903 ( .A1(n12008), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12009) );
  NAND2_X1 U14904 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12021) );
  AOI22_X1 U14905 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U14906 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U14907 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12011) );
  AOI22_X1 U14908 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12010) );
  NAND4_X1 U14909 ( .A1(n12013), .A2(n12012), .A3(n12011), .A4(n12010), .ZN(
        n12019) );
  AOI22_X1 U14910 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U14911 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U14912 ( .A1(n12559), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U14913 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12014) );
  NAND4_X1 U14914 ( .A1(n12017), .A2(n12016), .A3(n12015), .A4(n12014), .ZN(
        n12018) );
  NAND2_X1 U14915 ( .A1(n12132), .A2(n12038), .ZN(n12020) );
  NAND2_X1 U14916 ( .A1(n12024), .A2(n12023), .ZN(n12192) );
  NAND3_X1 U14917 ( .A1(n12036), .A2(n12192), .A3(n12080), .ZN(n12030) );
  INV_X1 U14918 ( .A(n12025), .ZN(n12027) );
  NAND2_X1 U14919 ( .A1(n12027), .A2(n12026), .ZN(n12037) );
  XNOR2_X1 U14920 ( .A(n12037), .B(n12038), .ZN(n12028) );
  NAND2_X1 U14921 ( .A1(n12028), .A2(n20841), .ZN(n12029) );
  NAND2_X1 U14922 ( .A1(n12030), .A2(n12029), .ZN(n16154) );
  OR2_X1 U14923 ( .A1(n16154), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12031) );
  NAND2_X1 U14924 ( .A1(n16154), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12032) );
  INV_X1 U14925 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12034) );
  NAND2_X1 U14926 ( .A1(n12132), .A2(n12047), .ZN(n12033) );
  OAI21_X1 U14927 ( .B1(n12034), .B2(n12120), .A(n12033), .ZN(n12035) );
  NAND2_X1 U14928 ( .A1(n12240), .A2(n12080), .ZN(n12042) );
  INV_X1 U14929 ( .A(n12037), .ZN(n12039) );
  NAND2_X1 U14930 ( .A1(n12039), .A2(n12038), .ZN(n12046) );
  XNOR2_X1 U14931 ( .A(n12046), .B(n12047), .ZN(n12040) );
  NAND2_X1 U14932 ( .A1(n12040), .A2(n20841), .ZN(n12041) );
  NAND2_X1 U14933 ( .A1(n12042), .A2(n12041), .ZN(n12043) );
  NAND2_X1 U14934 ( .A1(n12043), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14243) );
  AND2_X1 U14935 ( .A1(n12044), .A2(n12080), .ZN(n12045) );
  NAND2_X4 U14936 ( .A1(n12036), .A2(n12045), .ZN(n15138) );
  INV_X1 U14937 ( .A(n12046), .ZN(n12048) );
  NAND3_X1 U14938 ( .A1(n12048), .A2(n20841), .A3(n12047), .ZN(n12049) );
  NAND2_X1 U14939 ( .A1(n14264), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12051) );
  INV_X1 U14940 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16189) );
  NAND2_X1 U14941 ( .A1(n15138), .A2(n16189), .ZN(n12053) );
  INV_X1 U14942 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16181) );
  OR2_X1 U14943 ( .A1(n15138), .A2(n16181), .ZN(n14918) );
  NAND2_X1 U14944 ( .A1(n15138), .A2(n16181), .ZN(n12054) );
  INV_X1 U14945 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15134) );
  NAND2_X1 U14946 ( .A1(n15138), .A2(n15134), .ZN(n14936) );
  NAND2_X1 U14947 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12055) );
  NAND2_X1 U14948 ( .A1(n15138), .A2(n12055), .ZN(n14934) );
  INV_X1 U14949 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14922) );
  NAND2_X1 U14950 ( .A1(n15138), .A2(n14922), .ZN(n12056) );
  OR2_X1 U14951 ( .A1(n15138), .A2(n14922), .ZN(n12057) );
  INV_X1 U14952 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12058) );
  OR2_X1 U14953 ( .A1(n15138), .A2(n12058), .ZN(n15109) );
  XNOR2_X1 U14954 ( .A(n15138), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14909) );
  NAND2_X1 U14955 ( .A1(n15138), .A2(n12058), .ZN(n15108) );
  NAND2_X1 U14956 ( .A1(n14909), .A2(n15108), .ZN(n12059) );
  OAI21_X1 U14957 ( .B1(n15089), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15085), .ZN(n12064) );
  OR2_X1 U14958 ( .A1(n15138), .A2(n15134), .ZN(n14935) );
  NOR2_X1 U14959 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12060) );
  OR2_X1 U14960 ( .A1(n15138), .A2(n12060), .ZN(n14932) );
  NOR2_X1 U14961 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12062) );
  NOR2_X1 U14962 ( .A1(n15138), .A2(n12062), .ZN(n12063) );
  OR2_X1 U14963 ( .A1(n15138), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14896) );
  NAND2_X1 U14964 ( .A1(n15138), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12065) );
  NAND2_X1 U14965 ( .A1(n14896), .A2(n12065), .ZN(n14901) );
  INV_X1 U14966 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15045) );
  NAND2_X1 U14967 ( .A1(n10221), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12066) );
  INV_X1 U14968 ( .A(n14883), .ZN(n12071) );
  INV_X1 U14969 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15059) );
  INV_X1 U14970 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12068) );
  INV_X1 U14971 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12067) );
  AND2_X1 U14972 ( .A1(n10219), .A2(n12069), .ZN(n12070) );
  AND2_X1 U14973 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14997) );
  NAND2_X1 U14974 ( .A1(n14997), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14993) );
  NAND2_X1 U14975 ( .A1(n14816), .A2(n14993), .ZN(n12072) );
  INV_X1 U14976 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14996) );
  INV_X1 U14977 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15016) );
  NAND2_X1 U14978 ( .A1(n14996), .A2(n15016), .ZN(n14817) );
  AND2_X1 U14979 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14957) );
  AND2_X1 U14980 ( .A1(n15138), .A2(n14957), .ZN(n12073) );
  INV_X1 U14981 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13133) );
  NAND2_X1 U14982 ( .A1(n14808), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12078) );
  INV_X1 U14983 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14823) );
  INV_X1 U14984 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14989) );
  NAND2_X1 U14985 ( .A1(n14823), .A2(n14989), .ZN(n14979) );
  OR2_X1 U14986 ( .A1(n15138), .A2(n14979), .ZN(n12074) );
  INV_X1 U14987 ( .A(n14807), .ZN(n12076) );
  NAND2_X1 U14988 ( .A1(n12076), .A2(n12075), .ZN(n12077) );
  NAND2_X1 U14989 ( .A1(n12078), .A2(n12077), .ZN(n12079) );
  XNOR2_X1 U14990 ( .A(n12079), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14965) );
  NAND2_X1 U14991 ( .A1(n20547), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12091) );
  OAI21_X1 U14992 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20547), .A(
        n12091), .ZN(n12081) );
  INV_X1 U14993 ( .A(n12081), .ZN(n12085) );
  NAND2_X1 U14994 ( .A1(n12132), .A2(n12085), .ZN(n12082) );
  NAND2_X1 U14995 ( .A1(n12133), .A2(n12082), .ZN(n12088) );
  NAND2_X1 U14996 ( .A1(n12083), .A2(n13547), .ZN(n12084) );
  NAND2_X1 U14997 ( .A1(n12084), .A2(n14138), .ZN(n12104) );
  OAI211_X1 U14998 ( .C1(n13099), .C2(n12086), .A(n12104), .B(n12085), .ZN(
        n12087) );
  NAND2_X1 U14999 ( .A1(n12088), .A2(n12087), .ZN(n12100) );
  NOR2_X1 U15000 ( .A1(n12089), .A2(n9918), .ZN(n12090) );
  MUX2_X1 U15001 ( .A(n20517), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12093) );
  INV_X1 U15002 ( .A(n12091), .ZN(n12092) );
  XNOR2_X1 U15003 ( .A(n12093), .B(n12092), .ZN(n12970) );
  NAND2_X1 U15004 ( .A1(n12098), .A2(n14042), .ZN(n12123) );
  OAI211_X1 U15005 ( .C1(n12100), .C2(n12098), .A(n12970), .B(n12123), .ZN(
        n12108) );
  NAND2_X1 U15006 ( .A1(n12093), .A2(n12092), .ZN(n12095) );
  NAND2_X1 U15007 ( .A1(n20517), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12094) );
  NAND2_X1 U15008 ( .A1(n12095), .A2(n12094), .ZN(n12110) );
  MUX2_X1 U15009 ( .A(n12111), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12109) );
  XNOR2_X1 U15010 ( .A(n12110), .B(n12109), .ZN(n12969) );
  INV_X1 U15011 ( .A(n12969), .ZN(n12096) );
  NAND2_X1 U15012 ( .A1(n12132), .A2(n12096), .ZN(n12105) );
  NAND2_X1 U15013 ( .A1(n12124), .A2(n12969), .ZN(n12097) );
  NAND3_X1 U15014 ( .A1(n12105), .A2(n12104), .A3(n12097), .ZN(n12103) );
  INV_X1 U15015 ( .A(n12098), .ZN(n12099) );
  NOR2_X1 U15016 ( .A1(n12970), .A2(n12099), .ZN(n12101) );
  NAND2_X1 U15017 ( .A1(n12101), .A2(n12100), .ZN(n12102) );
  NOR2_X1 U15018 ( .A1(n12105), .A2(n12104), .ZN(n12106) );
  AOI21_X1 U15019 ( .B1(n12108), .B2(n12107), .A(n12106), .ZN(n12116) );
  NAND2_X1 U15020 ( .A1(n12110), .A2(n12109), .ZN(n12113) );
  NAND2_X1 U15021 ( .A1(n12111), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12112) );
  NAND2_X1 U15022 ( .A1(n12113), .A2(n12112), .ZN(n12119) );
  XNOR2_X1 U15023 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12118) );
  XNOR2_X1 U15024 ( .A(n12119), .B(n12118), .ZN(n12971) );
  INV_X1 U15025 ( .A(n12971), .ZN(n12114) );
  NOR2_X1 U15026 ( .A1(n12124), .A2(n12114), .ZN(n12115) );
  OAI22_X1 U15027 ( .A1(n12116), .A2(n12115), .B1(n12114), .B2(n12133), .ZN(
        n12122) );
  NOR2_X1 U15028 ( .A1(n11656), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12117) );
  AOI21_X1 U15029 ( .B1(n12119), .B2(n12118), .A(n12117), .ZN(n12131) );
  INV_X1 U15030 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20326) );
  NOR2_X1 U15031 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20326), .ZN(
        n12129) );
  AND2_X1 U15032 ( .A1(n12131), .A2(n12129), .ZN(n12972) );
  NAND2_X1 U15033 ( .A1(n12120), .A2(n12972), .ZN(n12121) );
  NAND2_X1 U15034 ( .A1(n12122), .A2(n12121), .ZN(n12128) );
  INV_X1 U15035 ( .A(n12123), .ZN(n12126) );
  NAND2_X1 U15036 ( .A1(n20326), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12130) );
  AOI21_X1 U15037 ( .B1(n12131), .B2(n12130), .A(n12129), .ZN(n12135) );
  INV_X1 U15038 ( .A(n12135), .ZN(n12974) );
  AND2_X1 U15039 ( .A1(n16001), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13564) );
  INV_X1 U15040 ( .A(n13564), .ZN(n20133) );
  AOI21_X1 U15041 ( .B1(n15153), .B2(n11788), .A(n12139), .ZN(n12140) );
  OR2_X1 U15042 ( .A1(n12994), .A2(n13099), .ZN(n15985) );
  INV_X1 U15043 ( .A(n12141), .ZN(n13217) );
  INV_X2 U15044 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20839) );
  NOR2_X1 U15045 ( .A1(n13217), .A2(n20839), .ZN(n12174) );
  INV_X1 U15046 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n12143) );
  NOR2_X1 U15047 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12643) );
  INV_X1 U15048 ( .A(n12636), .ZN(n14031) );
  XNOR2_X1 U15049 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14062) );
  AOI21_X1 U15050 ( .B1(n14031), .B2(n14062), .A(n12644), .ZN(n12142) );
  OAI21_X1 U15051 ( .B1(n12638), .B2(n12143), .A(n12142), .ZN(n12144) );
  AOI21_X1 U15052 ( .B1(n12174), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12144), .ZN(n12145) );
  NAND2_X1 U15053 ( .A1(n12644), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12167) );
  NAND2_X1 U15054 ( .A1(n12146), .A2(n12167), .ZN(n13654) );
  INV_X1 U15055 ( .A(n12147), .ZN(n12150) );
  INV_X1 U15056 ( .A(n12148), .ZN(n12149) );
  NAND2_X1 U15057 ( .A1(n12150), .A2(n12149), .ZN(n12151) );
  NAND2_X1 U15058 ( .A1(n15166), .A2(n12317), .ZN(n12156) );
  INV_X1 U15059 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n12153) );
  INV_X1 U15060 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14081) );
  OAI22_X1 U15061 ( .A1(n12638), .A2(n12153), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14081), .ZN(n12154) );
  AOI21_X1 U15062 ( .B1(n12174), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12154), .ZN(n12155) );
  NAND2_X1 U15063 ( .A1(n12156), .A2(n12155), .ZN(n13558) );
  NAND2_X1 U15064 ( .A1(n15167), .A2(n11811), .ZN(n12158) );
  NAND2_X1 U15065 ( .A1(n12158), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13609) );
  INV_X1 U15066 ( .A(n12174), .ZN(n12180) );
  NAND2_X1 U15067 ( .A1(n12645), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12161) );
  NAND2_X1 U15068 ( .A1(n20839), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12160) );
  OAI211_X1 U15069 ( .C1(n12180), .C2(n11802), .A(n12161), .B(n12160), .ZN(
        n12162) );
  AOI21_X1 U15070 ( .B1(n12159), .B2(n12317), .A(n12162), .ZN(n12163) );
  OR2_X1 U15071 ( .A1(n13609), .A2(n12163), .ZN(n13610) );
  INV_X1 U15072 ( .A(n12163), .ZN(n13611) );
  OR2_X1 U15073 ( .A1(n13611), .A2(n12636), .ZN(n12164) );
  NAND2_X1 U15074 ( .A1(n13610), .A2(n12164), .ZN(n13557) );
  NAND2_X1 U15075 ( .A1(n13558), .A2(n13557), .ZN(n13653) );
  INV_X1 U15076 ( .A(n13653), .ZN(n12165) );
  NAND2_X1 U15077 ( .A1(n12166), .A2(n12165), .ZN(n13656) );
  INV_X1 U15078 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n12172) );
  INV_X1 U15079 ( .A(n12168), .ZN(n12170) );
  INV_X1 U15080 ( .A(n12177), .ZN(n12169) );
  OAI21_X1 U15081 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12170), .A(
        n12169), .ZN(n14071) );
  AOI22_X1 U15082 ( .A1(n14031), .A2(n14071), .B1(n12644), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12171) );
  OAI21_X1 U15083 ( .B1(n12638), .B2(n12172), .A(n12171), .ZN(n12173) );
  AOI21_X1 U15084 ( .B1(n12174), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12173), .ZN(n12175) );
  NAND2_X1 U15085 ( .A1(n12176), .A2(n12317), .ZN(n12183) );
  OAI21_X1 U15086 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12177), .A(
        n12185), .ZN(n20297) );
  INV_X1 U15087 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16226) );
  INV_X1 U15088 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20840) );
  OAI21_X1 U15089 ( .B1(n20840), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20839), .ZN(n12179) );
  NAND2_X1 U15090 ( .A1(n12645), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12178) );
  OAI211_X1 U15091 ( .C1(n12180), .C2(n16226), .A(n12179), .B(n12178), .ZN(
        n12181) );
  OAI21_X1 U15092 ( .B1(n12636), .B2(n20297), .A(n12181), .ZN(n12182) );
  INV_X1 U15093 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n12188) );
  OAI21_X1 U15094 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n12186), .A(
        n12194), .ZN(n20201) );
  AOI22_X1 U15095 ( .A1(n12643), .A2(n20201), .B1(n12644), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12187) );
  OAI21_X1 U15096 ( .B1(n12638), .B2(n12188), .A(n12187), .ZN(n12189) );
  INV_X1 U15097 ( .A(n12189), .ZN(n12190) );
  NAND2_X1 U15098 ( .A1(n12192), .A2(n12317), .ZN(n12201) );
  INV_X1 U15099 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n12198) );
  INV_X1 U15100 ( .A(n12202), .ZN(n12234) );
  INV_X1 U15101 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12195) );
  NAND2_X1 U15102 ( .A1(n12195), .A2(n12194), .ZN(n12196) );
  NAND2_X1 U15103 ( .A1(n12234), .A2(n12196), .ZN(n20187) );
  AOI22_X1 U15104 ( .A1(n20187), .A2(n12643), .B1(n12644), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12197) );
  OAI21_X1 U15105 ( .B1(n12638), .B2(n12198), .A(n12197), .ZN(n12199) );
  INV_X1 U15106 ( .A(n12199), .ZN(n12200) );
  XNOR2_X1 U15107 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n12245), .ZN(
        n20161) );
  INV_X1 U15108 ( .A(n20161), .ZN(n12217) );
  AOI22_X1 U15109 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15110 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U15111 ( .A1(n12559), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U15112 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12203) );
  NAND4_X1 U15113 ( .A1(n12206), .A2(n12205), .A3(n12204), .A4(n12203), .ZN(
        n12212) );
  AOI22_X1 U15114 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15115 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12209) );
  AOI22_X1 U15116 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15117 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12207) );
  NAND4_X1 U15118 ( .A1(n12210), .A2(n12209), .A3(n12208), .A4(n12207), .ZN(
        n12211) );
  NOR2_X1 U15119 ( .A1(n12212), .A2(n12211), .ZN(n12215) );
  NAND2_X1 U15120 ( .A1(n12645), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12214) );
  NAND2_X1 U15121 ( .A1(n12644), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12213) );
  OAI211_X1 U15122 ( .C1(n12338), .C2(n12215), .A(n12214), .B(n12213), .ZN(
        n12216) );
  AOI21_X1 U15123 ( .B1(n12217), .B2(n14031), .A(n12216), .ZN(n14229) );
  INV_X1 U15124 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n14192) );
  XNOR2_X1 U15125 ( .A(n12232), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14267) );
  AOI22_X1 U15126 ( .A1(n14267), .A2(n14031), .B1(n12644), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12218) );
  OAI21_X1 U15127 ( .B1(n12638), .B2(n14192), .A(n12218), .ZN(n12219) );
  INV_X1 U15128 ( .A(n12219), .ZN(n12231) );
  AOI22_X1 U15129 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12223) );
  AOI22_X1 U15130 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12559), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U15131 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U15132 ( .A1(n12621), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12220) );
  NAND4_X1 U15133 ( .A1(n12223), .A2(n12222), .A3(n12221), .A4(n12220), .ZN(
        n12229) );
  AOI22_X1 U15134 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12498), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15135 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15136 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U15137 ( .A1(n11725), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12224) );
  NAND4_X1 U15138 ( .A1(n12227), .A2(n12226), .A3(n12225), .A4(n12224), .ZN(
        n12228) );
  OAI21_X1 U15139 ( .B1(n12229), .B2(n12228), .A(n12317), .ZN(n12230) );
  AND2_X1 U15140 ( .A1(n12231), .A2(n12230), .ZN(n14108) );
  NOR2_X1 U15141 ( .A1(n14229), .A2(n14108), .ZN(n12242) );
  INV_X1 U15142 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12238) );
  INV_X1 U15143 ( .A(n12232), .ZN(n12236) );
  INV_X1 U15144 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12233) );
  NAND2_X1 U15145 ( .A1(n12234), .A2(n12233), .ZN(n12235) );
  NAND2_X1 U15146 ( .A1(n12236), .A2(n12235), .ZN(n20178) );
  AOI22_X1 U15147 ( .A1(n20178), .A2(n12643), .B1(n12644), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12237) );
  OAI21_X1 U15148 ( .B1(n12638), .B2(n12238), .A(n12237), .ZN(n12239) );
  AOI21_X1 U15149 ( .B1(n12240), .B2(n12317), .A(n12239), .ZN(n14017) );
  INV_X1 U15150 ( .A(n14017), .ZN(n12241) );
  NAND2_X1 U15151 ( .A1(n12242), .A2(n12241), .ZN(n12243) );
  INV_X1 U15152 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12244) );
  INV_X1 U15153 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16113) );
  XNOR2_X1 U15154 ( .A(n12262), .B(n16113), .ZN(n16120) );
  OR2_X1 U15155 ( .A1(n16120), .A2(n12636), .ZN(n12261) );
  AOI22_X1 U15156 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U15157 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12498), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15158 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15159 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12246) );
  NAND4_X1 U15160 ( .A1(n12249), .A2(n12248), .A3(n12247), .A4(n12246), .ZN(
        n12255) );
  AOI22_X1 U15161 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15162 ( .A1(n12621), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15163 ( .A1(n12559), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U15164 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12250) );
  NAND4_X1 U15165 ( .A1(n12253), .A2(n12252), .A3(n12251), .A4(n12250), .ZN(
        n12254) );
  NOR2_X1 U15166 ( .A1(n12255), .A2(n12254), .ZN(n12258) );
  NAND2_X1 U15167 ( .A1(n12645), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12257) );
  NAND2_X1 U15168 ( .A1(n12644), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12256) );
  OAI211_X1 U15169 ( .C1(n12338), .C2(n12258), .A(n12257), .B(n12256), .ZN(
        n12259) );
  INV_X1 U15170 ( .A(n12259), .ZN(n12260) );
  NAND2_X1 U15171 ( .A1(n12261), .A2(n12260), .ZN(n14225) );
  INV_X1 U15172 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14301) );
  OAI21_X1 U15173 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12263), .A(
        n12301), .ZN(n16149) );
  AOI22_X1 U15174 ( .A1(n14031), .A2(n16149), .B1(n12644), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12264) );
  OAI21_X1 U15175 ( .B1(n12638), .B2(n14301), .A(n12264), .ZN(n14273) );
  INV_X1 U15176 ( .A(n14273), .ZN(n12265) );
  AOI22_X1 U15177 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U15178 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U15179 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U15180 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12266) );
  NAND4_X1 U15181 ( .A1(n12269), .A2(n12268), .A3(n12267), .A4(n12266), .ZN(
        n12275) );
  AOI22_X1 U15182 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U15183 ( .A1(n12559), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15184 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12271) );
  AOI22_X1 U15185 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12270) );
  NAND4_X1 U15186 ( .A1(n12273), .A2(n12272), .A3(n12271), .A4(n12270), .ZN(
        n12274) );
  OR2_X1 U15187 ( .A1(n12275), .A2(n12274), .ZN(n12276) );
  NAND2_X1 U15188 ( .A1(n12317), .A2(n12276), .ZN(n14299) );
  INV_X1 U15189 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16095) );
  XNOR2_X1 U15190 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12307), .ZN(
        n14941) );
  AOI22_X1 U15191 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12525), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12280) );
  AOI22_X1 U15192 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12279) );
  AOI22_X1 U15193 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12278) );
  AOI22_X1 U15194 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12277) );
  NAND4_X1 U15195 ( .A1(n12280), .A2(n12279), .A3(n12278), .A4(n12277), .ZN(
        n12286) );
  AOI22_X1 U15196 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12559), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12284) );
  AOI22_X1 U15197 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12283) );
  AOI22_X1 U15198 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12282) );
  AOI22_X1 U15199 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12281) );
  NAND4_X1 U15200 ( .A1(n12284), .A2(n12283), .A3(n12282), .A4(n12281), .ZN(
        n12285) );
  OR2_X1 U15201 ( .A1(n12286), .A2(n12285), .ZN(n12287) );
  AOI22_X1 U15202 ( .A1(n12317), .A2(n12287), .B1(n12644), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12289) );
  NAND2_X1 U15203 ( .A1(n12645), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12288) );
  OAI211_X1 U15204 ( .C1(n14941), .C2(n12636), .A(n12289), .B(n12288), .ZN(
        n14277) );
  INV_X1 U15205 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14330) );
  AOI22_X1 U15206 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12559), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15207 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12525), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U15208 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n9777), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U15209 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12290) );
  NAND4_X1 U15210 ( .A1(n12293), .A2(n12292), .A3(n12291), .A4(n12290), .ZN(
        n12299) );
  AOI22_X1 U15211 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U15212 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12296) );
  AOI22_X1 U15213 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n11725), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12295) );
  AOI22_X1 U15214 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12294) );
  NAND4_X1 U15215 ( .A1(n12297), .A2(n12296), .A3(n12295), .A4(n12294), .ZN(
        n12298) );
  OR2_X1 U15216 ( .A1(n12299), .A2(n12298), .ZN(n12300) );
  NAND2_X1 U15217 ( .A1(n12317), .A2(n12300), .ZN(n12304) );
  XNOR2_X1 U15218 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12301), .ZN(
        n16140) );
  INV_X1 U15219 ( .A(n16140), .ZN(n12302) );
  AOI22_X1 U15220 ( .A1(n12644), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n14031), .B2(n12302), .ZN(n12303) );
  OAI211_X1 U15221 ( .C1(n14330), .C2(n12638), .A(n12304), .B(n12303), .ZN(
        n14319) );
  NAND2_X1 U15222 ( .A1(n14277), .A2(n14319), .ZN(n12305) );
  INV_X1 U15223 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14282) );
  XNOR2_X1 U15224 ( .A(n12324), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14255) );
  NAND2_X1 U15225 ( .A1(n14255), .A2(n12643), .ZN(n12323) );
  INV_X1 U15226 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14291) );
  INV_X1 U15227 ( .A(n12644), .ZN(n12371) );
  INV_X1 U15228 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n14926) );
  OAI22_X1 U15229 ( .A1(n12638), .A2(n14291), .B1(n12371), .B2(n14926), .ZN(
        n12308) );
  INV_X1 U15230 ( .A(n12308), .ZN(n12321) );
  AOI22_X1 U15231 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U15232 ( .A1(n12621), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U15233 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12310) );
  AOI22_X1 U15234 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12309) );
  NAND4_X1 U15235 ( .A1(n12312), .A2(n12311), .A3(n12310), .A4(n12309), .ZN(
        n12319) );
  AOI22_X1 U15236 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12498), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12316) );
  AOI22_X1 U15237 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12315) );
  AOI22_X1 U15238 ( .A1(n12559), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12314) );
  AOI22_X1 U15239 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12313) );
  NAND4_X1 U15240 ( .A1(n12316), .A2(n12315), .A3(n12314), .A4(n12313), .ZN(
        n12318) );
  OAI21_X1 U15241 ( .B1(n12319), .B2(n12318), .A(n12317), .ZN(n12320) );
  AND2_X1 U15242 ( .A1(n12321), .A2(n12320), .ZN(n12322) );
  NAND2_X1 U15243 ( .A1(n12323), .A2(n12322), .ZN(n14251) );
  XNOR2_X1 U15244 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n12342), .ZN(
        n16083) );
  INV_X1 U15245 ( .A(n16083), .ZN(n16133) );
  AOI22_X1 U15246 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12328) );
  AOI22_X1 U15247 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U15248 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12326) );
  AOI22_X1 U15249 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12325) );
  NAND4_X1 U15250 ( .A1(n12328), .A2(n12327), .A3(n12326), .A4(n12325), .ZN(
        n12334) );
  AOI22_X1 U15251 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12332) );
  AOI22_X1 U15252 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12559), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12331) );
  AOI22_X1 U15253 ( .A1(n11725), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12330) );
  AOI22_X1 U15254 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12329) );
  NAND4_X1 U15255 ( .A1(n12332), .A2(n12331), .A3(n12330), .A4(n12329), .ZN(
        n12333) );
  NOR2_X1 U15256 ( .A1(n12334), .A2(n12333), .ZN(n12337) );
  NAND2_X1 U15257 ( .A1(n12645), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12336) );
  NAND2_X1 U15258 ( .A1(n12644), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12335) );
  OAI211_X1 U15259 ( .C1(n12338), .C2(n12337), .A(n12336), .B(n12335), .ZN(
        n12339) );
  AOI21_X1 U15260 ( .B1(n16133), .B2(n14031), .A(n12339), .ZN(n14333) );
  INV_X1 U15261 ( .A(n14333), .ZN(n12340) );
  INV_X1 U15262 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12341) );
  INV_X1 U15263 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14911) );
  XNOR2_X1 U15264 ( .A(n12359), .B(n14911), .ZN(n14913) );
  NAND2_X1 U15265 ( .A1(n14913), .A2(n12643), .ZN(n12358) );
  INV_X1 U15266 ( .A(n15153), .ZN(n12343) );
  NAND2_X1 U15267 ( .A1(n12343), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12614) );
  AOI22_X1 U15268 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U15269 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11831), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U15270 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12345) );
  AOI22_X1 U15271 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12559), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12344) );
  NAND4_X1 U15272 ( .A1(n12347), .A2(n12346), .A3(n12345), .A4(n12344), .ZN(
        n12353) );
  AOI22_X1 U15273 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U15274 ( .A1(n11725), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12350) );
  AOI22_X1 U15275 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12349) );
  AOI22_X1 U15276 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12348) );
  NAND4_X1 U15277 ( .A1(n12351), .A2(n12350), .A3(n12349), .A4(n12348), .ZN(
        n12352) );
  NOR2_X1 U15278 ( .A1(n12353), .A2(n12352), .ZN(n12356) );
  AOI21_X1 U15279 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14911), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12354) );
  AOI21_X1 U15280 ( .B1(n12645), .B2(P1_EAX_REG_16__SCAN_IN), .A(n12354), .ZN(
        n12355) );
  OAI21_X1 U15281 ( .B1(n12614), .B2(n12356), .A(n12355), .ZN(n12357) );
  NAND2_X1 U15282 ( .A1(n12358), .A2(n12357), .ZN(n14342) );
  XNOR2_X1 U15283 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12375), .ZN(
        n16128) );
  INV_X1 U15284 ( .A(n12614), .ZN(n12640) );
  AOI22_X1 U15285 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12363) );
  AOI22_X1 U15286 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12498), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U15287 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12559), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U15288 ( .A1(n11831), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12360) );
  NAND4_X1 U15289 ( .A1(n12363), .A2(n12362), .A3(n12361), .A4(n12360), .ZN(
        n12369) );
  AOI22_X1 U15290 ( .A1(n12627), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12367) );
  AOI22_X1 U15291 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12366) );
  AOI22_X1 U15292 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12365) );
  AOI22_X1 U15293 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12364) );
  NAND4_X1 U15294 ( .A1(n12367), .A2(n12366), .A3(n12365), .A4(n12364), .ZN(
        n12368) );
  OR2_X1 U15295 ( .A1(n12369), .A2(n12368), .ZN(n12373) );
  INV_X1 U15296 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14797) );
  INV_X1 U15297 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12370) );
  OAI22_X1 U15298 ( .A1(n12638), .A2(n14797), .B1(n12371), .B2(n12370), .ZN(
        n12372) );
  AOI21_X1 U15299 ( .B1(n12640), .B2(n12373), .A(n12372), .ZN(n12374) );
  OAI21_X1 U15300 ( .B1(n16128), .B2(n12636), .A(n12374), .ZN(n14671) );
  INV_X1 U15301 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16076) );
  INV_X1 U15302 ( .A(n12376), .ZN(n12378) );
  INV_X1 U15303 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12377) );
  NAND2_X1 U15304 ( .A1(n12378), .A2(n12377), .ZN(n12379) );
  NAND2_X1 U15305 ( .A1(n12430), .A2(n12379), .ZN(n16065) );
  AOI22_X1 U15306 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12383) );
  AOI22_X1 U15307 ( .A1(n12621), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12382) );
  AOI22_X1 U15308 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U15309 ( .A1(n12559), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12380) );
  NAND4_X1 U15310 ( .A1(n12383), .A2(n12382), .A3(n12381), .A4(n12380), .ZN(
        n12389) );
  AOI22_X1 U15311 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12498), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12387) );
  AOI22_X1 U15312 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12386) );
  AOI22_X1 U15313 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12385) );
  AOI22_X1 U15314 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12384) );
  NAND4_X1 U15315 ( .A1(n12387), .A2(n12386), .A3(n12385), .A4(n12384), .ZN(
        n12388) );
  NOR2_X1 U15316 ( .A1(n12389), .A2(n12388), .ZN(n12392) );
  OAI21_X1 U15317 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20840), .A(
        n20839), .ZN(n12391) );
  NAND2_X1 U15318 ( .A1(n12645), .A2(P1_EAX_REG_19__SCAN_IN), .ZN(n12390) );
  OAI211_X1 U15319 ( .C1(n12614), .C2(n12392), .A(n12391), .B(n12390), .ZN(
        n12393) );
  OAI21_X1 U15320 ( .B1(n16065), .B2(n12636), .A(n12393), .ZN(n14719) );
  XNOR2_X1 U15321 ( .A(n12394), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16079) );
  NAND2_X1 U15322 ( .A1(n16079), .A2(n12643), .ZN(n12409) );
  AOI22_X1 U15323 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12398) );
  AOI22_X1 U15324 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12397) );
  AOI22_X1 U15325 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12396) );
  AOI22_X1 U15326 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12395) );
  NAND4_X1 U15327 ( .A1(n12398), .A2(n12397), .A3(n12396), .A4(n12395), .ZN(
        n12404) );
  AOI22_X1 U15328 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12402) );
  AOI22_X1 U15329 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12401) );
  AOI22_X1 U15330 ( .A1(n12559), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12400) );
  AOI22_X1 U15331 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12399) );
  NAND4_X1 U15332 ( .A1(n12402), .A2(n12401), .A3(n12400), .A4(n12399), .ZN(
        n12403) );
  NOR2_X1 U15333 ( .A1(n12404), .A2(n12403), .ZN(n12407) );
  OAI21_X1 U15334 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n16076), .A(n12636), 
        .ZN(n12405) );
  AOI21_X1 U15335 ( .B1(n12645), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12405), .ZN(
        n12406) );
  OAI21_X1 U15336 ( .B1(n12614), .B2(n12407), .A(n12406), .ZN(n12408) );
  NAND2_X1 U15337 ( .A1(n12409), .A2(n12408), .ZN(n14788) );
  NOR2_X1 U15338 ( .A1(n14719), .A2(n14788), .ZN(n12410) );
  INV_X1 U15339 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14893) );
  INV_X1 U15340 ( .A(n12411), .ZN(n12413) );
  INV_X1 U15341 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12412) );
  NAND2_X1 U15342 ( .A1(n12413), .A2(n12412), .ZN(n12414) );
  NAND2_X1 U15343 ( .A1(n12464), .A2(n12414), .ZN(n16051) );
  AOI22_X1 U15344 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12418) );
  AOI22_X1 U15345 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U15346 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12416) );
  AOI22_X1 U15347 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12415) );
  NAND4_X1 U15348 ( .A1(n12418), .A2(n12417), .A3(n12416), .A4(n12415), .ZN(
        n12424) );
  AOI22_X1 U15349 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12422) );
  AOI22_X1 U15350 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U15351 ( .A1(n12559), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12420) );
  AOI22_X1 U15352 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12419) );
  NAND4_X1 U15353 ( .A1(n12422), .A2(n12421), .A3(n12420), .A4(n12419), .ZN(
        n12423) );
  OAI21_X1 U15354 ( .B1(n12424), .B2(n12423), .A(n12640), .ZN(n12427) );
  NAND2_X1 U15355 ( .A1(n12645), .A2(P1_EAX_REG_21__SCAN_IN), .ZN(n12426) );
  NAND2_X1 U15356 ( .A1(n20839), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12425) );
  NAND4_X1 U15357 ( .A1(n12427), .A2(n12636), .A3(n12426), .A4(n12425), .ZN(
        n12428) );
  NAND2_X1 U15358 ( .A1(n12429), .A2(n12428), .ZN(n14704) );
  XNOR2_X1 U15359 ( .A(n12430), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16056) );
  NAND2_X1 U15360 ( .A1(n16056), .A2(n12643), .ZN(n12445) );
  AOI22_X1 U15361 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12434) );
  AOI22_X1 U15362 ( .A1(n12621), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12559), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12433) );
  AOI22_X1 U15363 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11725), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U15364 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12431) );
  NAND4_X1 U15365 ( .A1(n12434), .A2(n12433), .A3(n12432), .A4(n12431), .ZN(
        n12440) );
  AOI22_X1 U15366 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11867), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U15367 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12498), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U15368 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U15369 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12435) );
  NAND4_X1 U15370 ( .A1(n12438), .A2(n12437), .A3(n12436), .A4(n12435), .ZN(
        n12439) );
  OAI21_X1 U15371 ( .B1(n12440), .B2(n12439), .A(n12640), .ZN(n12443) );
  NAND2_X1 U15372 ( .A1(n12645), .A2(P1_EAX_REG_20__SCAN_IN), .ZN(n12442) );
  NAND2_X1 U15373 ( .A1(n20839), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12441) );
  NAND4_X1 U15374 ( .A1(n12443), .A2(n12636), .A3(n12442), .A4(n12441), .ZN(
        n12444) );
  NAND2_X1 U15375 ( .A1(n12445), .A2(n12444), .ZN(n14711) );
  XNOR2_X1 U15376 ( .A(n12464), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14876) );
  NAND2_X1 U15377 ( .A1(n14876), .A2(n12643), .ZN(n12462) );
  AOI22_X1 U15378 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12451) );
  AOI22_X1 U15379 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12498), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12450) );
  AOI22_X1 U15380 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12449) );
  AOI22_X1 U15381 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12448) );
  NAND4_X1 U15382 ( .A1(n12451), .A2(n12450), .A3(n12449), .A4(n12448), .ZN(
        n12457) );
  AOI22_X1 U15383 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U15384 ( .A1(n11695), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U15385 ( .A1(n12621), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U15386 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12452) );
  NAND4_X1 U15387 ( .A1(n12455), .A2(n12454), .A3(n12453), .A4(n12452), .ZN(
        n12456) );
  NOR2_X1 U15388 ( .A1(n12457), .A2(n12456), .ZN(n12460) );
  INV_X1 U15389 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14878) );
  AOI21_X1 U15390 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14878), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12458) );
  AOI21_X1 U15391 ( .B1(n12645), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12458), .ZN(
        n12459) );
  OAI21_X1 U15392 ( .B1(n12614), .B2(n12460), .A(n12459), .ZN(n12461) );
  NAND2_X1 U15393 ( .A1(n12462), .A2(n12461), .ZN(n14661) );
  INV_X1 U15394 ( .A(n12466), .ZN(n12468) );
  INV_X1 U15395 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12467) );
  NAND2_X1 U15396 ( .A1(n12468), .A2(n12467), .ZN(n12469) );
  NAND2_X1 U15397 ( .A1(n12514), .A2(n12469), .ZN(n16026) );
  AOI22_X1 U15398 ( .A1(n12621), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12473) );
  AOI22_X1 U15399 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12498), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12472) );
  AOI22_X1 U15400 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12471) );
  AOI22_X1 U15401 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12470) );
  NAND4_X1 U15402 ( .A1(n12473), .A2(n12472), .A3(n12471), .A4(n12470), .ZN(
        n12479) );
  AOI22_X1 U15403 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12477) );
  AOI22_X1 U15404 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12559), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U15405 ( .A1(n11725), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U15406 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12474) );
  NAND4_X1 U15407 ( .A1(n12477), .A2(n12476), .A3(n12475), .A4(n12474), .ZN(
        n12478) );
  NOR2_X1 U15408 ( .A1(n12479), .A2(n12478), .ZN(n12496) );
  AOI22_X1 U15409 ( .A1(n12621), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U15410 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U15411 ( .A1(n12559), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12481) );
  AOI22_X1 U15412 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12480) );
  NAND4_X1 U15413 ( .A1(n12483), .A2(n12482), .A3(n12481), .A4(n12480), .ZN(
        n12489) );
  AOI22_X1 U15414 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12487) );
  AOI22_X1 U15415 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12498), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12486) );
  AOI22_X1 U15416 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12485) );
  AOI22_X1 U15417 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12484) );
  NAND4_X1 U15418 ( .A1(n12487), .A2(n12486), .A3(n12485), .A4(n12484), .ZN(
        n12488) );
  NOR2_X1 U15419 ( .A1(n12489), .A2(n12488), .ZN(n12497) );
  XNOR2_X1 U15420 ( .A(n12496), .B(n12497), .ZN(n12493) );
  INV_X1 U15421 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14761) );
  NAND2_X1 U15422 ( .A1(n20839), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12490) );
  OAI211_X1 U15423 ( .C1(n12638), .C2(n14761), .A(n12636), .B(n12490), .ZN(
        n12491) );
  INV_X1 U15424 ( .A(n12491), .ZN(n12492) );
  OAI21_X1 U15425 ( .B1(n12614), .B2(n12493), .A(n12492), .ZN(n12494) );
  XNOR2_X1 U15426 ( .A(n12514), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14867) );
  NAND2_X1 U15427 ( .A1(n14867), .A2(n14031), .ZN(n12513) );
  NOR2_X1 U15428 ( .A1(n12497), .A2(n12496), .ZN(n12520) );
  AOI22_X1 U15429 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12502) );
  AOI22_X1 U15430 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12501) );
  AOI22_X1 U15431 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12500) );
  AOI22_X1 U15432 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12499) );
  NAND4_X1 U15433 ( .A1(n12502), .A2(n12501), .A3(n12500), .A4(n12499), .ZN(
        n12508) );
  AOI22_X1 U15434 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12506) );
  AOI22_X1 U15435 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12505) );
  AOI22_X1 U15436 ( .A1(n11695), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12504) );
  AOI22_X1 U15437 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12503) );
  NAND4_X1 U15438 ( .A1(n12506), .A2(n12505), .A3(n12504), .A4(n12503), .ZN(
        n12507) );
  OR2_X1 U15439 ( .A1(n12508), .A2(n12507), .ZN(n12519) );
  XNOR2_X1 U15440 ( .A(n12520), .B(n12519), .ZN(n12511) );
  NAND2_X1 U15441 ( .A1(n12645), .A2(P1_EAX_REG_24__SCAN_IN), .ZN(n12510) );
  OAI21_X1 U15442 ( .B1(n20840), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n20839), .ZN(n12509) );
  OAI211_X1 U15443 ( .C1(n12511), .C2(n12614), .A(n12510), .B(n12509), .ZN(
        n12512) );
  NAND2_X1 U15444 ( .A1(n12513), .A2(n12512), .ZN(n14645) );
  INV_X1 U15445 ( .A(n12514), .ZN(n12515) );
  INV_X1 U15446 ( .A(n12516), .ZN(n12517) );
  INV_X1 U15447 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14634) );
  NAND2_X1 U15448 ( .A1(n12517), .A2(n14634), .ZN(n12518) );
  NAND2_X1 U15449 ( .A1(n12555), .A2(n12518), .ZN(n14856) );
  NAND2_X1 U15450 ( .A1(n12520), .A2(n12519), .ZN(n12538) );
  AOI22_X1 U15451 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11695), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12524) );
  AOI22_X1 U15452 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12523) );
  AOI22_X1 U15453 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12522) );
  AOI22_X1 U15454 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12521) );
  NAND4_X1 U15455 ( .A1(n12524), .A2(n12523), .A3(n12522), .A4(n12521), .ZN(
        n12531) );
  AOI22_X1 U15456 ( .A1(n12621), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12529) );
  AOI22_X1 U15457 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12498), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12528) );
  AOI22_X1 U15458 ( .A1(n11725), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12527) );
  AOI22_X1 U15459 ( .A1(n12525), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12526) );
  NAND4_X1 U15460 ( .A1(n12529), .A2(n12528), .A3(n12527), .A4(n12526), .ZN(
        n12530) );
  NOR2_X1 U15461 ( .A1(n12531), .A2(n12530), .ZN(n12539) );
  XNOR2_X1 U15462 ( .A(n12538), .B(n12539), .ZN(n12534) );
  OAI21_X1 U15463 ( .B1(n20840), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n20839), .ZN(n12533) );
  NAND2_X1 U15464 ( .A1(n12645), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n12532) );
  OAI211_X1 U15465 ( .C1(n12534), .C2(n12614), .A(n12533), .B(n12532), .ZN(
        n12535) );
  NAND2_X1 U15466 ( .A1(n12536), .A2(n12535), .ZN(n14628) );
  XNOR2_X1 U15467 ( .A(n12555), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14849) );
  NOR2_X1 U15468 ( .A1(n12539), .A2(n12538), .ZN(n12571) );
  AOI22_X1 U15469 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12543) );
  AOI22_X1 U15470 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12542) );
  AOI22_X1 U15471 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12541) );
  AOI22_X1 U15472 ( .A1(n11831), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12540) );
  NAND4_X1 U15473 ( .A1(n12543), .A2(n12542), .A3(n12541), .A4(n12540), .ZN(
        n12549) );
  AOI22_X1 U15474 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12547) );
  AOI22_X1 U15475 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12546) );
  AOI22_X1 U15476 ( .A1(n12559), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12545) );
  AOI22_X1 U15477 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12544) );
  NAND4_X1 U15478 ( .A1(n12547), .A2(n12546), .A3(n12545), .A4(n12544), .ZN(
        n12548) );
  OR2_X1 U15479 ( .A1(n12549), .A2(n12548), .ZN(n12570) );
  INV_X1 U15480 ( .A(n12570), .ZN(n12550) );
  XNOR2_X1 U15481 ( .A(n12571), .B(n12550), .ZN(n12553) );
  INV_X1 U15482 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14749) );
  NAND2_X1 U15483 ( .A1(n20839), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12551) );
  OAI211_X1 U15484 ( .C1(n12638), .C2(n14749), .A(n12636), .B(n12551), .ZN(
        n12552) );
  AOI21_X1 U15485 ( .B1(n12553), .B2(n12640), .A(n12552), .ZN(n12554) );
  AOI21_X1 U15486 ( .B1(n14849), .B2(n12643), .A(n12554), .ZN(n14615) );
  INV_X1 U15487 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14845) );
  INV_X1 U15488 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12556) );
  NAND2_X1 U15489 ( .A1(n12557), .A2(n12556), .ZN(n12558) );
  NAND2_X1 U15490 ( .A1(n12596), .A2(n12558), .ZN(n14838) );
  AOI22_X1 U15491 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12563) );
  AOI22_X1 U15492 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12559), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12562) );
  AOI22_X1 U15493 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12561) );
  AOI22_X1 U15494 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12560) );
  NAND4_X1 U15495 ( .A1(n12563), .A2(n12562), .A3(n12561), .A4(n12560), .ZN(
        n12569) );
  AOI22_X1 U15496 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11852), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12567) );
  AOI22_X1 U15497 ( .A1(n12621), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12566) );
  AOI22_X1 U15498 ( .A1(n11831), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12565) );
  AOI22_X1 U15499 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11940), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12564) );
  NAND4_X1 U15500 ( .A1(n12567), .A2(n12566), .A3(n12565), .A4(n12564), .ZN(
        n12568) );
  NOR2_X1 U15501 ( .A1(n12569), .A2(n12568), .ZN(n12577) );
  NAND2_X1 U15502 ( .A1(n12571), .A2(n12570), .ZN(n12576) );
  XNOR2_X1 U15503 ( .A(n12577), .B(n12576), .ZN(n12572) );
  NOR2_X1 U15504 ( .A1(n12572), .A2(n12614), .ZN(n12575) );
  INV_X1 U15505 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14744) );
  NAND2_X1 U15506 ( .A1(n20839), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12573) );
  OAI211_X1 U15507 ( .C1(n12638), .C2(n14744), .A(n12636), .B(n12573), .ZN(
        n12574) );
  OAI22_X1 U15508 ( .A1(n14838), .A2(n12636), .B1(n12575), .B2(n12574), .ZN(
        n14604) );
  XNOR2_X1 U15509 ( .A(n12596), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14825) );
  NAND2_X1 U15510 ( .A1(n14825), .A2(n14031), .ZN(n12594) );
  NOR2_X1 U15511 ( .A1(n12577), .A2(n12576), .ZN(n12611) );
  AOI22_X1 U15512 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12581) );
  AOI22_X1 U15513 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12580) );
  AOI22_X1 U15514 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12579) );
  AOI22_X1 U15515 ( .A1(n11831), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12578) );
  NAND4_X1 U15516 ( .A1(n12581), .A2(n12580), .A3(n12579), .A4(n12578), .ZN(
        n12588) );
  AOI22_X1 U15517 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12586) );
  AOI22_X1 U15518 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U15519 ( .A1(n12559), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12584) );
  AOI22_X1 U15520 ( .A1(n11852), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12583) );
  NAND4_X1 U15521 ( .A1(n12586), .A2(n12585), .A3(n12584), .A4(n12583), .ZN(
        n12587) );
  OR2_X1 U15522 ( .A1(n12588), .A2(n12587), .ZN(n12610) );
  XNOR2_X1 U15523 ( .A(n12611), .B(n12610), .ZN(n12592) );
  INV_X1 U15524 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14739) );
  NAND2_X1 U15525 ( .A1(n20839), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12589) );
  OAI211_X1 U15526 ( .C1(n12638), .C2(n14739), .A(n12636), .B(n12589), .ZN(
        n12590) );
  INV_X1 U15527 ( .A(n12590), .ZN(n12591) );
  OAI21_X1 U15528 ( .B1(n12592), .B2(n12614), .A(n12591), .ZN(n12593) );
  NAND2_X1 U15529 ( .A1(n12594), .A2(n12593), .ZN(n14591) );
  INV_X1 U15530 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14827) );
  NAND2_X1 U15531 ( .A1(n12597), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12648) );
  INV_X1 U15532 ( .A(n12597), .ZN(n12598) );
  INV_X1 U15533 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n21132) );
  NAND2_X1 U15534 ( .A1(n12598), .A2(n21132), .ZN(n12599) );
  NAND2_X1 U15535 ( .A1(n12648), .A2(n12599), .ZN(n14582) );
  AOI22_X1 U15536 ( .A1(n11831), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12621), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12603) );
  AOI22_X1 U15537 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12602) );
  AOI22_X1 U15538 ( .A1(n12559), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12601) );
  AOI22_X1 U15539 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12600) );
  NAND4_X1 U15540 ( .A1(n12603), .A2(n12602), .A3(n12601), .A4(n12600), .ZN(
        n12609) );
  AOI22_X1 U15541 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11852), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12607) );
  AOI22_X1 U15542 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12498), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12606) );
  AOI22_X1 U15543 ( .A1(n11867), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12605) );
  AOI22_X1 U15544 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12604) );
  NAND4_X1 U15545 ( .A1(n12607), .A2(n12606), .A3(n12605), .A4(n12604), .ZN(
        n12608) );
  NOR2_X1 U15546 ( .A1(n12609), .A2(n12608), .ZN(n12619) );
  NAND2_X1 U15547 ( .A1(n12611), .A2(n12610), .ZN(n12618) );
  XNOR2_X1 U15548 ( .A(n12619), .B(n12618), .ZN(n12615) );
  OAI21_X1 U15549 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n21132), .A(n12636), 
        .ZN(n12612) );
  AOI21_X1 U15550 ( .B1(n12645), .B2(P1_EAX_REG_29__SCAN_IN), .A(n12612), .ZN(
        n12613) );
  OAI21_X1 U15551 ( .B1(n12615), .B2(n12614), .A(n12613), .ZN(n12616) );
  NAND2_X1 U15552 ( .A1(n12617), .A2(n12616), .ZN(n14419) );
  XNOR2_X1 U15553 ( .A(n12648), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14812) );
  NOR2_X1 U15554 ( .A1(n12619), .A2(n12618), .ZN(n12635) );
  AOI22_X1 U15555 ( .A1(n12621), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12620), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12626) );
  AOI22_X1 U15556 ( .A1(n12559), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12622), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12625) );
  AOI22_X1 U15557 ( .A1(n11831), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12624) );
  AOI22_X1 U15558 ( .A1(n9777), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12582), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12623) );
  NAND4_X1 U15559 ( .A1(n12626), .A2(n12625), .A3(n12624), .A4(n12623), .ZN(
        n12633) );
  AOI22_X1 U15560 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11852), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U15561 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12498), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12630) );
  AOI22_X1 U15562 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12627), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12629) );
  AOI22_X1 U15563 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12628) );
  NAND4_X1 U15564 ( .A1(n12631), .A2(n12630), .A3(n12629), .A4(n12628), .ZN(
        n12632) );
  NOR2_X1 U15565 ( .A1(n12633), .A2(n12632), .ZN(n12634) );
  XNOR2_X1 U15566 ( .A(n12635), .B(n12634), .ZN(n12641) );
  INV_X1 U15567 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14731) );
  NAND2_X1 U15568 ( .A1(n20839), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12637) );
  OAI211_X1 U15569 ( .C1(n12638), .C2(n14731), .A(n12637), .B(n12636), .ZN(
        n12639) );
  AOI21_X1 U15570 ( .B1(n12641), .B2(n12640), .A(n12639), .ZN(n12642) );
  AOI21_X1 U15571 ( .B1(n14812), .B2(n12643), .A(n12642), .ZN(n14568) );
  AOI22_X1 U15572 ( .A1(n12645), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12644), .ZN(n12646) );
  INV_X1 U15573 ( .A(n12646), .ZN(n12647) );
  NAND2_X1 U15574 ( .A1(n9918), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16231) );
  NAND2_X1 U15575 ( .A1(n20839), .A2(n20526), .ZN(n20667) );
  NAND2_X1 U15576 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20809), .ZN(n13730) );
  INV_X1 U15577 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n21154) );
  INV_X1 U15578 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14559) );
  NAND2_X1 U15579 ( .A1(n12652), .A2(n20667), .ZN(n20845) );
  NAND2_X1 U15580 ( .A1(n20845), .A2(n9918), .ZN(n12650) );
  NAND2_X1 U15581 ( .A1(n9918), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15995) );
  NAND2_X1 U15582 ( .A1(n20840), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12651) );
  AND2_X1 U15583 ( .A1(n15995), .A2(n12651), .ZN(n13617) );
  INV_X2 U15584 ( .A(n20207), .ZN(n20299) );
  NAND2_X1 U15585 ( .A1(n20299), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14956) );
  NAND2_X1 U15586 ( .A1(n20287), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12653) );
  OAI211_X1 U15587 ( .C1(n14037), .C2(n20298), .A(n14956), .B(n12653), .ZN(
        n12654) );
  NOR2_X1 U15588 ( .A1(n16478), .A2(n16472), .ZN(n13436) );
  INV_X2 U15589 ( .A(n15319), .ZN(n15344) );
  NAND2_X1 U15590 ( .A1(n12655), .A2(n15341), .ZN(n12660) );
  NAND2_X1 U15591 ( .A1(n15344), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12657) );
  NAND2_X1 U15592 ( .A1(n12660), .A2(n12659), .ZN(P2_U2857) );
  AOI22_X1 U15593 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17277), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12677) );
  NOR2_X2 U15594 ( .A1(n12662), .A2(n18758), .ZN(n12749) );
  AOI22_X1 U15595 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17279), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12676) );
  NOR2_X1 U15596 ( .A1(n18758), .A2(n12666), .ZN(n12700) );
  INV_X1 U15597 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n21109) );
  NOR2_X1 U15598 ( .A1(n12662), .A2(n12667), .ZN(n12663) );
  AOI22_X1 U15599 ( .A1(n17303), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17305), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12664) );
  OAI21_X1 U15600 ( .B1(n21109), .B2(n10227), .A(n12664), .ZN(n12674) );
  INV_X1 U15601 ( .A(n17119), .ZN(n17262) );
  AOI22_X1 U15602 ( .A1(n9749), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12672) );
  INV_X4 U15603 ( .A(n13525), .ZN(n17247) );
  AOI22_X1 U15604 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12671) );
  NOR2_X2 U15605 ( .A1(n12667), .A2(n12666), .ZN(n13466) );
  AOI22_X1 U15606 ( .A1(n17267), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12670) );
  NOR2_X2 U15607 ( .A1(n18778), .A2(n12668), .ZN(n12838) );
  AOI22_X1 U15608 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n9758), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12669) );
  NAND4_X1 U15609 ( .A1(n12672), .A2(n12671), .A3(n12670), .A4(n12669), .ZN(
        n12673) );
  AOI211_X1 U15610 ( .C1(n9754), .C2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n12674), .B(n12673), .ZN(n12675) );
  NAND3_X1 U15611 ( .A1(n12677), .A2(n12676), .A3(n12675), .ZN(n16552) );
  AOI22_X1 U15612 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12687) );
  AOI22_X1 U15613 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12686) );
  INV_X1 U15614 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18337) );
  AOI22_X1 U15615 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12678) );
  OAI21_X1 U15616 ( .B1(n17019), .B2(n18337), .A(n12678), .ZN(n12684) );
  INV_X2 U15617 ( .A(n17233), .ZN(n17305) );
  AOI22_X1 U15618 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17305), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12682) );
  INV_X2 U15619 ( .A(n10227), .ZN(n17219) );
  AOI22_X1 U15620 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12681) );
  AOI22_X1 U15621 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12680) );
  AOI22_X1 U15622 ( .A1(n17248), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12679) );
  NAND4_X1 U15623 ( .A1(n12682), .A2(n12681), .A3(n12680), .A4(n12679), .ZN(
        n12683) );
  AOI211_X1 U15624 ( .C1(n17295), .C2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n12684), .B(n12683), .ZN(n12685) );
  NAND3_X1 U15625 ( .A1(n12687), .A2(n12686), .A3(n12685), .ZN(n12921) );
  AOI22_X1 U15626 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12699) );
  AOI22_X1 U15627 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12698) );
  INV_X1 U15628 ( .A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n20957) );
  AOI22_X1 U15629 ( .A1(n17303), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13466), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12689) );
  OAI21_X1 U15630 ( .B1(n12661), .B2(n20957), .A(n12689), .ZN(n12696) );
  AOI22_X1 U15631 ( .A1(n12833), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12690), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12694) );
  AOI22_X1 U15632 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13526), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12693) );
  AOI22_X1 U15633 ( .A1(n15901), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12692) );
  AOI22_X1 U15634 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12838), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12691) );
  NAND4_X1 U15635 ( .A1(n12694), .A2(n12693), .A3(n12692), .A4(n12691), .ZN(
        n12695) );
  AOI211_X1 U15636 ( .C1(n17295), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n12696), .B(n12695), .ZN(n12697) );
  NAND3_X1 U15637 ( .A1(n12699), .A2(n12698), .A3(n12697), .ZN(n12920) );
  AOI22_X1 U15638 ( .A1(n12749), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12700), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12703) );
  AOI22_X1 U15639 ( .A1(n12690), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13526), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12702) );
  AOI22_X1 U15640 ( .A1(n12838), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12704) );
  OAI21_X1 U15641 ( .B1(n12705), .B2(n20935), .A(n12704), .ZN(n12706) );
  INV_X1 U15642 ( .A(n12706), .ZN(n12713) );
  AOI22_X1 U15643 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9749), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12712) );
  AOI22_X1 U15644 ( .A1(n12750), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12707), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12711) );
  AOI22_X1 U15645 ( .A1(n12833), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13466), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12710) );
  AOI22_X1 U15646 ( .A1(n12688), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12708), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12709) );
  AOI22_X1 U15647 ( .A1(n12833), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12717) );
  AOI22_X1 U15648 ( .A1(n12749), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13466), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12716) );
  AOI22_X1 U15649 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12838), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12715) );
  AOI22_X1 U15650 ( .A1(n15901), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12714) );
  NAND4_X1 U15651 ( .A1(n12717), .A2(n12716), .A3(n12715), .A4(n12714), .ZN(
        n12723) );
  AOI22_X1 U15652 ( .A1(n12750), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12690), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U15653 ( .A1(n12688), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12720) );
  AOI22_X1 U15654 ( .A1(n12707), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12719) );
  AOI22_X1 U15655 ( .A1(n12700), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13526), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12718) );
  NAND4_X1 U15656 ( .A1(n12721), .A2(n12720), .A3(n12719), .A4(n12718), .ZN(
        n12722) );
  NAND2_X1 U15657 ( .A1(n17491), .A2(n12759), .ZN(n12763) );
  AOI22_X1 U15658 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17279), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12727) );
  AOI22_X1 U15659 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12726) );
  AOI22_X1 U15660 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17248), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12725) );
  AOI22_X1 U15661 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12724) );
  NAND4_X1 U15662 ( .A1(n12727), .A2(n12726), .A3(n12725), .A4(n12724), .ZN(
        n12733) );
  INV_X2 U15663 ( .A(n10227), .ZN(n17294) );
  AOI22_X1 U15664 ( .A1(n15901), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17294), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12731) );
  AOI22_X1 U15665 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12730) );
  AOI22_X1 U15666 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U15667 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12728) );
  NAND4_X1 U15668 ( .A1(n12731), .A2(n12730), .A3(n12729), .A4(n12728), .ZN(
        n12732) );
  INV_X1 U15669 ( .A(n17479), .ZN(n12932) );
  NAND2_X1 U15670 ( .A1(n12768), .A2(n12932), .ZN(n12744) );
  AOI22_X1 U15671 ( .A1(n15901), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12737) );
  AOI22_X1 U15672 ( .A1(n17303), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17294), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12736) );
  AOI22_X1 U15673 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12735) );
  AOI22_X1 U15674 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12734) );
  NAND4_X1 U15675 ( .A1(n12737), .A2(n12736), .A3(n12735), .A4(n12734), .ZN(
        n12743) );
  AOI22_X1 U15676 ( .A1(n9749), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U15677 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9754), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12740) );
  AOI22_X1 U15678 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12739) );
  AOI22_X1 U15679 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12738) );
  NAND4_X1 U15680 ( .A1(n12741), .A2(n12740), .A3(n12739), .A4(n12738), .ZN(
        n12742) );
  INV_X1 U15681 ( .A(n17472), .ZN(n12939) );
  NAND2_X1 U15682 ( .A1(n12771), .A2(n12939), .ZN(n12773) );
  NOR2_X4 U15683 ( .A1(n17468), .A2(n12773), .ZN(n17872) );
  INV_X1 U15684 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18097) );
  INV_X1 U15685 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18231) );
  XNOR2_X1 U15686 ( .A(n12744), .B(n12921), .ZN(n17907) );
  NAND2_X1 U15687 ( .A1(n12757), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12758) );
  AOI22_X1 U15688 ( .A1(n15901), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17294), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12747) );
  AOI22_X1 U15689 ( .A1(n12688), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12746) );
  INV_X1 U15690 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18312) );
  AOI22_X1 U15691 ( .A1(n12707), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12748) );
  OAI21_X1 U15692 ( .B1(n17019), .B2(n18312), .A(n12748), .ZN(n12756) );
  AOI22_X1 U15693 ( .A1(n12750), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12749), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12754) );
  AOI22_X1 U15694 ( .A1(n12838), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12753) );
  AOI22_X1 U15695 ( .A1(n13526), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13466), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12752) );
  AOI22_X1 U15696 ( .A1(n12833), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12751) );
  NAND4_X1 U15697 ( .A1(n12754), .A2(n12753), .A3(n12752), .A4(n12751), .ZN(
        n12755) );
  INV_X1 U15698 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18925) );
  NOR2_X1 U15699 ( .A1(n17960), .A2(n18925), .ZN(n17959) );
  NAND2_X1 U15700 ( .A1(n17959), .A2(n17951), .ZN(n17950) );
  NAND2_X1 U15701 ( .A1(n12758), .A2(n17950), .ZN(n17943) );
  XNOR2_X1 U15702 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12760), .ZN(
        n17944) );
  NAND2_X1 U15703 ( .A1(n17943), .A2(n17944), .ZN(n17942) );
  INV_X1 U15704 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18261) );
  XOR2_X1 U15705 ( .A(n12763), .B(n12762), .Z(n12766) );
  INV_X1 U15706 ( .A(n12766), .ZN(n12764) );
  NAND2_X1 U15707 ( .A1(n12766), .A2(n12765), .ZN(n12767) );
  NAND2_X1 U15708 ( .A1(n17927), .A2(n12767), .ZN(n17916) );
  INV_X1 U15709 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18243) );
  XNOR2_X1 U15710 ( .A(n12768), .B(n17479), .ZN(n12769) );
  XNOR2_X1 U15711 ( .A(n18243), .B(n12769), .ZN(n17917) );
  NAND2_X1 U15712 ( .A1(n17916), .A2(n17917), .ZN(n17915) );
  NAND2_X1 U15713 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12769), .ZN(
        n12770) );
  NAND2_X1 U15714 ( .A1(n17915), .A2(n12770), .ZN(n17906) );
  INV_X1 U15715 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18219) );
  XNOR2_X1 U15716 ( .A(n12771), .B(n17472), .ZN(n12772) );
  XNOR2_X1 U15717 ( .A(n18219), .B(n12772), .ZN(n17893) );
  NAND2_X1 U15718 ( .A1(n12776), .A2(n12775), .ZN(n12777) );
  INV_X1 U15719 ( .A(n12778), .ZN(n12782) );
  INV_X1 U15720 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n20868) );
  NAND2_X1 U15721 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18166) );
  INV_X1 U15722 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18169) );
  NOR2_X1 U15723 ( .A1(n18166), .A2(n18169), .ZN(n18151) );
  NAND2_X1 U15724 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18151), .ZN(
        n17784) );
  NOR2_X1 U15725 ( .A1(n20868), .A2(n17784), .ZN(n17771) );
  NAND2_X1 U15726 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17771), .ZN(
        n12953) );
  INV_X1 U15727 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18118) );
  NOR2_X1 U15728 ( .A1(n12953), .A2(n18118), .ZN(n16508) );
  INV_X1 U15729 ( .A(n12784), .ZN(n17694) );
  INV_X1 U15730 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18148) );
  INV_X1 U15731 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21139) );
  NAND4_X1 U15732 ( .A1(n18148), .A2(n20868), .A3(n21139), .A4(n18118), .ZN(
        n12783) );
  NAND3_X1 U15733 ( .A1(n18169), .A2(n12780), .A3(n12779), .ZN(n12781) );
  NOR2_X1 U15734 ( .A1(n17872), .A2(n17770), .ZN(n17804) );
  OAI221_X1 U15735 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17802), 
        .C1(n18097), .C2(n17694), .A(n17759), .ZN(n17748) );
  NOR2_X1 U15736 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17748), .ZN(
        n17747) );
  INV_X1 U15737 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18084) );
  NOR2_X1 U15738 ( .A1(n18097), .A2(n18084), .ZN(n18072) );
  INV_X1 U15739 ( .A(n18072), .ZN(n17744) );
  INV_X1 U15740 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21148) );
  NAND2_X1 U15741 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18049) );
  NOR2_X1 U15742 ( .A1(n21148), .A2(n18049), .ZN(n16560) );
  NAND2_X1 U15743 ( .A1(n16560), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17984) );
  INV_X1 U15744 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21092) );
  NAND2_X1 U15745 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18072), .ZN(
        n18029) );
  NOR2_X1 U15746 ( .A1(n18029), .A2(n17984), .ZN(n17682) );
  NAND2_X1 U15747 ( .A1(n17682), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17997) );
  NAND2_X1 U15748 ( .A1(n17802), .A2(n21092), .ZN(n17736) );
  NOR2_X1 U15749 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17736), .ZN(
        n12785) );
  INV_X1 U15750 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n20926) );
  NAND2_X1 U15751 ( .A1(n12785), .A2(n20926), .ZN(n17702) );
  NOR2_X1 U15752 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17702), .ZN(
        n17695) );
  INV_X1 U15753 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18043) );
  INV_X1 U15754 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n20898) );
  NAND3_X1 U15755 ( .A1(n17695), .A2(n18043), .A3(n20898), .ZN(n12786) );
  OAI21_X1 U15756 ( .B1(n12784), .B2(n17997), .A(n12786), .ZN(n12787) );
  INV_X1 U15757 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18014) );
  NAND2_X1 U15758 ( .A1(n17659), .A2(n18014), .ZN(n17658) );
  NAND2_X1 U15759 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17654), .ZN(
        n12791) );
  INV_X1 U15760 ( .A(n12791), .ZN(n12790) );
  INV_X1 U15761 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17995) );
  NAND2_X1 U15762 ( .A1(n17802), .A2(n17658), .ZN(n17653) );
  OAI21_X1 U15763 ( .B1(n12790), .B2(n12789), .A(n17653), .ZN(n17636) );
  NOR2_X1 U15764 ( .A1(n17636), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17635) );
  INV_X1 U15765 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17985) );
  OAI22_X1 U15766 ( .A1(n17872), .A2(n17635), .B1(n12791), .B2(n17985), .ZN(
        n12792) );
  INV_X1 U15767 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17606) );
  NOR2_X1 U15768 ( .A1(n17872), .A2(n12793), .ZN(n12795) );
  NAND2_X1 U15769 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16522) );
  INV_X1 U15770 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16536) );
  NOR2_X1 U15771 ( .A1(n16522), .A2(n16536), .ZN(n16539) );
  INV_X1 U15772 ( .A(n16539), .ZN(n16011) );
  INV_X1 U15773 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16012) );
  NOR2_X1 U15774 ( .A1(n16009), .A2(n16012), .ZN(n16008) );
  NOR2_X1 U15775 ( .A1(n12795), .A2(n16008), .ZN(n12799) );
  INV_X1 U15776 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18923) );
  AOI22_X1 U15777 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17802), .B1(
        n17872), .B2(n18923), .ZN(n12798) );
  NOR2_X1 U15778 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18923), .ZN(
        n16545) );
  NOR2_X1 U15779 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16012), .ZN(
        n16538) );
  OAI21_X1 U15780 ( .B1(n16545), .B2(n12796), .A(n12798), .ZN(n12797) );
  INV_X1 U15781 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18801) );
  INV_X1 U15782 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18798) );
  OAI22_X1 U15783 ( .A1(n18933), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18798), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12807) );
  NOR2_X1 U15784 ( .A1(n18940), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12913) );
  NOR2_X1 U15785 ( .A1(n21189), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12800) );
  OR2_X1 U15786 ( .A1(n12807), .A2(n12806), .ZN(n12801) );
  OAI21_X1 U15787 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18933), .A(
        n12801), .ZN(n12802) );
  OAI22_X1 U15788 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18801), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12802), .ZN(n12809) );
  NOR2_X1 U15789 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18801), .ZN(
        n12803) );
  NAND2_X1 U15790 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12802), .ZN(
        n12808) );
  AOI22_X1 U15791 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12809), .B1(
        n12803), .B2(n12808), .ZN(n12812) );
  AOI21_X1 U15792 ( .B1(n18940), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n12913), .ZN(n12917) );
  INV_X1 U15793 ( .A(n12917), .ZN(n12804) );
  NOR2_X1 U15794 ( .A1(n12914), .A2(n12804), .ZN(n12811) );
  OAI21_X1 U15795 ( .B1(n12807), .B2(n12806), .A(n12812), .ZN(n12805) );
  AOI21_X1 U15796 ( .B1(n12807), .B2(n12806), .A(n12805), .ZN(n12918) );
  INV_X1 U15797 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18754) );
  AND2_X1 U15798 ( .A1(n12808), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12810) );
  OAI22_X1 U15799 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18754), .B1(
        n12810), .B2(n12809), .ZN(n12915) );
  AOI211_X1 U15800 ( .C1(n12812), .C2(n12811), .A(n12918), .B(n12915), .ZN(
        n18745) );
  AOI22_X1 U15801 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12816) );
  AOI22_X1 U15802 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17277), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12815) );
  AOI22_X1 U15803 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12814) );
  AOI22_X1 U15804 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12813) );
  NAND4_X1 U15805 ( .A1(n12816), .A2(n12815), .A3(n12814), .A4(n12813), .ZN(
        n12822) );
  AOI22_X1 U15806 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12820) );
  AOI22_X1 U15807 ( .A1(n15901), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12819) );
  AOI22_X1 U15808 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12818) );
  AOI22_X1 U15809 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17248), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12817) );
  NAND4_X1 U15810 ( .A1(n12820), .A2(n12819), .A3(n12818), .A4(n12817), .ZN(
        n12821) );
  AOI22_X1 U15811 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12826) );
  AOI22_X1 U15812 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12825) );
  AOI22_X1 U15813 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12824) );
  AOI22_X1 U15814 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12823) );
  NAND4_X1 U15815 ( .A1(n12826), .A2(n12825), .A3(n12824), .A4(n12823), .ZN(
        n12832) );
  AOI22_X1 U15816 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12830) );
  AOI22_X1 U15817 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12829) );
  AOI22_X1 U15818 ( .A1(n17303), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12828) );
  AOI22_X1 U15819 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17305), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12827) );
  NAND4_X1 U15820 ( .A1(n12830), .A2(n12829), .A3(n12828), .A4(n12827), .ZN(
        n12831) );
  AOI22_X1 U15821 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17277), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12837) );
  AOI22_X1 U15822 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12836) );
  AOI22_X1 U15823 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9754), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12835) );
  AOI22_X1 U15824 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12834) );
  NAND4_X1 U15825 ( .A1(n12837), .A2(n12836), .A3(n12835), .A4(n12834), .ZN(
        n12844) );
  CLKBUF_X3 U15826 ( .A(n12838), .Z(n17304) );
  AOI22_X1 U15827 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12842) );
  AOI22_X1 U15828 ( .A1(n15901), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12841) );
  AOI22_X1 U15829 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12840) );
  AOI22_X1 U15830 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12839) );
  NAND4_X1 U15831 ( .A1(n12842), .A2(n12841), .A3(n12840), .A4(n12839), .ZN(
        n12843) );
  AOI22_X1 U15832 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17267), .ZN(n12848) );
  AOI22_X1 U15833 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17284), .ZN(n12847) );
  AOI22_X1 U15834 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n9758), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12846) );
  AOI22_X1 U15835 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17277), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12845) );
  AOI22_X1 U15836 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17301), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12852) );
  AOI22_X1 U15837 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12851) );
  AOI22_X1 U15838 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17278), .B1(
        n17305), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12850) );
  AOI22_X1 U15839 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17219), .B1(
        n9754), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12849) );
  NOR2_X1 U15840 ( .A1(n18323), .A2(n18348), .ZN(n12898) );
  AOI22_X1 U15841 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12856) );
  AOI22_X1 U15842 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17294), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12855) );
  AOI22_X1 U15843 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12854) );
  AOI22_X1 U15844 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12853) );
  NAND4_X1 U15845 ( .A1(n12856), .A2(n12855), .A3(n12854), .A4(n12853), .ZN(
        n12862) );
  AOI22_X1 U15846 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12860) );
  AOI22_X1 U15847 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12859) );
  AOI22_X1 U15848 ( .A1(n17303), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12858) );
  AOI22_X1 U15849 ( .A1(n15901), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12857) );
  NAND4_X1 U15850 ( .A1(n12860), .A2(n12859), .A3(n12858), .A4(n12857), .ZN(
        n12861) );
  AOI22_X1 U15851 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12872) );
  AOI22_X1 U15852 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12871) );
  INV_X1 U15853 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18321) );
  AOI22_X1 U15854 ( .A1(n15901), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17294), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12863) );
  OAI21_X1 U15855 ( .B1(n17119), .B2(n18321), .A(n12863), .ZN(n12869) );
  AOI22_X1 U15856 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17295), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12867) );
  AOI22_X1 U15857 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12866) );
  AOI22_X1 U15858 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12865) );
  AOI22_X1 U15859 ( .A1(n17303), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12864) );
  NAND4_X1 U15860 ( .A1(n12867), .A2(n12866), .A3(n12865), .A4(n12864), .ZN(
        n12868) );
  AOI211_X1 U15861 ( .C1(n9754), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n12869), .B(n12868), .ZN(n12870) );
  NAND3_X1 U15862 ( .A1(n12872), .A2(n12871), .A3(n12870), .ZN(n15929) );
  NOR2_X1 U15863 ( .A1(n18334), .A2(n15929), .ZN(n15932) );
  AOI22_X1 U15864 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9754), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12876) );
  AOI22_X1 U15865 ( .A1(n17303), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12875) );
  AOI22_X1 U15866 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12874) );
  AOI22_X1 U15867 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12873) );
  NAND4_X1 U15868 ( .A1(n12876), .A2(n12875), .A3(n12874), .A4(n12873), .ZN(
        n12882) );
  AOI22_X1 U15869 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12880) );
  AOI22_X1 U15870 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12879) );
  AOI22_X1 U15871 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12878) );
  AOI22_X1 U15872 ( .A1(n15901), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12877) );
  NAND4_X1 U15873 ( .A1(n12880), .A2(n12879), .A3(n12878), .A4(n12877), .ZN(
        n12881) );
  AOI22_X1 U15874 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17294), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U15875 ( .A1(n15901), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12889) );
  AOI22_X1 U15876 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12883) );
  OAI21_X1 U15877 ( .B1(n12661), .B2(n20962), .A(n12883), .ZN(n12888) );
  AOI22_X1 U15878 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17248), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12887) );
  AOI22_X1 U15879 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12886) );
  AOI22_X1 U15880 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12885) );
  AOI22_X1 U15881 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12884) );
  NOR2_X1 U15882 ( .A1(n18328), .A2(n17349), .ZN(n18761) );
  NAND3_X1 U15883 ( .A1(n12898), .A2(n15932), .A3(n18761), .ZN(n15923) );
  NAND2_X1 U15884 ( .A1(n18318), .A2(n18323), .ZN(n18764) );
  NAND2_X1 U15885 ( .A1(n17349), .A2(n18334), .ZN(n12896) );
  OAI21_X1 U15886 ( .B1(n18788), .B2(n18308), .A(n18328), .ZN(n12891) );
  OAI211_X1 U15887 ( .C1(n18788), .C2(n18328), .A(n12898), .B(n12891), .ZN(
        n12892) );
  INV_X1 U15888 ( .A(n12892), .ZN(n12893) );
  INV_X1 U15889 ( .A(n17349), .ZN(n18339) );
  NAND2_X1 U15890 ( .A1(n18339), .A2(n18328), .ZN(n12906) );
  INV_X1 U15891 ( .A(n18328), .ZN(n12895) );
  INV_X1 U15892 ( .A(n18334), .ZN(n17352) );
  NOR2_X1 U15893 ( .A1(n18764), .A2(n12896), .ZN(n13446) );
  NAND3_X1 U15894 ( .A1(n18313), .A2(n12902), .A3(n13446), .ZN(n12897) );
  NOR3_X1 U15895 ( .A1(n12898), .A2(n18313), .A3(n18774), .ZN(n12911) );
  INV_X1 U15896 ( .A(n15932), .ZN(n12900) );
  INV_X1 U15897 ( .A(n18788), .ZN(n16024) );
  NAND2_X1 U15898 ( .A1(n18313), .A2(n17500), .ZN(n12899) );
  AOI21_X1 U15899 ( .B1(n16024), .B2(n17431), .A(n12899), .ZN(n15916) );
  AOI21_X1 U15900 ( .B1(n12901), .B2(n12900), .A(n15916), .ZN(n12910) );
  INV_X1 U15901 ( .A(n12902), .ZN(n12909) );
  AOI21_X1 U15902 ( .B1(n18318), .B2(n18308), .A(n18788), .ZN(n12907) );
  NAND2_X1 U15903 ( .A1(n18308), .A2(n18959), .ZN(n12903) );
  NAND2_X1 U15904 ( .A1(n18318), .A2(n12903), .ZN(n15917) );
  AOI21_X1 U15905 ( .B1(n17431), .B2(n15928), .A(n18328), .ZN(n12904) );
  AOI21_X1 U15906 ( .B1(n15928), .B2(n15917), .A(n12904), .ZN(n12905) );
  OAI221_X1 U15907 ( .B1(n12907), .B2(n12906), .C1(n12907), .C2(n15928), .A(
        n12905), .ZN(n12908) );
  XNOR2_X1 U15908 ( .A(n12914), .B(n12913), .ZN(n12916) );
  INV_X1 U15909 ( .A(n18748), .ZN(n15931) );
  AOI21_X1 U15910 ( .B1(n12918), .B2(n12917), .A(n15931), .ZN(n18749) );
  NOR2_X1 U15911 ( .A1(n18313), .A2(n18308), .ZN(n13448) );
  NAND2_X1 U15912 ( .A1(n18926), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18821) );
  NOR2_X1 U15913 ( .A1(n18971), .A2(n18821), .ZN(n18957) );
  INV_X1 U15914 ( .A(n18957), .ZN(n18817) );
  NAND2_X1 U15915 ( .A1(n16547), .A2(n17873), .ZN(n12966) );
  NAND3_X1 U15916 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17994) );
  NOR2_X1 U15917 ( .A1(n17994), .A2(n17985), .ZN(n17973) );
  NAND2_X1 U15918 ( .A1(n17682), .A2(n17973), .ZN(n12954) );
  NAND2_X1 U15919 ( .A1(n12919), .A2(n12924), .ZN(n12923) );
  NAND2_X1 U15920 ( .A1(n12920), .A2(n12923), .ZN(n12931) );
  NOR2_X1 U15921 ( .A1(n17479), .A2(n12931), .ZN(n12922) );
  NAND2_X1 U15922 ( .A1(n12922), .A2(n12921), .ZN(n12938) );
  NOR2_X1 U15923 ( .A1(n17472), .A2(n12938), .ZN(n12943) );
  NAND2_X1 U15924 ( .A1(n12943), .A2(n16552), .ZN(n12944) );
  XNOR2_X1 U15925 ( .A(n17475), .B(n12922), .ZN(n12936) );
  AND2_X1 U15926 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12936), .ZN(
        n12937) );
  INV_X1 U15927 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18246) );
  XOR2_X1 U15928 ( .A(n12762), .B(n12923), .Z(n12929) );
  NOR2_X1 U15929 ( .A1(n18246), .A2(n12929), .ZN(n12930) );
  XOR2_X1 U15930 ( .A(n12919), .B(n12924), .Z(n12925) );
  NOR2_X1 U15931 ( .A1(n12925), .A2(n18261), .ZN(n12928) );
  XNOR2_X1 U15932 ( .A(n18261), .B(n12925), .ZN(n17941) );
  NOR2_X1 U15933 ( .A1(n12757), .A2(n18925), .ZN(n12927) );
  NAND3_X1 U15934 ( .A1(n17960), .A2(n12757), .A3(n18925), .ZN(n12926) );
  OAI221_X1 U15935 ( .B1(n12927), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n17960), .C2(n12757), .A(n12926), .ZN(n17940) );
  NOR2_X1 U15936 ( .A1(n17941), .A2(n17940), .ZN(n17939) );
  NOR2_X1 U15937 ( .A1(n12928), .A2(n17939), .ZN(n17931) );
  XNOR2_X1 U15938 ( .A(n18246), .B(n12929), .ZN(n17930) );
  NOR2_X1 U15939 ( .A1(n17931), .A2(n17930), .ZN(n17929) );
  NOR2_X1 U15940 ( .A1(n12930), .A2(n17929), .ZN(n12933) );
  XOR2_X1 U15941 ( .A(n12932), .B(n12931), .Z(n12934) );
  NOR2_X1 U15942 ( .A1(n12933), .A2(n12934), .ZN(n12935) );
  XNOR2_X1 U15943 ( .A(n12934), .B(n12933), .ZN(n17921) );
  XNOR2_X1 U15944 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n12936), .ZN(
        n17903) );
  XOR2_X1 U15945 ( .A(n12939), .B(n12938), .Z(n12941) );
  NOR2_X1 U15946 ( .A1(n12940), .A2(n12941), .ZN(n12942) );
  XNOR2_X1 U15947 ( .A(n12941), .B(n12940), .ZN(n17897) );
  NOR2_X1 U15948 ( .A1(n12942), .A2(n17896), .ZN(n12945) );
  XNOR2_X1 U15949 ( .A(n16552), .B(n12943), .ZN(n12946) );
  NAND2_X1 U15950 ( .A1(n12945), .A2(n12946), .ZN(n17883) );
  NAND2_X1 U15951 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17883), .ZN(
        n12948) );
  NOR2_X1 U15952 ( .A1(n12944), .A2(n12948), .ZN(n12950) );
  INV_X1 U15953 ( .A(n12944), .ZN(n12949) );
  OR2_X1 U15954 ( .A1(n12946), .A2(n12945), .ZN(n17884) );
  OAI21_X1 U15955 ( .B1(n12949), .B2(n12948), .A(n17884), .ZN(n12947) );
  AOI21_X1 U15956 ( .B1(n12949), .B2(n12948), .A(n12947), .ZN(n17869) );
  INV_X1 U15957 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18199) );
  NAND3_X1 U15958 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17967), .A3(
        n16539), .ZN(n12951) );
  XOR2_X1 U15959 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12951), .Z(
        n16550) );
  NOR2_X1 U15960 ( .A1(n17872), .A2(n12952), .ZN(n17828) );
  INV_X1 U15961 ( .A(n12953), .ZN(n18095) );
  INV_X1 U15962 ( .A(n12954), .ZN(n16509) );
  NAND2_X1 U15963 ( .A1(n18105), .A2(n16509), .ZN(n17605) );
  NOR2_X1 U15964 ( .A1(n17605), .A2(n16011), .ZN(n16515) );
  NAND2_X1 U15965 ( .A1(n16515), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12955) );
  XNOR2_X1 U15966 ( .A(n12955), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16546) );
  NAND2_X1 U15967 ( .A1(n16546), .A2(n17801), .ZN(n12963) );
  NOR2_X1 U15968 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21185) );
  INV_X1 U15969 ( .A(n21185), .ZN(n18928) );
  NAND2_X1 U15970 ( .A1(n18971), .A2(n18935), .ZN(n16665) );
  AND2_X1 U15971 ( .A1(n18928), .A2(n16665), .ZN(n18956) );
  OAI21_X4 U15972 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18956), .A(n9796), 
        .ZN(n17961) );
  NAND2_X1 U15973 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17922) );
  NOR2_X4 U15974 ( .A1(n18926), .A2(n17956), .ZN(n17800) );
  INV_X1 U15975 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17639) );
  INV_X1 U15976 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17879) );
  INV_X1 U15977 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16940) );
  NOR2_X1 U15978 ( .A1(n17841), .A2(n16940), .ZN(n16903) );
  NAND2_X1 U15979 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17810) );
  INV_X1 U15980 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17785) );
  INV_X1 U15981 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17752) );
  INV_X1 U15982 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17688) );
  INV_X1 U15983 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17672) );
  INV_X1 U15984 ( .A(n17610), .ZN(n17609) );
  INV_X1 U15985 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16749) );
  INV_X1 U15986 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16728) );
  NAND2_X1 U15987 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16524), .ZN(
        n12956) );
  INV_X1 U15988 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18897) );
  INV_X1 U15989 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18962) );
  NOR2_X1 U15990 ( .A1(n18897), .A2(n16866), .ZN(n16544) );
  NAND2_X1 U15991 ( .A1(n17608), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16526) );
  NOR2_X1 U15992 ( .A1(n16728), .A2(n16526), .ZN(n12957) );
  INV_X1 U15993 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17954) );
  NOR2_X1 U15994 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18971), .ZN(n17797) );
  NOR2_X1 U15995 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18935), .ZN(
        n21184) );
  INV_X1 U15996 ( .A(n21184), .ZN(n18937) );
  OAI221_X1 U15997 ( .B1(n18926), .B2(P3_STATE2_REG_2__SCAN_IN), .C1(
        P3_STATE2_REG_1__SCAN_IN), .C2(n18971), .A(n18937), .ZN(n18306) );
  NAND2_X1 U15998 ( .A1(n18962), .A2(n18306), .ZN(n18612) );
  INV_X1 U15999 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16685) );
  NOR3_X1 U16000 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n16685), .ZN(n18663) );
  NAND2_X1 U16001 ( .A1(n18518), .A2(n18663), .ZN(n18340) );
  OAI21_X2 U16002 ( .B1(n17954), .B2(n17749), .A(n18349), .ZN(n17774) );
  NAND2_X1 U16003 ( .A1(n12957), .A2(n17774), .ZN(n16512) );
  INV_X1 U16004 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16716) );
  XOR2_X1 U16005 ( .A(n16716), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n12960) );
  NOR2_X1 U16006 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17749), .ZN(
        n16525) );
  INV_X1 U16007 ( .A(n18340), .ZN(n18692) );
  INV_X1 U16008 ( .A(n12957), .ZN(n12958) );
  AOI22_X1 U16009 ( .A1(n18692), .A2(n12958), .B1(n17797), .B2(n9860), .ZN(
        n12959) );
  NAND2_X1 U16010 ( .A1(n12959), .A2(n17961), .ZN(n16527) );
  NOR2_X1 U16011 ( .A1(n16525), .A2(n16527), .ZN(n16511) );
  OAI22_X1 U16012 ( .A1(n16512), .A2(n12960), .B1(n16511), .B2(n16716), .ZN(
        n12961) );
  AOI211_X1 U16013 ( .C1(n17800), .C2(n10031), .A(n16544), .B(n12961), .ZN(
        n12962) );
  INV_X1 U16014 ( .A(n12964), .ZN(n12965) );
  NAND2_X1 U16015 ( .A1(n12966), .A2(n12965), .ZN(P3_U2799) );
  NAND2_X1 U16016 ( .A1(n12967), .A2(n9806), .ZN(n12968) );
  XNOR2_X1 U16017 ( .A(n12968), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14424) );
  OR4_X1 U16018 ( .A1(n12972), .A2(n12971), .A3(n12970), .A4(n12969), .ZN(
        n12973) );
  NAND2_X1 U16019 ( .A1(n12974), .A2(n12973), .ZN(n13369) );
  NAND2_X1 U16020 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20846) );
  INV_X1 U16021 ( .A(n20846), .ZN(n20732) );
  OR2_X1 U16022 ( .A1(n13369), .A2(n20732), .ZN(n13212) );
  INV_X1 U16023 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20738) );
  NAND2_X1 U16024 ( .A1(n12975), .A2(n20738), .ZN(n16017) );
  AND2_X1 U16025 ( .A1(n14042), .A2(n16017), .ZN(n12976) );
  OR2_X1 U16026 ( .A1(n13212), .A2(n12976), .ZN(n12983) );
  NAND2_X1 U16027 ( .A1(n14138), .A2(n16017), .ZN(n14041) );
  NAND2_X1 U16028 ( .A1(n14041), .A2(n20846), .ZN(n12978) );
  OAI211_X1 U16029 ( .C1(n12977), .C2(n12978), .A(n13547), .B(n13217), .ZN(
        n12979) );
  INV_X1 U16030 ( .A(n12979), .ZN(n12980) );
  OR2_X1 U16031 ( .A1(n13429), .A2(n12980), .ZN(n12982) );
  MUX2_X1 U16032 ( .A(n12983), .B(n12982), .S(n12981), .Z(n12991) );
  NOR2_X1 U16033 ( .A1(n13923), .A2(n14138), .ZN(n13113) );
  INV_X1 U16034 ( .A(n12984), .ZN(n12989) );
  NOR2_X1 U16035 ( .A1(n13113), .A2(n11788), .ZN(n12985) );
  NAND2_X1 U16036 ( .A1(n12986), .A2(n12985), .ZN(n13098) );
  INV_X1 U16037 ( .A(n12994), .ZN(n12987) );
  NAND2_X1 U16038 ( .A1(n13098), .A2(n12987), .ZN(n12988) );
  AND2_X1 U16039 ( .A1(n12989), .A2(n12988), .ZN(n13408) );
  AOI21_X1 U16040 ( .B1(n13429), .B2(n13113), .A(n13408), .ZN(n12990) );
  NAND2_X1 U16041 ( .A1(n12991), .A2(n12990), .ZN(n12992) );
  OR2_X1 U16042 ( .A1(n12994), .A2(n14038), .ZN(n13421) );
  AND2_X1 U16043 ( .A1(n13421), .A2(n15985), .ZN(n13367) );
  OAI211_X1 U16044 ( .C1(n11786), .C2(n12997), .A(n11801), .B(n13367), .ZN(
        n12995) );
  NAND2_X1 U16045 ( .A1(n13361), .A2(n14138), .ZN(n15998) );
  OAI21_X1 U16046 ( .B1(n12997), .B2(n12996), .A(n15998), .ZN(n12998) );
  INV_X1 U16047 ( .A(n13061), .ZN(n13091) );
  NAND2_X1 U16048 ( .A1(n13064), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12999) );
  OAI211_X1 U16049 ( .C1(n14540), .C2(P1_EBX_REG_1__SCAN_IN), .A(n9772), .B(
        n12999), .ZN(n13000) );
  NAND2_X1 U16050 ( .A1(n13001), .A2(n13000), .ZN(n13005) );
  INV_X1 U16051 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13002) );
  OR2_X1 U16052 ( .A1(n9772), .A2(n13002), .ZN(n13004) );
  NAND2_X1 U16053 ( .A1(n13091), .A2(n13002), .ZN(n13003) );
  NAND2_X1 U16054 ( .A1(n13004), .A2(n13003), .ZN(n13658) );
  XNOR2_X1 U16055 ( .A(n13005), .B(n13658), .ZN(n13566) );
  AOI21_X1 U16056 ( .B1(n13566), .B2(n13560), .A(n13005), .ZN(n13651) );
  MUX2_X1 U16057 ( .A(n13080), .B(n13064), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n13008) );
  OR2_X1 U16058 ( .A1(n9773), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13007) );
  MUX2_X1 U16059 ( .A(n13090), .B(n9772), .S(P1_EBX_REG_3__SCAN_IN), .Z(n13011) );
  OR2_X1 U16060 ( .A1(n9772), .A2(n13560), .ZN(n13058) );
  NAND2_X1 U16061 ( .A1(n14540), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13009) );
  AND2_X1 U16062 ( .A1(n13058), .A2(n13009), .ZN(n13010) );
  NAND2_X1 U16063 ( .A1(n13011), .A2(n13010), .ZN(n13774) );
  MUX2_X1 U16064 ( .A(n13080), .B(n13064), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n13012) );
  OAI21_X1 U16065 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n9773), .A(
        n13012), .ZN(n13828) );
  INV_X1 U16066 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20195) );
  NAND2_X1 U16067 ( .A1(n13056), .A2(n20195), .ZN(n13016) );
  NAND2_X1 U16068 ( .A1(n9772), .A2(n13109), .ZN(n13014) );
  NAND2_X1 U16069 ( .A1(n13560), .A2(n20195), .ZN(n13013) );
  NAND3_X1 U16070 ( .A1(n13014), .A2(n13013), .A3(n13064), .ZN(n13015) );
  OR2_X1 U16071 ( .A1(n13080), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n13019) );
  NAND2_X1 U16072 ( .A1(n13064), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13017) );
  OAI211_X1 U16073 ( .C1(n14540), .C2(P1_EBX_REG_6__SCAN_IN), .A(n9772), .B(
        n13017), .ZN(n13018) );
  NAND2_X1 U16074 ( .A1(n13019), .A2(n13018), .ZN(n16206) );
  INV_X1 U16075 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16199) );
  NAND2_X1 U16076 ( .A1(n9772), .A2(n16199), .ZN(n13021) );
  INV_X1 U16077 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20171) );
  NAND2_X1 U16078 ( .A1(n13560), .A2(n20171), .ZN(n13020) );
  NAND3_X1 U16079 ( .A1(n13021), .A2(n13020), .A3(n13064), .ZN(n13022) );
  OAI21_X1 U16080 ( .B1(P1_EBX_REG_7__SCAN_IN), .B2(n13090), .A(n13022), .ZN(
        n14019) );
  OR2_X1 U16081 ( .A1(n13080), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n13025) );
  NAND2_X1 U16082 ( .A1(n13064), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13023) );
  OAI211_X1 U16083 ( .C1(n14540), .C2(P1_EBX_REG_8__SCAN_IN), .A(n9772), .B(
        n13023), .ZN(n13024) );
  NAND2_X1 U16084 ( .A1(n13025), .A2(n13024), .ZN(n14113) );
  INV_X1 U16085 ( .A(n9772), .ZN(n13055) );
  MUX2_X1 U16086 ( .A(n13056), .B(n13055), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n13028) );
  NAND2_X1 U16087 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n14540), .ZN(
        n13026) );
  NAND2_X1 U16088 ( .A1(n13058), .A2(n13026), .ZN(n13027) );
  NOR2_X1 U16089 ( .A1(n13028), .A2(n13027), .ZN(n14232) );
  MUX2_X1 U16090 ( .A(n13080), .B(n13064), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n13030) );
  OR2_X1 U16091 ( .A1(n9773), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13029) );
  AND2_X1 U16092 ( .A1(n13030), .A2(n13029), .ZN(n14221) );
  MUX2_X1 U16093 ( .A(n13090), .B(n9772), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13033) );
  NAND2_X1 U16094 ( .A1(n14540), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13031) );
  AND2_X1 U16095 ( .A1(n13058), .A2(n13031), .ZN(n13032) );
  NAND2_X1 U16096 ( .A1(n13033), .A2(n13032), .ZN(n14302) );
  MUX2_X1 U16097 ( .A(n13080), .B(n13064), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n13035) );
  OR2_X1 U16098 ( .A1(n9773), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13034) );
  NAND2_X1 U16099 ( .A1(n13035), .A2(n13034), .ZN(n14325) );
  MUX2_X1 U16100 ( .A(n13080), .B(n13064), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n13037) );
  OR2_X1 U16101 ( .A1(n9773), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13036) );
  AND2_X1 U16102 ( .A1(n13037), .A2(n13036), .ZN(n14256) );
  INV_X1 U16103 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n13038) );
  NAND2_X1 U16104 ( .A1(n13056), .A2(n13038), .ZN(n13042) );
  NAND2_X1 U16105 ( .A1(n9772), .A2(n16181), .ZN(n13040) );
  NAND2_X1 U16106 ( .A1(n13560), .A2(n13038), .ZN(n13039) );
  NAND3_X1 U16107 ( .A1(n13040), .A2(n13039), .A3(n13064), .ZN(n13041) );
  NAND2_X1 U16108 ( .A1(n13042), .A2(n13041), .ZN(n14278) );
  NAND2_X1 U16109 ( .A1(n14256), .A2(n14278), .ZN(n13043) );
  MUX2_X1 U16110 ( .A(n13056), .B(n13055), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n13046) );
  NAND2_X1 U16111 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n14540), .ZN(
        n13044) );
  NAND2_X1 U16112 ( .A1(n13058), .A2(n13044), .ZN(n13045) );
  NOR2_X1 U16113 ( .A1(n13046), .A2(n13045), .ZN(n14344) );
  MUX2_X1 U16114 ( .A(n13080), .B(n13064), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n13048) );
  OR2_X1 U16115 ( .A1(n9773), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13047) );
  NAND2_X1 U16116 ( .A1(n13048), .A2(n13047), .ZN(n14345) );
  INV_X1 U16117 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15090) );
  NAND2_X1 U16118 ( .A1(n9772), .A2(n15090), .ZN(n13050) );
  INV_X1 U16119 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14727) );
  NAND2_X1 U16120 ( .A1(n13560), .A2(n14727), .ZN(n13049) );
  NAND3_X1 U16121 ( .A1(n13050), .A2(n13049), .A3(n13064), .ZN(n13051) );
  OAI21_X1 U16122 ( .B1(P1_EBX_REG_17__SCAN_IN), .B2(n13090), .A(n13051), .ZN(
        n14677) );
  OR2_X1 U16123 ( .A1(n13080), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n13054) );
  NAND2_X1 U16124 ( .A1(n13064), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13052) );
  OAI211_X1 U16125 ( .C1(n14540), .C2(P1_EBX_REG_18__SCAN_IN), .A(n9772), .B(
        n13052), .ZN(n13053) );
  NAND2_X1 U16126 ( .A1(n13054), .A2(n13053), .ZN(n15076) );
  MUX2_X1 U16127 ( .A(n13056), .B(n13055), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n13060) );
  NAND2_X1 U16128 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n14540), .ZN(
        n13057) );
  NAND2_X1 U16129 ( .A1(n13058), .A2(n13057), .ZN(n13059) );
  NOR2_X1 U16130 ( .A1(n13060), .A2(n13059), .ZN(n14722) );
  MUX2_X1 U16131 ( .A(n13080), .B(n13064), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n13063) );
  OR2_X1 U16132 ( .A1(n9773), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13062) );
  NAND2_X1 U16133 ( .A1(n13063), .A2(n13062), .ZN(n14713) );
  NAND2_X1 U16134 ( .A1(n9772), .A2(n15045), .ZN(n13066) );
  INV_X1 U16135 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14708) );
  NAND2_X1 U16136 ( .A1(n13560), .A2(n14708), .ZN(n13065) );
  NAND3_X1 U16137 ( .A1(n13066), .A2(n13065), .A3(n13064), .ZN(n13067) );
  OAI21_X1 U16138 ( .B1(P1_EBX_REG_21__SCAN_IN), .B2(n13090), .A(n13067), .ZN(
        n14706) );
  MUX2_X1 U16139 ( .A(n13080), .B(n13064), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n13069) );
  OR2_X1 U16140 ( .A1(n9773), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13068) );
  NAND2_X1 U16141 ( .A1(n13069), .A2(n13068), .ZN(n14663) );
  MUX2_X1 U16142 ( .A(n13090), .B(n9772), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n13071) );
  NAND2_X1 U16143 ( .A1(n14540), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13070) );
  NAND2_X1 U16144 ( .A1(n13071), .A2(n13070), .ZN(n14698) );
  MUX2_X1 U16145 ( .A(n13080), .B(n13064), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n13073) );
  OR2_X1 U16146 ( .A1(n9773), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13072) );
  AND2_X1 U16147 ( .A1(n13073), .A2(n13072), .ZN(n14648) );
  NAND2_X1 U16148 ( .A1(n14698), .A2(n14648), .ZN(n13074) );
  NAND2_X1 U16149 ( .A1(n9772), .A2(n14996), .ZN(n13075) );
  OAI211_X1 U16150 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n14540), .A(n13075), .B(
        n13064), .ZN(n13076) );
  OAI21_X1 U16151 ( .B1(P1_EBX_REG_25__SCAN_IN), .B2(n13090), .A(n13076), .ZN(
        n14630) );
  OR2_X1 U16152 ( .A1(n13080), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n13079) );
  NAND2_X1 U16153 ( .A1(n13064), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13077) );
  OAI211_X1 U16154 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n14540), .A(n9772), .B(
        n13077), .ZN(n13078) );
  NAND2_X1 U16155 ( .A1(n13079), .A2(n13078), .ZN(n14620) );
  MUX2_X1 U16156 ( .A(n13080), .B(n13064), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n13082) );
  OR2_X1 U16157 ( .A1(n9773), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13081) );
  AND2_X1 U16158 ( .A1(n13082), .A2(n13081), .ZN(n14592) );
  NAND2_X1 U16159 ( .A1(n9772), .A2(n14989), .ZN(n13085) );
  OR2_X1 U16160 ( .A1(n14540), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n13084) );
  NAND3_X1 U16161 ( .A1(n13085), .A2(n13064), .A3(n13084), .ZN(n13086) );
  OAI21_X1 U16162 ( .B1(P1_EBX_REG_27__SCAN_IN), .B2(n13090), .A(n13086), .ZN(
        n14605) );
  NAND2_X1 U16163 ( .A1(n14592), .A2(n14605), .ZN(n13087) );
  OR2_X1 U16164 ( .A1(n9773), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13089) );
  OR2_X1 U16165 ( .A1(n14540), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n13088) );
  NAND2_X1 U16166 ( .A1(n13089), .A2(n13088), .ZN(n14569) );
  OAI22_X1 U16167 ( .A1(n14569), .A2(n13091), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n13090), .ZN(n13092) );
  NOR2_X1 U16168 ( .A1(n14593), .A2(n13092), .ZN(n13093) );
  NAND2_X1 U16169 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20303) );
  NOR3_X1 U16170 ( .A1(n20320), .A2(n9923), .A3(n20303), .ZN(n14241) );
  NAND2_X1 U16171 ( .A1(n13095), .A2(n14042), .ZN(n13096) );
  AND3_X1 U16172 ( .A1(n13098), .A2(n13097), .A3(n13096), .ZN(n13420) );
  INV_X1 U16173 ( .A(n14044), .ZN(n13100) );
  AND2_X1 U16174 ( .A1(n13100), .A2(n13099), .ZN(n13101) );
  OR2_X1 U16175 ( .A1(n13102), .A2(n13101), .ZN(n13112) );
  INV_X1 U16176 ( .A(n13112), .ZN(n13106) );
  MUX2_X1 U16177 ( .A(n13103), .B(n12981), .S(n13547), .Z(n13104) );
  NAND4_X1 U16178 ( .A1(n13420), .A2(n13106), .A3(n13105), .A4(n13104), .ZN(
        n13107) );
  INV_X1 U16179 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13642) );
  AND2_X1 U16180 ( .A1(n12984), .A2(n14042), .ZN(n15150) );
  NAND2_X1 U16181 ( .A1(n13120), .A2(n15150), .ZN(n16175) );
  NAND2_X1 U16182 ( .A1(n13108), .A2(n16175), .ZN(n20321) );
  NAND2_X1 U16183 ( .A1(n14241), .A2(n20321), .ZN(n14238) );
  NAND2_X1 U16184 ( .A1(n13110), .A2(n12977), .ZN(n13111) );
  NOR2_X1 U16185 ( .A1(n13112), .A2(n13111), .ZN(n13418) );
  AOI21_X1 U16186 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13790) );
  NOR2_X1 U16187 ( .A1(n13790), .A2(n20303), .ZN(n16217) );
  NAND2_X1 U16188 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n16217), .ZN(
        n14239) );
  NOR2_X1 U16189 ( .A1(n20314), .A2(n14239), .ZN(n15051) );
  INV_X1 U16190 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16190) );
  NAND3_X1 U16191 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14309) );
  NOR3_X1 U16192 ( .A1(n16190), .A2(n16189), .A3(n14309), .ZN(n15125) );
  NAND2_X1 U16193 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15125), .ZN(
        n15131) );
  NOR2_X1 U16194 ( .A1(n15134), .A2(n15131), .ZN(n15052) );
  NAND2_X1 U16195 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15052), .ZN(
        n13118) );
  INV_X1 U16196 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15084) );
  NOR4_X1 U16197 ( .A1(n12058), .A2(n14922), .A3(n15090), .A4(n15084), .ZN(
        n15074) );
  INV_X1 U16198 ( .A(n15074), .ZN(n15079) );
  NOR2_X1 U16199 ( .A1(n12068), .A2(n15079), .ZN(n13119) );
  AND2_X1 U16200 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15020) );
  INV_X1 U16201 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14998) );
  NOR2_X1 U16202 ( .A1(n14993), .A2(n14998), .ZN(n13114) );
  NAND3_X1 U16203 ( .A1(n14990), .A2(n14957), .A3(n13133), .ZN(n13116) );
  INV_X1 U16204 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21141) );
  NOR2_X1 U16205 ( .A1(n20207), .A2(n21141), .ZN(n14420) );
  INV_X1 U16206 ( .A(n14420), .ZN(n13115) );
  OAI211_X1 U16207 ( .C1(n16218), .C2(n14690), .A(n13116), .B(n13115), .ZN(
        n13117) );
  INV_X1 U16208 ( .A(n13117), .ZN(n13134) );
  NAND2_X1 U16209 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14241), .ZN(
        n14310) );
  INV_X1 U16210 ( .A(n14310), .ZN(n15126) );
  NAND2_X1 U16211 ( .A1(n15126), .A2(n15052), .ZN(n16176) );
  NOR2_X1 U16212 ( .A1(n16181), .A2(n16176), .ZN(n15071) );
  AOI21_X1 U16213 ( .B1(n15071), .B2(n13119), .A(n15124), .ZN(n13122) );
  NOR2_X1 U16214 ( .A1(n14239), .A2(n13118), .ZN(n15070) );
  AOI21_X1 U16215 ( .B1(n13119), .B2(n15070), .A(n20314), .ZN(n13121) );
  OAI22_X1 U16216 ( .A1(n20299), .A2(n13120), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n15050), .ZN(n15073) );
  NOR3_X1 U16217 ( .A1(n13122), .A2(n13121), .A3(n15073), .ZN(n15063) );
  NAND2_X1 U16218 ( .A1(n15063), .A2(n10221), .ZN(n13125) );
  INV_X1 U16219 ( .A(n15073), .ZN(n13123) );
  AND2_X1 U16220 ( .A1(n15100), .A2(n13123), .ZN(n14313) );
  INV_X1 U16221 ( .A(n14313), .ZN(n13124) );
  NAND2_X1 U16222 ( .A1(n13125), .A2(n13124), .ZN(n15041) );
  OR2_X1 U16223 ( .A1(n15100), .A2(n15020), .ZN(n13126) );
  NAND2_X1 U16224 ( .A1(n15041), .A2(n13126), .ZN(n15029) );
  NOR2_X1 U16225 ( .A1(n20314), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13127) );
  NAND2_X1 U16226 ( .A1(n20314), .A2(n16175), .ZN(n13128) );
  NAND2_X1 U16227 ( .A1(n13128), .A2(n14993), .ZN(n13129) );
  OAI21_X1 U16228 ( .B1(n14997), .B2(n15050), .A(n13129), .ZN(n13130) );
  NAND2_X1 U16229 ( .A1(n15004), .A2(n15100), .ZN(n14962) );
  NAND3_X1 U16230 ( .A1(n15004), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13131) );
  NAND2_X1 U16231 ( .A1(n14962), .A2(n13131), .ZN(n14987) );
  INV_X1 U16232 ( .A(n14957), .ZN(n14980) );
  NAND2_X1 U16233 ( .A1(n14962), .A2(n14980), .ZN(n13132) );
  AND2_X1 U16234 ( .A1(n14987), .A2(n13132), .ZN(n14961) );
  AND2_X1 U16235 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13135) );
  NAND2_X1 U16236 ( .A1(n13176), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13173) );
  NAND2_X1 U16237 ( .A1(n13174), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13171) );
  INV_X1 U16238 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19123) );
  INV_X1 U16239 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16358) );
  INV_X1 U16240 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16347) );
  NAND2_X1 U16241 ( .A1(n13168), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13165) );
  INV_X1 U16242 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16340) );
  NAND2_X1 U16243 ( .A1(n13166), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13162) );
  INV_X1 U16244 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13164) );
  NAND2_X1 U16245 ( .A1(n13163), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13161) );
  INV_X1 U16246 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14411) );
  INV_X1 U16247 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15495) );
  INV_X1 U16248 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15501) );
  AND2_X1 U16249 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n13151) );
  INV_X1 U16250 ( .A(n13151), .ZN(n13136) );
  NOR2_X1 U16251 ( .A1(n15501), .A2(n13136), .ZN(n13149) );
  AND2_X1 U16252 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n13149), .ZN(
        n13147) );
  INV_X1 U16253 ( .A(n13147), .ZN(n13137) );
  NOR2_X1 U16254 ( .A1(n15495), .A2(n13137), .ZN(n13138) );
  AND2_X1 U16255 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13142) );
  AND2_X1 U16256 ( .A1(n13142), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13139) );
  INV_X1 U16257 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n21126) );
  INV_X1 U16258 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15468) );
  NAND2_X1 U16259 ( .A1(n13144), .A2(n13142), .ZN(n13145) );
  AOI21_X1 U16260 ( .B1(n15468), .B2(n13145), .A(n13143), .ZN(n16253) );
  INV_X1 U16261 ( .A(n13144), .ZN(n13183) );
  AND2_X1 U16262 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n13144), .ZN(
        n13182) );
  OAI21_X1 U16263 ( .B1(n13182), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n13145), .ZN(n14484) );
  INV_X1 U16264 ( .A(n14484), .ZN(n13285) );
  NAND2_X1 U16265 ( .A1(n13146), .A2(n13147), .ZN(n13150) );
  AOI21_X1 U16266 ( .B1(n15495), .B2(n13150), .A(n13148), .ZN(n16284) );
  AND2_X1 U16267 ( .A1(n13146), .A2(n13149), .ZN(n13152) );
  OAI21_X1 U16268 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n13152), .A(
        n13150), .ZN(n16327) );
  INV_X1 U16269 ( .A(n16327), .ZN(n16300) );
  NAND2_X1 U16270 ( .A1(n13146), .A2(n13151), .ZN(n13153) );
  AOI21_X1 U16271 ( .B1(n13153), .B2(n15501), .A(n13152), .ZN(n16307) );
  AND2_X1 U16272 ( .A1(n13146), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13155) );
  OAI21_X1 U16273 ( .B1(n13155), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n13153), .ZN(n15515) );
  INV_X1 U16274 ( .A(n15515), .ZN(n15953) );
  NOR2_X1 U16275 ( .A1(n13146), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13154) );
  NOR2_X1 U16276 ( .A1(n13155), .A2(n13154), .ZN(n14524) );
  INV_X1 U16277 ( .A(n13146), .ZN(n13160) );
  INV_X1 U16278 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n13158) );
  INV_X1 U16279 ( .A(n13156), .ZN(n13157) );
  NAND2_X1 U16280 ( .A1(n13158), .A2(n13157), .ZN(n13159) );
  NAND2_X1 U16281 ( .A1(n13160), .A2(n13159), .ZN(n15529) );
  INV_X1 U16282 ( .A(n15529), .ZN(n19001) );
  AOI21_X1 U16283 ( .B1(n13161), .B2(n14411), .A(n13156), .ZN(n19012) );
  AOI21_X1 U16284 ( .B1(n13164), .B2(n13162), .A(n13163), .ZN(n19036) );
  AOI21_X1 U16285 ( .B1(n16340), .B2(n13165), .A(n13166), .ZN(n19065) );
  AOI21_X1 U16286 ( .B1(n16347), .B2(n13167), .A(n13168), .ZN(n19086) );
  AOI21_X1 U16287 ( .B1(n16358), .B2(n13169), .A(n13170), .ZN(n19108) );
  AOI21_X1 U16288 ( .B1(n19123), .B2(n13171), .A(n13172), .ZN(n19127) );
  AOI21_X1 U16289 ( .B1(n19145), .B2(n13173), .A(n13174), .ZN(n19149) );
  INV_X1 U16290 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16383) );
  NAND2_X1 U16291 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n13175), .ZN(
        n13178) );
  AOI21_X1 U16292 ( .B1(n16383), .B2(n13178), .A(n13176), .ZN(n19175) );
  INV_X1 U16293 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20858) );
  NOR2_X1 U16294 ( .A1(n20858), .A2(n13177), .ZN(n13179) );
  AOI21_X1 U16295 ( .B1(n20858), .B2(n13177), .A(n13179), .ZN(n13867) );
  INV_X1 U16296 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19389) );
  AOI22_X1 U16297 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19399), .B1(n19389), 
        .B2(n20119), .ZN(n19197) );
  AOI22_X1 U16298 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19398), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20119), .ZN(n13715) );
  NOR2_X1 U16299 ( .A1(n19197), .A2(n13715), .ZN(n13714) );
  OAI21_X1 U16300 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n13177), .ZN(n13627) );
  NAND2_X1 U16301 ( .A1(n13714), .A2(n13627), .ZN(n13570) );
  NOR2_X1 U16302 ( .A1(n13867), .A2(n13570), .ZN(n19188) );
  OAI21_X1 U16303 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13179), .A(
        n13178), .ZN(n19373) );
  NAND2_X1 U16304 ( .A1(n19188), .A2(n19373), .ZN(n19172) );
  OAI21_X1 U16305 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13176), .A(
        n13173), .ZN(n19160) );
  NAND2_X1 U16306 ( .A1(n19159), .A2(n19160), .ZN(n19147) );
  NOR2_X1 U16307 ( .A1(n19149), .A2(n19147), .ZN(n19135) );
  OAI21_X1 U16308 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13174), .A(
        n13171), .ZN(n19136) );
  NAND2_X1 U16309 ( .A1(n19135), .A2(n19136), .ZN(n19125) );
  NOR2_X1 U16310 ( .A1(n19127), .A2(n19125), .ZN(n19115) );
  OAI21_X1 U16311 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13172), .A(
        n13169), .ZN(n19116) );
  NAND2_X1 U16312 ( .A1(n19115), .A2(n19116), .ZN(n19104) );
  NOR2_X1 U16313 ( .A1(n19108), .A2(n19104), .ZN(n19091) );
  OAI21_X1 U16314 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n13170), .A(
        n13167), .ZN(n19092) );
  NAND2_X1 U16315 ( .A1(n19091), .A2(n19092), .ZN(n19084) );
  NOR2_X1 U16316 ( .A1(n19086), .A2(n19084), .ZN(n19074) );
  OAI21_X1 U16317 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n13168), .A(
        n13165), .ZN(n19075) );
  NAND2_X1 U16318 ( .A1(n19074), .A2(n19075), .ZN(n19063) );
  OAI21_X1 U16319 ( .B1(n19065), .B2(n19063), .A(n13180), .ZN(n19050) );
  OAI21_X1 U16320 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n13166), .A(
        n13162), .ZN(n19051) );
  OAI21_X1 U16321 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n13163), .A(
        n13161), .ZN(n15544) );
  INV_X1 U16322 ( .A(n15544), .ZN(n19025) );
  NOR2_X1 U16323 ( .A1(n19012), .A2(n19011), .ZN(n19010) );
  NOR2_X1 U16324 ( .A1(n10058), .A2(n13240), .ZN(n15951) );
  NOR2_X1 U16325 ( .A1(n15953), .A2(n15951), .ZN(n15952) );
  NOR2_X1 U16326 ( .A1(n10058), .A2(n16299), .ZN(n16283) );
  NOR2_X1 U16327 ( .A1(n16284), .A2(n16283), .ZN(n16282) );
  NOR2_X2 U16328 ( .A1(n16282), .A2(n10058), .ZN(n16272) );
  OAI21_X1 U16329 ( .B1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n13148), .A(
        n13183), .ZN(n15484) );
  INV_X1 U16330 ( .A(n15484), .ZN(n16273) );
  INV_X1 U16332 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16261) );
  AOI21_X1 U16333 ( .B1(n13183), .B2(n16261), .A(n13182), .ZN(n16260) );
  NOR2_X1 U16334 ( .A1(n10058), .A2(n13284), .ZN(n16254) );
  XNOR2_X1 U16336 ( .A(n13143), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16246) );
  XNOR2_X1 U16337 ( .A(n13184), .B(n16246), .ZN(n13185) );
  NAND2_X1 U16338 ( .A1(n13185), .A2(n19198), .ZN(n13205) );
  AND2_X1 U16339 ( .A1(n15876), .A2(n20123), .ZN(n13313) );
  AND3_X1 U16340 ( .A1(n13186), .A2(n16502), .A3(n13313), .ZN(n13301) );
  AND2_X2 U16341 ( .A1(n13301), .A2(n19422), .ZN(n19362) );
  NOR2_X1 U16342 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13433), .ZN(n16501) );
  NOR2_X1 U16343 ( .A1(n19422), .A2(n20114), .ZN(n13187) );
  INV_X1 U16344 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20107) );
  INV_X1 U16345 ( .A(n16501), .ZN(n13188) );
  NAND2_X1 U16346 ( .A1(n19362), .A2(n13188), .ZN(n16242) );
  NAND2_X1 U16347 ( .A1(n20107), .A2(n20118), .ZN(n13189) );
  NAND2_X1 U16348 ( .A1(n13301), .A2(n13189), .ZN(n13193) );
  OR2_X1 U16349 ( .A1(n13193), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n13190) );
  NAND2_X1 U16350 ( .A1(n16242), .A2(n13190), .ZN(n19167) );
  INV_X1 U16351 ( .A(n13191), .ZN(n13200) );
  NAND2_X1 U16352 ( .A1(n9748), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n13192) );
  NOR2_X1 U16353 ( .A1(n16473), .A2(n9755), .ZN(n13296) );
  INV_X1 U16354 ( .A(n13296), .ZN(n13194) );
  OR2_X1 U16355 ( .A1(n10859), .A2(n13194), .ZN(n20120) );
  INV_X1 U16356 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20113) );
  NAND2_X1 U16357 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20113), .ZN(n15871) );
  NOR2_X1 U16358 ( .A1(n13195), .A2(n15871), .ZN(n16459) );
  INV_X1 U16359 ( .A(n19365), .ZN(n13196) );
  OR2_X1 U16360 ( .A1(n19185), .A2(n19198), .ZN(n13197) );
  NOR2_X1 U16361 ( .A1(n16459), .A2(n13197), .ZN(n13198) );
  NAND2_X1 U16362 ( .A1(n20120), .A2(n13198), .ZN(n19154) );
  NOR2_X1 U16363 ( .A1(n19204), .A2(n19879), .ZN(n19211) );
  AOI22_X1 U16364 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19166), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19204), .ZN(n13199) );
  OAI21_X1 U16365 ( .B1(n13200), .B2(n19169), .A(n13199), .ZN(n13201) );
  AOI21_X1 U16366 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n19167), .A(n13201), .ZN(
        n13202) );
  OAI21_X1 U16367 ( .B1(n15630), .B2(n19199), .A(n13202), .ZN(n13203) );
  NAND2_X1 U16368 ( .A1(n13205), .A2(n13204), .ZN(P2_U2825) );
  INV_X1 U16369 ( .A(n13206), .ZN(n13207) );
  NAND2_X1 U16370 ( .A1(n13207), .A2(n20846), .ZN(n13208) );
  INV_X1 U16371 ( .A(n13209), .ZN(n13210) );
  NAND4_X1 U16372 ( .A1(n13210), .A2(n11786), .A3(n13854), .A4(n13687), .ZN(
        n13559) );
  OR2_X1 U16373 ( .A1(n13211), .A2(n13212), .ZN(n13409) );
  OAI21_X1 U16374 ( .B1(n14038), .B2(n13559), .A(n13409), .ZN(n13213) );
  INV_X1 U16375 ( .A(n13213), .ZN(n13214) );
  OAI21_X1 U16376 ( .B1(n13429), .B2(n13404), .A(n13214), .ZN(n13215) );
  AND2_X1 U16377 ( .A1(n14762), .A2(n13854), .ZN(n13216) );
  NAND2_X1 U16378 ( .A1(n14545), .A2(n13216), .ZN(n13233) );
  NOR4_X1 U16379 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n13221) );
  NOR4_X1 U16380 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13220) );
  NOR4_X1 U16381 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n13219) );
  NOR4_X1 U16382 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13218) );
  AND4_X1 U16383 ( .A1(n13221), .A2(n13220), .A3(n13219), .A4(n13218), .ZN(
        n13226) );
  NOR4_X1 U16384 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_3__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n13224) );
  NOR4_X1 U16385 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n13223) );
  NOR4_X1 U16386 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P1_ADDRESS_REG_27__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_25__SCAN_IN), .ZN(n13222) );
  INV_X1 U16387 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20748) );
  AND4_X1 U16388 ( .A1(n13224), .A2(n13223), .A3(n13222), .A4(n20748), .ZN(
        n13225) );
  NAND2_X1 U16389 ( .A1(n13226), .A2(n13225), .ZN(n13227) );
  INV_X1 U16390 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16571) );
  NOR2_X1 U16391 ( .A1(n14793), .A2(n16571), .ZN(n13231) );
  NOR2_X2 U16392 ( .A1(n13228), .A2(n14327), .ZN(n14802) );
  AOI22_X1 U16393 ( .A1(n14802), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14789), .ZN(n13229) );
  NOR2_X1 U16394 ( .A1(n13231), .A2(n13230), .ZN(n13232) );
  NAND2_X1 U16395 ( .A1(n13233), .A2(n13232), .ZN(P1_U2873) );
  INV_X1 U16396 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20837) );
  NOR3_X1 U16397 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20837), .ZN(n13235) );
  NOR4_X1 U16398 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13234) );
  NAND4_X1 U16399 ( .A1(n14327), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13235), .A4(
        n13234), .ZN(U214) );
  NOR2_X1 U16400 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13237) );
  NOR4_X1 U16401 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13236) );
  NAND4_X1 U16402 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13237), .A4(n13236), .ZN(n13238) );
  NOR2_X1 U16403 ( .A1(n15878), .A2(n13238), .ZN(n16570) );
  NAND2_X1 U16404 ( .A1(n16570), .A2(U214), .ZN(U212) );
  NOR2_X1 U16405 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13238), .ZN(n16655)
         );
  INV_X1 U16406 ( .A(n19198), .ZN(n19972) );
  AOI211_X1 U16407 ( .C1(n14524), .C2(n13239), .A(n13240), .B(n19972), .ZN(
        n13250) );
  INV_X1 U16408 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14526) );
  INV_X1 U16409 ( .A(n19211), .ZN(n19144) );
  INV_X1 U16410 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20027) );
  OAI22_X1 U16411 ( .A1(n14526), .A2(n19144), .B1(n20027), .B2(n19154), .ZN(
        n13249) );
  INV_X1 U16412 ( .A(n19167), .ZN(n19207) );
  OAI22_X1 U16413 ( .A1(n13241), .A2(n19169), .B1(n11610), .B2(n19207), .ZN(
        n13248) );
  AND2_X1 U16414 ( .A1(n15315), .A2(n13242), .ZN(n13243) );
  OR2_X1 U16415 ( .A1(n13243), .A2(n15301), .ZN(n15309) );
  NAND2_X1 U16416 ( .A1(n13244), .A2(n13245), .ZN(n13246) );
  OAI22_X1 U16417 ( .A1(n15309), .A2(n19199), .B1(n9821), .B2(n19182), .ZN(
        n13247) );
  OR4_X1 U16418 ( .A1(n13250), .A2(n13249), .A3(n13248), .A4(n13247), .ZN(
        P2_U2834) );
  INV_X1 U16419 ( .A(n13251), .ZN(n19392) );
  MUX2_X1 U16420 ( .A(n15815), .B(n19392), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13263) );
  OAI21_X1 U16421 ( .B1(n13253), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13252), .ZN(n19386) );
  OAI22_X1 U16422 ( .A1(n16411), .A2(n19200), .B1(n19406), .B2(n19386), .ZN(
        n13262) );
  OAI21_X1 U16423 ( .B1(n19201), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13395), .ZN(n19378) );
  INV_X1 U16424 ( .A(n13254), .ZN(n13257) );
  INV_X1 U16425 ( .A(n13255), .ZN(n13256) );
  NAND2_X1 U16426 ( .A1(n13257), .A2(n13256), .ZN(n13259) );
  AND2_X1 U16427 ( .A1(n13259), .A2(n13258), .ZN(n19273) );
  NAND2_X1 U16428 ( .A1(n19391), .A2(n19273), .ZN(n13260) );
  INV_X1 U16429 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18993) );
  NAND2_X1 U16430 ( .A1(n19365), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n19377) );
  OAI211_X1 U16431 ( .C1(n19395), .C2(n19378), .A(n13260), .B(n19377), .ZN(
        n13261) );
  OR3_X1 U16432 ( .A1(n13263), .A2(n13262), .A3(n13261), .ZN(P2_U3046) );
  NOR2_X1 U16433 ( .A1(n14426), .A2(n13264), .ZN(n13872) );
  NOR2_X1 U16434 ( .A1(n14427), .A2(n13266), .ZN(n13268) );
  OAI21_X1 U16435 ( .B1(n14426), .B2(n13266), .A(n13265), .ZN(n13267) );
  MUX2_X1 U16436 ( .A(n13268), .B(n13267), .S(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n13282) );
  OR2_X1 U16437 ( .A1(n13270), .A2(n13269), .ZN(n13272) );
  AND2_X1 U16438 ( .A1(n13272), .A2(n13271), .ZN(n13889) );
  INV_X1 U16439 ( .A(n13889), .ZN(n20074) );
  AND2_X1 U16440 ( .A1(n19185), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n13386) );
  OAI21_X1 U16441 ( .B1(n13275), .B2(n13274), .A(n13273), .ZN(n13381) );
  OAI21_X1 U16442 ( .B1(n13278), .B2(n13277), .A(n13276), .ZN(n13384) );
  OAI22_X1 U16443 ( .A1(n19395), .A2(n13381), .B1(n13384), .B2(n19406), .ZN(
        n13279) );
  AOI211_X1 U16444 ( .C1(n19391), .C2(n20074), .A(n13386), .B(n13279), .ZN(
        n13280) );
  OAI21_X1 U16445 ( .B1(n13588), .B2(n16411), .A(n13280), .ZN(n13281) );
  OR3_X1 U16446 ( .A1(n13872), .A2(n13282), .A3(n13281), .ZN(P2_U3044) );
  AOI211_X1 U16447 ( .C1(n13285), .C2(n13283), .A(n13284), .B(n19972), .ZN(
        n13295) );
  INV_X1 U16448 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13286) );
  OAI22_X1 U16449 ( .A1(n13287), .A2(n19169), .B1(n13286), .B2(n19144), .ZN(
        n13294) );
  OAI22_X1 U16450 ( .A1(n19207), .A2(n11633), .B1(n20041), .B2(n19154), .ZN(
        n13293) );
  NAND2_X1 U16451 ( .A1(n13288), .A2(n13289), .ZN(n13290) );
  NAND2_X1 U16452 ( .A1(n15241), .A2(n13290), .ZN(n15258) );
  OAI22_X1 U16453 ( .A1(n15258), .A2(n19199), .B1(n15359), .B2(n19182), .ZN(
        n13292) );
  OR4_X1 U16454 ( .A1(n13295), .A2(n13294), .A3(n13293), .A4(n13292), .ZN(
        P2_U2827) );
  INV_X1 U16455 ( .A(n10850), .ZN(n13297) );
  NAND2_X1 U16456 ( .A1(n13297), .A2(n13296), .ZN(n13729) );
  INV_X1 U16457 ( .A(n13729), .ZN(n19210) );
  INV_X1 U16458 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n20128) );
  AND2_X1 U16459 ( .A1(n20064), .A2(n13298), .ZN(n14534) );
  INV_X1 U16460 ( .A(n14534), .ZN(n13300) );
  INV_X1 U16461 ( .A(n13301), .ZN(n13299) );
  OAI211_X1 U16462 ( .C1(n19210), .C2(n20128), .A(n13300), .B(n13299), .ZN(
        P2_U2814) );
  OAI21_X1 U16463 ( .B1(n19422), .B2(n20118), .A(n13301), .ZN(n13356) );
  AOI22_X1 U16464 ( .A1(P2_EAX_REG_26__SCAN_IN), .A2(n19362), .B1(n13356), 
        .B2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13304) );
  INV_X1 U16465 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16603) );
  OR2_X1 U16466 ( .A1(n15878), .A2(n16603), .ZN(n13303) );
  NAND2_X1 U16467 ( .A1(n15878), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13302) );
  AND2_X1 U16468 ( .A1(n13303), .A2(n13302), .ZN(n19232) );
  INV_X1 U16469 ( .A(n19232), .ZN(n15374) );
  NAND2_X1 U16470 ( .A1(n19357), .A2(n15374), .ZN(n13327) );
  NAND2_X1 U16471 ( .A1(n13304), .A2(n13327), .ZN(P2_U2962) );
  AOI22_X1 U16472 ( .A1(P2_EAX_REG_23__SCAN_IN), .A2(n19362), .B1(n13356), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13305) );
  INV_X1 U16473 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16607) );
  INV_X1 U16474 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18345) );
  AOI22_X1 U16475 ( .A1(n15880), .A2(n16607), .B1(n18345), .B2(n15878), .ZN(
        n19240) );
  NAND2_X1 U16476 ( .A1(n19357), .A2(n19240), .ZN(n13329) );
  NAND2_X1 U16477 ( .A1(n13305), .A2(n13329), .ZN(P2_U2959) );
  AOI22_X1 U16478 ( .A1(P2_EAX_REG_25__SCAN_IN), .A2(n19362), .B1(n13356), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13308) );
  INV_X1 U16479 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n14207) );
  OR2_X1 U16480 ( .A1(n15878), .A2(n14207), .ZN(n13307) );
  NAND2_X1 U16481 ( .A1(n15878), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13306) );
  AND2_X1 U16482 ( .A1(n13307), .A2(n13306), .ZN(n19236) );
  INV_X1 U16483 ( .A(n19236), .ZN(n15384) );
  NAND2_X1 U16484 ( .A1(n19357), .A2(n15384), .ZN(n13350) );
  NAND2_X1 U16485 ( .A1(n13308), .A2(n13350), .ZN(P2_U2961) );
  INV_X1 U16486 ( .A(n13309), .ZN(n13312) );
  NOR3_X1 U16487 ( .A1(n13312), .A2(n13311), .A3(n13310), .ZN(n16479) );
  NOR2_X1 U16488 ( .A1(n16479), .A2(n9755), .ZN(n20104) );
  NAND2_X1 U16489 ( .A1(n13314), .A2(n13313), .ZN(n13380) );
  OAI21_X1 U16490 ( .B1(n21077), .B2(n20104), .A(n13380), .ZN(P2_U2819) );
  AOI22_X1 U16491 ( .A1(P2_EAX_REG_21__SCAN_IN), .A2(n19362), .B1(n13356), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13315) );
  AOI22_X1 U16492 ( .A1(n15880), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13340), .ZN(n19439) );
  INV_X1 U16493 ( .A(n19439), .ZN(n15408) );
  NAND2_X1 U16494 ( .A1(n19357), .A2(n15408), .ZN(n13325) );
  NAND2_X1 U16495 ( .A1(n13315), .A2(n13325), .ZN(P2_U2957) );
  INV_X1 U16496 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n20917) );
  NAND2_X1 U16497 ( .A1(n15878), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13317) );
  INV_X1 U16498 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n21125) );
  OR2_X1 U16499 ( .A1(n15878), .A2(n21125), .ZN(n13316) );
  NAND2_X1 U16500 ( .A1(n13317), .A2(n13316), .ZN(n19229) );
  NAND2_X1 U16501 ( .A1(n19357), .A2(n19229), .ZN(n13320) );
  NAND2_X1 U16502 ( .A1(n19361), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13318) );
  OAI211_X1 U16503 ( .C1(n19283), .C2(n20917), .A(n13320), .B(n13318), .ZN(
        P2_U2978) );
  INV_X1 U16504 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n21123) );
  NAND2_X1 U16505 ( .A1(n19361), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13319) );
  OAI211_X1 U16506 ( .C1(n19283), .C2(n21123), .A(n13320), .B(n13319), .ZN(
        P2_U2963) );
  AOI22_X1 U16507 ( .A1(P2_EAX_REG_17__SCAN_IN), .A2(n19362), .B1(n19361), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13321) );
  AOI22_X1 U16508 ( .A1(n15880), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13340), .ZN(n19423) );
  INV_X1 U16509 ( .A(n19423), .ZN(n15439) );
  NAND2_X1 U16510 ( .A1(n19357), .A2(n15439), .ZN(n13348) );
  NAND2_X1 U16511 ( .A1(n13321), .A2(n13348), .ZN(P2_U2953) );
  AOI22_X1 U16512 ( .A1(P2_EAX_REG_0__SCAN_IN), .A2(n19362), .B1(n19361), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n13323) );
  AOI22_X1 U16513 ( .A1(n15880), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13340), .ZN(n13322) );
  INV_X1 U16514 ( .A(n13322), .ZN(n19281) );
  NAND2_X1 U16515 ( .A1(n19357), .A2(n19281), .ZN(n13342) );
  NAND2_X1 U16516 ( .A1(n13323), .A2(n13342), .ZN(P2_U2967) );
  AOI22_X1 U16517 ( .A1(P2_EAX_REG_3__SCAN_IN), .A2(n19362), .B1(n19361), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13324) );
  AOI22_X1 U16518 ( .A1(n15880), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13340), .ZN(n19432) );
  INV_X1 U16519 ( .A(n19432), .ZN(n15422) );
  NAND2_X1 U16520 ( .A1(n19357), .A2(n15422), .ZN(n13354) );
  NAND2_X1 U16521 ( .A1(n13324), .A2(n13354), .ZN(P2_U2970) );
  AOI22_X1 U16522 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19362), .B1(n19361), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n13326) );
  NAND2_X1 U16523 ( .A1(n13326), .A2(n13325), .ZN(P2_U2972) );
  AOI22_X1 U16524 ( .A1(n19362), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n19361), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13328) );
  NAND2_X1 U16525 ( .A1(n13328), .A2(n13327), .ZN(P2_U2977) );
  AOI22_X1 U16526 ( .A1(P2_EAX_REG_7__SCAN_IN), .A2(n19362), .B1(n19361), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n13330) );
  NAND2_X1 U16527 ( .A1(n13330), .A2(n13329), .ZN(P2_U2974) );
  AOI22_X1 U16528 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19362), .B1(n19361), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13333) );
  INV_X1 U16529 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n14328) );
  OR2_X1 U16530 ( .A1(n15878), .A2(n14328), .ZN(n13332) );
  NAND2_X1 U16531 ( .A1(n15878), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13331) );
  AND2_X1 U16532 ( .A1(n13332), .A2(n13331), .ZN(n19228) );
  INV_X1 U16533 ( .A(n19228), .ZN(n15356) );
  NAND2_X1 U16534 ( .A1(n19357), .A2(n15356), .ZN(n13334) );
  NAND2_X1 U16535 ( .A1(n13333), .A2(n13334), .ZN(P2_U2979) );
  AOI22_X1 U16536 ( .A1(P2_EAX_REG_28__SCAN_IN), .A2(n19362), .B1(n19361), 
        .B2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13335) );
  NAND2_X1 U16537 ( .A1(n13335), .A2(n13334), .ZN(P2_U2964) );
  AOI22_X1 U16538 ( .A1(n19362), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n19361), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13337) );
  AOI22_X1 U16539 ( .A1(n15880), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n15878), .ZN(n19443) );
  INV_X1 U16540 ( .A(n19443), .ZN(n13336) );
  NAND2_X1 U16541 ( .A1(n19357), .A2(n13336), .ZN(n13352) );
  NAND2_X1 U16542 ( .A1(n13337), .A2(n13352), .ZN(P2_U2958) );
  AOI22_X1 U16543 ( .A1(n19362), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n19361), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13338) );
  INV_X1 U16544 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16613) );
  INV_X1 U16545 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18327) );
  OAI22_X1 U16546 ( .A1(n15878), .A2(n16613), .B1(n18327), .B2(n15880), .ZN(
        n19436) );
  NAND2_X1 U16547 ( .A1(n19357), .A2(n19436), .ZN(n13357) );
  NAND2_X1 U16548 ( .A1(n13338), .A2(n13357), .ZN(P2_U2956) );
  AOI22_X1 U16549 ( .A1(n19362), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n13356), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13339) );
  AOI22_X1 U16550 ( .A1(n15880), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n15878), .ZN(n19237) );
  INV_X1 U16551 ( .A(n19237), .ZN(n15392) );
  NAND2_X1 U16552 ( .A1(n19357), .A2(n15392), .ZN(n13344) );
  NAND2_X1 U16553 ( .A1(n13339), .A2(n13344), .ZN(P2_U2960) );
  AOI22_X1 U16554 ( .A1(n19362), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n19361), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13341) );
  AOI22_X1 U16555 ( .A1(n15880), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13340), .ZN(n19427) );
  INV_X1 U16556 ( .A(n19427), .ZN(n15433) );
  NAND2_X1 U16557 ( .A1(n19357), .A2(n15433), .ZN(n13346) );
  NAND2_X1 U16558 ( .A1(n13341), .A2(n13346), .ZN(P2_U2954) );
  AOI22_X1 U16559 ( .A1(n19362), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n19361), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13343) );
  NAND2_X1 U16560 ( .A1(n13343), .A2(n13342), .ZN(P2_U2952) );
  AOI22_X1 U16561 ( .A1(n19362), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n19361), .B2(
        P2_LWORD_REG_8__SCAN_IN), .ZN(n13345) );
  NAND2_X1 U16562 ( .A1(n13345), .A2(n13344), .ZN(P2_U2975) );
  AOI22_X1 U16563 ( .A1(P2_EAX_REG_2__SCAN_IN), .A2(n19362), .B1(n19361), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13347) );
  NAND2_X1 U16564 ( .A1(n13347), .A2(n13346), .ZN(P2_U2969) );
  AOI22_X1 U16565 ( .A1(P2_EAX_REG_1__SCAN_IN), .A2(n19362), .B1(n19361), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13349) );
  NAND2_X1 U16566 ( .A1(n13349), .A2(n13348), .ZN(P2_U2968) );
  AOI22_X1 U16567 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(n19362), .B1(n19361), .B2(
        P2_LWORD_REG_9__SCAN_IN), .ZN(n13351) );
  NAND2_X1 U16568 ( .A1(n13351), .A2(n13350), .ZN(P2_U2976) );
  AOI22_X1 U16569 ( .A1(P2_EAX_REG_6__SCAN_IN), .A2(n19362), .B1(n19361), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n13353) );
  NAND2_X1 U16570 ( .A1(n13353), .A2(n13352), .ZN(P2_U2973) );
  AOI22_X1 U16571 ( .A1(P2_EAX_REG_19__SCAN_IN), .A2(n19362), .B1(n19361), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13355) );
  NAND2_X1 U16572 ( .A1(n13355), .A2(n13354), .ZN(P2_U2955) );
  AOI22_X1 U16573 ( .A1(P2_EAX_REG_4__SCAN_IN), .A2(n19362), .B1(n13356), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n13358) );
  NAND2_X1 U16574 ( .A1(n13358), .A2(n13357), .ZN(P2_U2971) );
  AOI22_X1 U16575 ( .A1(n15880), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15878), .ZN(n19220) );
  INV_X1 U16576 ( .A(n19357), .ZN(n13360) );
  AOI22_X1 U16577 ( .A1(n19362), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n19361), 
        .B2(P2_LWORD_REG_15__SCAN_IN), .ZN(n13359) );
  OAI21_X1 U16578 ( .B1(n19220), .B2(n13360), .A(n13359), .ZN(P2_U2982) );
  INV_X1 U16579 ( .A(n13361), .ZN(n13390) );
  INV_X1 U16580 ( .A(n13369), .ZN(n13362) );
  NAND2_X1 U16581 ( .A1(n12984), .A2(n13362), .ZN(n13391) );
  AOI22_X1 U16582 ( .A1(n13429), .A2(n14038), .B1(n13390), .B2(n13391), .ZN(
        n20132) );
  NAND3_X1 U16583 ( .A1(n14038), .A2(n14540), .A3(n16017), .ZN(n13363) );
  NAND2_X1 U16584 ( .A1(n13363), .A2(n20846), .ZN(n20838) );
  NAND2_X1 U16585 ( .A1(n20132), .A2(n20838), .ZN(n15987) );
  AND2_X1 U16586 ( .A1(n15987), .A2(n13564), .ZN(n20141) );
  INV_X1 U16587 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13376) );
  INV_X1 U16588 ( .A(n13422), .ZN(n13372) );
  NAND3_X1 U16589 ( .A1(n13364), .A2(n13365), .A3(n13547), .ZN(n13366) );
  NAND2_X1 U16590 ( .A1(n13367), .A2(n13366), .ZN(n13368) );
  NAND2_X1 U16591 ( .A1(n13429), .A2(n13368), .ZN(n13371) );
  NAND2_X1 U16592 ( .A1(n12984), .A2(n13369), .ZN(n13370) );
  OAI211_X1 U16593 ( .C1(n13429), .C2(n13372), .A(n13371), .B(n13370), .ZN(
        n13373) );
  NAND2_X1 U16594 ( .A1(n13373), .A2(n14360), .ZN(n15984) );
  INV_X1 U16595 ( .A(n15984), .ZN(n13374) );
  NAND2_X1 U16596 ( .A1(n20141), .A2(n13374), .ZN(n13375) );
  OAI21_X1 U16597 ( .B1(n20141), .B2(n13376), .A(n13375), .ZN(P1_U3484) );
  NOR2_X1 U16598 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13840) );
  OR2_X1 U16599 ( .A1(n20064), .A2(n13840), .ZN(n20077) );
  NAND2_X1 U16600 ( .A1(n20077), .A2(n20119), .ZN(n13377) );
  NAND2_X1 U16601 ( .A1(n20107), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13378) );
  NAND2_X1 U16602 ( .A1(n13379), .A2(n13378), .ZN(n19375) );
  INV_X1 U16603 ( .A(n13380), .ZN(n13382) );
  NAND2_X1 U16604 ( .A1(n13382), .A2(n9748), .ZN(n19379) );
  INV_X1 U16605 ( .A(n19379), .ZN(n16379) );
  INV_X1 U16606 ( .A(n13381), .ZN(n13387) );
  NAND2_X1 U16607 ( .A1(n13382), .A2(n19422), .ZN(n19385) );
  INV_X1 U16608 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13383) );
  OAI22_X1 U16609 ( .A1(n19385), .A2(n13384), .B1(n16382), .B2(n13383), .ZN(
        n13385) );
  AOI211_X1 U16610 ( .C1(n16379), .C2(n13387), .A(n13386), .B(n13385), .ZN(
        n13389) );
  AND2_X1 U16611 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20078) );
  NAND2_X1 U16612 ( .A1(n15847), .A2(n19382), .ZN(n13388) );
  OAI211_X1 U16613 ( .C1(n13627), .C2(n19374), .A(n13389), .B(n13388), .ZN(
        P2_U3012) );
  NOR2_X1 U16614 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20667), .ZN(n14564) );
  NOR2_X1 U16615 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(n14564), .ZN(n13394)
         );
  NAND2_X1 U16616 ( .A1(n20844), .A2(n13392), .ZN(n13393) );
  OAI21_X1 U16617 ( .B1(n20844), .B2(n13394), .A(n13393), .ZN(P1_U3487) );
  INV_X1 U16618 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13402) );
  XNOR2_X1 U16619 ( .A(n13395), .B(n19398), .ZN(n13396) );
  XNOR2_X1 U16620 ( .A(n13722), .B(n13396), .ZN(n19394) );
  NAND2_X1 U16621 ( .A1(n19365), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n19403) );
  OAI21_X1 U16622 ( .B1(n19379), .B2(n19394), .A(n19403), .ZN(n13401) );
  OR2_X1 U16623 ( .A1(n13397), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13399) );
  NAND2_X1 U16624 ( .A1(n13399), .A2(n13398), .ZN(n19405) );
  OAI22_X1 U16625 ( .A1(n19385), .A2(n19405), .B1(n16382), .B2(n13402), .ZN(
        n13400) );
  AOI211_X1 U16626 ( .C1(n16370), .C2(n13402), .A(n13401), .B(n13400), .ZN(
        n13403) );
  OAI21_X1 U16627 ( .B1(n13602), .B2(n14529), .A(n13403), .ZN(P2_U3013) );
  NAND2_X1 U16628 ( .A1(n13429), .A2(n13422), .ZN(n13563) );
  NAND2_X1 U16629 ( .A1(n13421), .A2(n12977), .ZN(n13406) );
  OAI21_X1 U16630 ( .B1(n20732), .B2(n16017), .A(n13404), .ZN(n13405) );
  OAI21_X1 U16631 ( .B1(n15150), .B2(n13406), .A(n13405), .ZN(n13407) );
  OR2_X1 U16632 ( .A1(n13429), .A2(n13407), .ZN(n13414) );
  INV_X1 U16633 ( .A(n13408), .ZN(n13410) );
  OAI211_X1 U16634 ( .C1(n14044), .C2(n13411), .A(n13410), .B(n13409), .ZN(
        n13412) );
  INV_X1 U16635 ( .A(n13412), .ZN(n13413) );
  NAND3_X1 U16636 ( .A1(n13563), .A2(n13414), .A3(n13413), .ZN(n13694) );
  NOR2_X1 U16637 ( .A1(n20839), .A2(n20727), .ZN(n16233) );
  INV_X1 U16638 ( .A(n16233), .ZN(n16237) );
  NOR2_X1 U16639 ( .A1(n9918), .A2(n16237), .ZN(n13702) );
  AOI22_X1 U16640 ( .A1(n13564), .A2(n13694), .B1(P1_FLUSH_REG_SCAN_IN), .B2(
        n13702), .ZN(n16228) );
  OAI21_X1 U16641 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n20526), .A(n16228), 
        .ZN(n20807) );
  INV_X1 U16642 ( .A(n20807), .ZN(n14502) );
  INV_X1 U16643 ( .A(n13415), .ZN(n14046) );
  INV_X1 U16644 ( .A(n13416), .ZN(n13417) );
  AND2_X1 U16645 ( .A1(n13418), .A2(n13417), .ZN(n13419) );
  NAND3_X1 U16646 ( .A1(n13420), .A2(n13419), .A3(n13211), .ZN(n15155) );
  INV_X1 U16647 ( .A(n15155), .ZN(n14499) );
  INV_X1 U16648 ( .A(n13421), .ZN(n13423) );
  OR2_X1 U16649 ( .A1(n13423), .A2(n13422), .ZN(n13684) );
  INV_X1 U16650 ( .A(n13424), .ZN(n15151) );
  NAND2_X1 U16651 ( .A1(n15151), .A2(n9930), .ZN(n13679) );
  NAND2_X1 U16652 ( .A1(n13424), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13685) );
  AND2_X1 U16653 ( .A1(n13679), .A2(n13685), .ZN(n13430) );
  INV_X1 U16654 ( .A(n13430), .ZN(n13426) );
  XNOR2_X1 U16655 ( .A(n9930), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13425) );
  AOI22_X1 U16656 ( .A1(n13684), .A2(n13426), .B1(n15150), .B2(n13425), .ZN(
        n13428) );
  NAND3_X1 U16657 ( .A1(n14499), .A2(n13687), .A3(n13430), .ZN(n13427) );
  OAI211_X1 U16658 ( .C1(n13415), .C2(n14499), .A(n13428), .B(n13427), .ZN(
        n13695) );
  NOR2_X1 U16659 ( .A1(n20727), .A2(n13642), .ZN(n15159) );
  INV_X1 U16660 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n20945) );
  AOI22_X1 U16661 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n9923), .B2(n20945), .ZN(
        n15157) );
  AOI222_X1 U16662 ( .A1(n13695), .A2(n20804), .B1(n15159), .B2(n15157), .C1(
        n13430), .C2(n20803), .ZN(n13432) );
  NAND2_X1 U16663 ( .A1(n14502), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13431) );
  OAI21_X1 U16664 ( .B1(n14502), .B2(n13432), .A(n13431), .ZN(P1_U3472) );
  NOR2_X1 U16665 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19879), .ZN(n16506) );
  OR2_X1 U16666 ( .A1(n10850), .A2(n13433), .ZN(n13439) );
  INV_X1 U16667 ( .A(n13434), .ZN(n13435) );
  NOR2_X1 U16668 ( .A1(n13436), .A2(n13435), .ZN(n13437) );
  OAI211_X1 U16669 ( .C1(n13439), .C2(n19285), .A(n13438), .B(n13437), .ZN(
        n16488) );
  INV_X1 U16670 ( .A(n16488), .ZN(n16483) );
  AND2_X1 U16671 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20089) );
  NAND2_X1 U16672 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20089), .ZN(n16500) );
  OAI22_X1 U16673 ( .A1(n16483), .A2(n9755), .B1(n21077), .B2(n16500), .ZN(
        n13440) );
  NOR2_X1 U16674 ( .A1(n16506), .A2(n13440), .ZN(n15862) );
  INV_X1 U16675 ( .A(n15862), .ZN(n13445) );
  INV_X1 U16676 ( .A(n13840), .ZN(n20061) );
  NAND2_X1 U16677 ( .A1(n19422), .A2(n13441), .ZN(n13442) );
  OR2_X1 U16678 ( .A1(n10850), .A2(n13442), .ZN(n16480) );
  OR3_X1 U16679 ( .A1(n15862), .A2(n20061), .A3(n16480), .ZN(n13443) );
  OAI21_X1 U16680 ( .B1(n13445), .B2(n13444), .A(n13443), .ZN(P2_U3595) );
  INV_X1 U16681 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n20963) );
  INV_X1 U16682 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17096) );
  NOR2_X1 U16683 ( .A1(n20963), .A2(n17096), .ZN(n13538) );
  INV_X1 U16684 ( .A(n18745), .ZN(n15924) );
  NAND3_X1 U16685 ( .A1(n18328), .A2(n18348), .A3(n13446), .ZN(n13447) );
  OAI21_X1 U16686 ( .B1(n15923), .B2(n15924), .A(n13447), .ZN(n16021) );
  NAND3_X1 U16687 ( .A1(n16021), .A2(n13448), .A3(n18957), .ZN(n14375) );
  NAND2_X1 U16688 ( .A1(n18348), .A2(n17346), .ZN(n17341) );
  INV_X2 U16689 ( .A(n17343), .ZN(n17338) );
  INV_X1 U16690 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17158) );
  INV_X1 U16691 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16838) );
  INV_X1 U16692 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17200) );
  INV_X1 U16693 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16914) );
  INV_X1 U16694 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n13450) );
  INV_X1 U16695 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n20960) );
  NAND2_X1 U16696 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17334) );
  NOR2_X1 U16697 ( .A1(n20960), .A2(n17334), .ZN(n17327) );
  NAND3_X1 U16698 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17327), .ZN(n17318) );
  INV_X1 U16699 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16937) );
  INV_X1 U16700 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17274) );
  INV_X1 U16701 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17319) );
  NAND2_X1 U16702 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .ZN(n17317) );
  NOR4_X1 U16703 ( .A1(n16937), .A2(n17274), .A3(n17319), .A4(n17317), .ZN(
        n13449) );
  NAND3_X1 U16704 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(n13449), .ZN(n14376) );
  NOR4_X1 U16705 ( .A1(n16914), .A2(n13450), .A3(n17318), .A4(n14376), .ZN(
        n13451) );
  NAND4_X1 U16706 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(P3_EBX_REG_14__SCAN_IN), .A4(n13451), .ZN(n17199) );
  NOR2_X1 U16707 ( .A1(n17200), .A2(n17199), .ZN(n17185) );
  NAND3_X1 U16708 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17346), .A3(n17185), 
        .ZN(n17173) );
  NOR2_X1 U16709 ( .A1(n16838), .A2(n17173), .ZN(n17172) );
  NAND2_X1 U16710 ( .A1(n18348), .A2(n17172), .ZN(n17157) );
  NOR2_X1 U16711 ( .A1(n17158), .A2(n17157), .ZN(n17143) );
  NAND2_X1 U16712 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17143), .ZN(n17131) );
  NAND4_X1 U16713 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(P3_EBX_REG_23__SCAN_IN), .A4(P3_EBX_REG_22__SCAN_IN), .ZN(n13537)
         );
  NOR2_X1 U16714 ( .A1(n17131), .A2(n13537), .ZN(n17106) );
  NAND2_X1 U16715 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17106), .ZN(n17097) );
  NAND2_X1 U16716 ( .A1(n17338), .A2(n17097), .ZN(n17095) );
  OAI21_X1 U16717 ( .B1(n13538), .B2(n17341), .A(n17095), .ZN(n17089) );
  AOI22_X1 U16718 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13455) );
  AOI22_X1 U16719 ( .A1(n12749), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13454) );
  AOI22_X1 U16720 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13453) );
  AOI22_X1 U16721 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13452) );
  NAND4_X1 U16722 ( .A1(n13455), .A2(n13454), .A3(n13453), .A4(n13452), .ZN(
        n13461) );
  AOI22_X1 U16723 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13459) );
  AOI22_X1 U16724 ( .A1(n17267), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13458) );
  AOI22_X1 U16725 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17277), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13457) );
  AOI22_X1 U16726 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17305), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13456) );
  NAND4_X1 U16727 ( .A1(n13459), .A2(n13458), .A3(n13457), .A4(n13456), .ZN(
        n13460) );
  NOR2_X1 U16728 ( .A1(n13461), .A2(n13460), .ZN(n13536) );
  AOI22_X1 U16729 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13465) );
  AOI22_X1 U16730 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9754), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13464) );
  AOI22_X1 U16731 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13463) );
  AOI22_X1 U16732 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13462) );
  NAND4_X1 U16733 ( .A1(n13465), .A2(n13464), .A3(n13463), .A4(n13462), .ZN(
        n13472) );
  AOI22_X1 U16734 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17294), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13470) );
  AOI22_X1 U16735 ( .A1(n17305), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13469) );
  AOI22_X1 U16736 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13468) );
  AOI22_X1 U16737 ( .A1(n12749), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13467) );
  NAND4_X1 U16738 ( .A1(n13470), .A2(n13469), .A3(n13468), .A4(n13467), .ZN(
        n13471) );
  NOR2_X1 U16739 ( .A1(n13472), .A2(n13471), .ZN(n17093) );
  AOI22_X1 U16740 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17305), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13476) );
  AOI22_X1 U16741 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13475) );
  AOI22_X1 U16742 ( .A1(n17248), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13474) );
  AOI22_X1 U16743 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13473) );
  NAND4_X1 U16744 ( .A1(n13476), .A2(n13475), .A3(n13474), .A4(n13473), .ZN(
        n13482) );
  AOI22_X1 U16745 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17294), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13480) );
  AOI22_X1 U16746 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13479) );
  AOI22_X1 U16747 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13478) );
  AOI22_X1 U16748 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13477) );
  NAND4_X1 U16749 ( .A1(n13480), .A2(n13479), .A3(n13478), .A4(n13477), .ZN(
        n13481) );
  NOR2_X1 U16750 ( .A1(n13482), .A2(n13481), .ZN(n17103) );
  AOI22_X1 U16751 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13486) );
  AOI22_X1 U16752 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13485) );
  AOI22_X1 U16753 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13484) );
  AOI22_X1 U16754 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13483) );
  NAND4_X1 U16755 ( .A1(n13486), .A2(n13485), .A3(n13484), .A4(n13483), .ZN(
        n13492) );
  AOI22_X1 U16756 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13490) );
  AOI22_X1 U16757 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13489) );
  AOI22_X1 U16758 ( .A1(n17248), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17305), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13488) );
  AOI22_X1 U16759 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13487) );
  NAND4_X1 U16760 ( .A1(n13490), .A2(n13489), .A3(n13488), .A4(n13487), .ZN(
        n13491) );
  NOR2_X1 U16761 ( .A1(n13492), .A2(n13491), .ZN(n17113) );
  AOI22_X1 U16762 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17262), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n17284), .ZN(n13496) );
  AOI22_X1 U16763 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17295), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13495) );
  AOI22_X1 U16764 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17277), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13494) );
  AOI22_X1 U16765 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n9758), .ZN(n13493) );
  NAND4_X1 U16766 ( .A1(n13496), .A2(n13495), .A3(n13494), .A4(n13493), .ZN(
        n13502) );
  AOI22_X1 U16767 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17302), .ZN(n13500) );
  AOI22_X1 U16768 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17219), .ZN(n13499) );
  AOI22_X1 U16769 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17305), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17278), .ZN(n13498) );
  AOI22_X1 U16770 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17267), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n17304), .ZN(n13497) );
  NAND4_X1 U16771 ( .A1(n13500), .A2(n13499), .A3(n13498), .A4(n13497), .ZN(
        n13501) );
  NOR2_X1 U16772 ( .A1(n13502), .A2(n13501), .ZN(n17114) );
  NOR2_X1 U16773 ( .A1(n17113), .A2(n17114), .ZN(n17112) );
  AOI22_X1 U16774 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13513) );
  AOI22_X1 U16775 ( .A1(n17248), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13512) );
  AOI22_X1 U16776 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13503) );
  OAI21_X1 U16777 ( .B1(n13504), .B2(n20935), .A(n13503), .ZN(n13510) );
  AOI22_X1 U16778 ( .A1(n17305), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13508) );
  AOI22_X1 U16779 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17294), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13507) );
  AOI22_X1 U16780 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13506) );
  AOI22_X1 U16781 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13505) );
  NAND4_X1 U16782 ( .A1(n13508), .A2(n13507), .A3(n13506), .A4(n13505), .ZN(
        n13509) );
  AOI211_X1 U16783 ( .C1(n9754), .C2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n13510), .B(n13509), .ZN(n13511) );
  NAND3_X1 U16784 ( .A1(n13513), .A2(n13512), .A3(n13511), .ZN(n17108) );
  NAND2_X1 U16785 ( .A1(n17112), .A2(n17108), .ZN(n17107) );
  NOR2_X1 U16786 ( .A1(n17103), .A2(n17107), .ZN(n17102) );
  AOI22_X1 U16787 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17294), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13523) );
  AOI22_X1 U16788 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13522) );
  AOI22_X1 U16789 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13514) );
  OAI21_X1 U16790 ( .B1(n17119), .B2(n20957), .A(n13514), .ZN(n13520) );
  AOI22_X1 U16791 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13518) );
  AOI22_X1 U16792 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13517) );
  AOI22_X1 U16793 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13516) );
  AOI22_X1 U16794 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17305), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13515) );
  NAND4_X1 U16795 ( .A1(n13518), .A2(n13517), .A3(n13516), .A4(n13515), .ZN(
        n13519) );
  AOI211_X1 U16796 ( .C1(n9754), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n13520), .B(n13519), .ZN(n13521) );
  NAND3_X1 U16797 ( .A1(n13523), .A2(n13522), .A3(n13521), .ZN(n17099) );
  NAND2_X1 U16798 ( .A1(n17102), .A2(n17099), .ZN(n17098) );
  NOR2_X1 U16799 ( .A1(n17093), .A2(n17098), .ZN(n17092) );
  AOI22_X1 U16800 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13535) );
  AOI22_X1 U16801 ( .A1(n17305), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13534) );
  AOI22_X1 U16802 ( .A1(n12749), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13524) );
  OAI21_X1 U16803 ( .B1(n13525), .B2(n18337), .A(n13524), .ZN(n13532) );
  AOI22_X1 U16804 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13530) );
  AOI22_X1 U16805 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13529) );
  AOI22_X1 U16806 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13528) );
  AOI22_X1 U16807 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13527) );
  NAND4_X1 U16808 ( .A1(n13530), .A2(n13529), .A3(n13528), .A4(n13527), .ZN(
        n13531) );
  AOI211_X1 U16809 ( .C1(n17296), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n13532), .B(n13531), .ZN(n13533) );
  NAND3_X1 U16810 ( .A1(n13535), .A2(n13534), .A3(n13533), .ZN(n17088) );
  NAND2_X1 U16811 ( .A1(n17092), .A2(n17088), .ZN(n17087) );
  NOR2_X1 U16812 ( .A1(n13536), .A2(n17087), .ZN(n17083) );
  AOI21_X1 U16813 ( .B1(n13536), .B2(n17087), .A(n17083), .ZN(n17357) );
  AOI22_X1 U16814 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17089), .B1(n17357), 
        .B2(n17343), .ZN(n13543) );
  INV_X1 U16815 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n13541) );
  INV_X1 U16816 ( .A(n13537), .ZN(n13539) );
  NAND4_X1 U16817 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n13539), .A4(n13538), .ZN(n14381) );
  INV_X1 U16818 ( .A(n14381), .ZN(n13540) );
  NAND3_X1 U16819 ( .A1(n17143), .A2(n13541), .A3(n13540), .ZN(n13542) );
  NAND2_X1 U16820 ( .A1(n13543), .A2(n13542), .ZN(P3_U2674) );
  INV_X1 U16821 ( .A(n15998), .ZN(n13544) );
  NOR2_X1 U16822 ( .A1(n15150), .A2(n13544), .ZN(n13545) );
  NAND2_X1 U16823 ( .A1(n20228), .A2(n13547), .ZN(n13674) );
  OR2_X1 U16824 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16237), .ZN(n20230) );
  INV_X2 U16825 ( .A(n20230), .ZN(n20847) );
  AOI22_X1 U16826 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20847), .B1(n20239), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13548) );
  OAI21_X1 U16827 ( .B1(n14749), .B2(n13674), .A(n13548), .ZN(P1_U2910) );
  INV_X1 U16828 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13550) );
  AOI22_X1 U16829 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20847), .B1(n20239), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13549) );
  OAI21_X1 U16830 ( .B1(n13550), .B2(n13674), .A(n13549), .ZN(P1_U2912) );
  INV_X1 U16831 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n20882) );
  AOI22_X1 U16832 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20847), .B1(n20239), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13551) );
  OAI21_X1 U16833 ( .B1(n20882), .B2(n13674), .A(n13551), .ZN(P1_U2911) );
  INV_X1 U16834 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13553) );
  AOI22_X1 U16835 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n20239), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20847), .ZN(n13552) );
  OAI21_X1 U16836 ( .B1(n13553), .B2(n13674), .A(n13552), .ZN(P1_U2918) );
  AOI22_X1 U16837 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20847), .B1(n20239), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13554) );
  OAI21_X1 U16838 ( .B1(n14739), .B2(n13674), .A(n13554), .ZN(P1_U2908) );
  INV_X1 U16839 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13556) );
  AOI22_X1 U16840 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20847), .B1(n20239), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13555) );
  OAI21_X1 U16841 ( .B1(n13556), .B2(n13674), .A(n13555), .ZN(P1_U2907) );
  OAI21_X1 U16842 ( .B1(n13558), .B2(n13557), .A(n13653), .ZN(n14083) );
  INV_X1 U16843 ( .A(n13559), .ZN(n13561) );
  NAND2_X1 U16844 ( .A1(n13561), .A2(n13560), .ZN(n13562) );
  NAND2_X1 U16845 ( .A1(n13563), .A2(n13562), .ZN(n13565) );
  NAND2_X1 U16846 ( .A1(n20227), .A2(n14360), .ZN(n14701) );
  XNOR2_X1 U16847 ( .A(n13566), .B(n14540), .ZN(n14078) );
  INV_X1 U16848 ( .A(n14078), .ZN(n13645) );
  AOI22_X1 U16849 ( .A1(n20222), .A2(n13645), .B1(n14716), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13567) );
  OAI21_X1 U16850 ( .B1(n14083), .B2(n14701), .A(n13567), .ZN(P1_U2871) );
  NAND2_X1 U16851 ( .A1(n19173), .A2(n13570), .ZN(n13571) );
  XNOR2_X1 U16852 ( .A(n13867), .B(n13571), .ZN(n13572) );
  NAND2_X1 U16853 ( .A1(n13572), .A2(n19198), .ZN(n13583) );
  NAND2_X1 U16854 ( .A1(n13574), .A2(n13573), .ZN(n13576) );
  INV_X1 U16855 ( .A(n13891), .ZN(n13575) );
  NAND2_X1 U16856 ( .A1(n13576), .A2(n13575), .ZN(n13890) );
  OAI22_X1 U16857 ( .A1(n20858), .A2(n19144), .B1(n19182), .B2(n13890), .ZN(
        n13578) );
  INV_X1 U16858 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19998) );
  NOR2_X1 U16859 ( .A1(n19154), .A2(n19998), .ZN(n13577) );
  AOI211_X1 U16860 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n19167), .A(n13578), .B(
        n13577), .ZN(n13579) );
  OAI21_X1 U16861 ( .B1(n13580), .B2(n19169), .A(n13579), .ZN(n13581) );
  AOI21_X1 U16862 ( .B1(n15861), .B2(n19187), .A(n13581), .ZN(n13582) );
  OAI211_X1 U16863 ( .C1(n15893), .C2(n13729), .A(n13583), .B(n13582), .ZN(
        P2_U2852) );
  MUX2_X1 U16864 ( .A(n10394), .B(n13588), .S(n15319), .Z(n13589) );
  OAI21_X1 U16865 ( .B1(n20072), .B2(n15337), .A(n13589), .ZN(P2_U2885) );
  MUX2_X1 U16866 ( .A(n13590), .B(n11084), .S(n15319), .Z(n13591) );
  OAI21_X1 U16867 ( .B1(n15893), .B2(n15337), .A(n13591), .ZN(P2_U2884) );
  OAI21_X1 U16868 ( .B1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B2(
        P2_STATE2_REG_3__SCAN_IN), .A(n13592), .ZN(n13594) );
  AND2_X1 U16869 ( .A1(n13594), .A2(n13593), .ZN(n13595) );
  MUX2_X1 U16870 ( .A(n19200), .B(n11203), .S(n9778), .Z(n13597) );
  OAI21_X1 U16871 ( .B1(n20086), .B2(n15337), .A(n13597), .ZN(P2_U2887) );
  OR2_X1 U16872 ( .A1(n13600), .A2(n13599), .ZN(n13601) );
  MUX2_X1 U16873 ( .A(n13724), .B(n13602), .S(n15319), .Z(n13603) );
  OAI21_X1 U16874 ( .B1(n19407), .B2(n15337), .A(n13603), .ZN(P2_U2886) );
  AND2_X1 U16875 ( .A1(n13604), .A2(n20732), .ZN(n13605) );
  OR2_X1 U16876 ( .A1(n20257), .A2(n14042), .ZN(n13793) );
  INV_X1 U16877 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14338) );
  NOR2_X2 U16878 ( .A1(n20257), .A2(n14138), .ZN(n20269) );
  INV_X1 U16879 ( .A(n20269), .ZN(n13608) );
  INV_X1 U16880 ( .A(DATAI_15_), .ZN(n13607) );
  INV_X1 U16881 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13606) );
  MUX2_X1 U16882 ( .A(n13607), .B(n13606), .S(n14327), .Z(n14336) );
  INV_X1 U16883 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20231) );
  OAI222_X1 U16884 ( .A1(n13793), .A2(n14338), .B1(n13608), .B2(n14336), .C1(
        n13802), .C2(n20231), .ZN(P1_U2967) );
  INV_X1 U16885 ( .A(n13609), .ZN(n13612) );
  OAI21_X1 U16886 ( .B1(n13612), .B2(n13611), .A(n13610), .ZN(n14090) );
  INV_X1 U16887 ( .A(n13613), .ZN(n13615) );
  AOI21_X1 U16888 ( .B1(n13615), .B2(n13642), .A(n13614), .ZN(n13753) );
  AND2_X1 U16889 ( .A1(n20299), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13757) );
  INV_X1 U16890 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13616) );
  AOI21_X1 U16891 ( .B1(n14950), .B2(n13617), .A(n13616), .ZN(n13618) );
  AOI211_X1 U16892 ( .C1(n13753), .C2(n20294), .A(n13757), .B(n13618), .ZN(
        n13619) );
  OAI21_X1 U16893 ( .B1(n14954), .B2(n14090), .A(n13619), .ZN(P1_U2999) );
  NAND2_X1 U16894 ( .A1(n13620), .A2(n14507), .ZN(n13622) );
  INV_X1 U16895 ( .A(n13637), .ZN(n13621) );
  NAND2_X1 U16896 ( .A1(n13622), .A2(n13621), .ZN(n19165) );
  NOR2_X1 U16897 ( .A1(n14505), .A2(n10538), .ZN(n13624) );
  OAI211_X1 U16898 ( .C1(n13624), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15341), .B(n13623), .ZN(n13626) );
  NAND2_X1 U16899 ( .A1(n15344), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13625) );
  OAI211_X1 U16900 ( .C1(n19165), .C2(n9778), .A(n13626), .B(n13625), .ZN(
        P2_U2881) );
  NOR2_X1 U16901 ( .A1(n10058), .A2(n13714), .ZN(n13628) );
  XNOR2_X1 U16902 ( .A(n13628), .B(n13627), .ZN(n13629) );
  NAND2_X1 U16903 ( .A1(n13629), .A2(n19198), .ZN(n13636) );
  OAI22_X1 U16904 ( .A1(n19207), .A2(n10394), .B1(n13889), .B2(n19182), .ZN(
        n13631) );
  INV_X1 U16905 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19996) );
  NOR2_X1 U16906 ( .A1(n19154), .A2(n19996), .ZN(n13630) );
  AOI211_X1 U16907 ( .C1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .C2(n19211), .A(
        n13631), .B(n13630), .ZN(n13632) );
  OAI21_X1 U16908 ( .B1(n13633), .B2(n19169), .A(n13632), .ZN(n13634) );
  AOI21_X1 U16909 ( .B1(n15847), .B2(n19187), .A(n13634), .ZN(n13635) );
  OAI211_X1 U16910 ( .C1(n13729), .C2(n20072), .A(n13636), .B(n13635), .ZN(
        P2_U2853) );
  XOR2_X1 U16911 ( .A(n13623), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13641)
         );
  OR2_X1 U16912 ( .A1(n13638), .A2(n13637), .ZN(n13639) );
  NAND2_X1 U16913 ( .A1(n13639), .A2(n13761), .ZN(n19153) );
  MUX2_X1 U16914 ( .A(n19153), .B(n11555), .S(n9778), .Z(n13640) );
  OAI21_X1 U16915 ( .B1(n13641), .B2(n15337), .A(n13640), .ZN(P2_U2880) );
  INV_X1 U16916 ( .A(n20314), .ZN(n15129) );
  AOI21_X1 U16917 ( .B1(n15129), .B2(n13642), .A(n15073), .ZN(n13754) );
  NAND2_X1 U16918 ( .A1(n20299), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n13738) );
  OAI21_X1 U16919 ( .B1(n13754), .B2(n9923), .A(n13738), .ZN(n13644) );
  AOI211_X1 U16920 ( .C1(n13642), .C2(n16175), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n15100), .ZN(n13643) );
  AOI211_X1 U16921 ( .C1(n13645), .C2(n20312), .A(n13644), .B(n13643), .ZN(
        n13649) );
  OR2_X1 U16922 ( .A1(n13646), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13740) );
  NAND3_X1 U16923 ( .A1(n13740), .A2(n13647), .A3(n20318), .ZN(n13648) );
  NAND2_X1 U16924 ( .A1(n13649), .A2(n13648), .ZN(P1_U3030) );
  NOR2_X1 U16925 ( .A1(n13651), .A2(n13650), .ZN(n13652) );
  OR2_X1 U16926 ( .A1(n13775), .A2(n13652), .ZN(n20308) );
  INV_X1 U16927 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13657) );
  NAND2_X1 U16928 ( .A1(n13654), .A2(n13653), .ZN(n13655) );
  AND2_X1 U16929 ( .A1(n13656), .A2(n13655), .ZN(n14039) );
  INV_X1 U16930 ( .A(n14039), .ZN(n13930) );
  OAI222_X1 U16931 ( .A1(n20308), .A2(n14725), .B1(n20227), .B2(n13657), .C1(
        n13930), .C2(n14730), .ZN(P1_U2870) );
  INV_X1 U16932 ( .A(n13658), .ZN(n13660) );
  OR2_X1 U16933 ( .A1(n9773), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13659) );
  NAND2_X1 U16934 ( .A1(n13660), .A2(n13659), .ZN(n14085) );
  OAI222_X1 U16935 ( .A1(n14085), .A2(n14725), .B1(n13002), .B2(n20227), .C1(
        n14090), .C2(n14730), .ZN(P1_U2872) );
  AOI22_X1 U16936 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13661) );
  OAI21_X1 U16937 ( .B1(n14761), .B2(n13674), .A(n13661), .ZN(P1_U2913) );
  INV_X1 U16938 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13663) );
  AOI22_X1 U16939 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13662) );
  OAI21_X1 U16940 ( .B1(n13663), .B2(n13674), .A(n13662), .ZN(P1_U2920) );
  INV_X1 U16941 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13665) );
  AOI22_X1 U16942 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13664) );
  OAI21_X1 U16943 ( .B1(n13665), .B2(n13674), .A(n13664), .ZN(P1_U2916) );
  INV_X1 U16944 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13667) );
  AOI22_X1 U16945 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13666) );
  OAI21_X1 U16946 ( .B1(n13667), .B2(n13674), .A(n13666), .ZN(P1_U2915) );
  INV_X1 U16947 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14782) );
  AOI22_X1 U16948 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13668) );
  OAI21_X1 U16949 ( .B1(n14782), .B2(n13674), .A(n13668), .ZN(P1_U2917) );
  AOI22_X1 U16950 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13669) );
  OAI21_X1 U16951 ( .B1(n14744), .B2(n13674), .A(n13669), .ZN(P1_U2909) );
  AOI22_X1 U16952 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13670) );
  OAI21_X1 U16953 ( .B1(n14731), .B2(n13674), .A(n13670), .ZN(P1_U2906) );
  INV_X1 U16954 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13672) );
  AOI22_X1 U16955 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13671) );
  OAI21_X1 U16956 ( .B1(n13672), .B2(n13674), .A(n13671), .ZN(P1_U2914) );
  AOI22_X1 U16957 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13673) );
  OAI21_X1 U16958 ( .B1(n14797), .B2(n13674), .A(n13673), .ZN(P1_U2919) );
  NOR2_X1 U16959 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20727), .ZN(n13696) );
  INV_X1 U16960 ( .A(n13694), .ZN(n15972) );
  INV_X1 U16961 ( .A(n13901), .ZN(n13968) );
  OR2_X1 U16962 ( .A1(n11931), .A2(n13968), .ZN(n13675) );
  XNOR2_X1 U16963 ( .A(n13675), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20212) );
  INV_X1 U16964 ( .A(n13211), .ZN(n13676) );
  AND2_X1 U16965 ( .A1(n20212), .A2(n13676), .ZN(n16225) );
  OAI21_X1 U16966 ( .B1(n16225), .B2(n15972), .A(n20727), .ZN(n13677) );
  AOI21_X1 U16967 ( .B1(n15972), .B2(n16226), .A(n13677), .ZN(n13678) );
  AOI21_X1 U16968 ( .B1(n13696), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13678), .ZN(n15992) );
  NAND2_X1 U16969 ( .A1(n20815), .A2(n15155), .ZN(n13691) );
  XNOR2_X1 U16970 ( .A(n13679), .B(n11656), .ZN(n13683) );
  NAND2_X1 U16971 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13680) );
  AOI22_X1 U16972 ( .A1(n13681), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n11656), .B2(n13680), .ZN(n13682) );
  AOI22_X1 U16973 ( .A1(n13684), .A2(n13683), .B1(n15150), .B2(n13682), .ZN(
        n13689) );
  NAND2_X1 U16974 ( .A1(n13685), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13686) );
  NAND2_X1 U16975 ( .A1(n11866), .A2(n13686), .ZN(n20802) );
  NAND3_X1 U16976 ( .A1(n14499), .A2(n13687), .A3(n20802), .ZN(n13688) );
  AND2_X1 U16977 ( .A1(n13689), .A2(n13688), .ZN(n13690) );
  NAND2_X1 U16978 ( .A1(n13691), .A2(n13690), .ZN(n20805) );
  NAND2_X1 U16979 ( .A1(n20805), .A2(n13694), .ZN(n13693) );
  OR2_X1 U16980 ( .A1(n13694), .A2(n11656), .ZN(n13692) );
  NAND2_X1 U16981 ( .A1(n13693), .A2(n13692), .ZN(n15979) );
  NAND2_X1 U16982 ( .A1(n15979), .A2(n20727), .ZN(n13699) );
  NAND2_X1 U16983 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13696), .ZN(
        n13698) );
  MUX2_X1 U16984 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13695), .S(
        n13694), .Z(n15974) );
  AOI22_X1 U16985 ( .A1(n13696), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15974), .B2(n20727), .ZN(n13697) );
  AOI21_X1 U16986 ( .B1(n13699), .B2(n13698), .A(n13697), .ZN(n15989) );
  INV_X1 U16987 ( .A(n13700), .ZN(n15152) );
  NAND2_X1 U16988 ( .A1(n15989), .A2(n15152), .ZN(n13701) );
  NAND2_X1 U16989 ( .A1(n15992), .A2(n13701), .ZN(n13735) );
  OAI21_X1 U16990 ( .B1(n13735), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13702), .ZN(
        n13703) );
  NOR2_X1 U16991 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16229) );
  NAND2_X1 U16992 ( .A1(n13703), .A2(n15174), .ZN(n20823) );
  NOR2_X1 U16993 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20727), .ZN(n20813) );
  AOI21_X1 U16994 ( .B1(n15166), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20667), 
        .ZN(n20598) );
  OAI21_X1 U16995 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15166), .A(n20598), 
        .ZN(n13705) );
  OAI21_X1 U16996 ( .B1(n20813), .B2(n20518), .A(n13705), .ZN(n13706) );
  NAND2_X1 U16997 ( .A1(n20823), .A2(n13706), .ZN(n13707) );
  OAI21_X1 U16998 ( .B1(n20823), .B2(n20517), .A(n13707), .ZN(P1_U3477) );
  OAI21_X1 U16999 ( .B1(n13708), .B2(n13710), .A(n13709), .ZN(n20316) );
  NAND2_X1 U17000 ( .A1(n20299), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n20309) );
  NAND2_X1 U17001 ( .A1(n20287), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13711) );
  OAI211_X1 U17002 ( .C1(n20298), .C2(n14062), .A(n20309), .B(n13711), .ZN(
        n13712) );
  AOI21_X1 U17003 ( .B1(n14039), .B2(n20293), .A(n13712), .ZN(n13713) );
  OAI21_X1 U17004 ( .B1(n20139), .B2(n20316), .A(n13713), .ZN(P1_U2997) );
  AOI211_X1 U17005 ( .C1(n19197), .C2(n13715), .A(n10058), .B(n13714), .ZN(
        n13830) );
  NOR2_X1 U17006 ( .A1(n19972), .A2(n19173), .ZN(n19107) );
  AOI22_X1 U17007 ( .A1(n13830), .A2(n19198), .B1(n19107), .B2(n13402), .ZN(
        n13728) );
  INV_X1 U17008 ( .A(n13716), .ZN(n13719) );
  INV_X1 U17009 ( .A(n13717), .ZN(n13718) );
  NAND2_X1 U17010 ( .A1(n13719), .A2(n13718), .ZN(n13720) );
  NAND2_X1 U17011 ( .A1(n13721), .A2(n13720), .ZN(n20083) );
  INV_X1 U17012 ( .A(n20083), .ZN(n13888) );
  OAI22_X1 U17013 ( .A1(n13888), .A2(n19182), .B1(n13722), .B2(n19169), .ZN(
        n13726) );
  AOI22_X1 U17014 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19166), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n19204), .ZN(n13723) );
  OAI21_X1 U17015 ( .B1(n19207), .B2(n13724), .A(n13723), .ZN(n13725) );
  AOI211_X1 U17016 ( .C1(n19187), .C2(n11087), .A(n13726), .B(n13725), .ZN(
        n13727) );
  OAI211_X1 U17017 ( .C1(n19407), .C2(n13729), .A(n13728), .B(n13727), .ZN(
        P2_U2854) );
  NOR2_X1 U17018 ( .A1(n13415), .A2(n20813), .ZN(n13733) );
  INV_X1 U17019 ( .A(n13730), .ZN(n20810) );
  AND2_X1 U17020 ( .A1(n15166), .A2(n20810), .ZN(n20816) );
  MUX2_X1 U17021 ( .A(n20598), .B(n20816), .S(n13731), .Z(n13732) );
  OAI21_X1 U17022 ( .B1(n13733), .B2(n13732), .A(n20823), .ZN(n13734) );
  OAI21_X1 U17023 ( .B1(n12111), .B2(n20823), .A(n13734), .ZN(P1_U3476) );
  NOR2_X1 U17024 ( .A1(n13735), .A2(n16237), .ZN(n15999) );
  INV_X1 U17025 ( .A(n12159), .ZN(n20393) );
  OAI22_X1 U17026 ( .A1(n15167), .A2(n20667), .B1(n20393), .B2(n20813), .ZN(
        n13736) );
  OAI21_X1 U17027 ( .B1(n15999), .B2(n13736), .A(n20823), .ZN(n13737) );
  OAI21_X1 U17028 ( .B1(n20823), .B2(n20547), .A(n13737), .ZN(P1_U3478) );
  OAI21_X1 U17029 ( .B1(n14950), .B2(n14081), .A(n13738), .ZN(n13739) );
  AOI21_X1 U17030 ( .B1(n16141), .B2(n14081), .A(n13739), .ZN(n13742) );
  NAND3_X1 U17031 ( .A1(n13740), .A2(n13647), .A3(n20294), .ZN(n13741) );
  OAI211_X1 U17032 ( .C1(n14083), .C2(n14954), .A(n13742), .B(n13741), .ZN(
        P1_U2998) );
  OR2_X1 U17033 ( .A1(n19200), .A2(n13832), .ZN(n13748) );
  NAND2_X1 U17034 ( .A1(n9896), .A2(n13744), .ZN(n13836) );
  MUX2_X1 U17035 ( .A(n10381), .B(n13836), .S(n13745), .Z(n13746) );
  INV_X1 U17036 ( .A(n13746), .ZN(n13747) );
  NAND2_X1 U17037 ( .A1(n13748), .A2(n13747), .ZN(n16461) );
  OAI22_X1 U17038 ( .A1(n19173), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19197), .B2(n10058), .ZN(n13831) );
  AOI222_X1 U17039 ( .A1(n16461), .A2(n13840), .B1(n13750), .B2(n15835), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n13831), .ZN(n13752) );
  NAND2_X1 U17040 ( .A1(n15862), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13751) );
  OAI21_X1 U17041 ( .B1(n13752), .B2(n15862), .A(n13751), .ZN(P2_U3601) );
  INV_X1 U17042 ( .A(n13753), .ZN(n13760) );
  INV_X1 U17043 ( .A(n14085), .ZN(n13758) );
  NOR2_X1 U17044 ( .A1(n15129), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13755) );
  AOI22_X1 U17045 ( .A1(n13755), .A2(n15050), .B1(n13754), .B2(n16175), .ZN(
        n13756) );
  AOI211_X1 U17046 ( .C1(n13758), .C2(n20312), .A(n13757), .B(n13756), .ZN(
        n13759) );
  OAI21_X1 U17047 ( .B1(n15137), .B2(n13760), .A(n13759), .ZN(P1_U3031) );
  NAND2_X1 U17048 ( .A1(n13762), .A2(n13761), .ZN(n13764) );
  AND2_X1 U17049 ( .A1(n13764), .A2(n10097), .ZN(n19139) );
  INV_X1 U17050 ( .A(n19139), .ZN(n13770) );
  OAI211_X1 U17051 ( .C1(n13767), .C2(n13766), .A(n13765), .B(n15341), .ZN(
        n13769) );
  NAND2_X1 U17052 ( .A1(n15344), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13768) );
  OAI211_X1 U17053 ( .C1(n13770), .C2(n15344), .A(n13769), .B(n13768), .ZN(
        P2_U2879) );
  OR2_X1 U17054 ( .A1(n13772), .A2(n13771), .ZN(n13773) );
  NAND2_X1 U17055 ( .A1(n13823), .A2(n13773), .ZN(n14075) );
  INV_X1 U17056 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13777) );
  OR2_X1 U17057 ( .A1(n13775), .A2(n13774), .ZN(n13776) );
  NAND2_X1 U17058 ( .A1(n13827), .A2(n13776), .ZN(n14070) );
  OAI222_X1 U17059 ( .A1(n14075), .A2(n14701), .B1(n20227), .B2(n13777), .C1(
        n14070), .C2(n14725), .ZN(P1_U2869) );
  XNOR2_X1 U17060 ( .A(n13765), .B(n13778), .ZN(n13783) );
  NOR2_X1 U17061 ( .A1(n13780), .A2(n13763), .ZN(n13781) );
  OR2_X1 U17062 ( .A1(n13779), .A2(n13781), .ZN(n19131) );
  MUX2_X1 U17063 ( .A(n19131), .B(n11564), .S(n9778), .Z(n13782) );
  OAI21_X1 U17064 ( .B1(n13783), .B2(n15337), .A(n13782), .ZN(P2_U2878) );
  OAI21_X1 U17065 ( .B1(n13784), .B2(n13786), .A(n13785), .ZN(n13814) );
  NAND2_X1 U17066 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13787) );
  INV_X1 U17067 ( .A(n20321), .ZN(n15018) );
  OAI22_X1 U17068 ( .A1(n13790), .A2(n20314), .B1(n13787), .B2(n15018), .ZN(
        n20304) );
  INV_X1 U17069 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20749) );
  OAI22_X1 U17070 ( .A1(n16218), .A2(n14070), .B1(n20749), .B2(n20207), .ZN(
        n13788) );
  AOI21_X1 U17071 ( .B1(n20304), .B2(n13789), .A(n13788), .ZN(n13792) );
  INV_X1 U17072 ( .A(n15124), .ZN(n14311) );
  AOI21_X1 U17073 ( .B1(n9923), .B2(n14311), .A(n15073), .ZN(n20313) );
  NAND2_X1 U17074 ( .A1(n15129), .A2(n13790), .ZN(n20323) );
  OAI211_X1 U17075 ( .C1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n15124), .A(
        n20313), .B(n20323), .ZN(n20301) );
  NAND2_X1 U17076 ( .A1(n20301), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13791) );
  OAI211_X1 U17077 ( .C1(n13814), .C2(n15137), .A(n13792), .B(n13791), .ZN(
        P1_U3028) );
  AOI22_X1 U17078 ( .A1(n20281), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20284), .ZN(n13797) );
  NAND2_X1 U17079 ( .A1(n13927), .A2(DATAI_4_), .ZN(n13795) );
  NAND2_X1 U17080 ( .A1(n14327), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13794) );
  AND2_X1 U17081 ( .A1(n13795), .A2(n13794), .ZN(n14777) );
  INV_X1 U17082 ( .A(n14777), .ZN(n13796) );
  NAND2_X1 U17083 ( .A1(n20269), .A2(n13796), .ZN(n14217) );
  NAND2_X1 U17084 ( .A1(n13797), .A2(n14217), .ZN(P1_U2956) );
  AOI22_X1 U17085 ( .A1(n20281), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20284), .ZN(n13801) );
  NAND2_X1 U17086 ( .A1(n13927), .A2(DATAI_6_), .ZN(n13799) );
  NAND2_X1 U17087 ( .A1(n14327), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13798) );
  AND2_X1 U17088 ( .A1(n13799), .A2(n13798), .ZN(n14767) );
  INV_X1 U17089 ( .A(n14767), .ZN(n13800) );
  NAND2_X1 U17090 ( .A1(n20269), .A2(n13800), .ZN(n14211) );
  NAND2_X1 U17091 ( .A1(n13801), .A2(n14211), .ZN(P1_U2958) );
  INV_X1 U17092 ( .A(n13802), .ZN(n20284) );
  AOI22_X1 U17093 ( .A1(n20281), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20284), .ZN(n13805) );
  NAND2_X1 U17094 ( .A1(n14327), .A2(n16607), .ZN(n13803) );
  OAI21_X1 U17095 ( .B1(n14327), .B2(DATAI_7_), .A(n13803), .ZN(n14763) );
  INV_X1 U17096 ( .A(n14763), .ZN(n13804) );
  NAND2_X1 U17097 ( .A1(n20269), .A2(n13804), .ZN(n14205) );
  NAND2_X1 U17098 ( .A1(n13805), .A2(n14205), .ZN(P1_U2959) );
  AOI22_X1 U17099 ( .A1(n20281), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20284), .ZN(n13809) );
  NAND2_X1 U17100 ( .A1(n13927), .A2(DATAI_5_), .ZN(n13807) );
  NAND2_X1 U17101 ( .A1(n14327), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13806) );
  AND2_X1 U17102 ( .A1(n13807), .A2(n13806), .ZN(n14772) );
  INV_X1 U17103 ( .A(n14772), .ZN(n13808) );
  NAND2_X1 U17104 ( .A1(n20269), .A2(n13808), .ZN(n14213) );
  NAND2_X1 U17105 ( .A1(n13809), .A2(n14213), .ZN(P1_U2957) );
  INV_X1 U17106 ( .A(n14075), .ZN(n13812) );
  AOI22_X1 U17107 ( .A1(n20287), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20299), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n13810) );
  OAI21_X1 U17108 ( .B1(n20298), .B2(n14071), .A(n13810), .ZN(n13811) );
  AOI21_X1 U17109 ( .B1(n13812), .B2(n20293), .A(n13811), .ZN(n13813) );
  OAI21_X1 U17110 ( .B1(n13814), .B2(n20139), .A(n13813), .ZN(P1_U2996) );
  NOR2_X1 U17111 ( .A1(n13816), .A2(n13817), .ZN(n13818) );
  OR2_X1 U17112 ( .A1(n13815), .A2(n13818), .ZN(n16162) );
  NAND2_X1 U17113 ( .A1(n13825), .A2(n13819), .ZN(n13820) );
  NAND2_X1 U17114 ( .A1(n16207), .A2(n13820), .ZN(n20190) );
  INV_X1 U17115 ( .A(n20190), .ZN(n13821) );
  AOI22_X1 U17116 ( .A1(n20222), .A2(n13821), .B1(n14716), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n13822) );
  OAI21_X1 U17117 ( .B1(n16162), .B2(n14701), .A(n13822), .ZN(P1_U2867) );
  XOR2_X1 U17118 ( .A(n13824), .B(n13823), .Z(n20292) );
  INV_X1 U17119 ( .A(n20292), .ZN(n14228) );
  INV_X1 U17120 ( .A(n13825), .ZN(n13826) );
  AOI21_X1 U17121 ( .B1(n13828), .B2(n13827), .A(n13826), .ZN(n20300) );
  AOI22_X1 U17122 ( .A1(n20222), .A2(n20300), .B1(n14716), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n13829) );
  OAI21_X1 U17123 ( .B1(n14228), .B2(n14701), .A(n13829), .ZN(P1_U2868) );
  AOI21_X1 U17124 ( .B1(n10058), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n13830), .ZN(n15849) );
  NOR2_X1 U17125 ( .A1(n13298), .A2(n13831), .ZN(n15836) );
  INV_X1 U17126 ( .A(n13832), .ZN(n15860) );
  NAND2_X1 U17127 ( .A1(n11087), .A2(n15860), .ZN(n13839) );
  NOR2_X1 U17128 ( .A1(n13833), .A2(n13834), .ZN(n13835) );
  AOI22_X1 U17129 ( .A1(n13837), .A2(n10381), .B1(n13836), .B2(n13835), .ZN(
        n13838) );
  NAND2_X1 U17130 ( .A1(n13839), .A2(n13838), .ZN(n16465) );
  AOI222_X1 U17131 ( .A1(n20079), .A2(n15835), .B1(n15849), .B2(n15836), .C1(
        n16465), .C2(n13840), .ZN(n13842) );
  NAND2_X1 U17132 ( .A1(n15862), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13841) );
  OAI21_X1 U17133 ( .B1(n13842), .B2(n15862), .A(n13841), .ZN(P2_U3600) );
  NAND3_X1 U17134 ( .A1(n20825), .A2(n12111), .A3(n20517), .ZN(n20328) );
  INV_X1 U17135 ( .A(n20328), .ZN(n13845) );
  INV_X1 U17136 ( .A(n20391), .ZN(n20394) );
  INV_X1 U17137 ( .A(n13843), .ZN(n20548) );
  NOR2_X1 U17138 ( .A1(n20547), .A2(n20328), .ZN(n20366) );
  AOI21_X1 U17139 ( .B1(n9847), .B2(n20548), .A(n20366), .ZN(n13848) );
  OAI211_X1 U17140 ( .C1(n20394), .C2(n20840), .A(n13848), .B(n20809), .ZN(
        n13844) );
  OAI211_X1 U17141 ( .C1(n13845), .C2(n20809), .A(n13844), .B(n20673), .ZN(
        n20369) );
  INV_X1 U17142 ( .A(n20369), .ZN(n13860) );
  INV_X1 U17143 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13853) );
  INV_X1 U17144 ( .A(n20372), .ZN(n13857) );
  NOR2_X2 U17145 ( .A1(n14954), .A2(n13927), .ZN(n15176) );
  NOR2_X2 U17146 ( .A1(n14327), .A2(n14954), .ZN(n15177) );
  AOI22_X1 U17147 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n15176), .B1(DATAI_26_), 
        .B2(n15177), .ZN(n20691) );
  INV_X1 U17148 ( .A(n20691), .ZN(n20651) );
  NOR2_X1 U17149 ( .A1(n15166), .A2(n15167), .ZN(n13948) );
  NAND2_X1 U17150 ( .A1(n13927), .A2(DATAI_2_), .ZN(n13847) );
  NAND2_X1 U17151 ( .A1(n14327), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13846) );
  AND2_X1 U17152 ( .A1(n13847), .A2(n13846), .ZN(n14195) );
  NOR2_X2 U17153 ( .A1(n14195), .A2(n15174), .ZN(n20687) );
  OAI22_X1 U17154 ( .A1(n13848), .A2(n20667), .B1(n20328), .B2(n20839), .ZN(
        n20367) );
  NOR2_X2 U17155 ( .A1(n15178), .A2(n12981), .ZN(n20686) );
  AOI22_X1 U17156 ( .A1(n20687), .A2(n20367), .B1(n20686), .B2(n20366), .ZN(
        n13850) );
  OAI21_X1 U17157 ( .B1(n20654), .B2(n20385), .A(n13850), .ZN(n13851) );
  AOI21_X1 U17158 ( .B1(n13857), .B2(n20651), .A(n13851), .ZN(n13852) );
  OAI21_X1 U17159 ( .B1(n13860), .B2(n13853), .A(n13852), .ZN(P1_U3043) );
  INV_X1 U17160 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13859) );
  AOI22_X1 U17161 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n15176), .B1(DATAI_31_), 
        .B2(n15177), .ZN(n20726) );
  INV_X1 U17162 ( .A(n20726), .ZN(n20587) );
  AOI22_X1 U17163 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n15176), .B1(DATAI_23_), 
        .B2(n15177), .ZN(n20593) );
  NOR2_X2 U17164 ( .A1(n14763), .A2(n15174), .ZN(n20719) );
  NOR2_X2 U17165 ( .A1(n15178), .A2(n13854), .ZN(n20716) );
  AOI22_X1 U17166 ( .A1(n20719), .A2(n20367), .B1(n20716), .B2(n20366), .ZN(
        n13855) );
  OAI21_X1 U17167 ( .B1(n20593), .B2(n20385), .A(n13855), .ZN(n13856) );
  AOI21_X1 U17168 ( .B1(n13857), .B2(n20587), .A(n13856), .ZN(n13858) );
  OAI21_X1 U17169 ( .B1(n13860), .B2(n13859), .A(n13858), .ZN(P1_U3048) );
  NAND2_X1 U17170 ( .A1(n13862), .A2(n13861), .ZN(n13864) );
  XNOR2_X1 U17171 ( .A(n13864), .B(n13863), .ZN(n13882) );
  NOR2_X1 U17172 ( .A1(n13196), .A2(n19998), .ZN(n13876) );
  NOR2_X1 U17173 ( .A1(n16382), .A2(n20858), .ZN(n13866) );
  AOI211_X1 U17174 ( .C1(n13867), .C2(n16370), .A(n13876), .B(n13866), .ZN(
        n13868) );
  OAI21_X1 U17175 ( .B1(n11084), .B2(n14529), .A(n13868), .ZN(n13869) );
  AOI21_X1 U17176 ( .B1(n13880), .B2(n16378), .A(n13869), .ZN(n13870) );
  OAI21_X1 U17177 ( .B1(n13882), .B2(n9780), .A(n13870), .ZN(P2_U3011) );
  NAND2_X1 U17178 ( .A1(n13873), .A2(n15815), .ZN(n13874) );
  NOR2_X1 U17179 ( .A1(n13872), .A2(n13871), .ZN(n14004) );
  OAI22_X1 U17180 ( .A1(n13875), .A2(n13874), .B1(n14004), .B2(n13873), .ZN(
        n13879) );
  INV_X1 U17181 ( .A(n13890), .ZN(n20065) );
  AOI21_X1 U17182 ( .B1(n19391), .B2(n20065), .A(n13876), .ZN(n13877) );
  OAI21_X1 U17183 ( .B1(n11084), .B2(n16411), .A(n13877), .ZN(n13878) );
  AOI211_X1 U17184 ( .C1(n13880), .C2(n16450), .A(n13879), .B(n13878), .ZN(
        n13881) );
  OAI21_X1 U17185 ( .B1(n13882), .B2(n19395), .A(n13881), .ZN(P2_U3043) );
  INV_X1 U17186 ( .A(n13884), .ZN(n13885) );
  NAND2_X1 U17187 ( .A1(n13883), .A2(n13885), .ZN(n13886) );
  OAI21_X1 U17188 ( .B1(n13887), .B2(n13886), .A(n14505), .ZN(n19186) );
  XNOR2_X1 U17189 ( .A(n20079), .B(n20083), .ZN(n19265) );
  AND2_X1 U17190 ( .A1(n19274), .A2(n19273), .ZN(n19277) );
  NOR2_X1 U17191 ( .A1(n19265), .A2(n19277), .ZN(n19264) );
  AOI21_X1 U17192 ( .B1(n13888), .B2(n19407), .A(n19264), .ZN(n19257) );
  XNOR2_X1 U17193 ( .A(n20072), .B(n13889), .ZN(n19258) );
  NOR2_X1 U17194 ( .A1(n19257), .A2(n19258), .ZN(n19256) );
  AOI21_X1 U17195 ( .B1(n13889), .B2(n20072), .A(n19256), .ZN(n19251) );
  XNOR2_X1 U17196 ( .A(n15893), .B(n13890), .ZN(n19252) );
  NOR2_X1 U17197 ( .A1(n19251), .A2(n19252), .ZN(n19250) );
  INV_X1 U17198 ( .A(n15893), .ZN(n20066) );
  NOR2_X1 U17199 ( .A1(n20066), .A2(n20065), .ZN(n13894) );
  OR2_X1 U17200 ( .A1(n13892), .A2(n13891), .ZN(n13893) );
  NAND2_X1 U17201 ( .A1(n13893), .A2(n16445), .ZN(n19181) );
  OAI21_X1 U17202 ( .B1(n19250), .B2(n13894), .A(n19181), .ZN(n19247) );
  XOR2_X1 U17203 ( .A(n19186), .B(n19247), .Z(n13900) );
  INV_X1 U17204 ( .A(n19181), .ZN(n13895) );
  AOI22_X1 U17205 ( .A1(n19263), .A2(n13895), .B1(n19262), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n13899) );
  INV_X1 U17206 ( .A(n16315), .ZN(n15402) );
  INV_X1 U17207 ( .A(n13896), .ZN(n13897) );
  NAND2_X1 U17208 ( .A1(n15402), .A2(n13897), .ZN(n19280) );
  NAND2_X1 U17209 ( .A1(n19280), .A2(n19436), .ZN(n13898) );
  OAI211_X1 U17210 ( .C1(n13900), .C2(n19275), .A(n13899), .B(n13898), .ZN(
        P2_U2915) );
  NAND3_X1 U17211 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20825), .A3(
        n20517), .ZN(n20434) );
  INV_X1 U17212 ( .A(n20434), .ZN(n13903) );
  NOR2_X1 U17213 ( .A1(n13415), .A2(n13901), .ZN(n20487) );
  NOR2_X1 U17214 ( .A1(n20547), .A2(n20434), .ZN(n20468) );
  AOI21_X1 U17215 ( .B1(n20487), .B2(n20548), .A(n20468), .ZN(n13906) );
  OAI211_X1 U17216 ( .C1(n14161), .C2(n20840), .A(n13906), .B(n20809), .ZN(
        n13902) );
  OAI211_X1 U17217 ( .C1(n13903), .C2(n20809), .A(n20673), .B(n13902), .ZN(
        n20470) );
  INV_X1 U17218 ( .A(n20470), .ZN(n13999) );
  INV_X1 U17219 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13910) );
  INV_X1 U17220 ( .A(n20516), .ZN(n13904) );
  INV_X1 U17221 ( .A(n13948), .ZN(n13905) );
  INV_X1 U17222 ( .A(n20481), .ZN(n14184) );
  OAI22_X1 U17223 ( .A1(n13906), .A2(n20667), .B1(n20434), .B2(n20839), .ZN(
        n20469) );
  AOI22_X1 U17224 ( .A1(n20687), .A2(n20469), .B1(n20686), .B2(n20468), .ZN(
        n13907) );
  OAI21_X1 U17225 ( .B1(n20654), .B2(n14184), .A(n13907), .ZN(n13908) );
  AOI21_X1 U17226 ( .B1(n20457), .B2(n20651), .A(n13908), .ZN(n13909) );
  OAI21_X1 U17227 ( .B1(n13999), .B2(n13910), .A(n13909), .ZN(P1_U3075) );
  INV_X1 U17228 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13914) );
  AOI22_X1 U17229 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n15176), .B1(DATAI_29_), 
        .B2(n15177), .ZN(n20709) );
  INV_X1 U17230 ( .A(n20709), .ZN(n20614) );
  AOI22_X1 U17231 ( .A1(DATAI_21_), .A2(n15177), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n15176), .ZN(n20617) );
  NOR2_X2 U17232 ( .A1(n14772), .A2(n15174), .ZN(n20705) );
  NOR2_X2 U17233 ( .A1(n15178), .A2(n12083), .ZN(n20704) );
  AOI22_X1 U17234 ( .A1(n20705), .A2(n20469), .B1(n20704), .B2(n20468), .ZN(
        n13911) );
  OAI21_X1 U17235 ( .B1(n20617), .B2(n14184), .A(n13911), .ZN(n13912) );
  AOI21_X1 U17236 ( .B1(n20457), .B2(n20614), .A(n13912), .ZN(n13913) );
  OAI21_X1 U17237 ( .B1(n13999), .B2(n13914), .A(n13913), .ZN(P1_U3078) );
  INV_X1 U17238 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13922) );
  AOI22_X1 U17239 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n15176), .B1(DATAI_27_), 
        .B2(n15177), .ZN(n20697) );
  INV_X1 U17240 ( .A(n20697), .ZN(n20608) );
  AOI22_X1 U17241 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n15176), .B1(DATAI_19_), 
        .B2(n15177), .ZN(n20611) );
  NAND2_X1 U17242 ( .A1(n13927), .A2(DATAI_3_), .ZN(n13916) );
  NAND2_X1 U17243 ( .A1(n14327), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13915) );
  AND2_X1 U17244 ( .A1(n13916), .A2(n13915), .ZN(n14783) );
  NOR2_X2 U17245 ( .A1(n14783), .A2(n15174), .ZN(n20693) );
  INV_X1 U17246 ( .A(n15178), .ZN(n13918) );
  NAND2_X1 U17247 ( .A1(n13918), .A2(n13917), .ZN(n20410) );
  AOI22_X1 U17248 ( .A1(n20693), .A2(n20469), .B1(n20692), .B2(n20468), .ZN(
        n13919) );
  OAI21_X1 U17249 ( .B1(n20611), .B2(n14184), .A(n13919), .ZN(n13920) );
  AOI21_X1 U17250 ( .B1(n20457), .B2(n20608), .A(n13920), .ZN(n13921) );
  OAI21_X1 U17251 ( .B1(n13999), .B2(n13922), .A(n13921), .ZN(P1_U3076) );
  NAND2_X1 U17252 ( .A1(n13923), .A2(n14360), .ZN(n13924) );
  NAND2_X2 U17253 ( .A1(n14762), .A2(n13924), .ZN(n14805) );
  INV_X1 U17254 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n21053) );
  NAND2_X1 U17255 ( .A1(n13927), .A2(DATAI_0_), .ZN(n13926) );
  NAND2_X1 U17256 ( .A1(n14327), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13925) );
  AND2_X1 U17257 ( .A1(n13926), .A2(n13925), .ZN(n15175) );
  OAI222_X1 U17258 ( .A1(n14805), .A2(n14090), .B1(n14762), .B2(n21053), .C1(
        n14337), .C2(n15175), .ZN(P1_U2904) );
  OAI222_X1 U17259 ( .A1(n14805), .A2(n16162), .B1(n14762), .B2(n12188), .C1(
        n14337), .C2(n14772), .ZN(P1_U2899) );
  NAND2_X1 U17260 ( .A1(n13927), .A2(DATAI_1_), .ZN(n13929) );
  NAND2_X1 U17261 ( .A1(n14327), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13928) );
  AND2_X1 U17262 ( .A1(n13929), .A2(n13928), .ZN(n14798) );
  OAI222_X1 U17263 ( .A1(n14805), .A2(n14083), .B1(n14762), .B2(n12153), .C1(
        n14337), .C2(n14798), .ZN(P1_U2903) );
  OAI222_X1 U17264 ( .A1(n14805), .A2(n14075), .B1(n14762), .B2(n12172), .C1(
        n14337), .C2(n14783), .ZN(P1_U2901) );
  OAI222_X1 U17265 ( .A1(n14805), .A2(n13930), .B1(n14762), .B2(n12143), .C1(
        n14337), .C2(n14195), .ZN(P1_U2902) );
  XNOR2_X1 U17266 ( .A(n13931), .B(n14094), .ZN(n13937) );
  OR2_X1 U17267 ( .A1(n13944), .A2(n13932), .ZN(n13934) );
  NAND2_X1 U17268 ( .A1(n13934), .A2(n13933), .ZN(n19111) );
  MUX2_X1 U17269 ( .A(n19111), .B(n13935), .S(n9778), .Z(n13936) );
  OAI21_X1 U17270 ( .B1(n13937), .B2(n15337), .A(n13936), .ZN(P2_U2876) );
  INV_X1 U17271 ( .A(n13938), .ZN(n13941) );
  INV_X1 U17272 ( .A(n13931), .ZN(n13939) );
  OAI211_X1 U17273 ( .C1(n13941), .C2(n13940), .A(n13939), .B(n15341), .ZN(
        n13946) );
  NOR2_X1 U17274 ( .A1(n13779), .A2(n13942), .ZN(n13943) );
  NAND2_X1 U17275 ( .A1(n9846), .A2(n15319), .ZN(n13945) );
  OAI211_X1 U17276 ( .C1(n15319), .C2(n11570), .A(n13946), .B(n13945), .ZN(
        P2_U2877) );
  INV_X1 U17277 ( .A(n13731), .ZN(n13947) );
  OAI21_X1 U17278 ( .B1(n20618), .B2(n20588), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13949) );
  NAND2_X1 U17279 ( .A1(n13949), .A2(n20809), .ZN(n13955) );
  AND2_X1 U17280 ( .A1(n20815), .A2(n13415), .ZN(n20595) );
  INV_X1 U17281 ( .A(n20518), .ZN(n20437) );
  AND2_X1 U17282 ( .A1(n20595), .A2(n20437), .ZN(n13952) );
  NAND3_X1 U17283 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n12111), .ZN(n20596) );
  NOR2_X1 U17284 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20596), .ZN(
        n20586) );
  OR2_X1 U17285 ( .A1(n20332), .A2(n20825), .ZN(n13974) );
  NAND2_X1 U17286 ( .A1(n13974), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13971) );
  OAI21_X1 U17287 ( .B1(n20526), .B2(n20586), .A(n13971), .ZN(n13950) );
  INV_X1 U17288 ( .A(n13950), .ZN(n13951) );
  NAND2_X1 U17289 ( .A1(n13953), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20432) );
  OAI211_X1 U17290 ( .C1(n13955), .C2(n13952), .A(n13951), .B(n20525), .ZN(
        n20590) );
  INV_X1 U17291 ( .A(n20590), .ZN(n13964) );
  INV_X1 U17292 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13959) );
  INV_X1 U17293 ( .A(n13952), .ZN(n13954) );
  OR2_X1 U17294 ( .A1(n13953), .A2(n20839), .ZN(n20520) );
  OAI22_X1 U17295 ( .A1(n13955), .A2(n13954), .B1(n20520), .B2(n13974), .ZN(
        n20589) );
  AOI22_X1 U17296 ( .A1(n20588), .A2(n20651), .B1(n20586), .B2(n20686), .ZN(
        n13956) );
  OAI21_X1 U17297 ( .B1(n20654), .B2(n20627), .A(n13956), .ZN(n13957) );
  AOI21_X1 U17298 ( .B1(n20589), .B2(n20687), .A(n13957), .ZN(n13958) );
  OAI21_X1 U17299 ( .B1(n13964), .B2(n13959), .A(n13958), .ZN(P1_U3115) );
  INV_X1 U17300 ( .A(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13963) );
  AOI22_X1 U17301 ( .A1(n20588), .A2(n20608), .B1(n20586), .B2(n20692), .ZN(
        n13960) );
  OAI21_X1 U17302 ( .B1(n20611), .B2(n20627), .A(n13960), .ZN(n13961) );
  AOI21_X1 U17303 ( .B1(n20589), .B2(n20693), .A(n13961), .ZN(n13962) );
  OAI21_X1 U17304 ( .B1(n13964), .B2(n13963), .A(n13962), .ZN(P1_U3116) );
  INV_X1 U17305 ( .A(n20672), .ZN(n13966) );
  INV_X1 U17306 ( .A(n20725), .ZN(n13967) );
  OAI21_X1 U17307 ( .B1(n20658), .B2(n13967), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13969) );
  NOR2_X1 U17308 ( .A1(n13415), .A2(n13968), .ZN(n20665) );
  NAND2_X1 U17309 ( .A1(n20665), .A2(n20437), .ZN(n13973) );
  AOI21_X1 U17310 ( .B1(n13969), .B2(n13973), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n13972) );
  NOR2_X1 U17311 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20666), .ZN(
        n20655) );
  NAND2_X1 U17312 ( .A1(n20520), .A2(n13970), .ZN(n15171) );
  OR2_X1 U17313 ( .A1(n13973), .A2(n20667), .ZN(n13978) );
  INV_X1 U17314 ( .A(n20432), .ZN(n13976) );
  INV_X1 U17315 ( .A(n13974), .ZN(n13975) );
  NAND2_X1 U17316 ( .A1(n13976), .A2(n13975), .ZN(n13977) );
  NAND2_X1 U17317 ( .A1(n13978), .A2(n13977), .ZN(n20656) );
  AOI22_X1 U17318 ( .A1(n20719), .A2(n20656), .B1(n20716), .B2(n20655), .ZN(
        n13980) );
  NAND2_X1 U17319 ( .A1(n20658), .A2(n20587), .ZN(n13979) );
  OAI211_X1 U17320 ( .C1(n20593), .C2(n20725), .A(n13980), .B(n13979), .ZN(
        n13981) );
  AOI21_X1 U17321 ( .B1(n20659), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n13981), .ZN(n13982) );
  INV_X1 U17322 ( .A(n13982), .ZN(P1_U3152) );
  AOI22_X1 U17323 ( .A1(DATAI_20_), .A2(n15177), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n15176), .ZN(n20581) );
  NOR2_X2 U17324 ( .A1(n14777), .A2(n15174), .ZN(n20699) );
  NOR2_X2 U17325 ( .A1(n15178), .A2(n11786), .ZN(n20698) );
  AOI22_X1 U17326 ( .A1(n20699), .A2(n20656), .B1(n20655), .B2(n20698), .ZN(
        n13984) );
  AOI22_X1 U17327 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n15176), .B1(DATAI_28_), 
        .B2(n15177), .ZN(n20703) );
  INV_X1 U17328 ( .A(n20703), .ZN(n20578) );
  NAND2_X1 U17329 ( .A1(n20658), .A2(n20578), .ZN(n13983) );
  OAI211_X1 U17330 ( .C1(n20581), .C2(n20725), .A(n13984), .B(n13983), .ZN(
        n13985) );
  AOI21_X1 U17331 ( .B1(n20659), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n13985), .ZN(n13986) );
  INV_X1 U17332 ( .A(n13986), .ZN(P1_U3149) );
  AOI22_X1 U17333 ( .A1(n20693), .A2(n20656), .B1(n20692), .B2(n20655), .ZN(
        n13988) );
  NAND2_X1 U17334 ( .A1(n20658), .A2(n20608), .ZN(n13987) );
  OAI211_X1 U17335 ( .C1(n20611), .C2(n20725), .A(n13988), .B(n13987), .ZN(
        n13989) );
  AOI21_X1 U17336 ( .B1(n20659), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n13989), .ZN(n13990) );
  INV_X1 U17337 ( .A(n13990), .ZN(P1_U3148) );
  AOI22_X1 U17338 ( .A1(n20705), .A2(n20656), .B1(n20704), .B2(n20655), .ZN(
        n13992) );
  NAND2_X1 U17339 ( .A1(n20658), .A2(n20614), .ZN(n13991) );
  OAI211_X1 U17340 ( .C1(n20617), .C2(n20725), .A(n13992), .B(n13991), .ZN(
        n13993) );
  AOI21_X1 U17341 ( .B1(n20659), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n13993), .ZN(n13994) );
  INV_X1 U17342 ( .A(n13994), .ZN(P1_U3150) );
  INV_X1 U17343 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13998) );
  AOI22_X1 U17344 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n15176), .B1(DATAI_30_), 
        .B2(n15177), .ZN(n20715) );
  INV_X1 U17345 ( .A(n20715), .ZN(n20657) );
  AOI22_X1 U17346 ( .A1(DATAI_22_), .A2(n15177), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n15176), .ZN(n20662) );
  NOR2_X2 U17347 ( .A1(n14767), .A2(n15174), .ZN(n20711) );
  NOR2_X2 U17348 ( .A1(n15178), .A2(n11811), .ZN(n20710) );
  AOI22_X1 U17349 ( .A1(n20711), .A2(n20469), .B1(n20710), .B2(n20468), .ZN(
        n13995) );
  OAI21_X1 U17350 ( .B1(n20662), .B2(n14184), .A(n13995), .ZN(n13996) );
  AOI21_X1 U17351 ( .B1(n20457), .B2(n20657), .A(n13996), .ZN(n13997) );
  OAI21_X1 U17352 ( .B1(n13999), .B2(n13998), .A(n13997), .ZN(P1_U3079) );
  XNOR2_X1 U17353 ( .A(n14001), .B(n14000), .ZN(n19367) );
  OAI21_X1 U17354 ( .B1(n14002), .B2(n20857), .A(n14003), .ZN(n19366) );
  OAI21_X1 U17355 ( .B1(n19396), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n14004), .ZN(n16447) );
  INV_X1 U17356 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19999) );
  NOR2_X1 U17357 ( .A1(n19999), .A2(n13196), .ZN(n14005) );
  AOI221_X1 U17358 ( .B1(n16454), .B2(n20857), .C1(n16447), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n14005), .ZN(n14010) );
  AOI21_X1 U17359 ( .B1(n14008), .B2(n14007), .A(n14006), .ZN(n19370) );
  NAND2_X1 U17360 ( .A1(n19370), .A2(n19402), .ZN(n14009) );
  OAI211_X1 U17361 ( .C1(n16433), .C2(n19181), .A(n14010), .B(n14009), .ZN(
        n14011) );
  AOI21_X1 U17362 ( .B1(n19366), .B2(n16450), .A(n14011), .ZN(n14012) );
  OAI21_X1 U17363 ( .B1(n19395), .B2(n19367), .A(n14012), .ZN(P2_U3042) );
  OR2_X1 U17364 ( .A1(n13815), .A2(n14014), .ZN(n14015) );
  INV_X1 U17365 ( .A(n20224), .ZN(n14016) );
  OAI222_X1 U17366 ( .A1(n14805), .A2(n14016), .B1(n14762), .B2(n12198), .C1(
        n14337), .C2(n14767), .ZN(P1_U2898) );
  OR2_X1 U17367 ( .A1(n14013), .A2(n14017), .ZN(n14109) );
  NAND2_X1 U17368 ( .A1(n14013), .A2(n14017), .ZN(n14018) );
  AND2_X1 U17369 ( .A1(n14109), .A2(n14018), .ZN(n20174) );
  INV_X1 U17370 ( .A(n20174), .ZN(n14030) );
  OR2_X1 U17371 ( .A1(n16209), .A2(n14019), .ZN(n14020) );
  NAND2_X1 U17372 ( .A1(n14114), .A2(n14020), .ZN(n20167) );
  INV_X1 U17373 ( .A(n20167), .ZN(n14021) );
  AOI22_X1 U17374 ( .A1(n20222), .A2(n14021), .B1(n14716), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n14022) );
  OAI21_X1 U17375 ( .B1(n14030), .B2(n14701), .A(n14022), .ZN(P1_U2865) );
  XNOR2_X1 U17376 ( .A(n14023), .B(n14098), .ZN(n14029) );
  OAI21_X1 U17377 ( .B1(n14026), .B2(n14024), .A(n14025), .ZN(n19090) );
  INV_X1 U17378 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n14027) );
  MUX2_X1 U17379 ( .A(n19090), .B(n14027), .S(n9778), .Z(n14028) );
  OAI21_X1 U17380 ( .B1(n14029), .B2(n15337), .A(n14028), .ZN(P2_U2874) );
  OAI222_X1 U17381 ( .A1(n14030), .A2(n14805), .B1(n14762), .B2(n12238), .C1(
        n14763), .C2(n14337), .ZN(P1_U2897) );
  NAND2_X1 U17382 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n16229), .ZN(n16002) );
  NAND2_X1 U17383 ( .A1(n14031), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14032) );
  MUX2_X1 U17384 ( .A(n16002), .B(n14032), .S(n9918), .Z(n14033) );
  INV_X1 U17385 ( .A(n14033), .ZN(n14034) );
  NAND2_X1 U17386 ( .A1(n14112), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14036) );
  INV_X1 U17387 ( .A(n14036), .ZN(n14035) );
  INV_X1 U17388 ( .A(n20844), .ZN(n14045) );
  OAI21_X1 U17389 ( .B1(n14038), .B2(n14045), .A(n16117), .ZN(n20218) );
  NAND2_X1 U17390 ( .A1(n20218), .A2(n14039), .ZN(n14061) );
  NAND2_X1 U17391 ( .A1(n20846), .A2(n20840), .ZN(n14054) );
  INV_X1 U17392 ( .A(n14054), .ZN(n14040) );
  AND2_X1 U17393 ( .A1(n14041), .A2(n14040), .ZN(n15993) );
  AND2_X1 U17394 ( .A1(n14042), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14055) );
  NOR2_X1 U17395 ( .A1(n15993), .A2(n14055), .ZN(n14043) );
  NOR2_X1 U17396 ( .A1(n14045), .A2(n14044), .ZN(n20213) );
  NAND2_X1 U17397 ( .A1(n20213), .A2(n14046), .ZN(n14053) );
  INV_X1 U17398 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n14048) );
  OR3_X1 U17399 ( .A1(n14048), .A2(n20203), .A3(P1_REIP_REG_2__SCAN_IN), .ZN(
        n14052) );
  NAND2_X1 U17400 ( .A1(n20193), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14051) );
  OAI21_X1 U17401 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20203), .A(n14112), .ZN(
        n14049) );
  NAND2_X1 U17402 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n14049), .ZN(n14050) );
  NAND4_X1 U17403 ( .A1(n14053), .A2(n14052), .A3(n14051), .A4(n14050), .ZN(
        n14059) );
  NAND2_X1 U17404 ( .A1(n14055), .A2(n14054), .ZN(n14056) );
  NOR2_X2 U17405 ( .A1(n14057), .A2(n14056), .ZN(n20205) );
  NOR2_X1 U17406 ( .A1(n20191), .A2(n20308), .ZN(n14058) );
  AOI211_X1 U17407 ( .C1(n20206), .C2(P1_EBX_REG_2__SCAN_IN), .A(n14059), .B(
        n14058), .ZN(n14060) );
  OAI211_X1 U17408 ( .C1(n20216), .C2(n14062), .A(n14061), .B(n14060), .ZN(
        P1_U2838) );
  INV_X1 U17409 ( .A(n20218), .ZN(n14091) );
  INV_X1 U17410 ( .A(n20203), .ZN(n14063) );
  NAND4_X1 U17411 ( .A1(n14063), .A2(P1_REIP_REG_1__SCAN_IN), .A3(
        P1_REIP_REG_2__SCAN_IN), .A4(n20749), .ZN(n14066) );
  OAI221_X1 U17412 ( .B1(n20203), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n20203), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n14112), .ZN(n14064) );
  NAND2_X1 U17413 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n14064), .ZN(n14065) );
  OAI211_X1 U17414 ( .C1(n20210), .C2(n14067), .A(n14066), .B(n14065), .ZN(
        n14068) );
  AOI21_X1 U17415 ( .B1(P1_EBX_REG_3__SCAN_IN), .B2(n20206), .A(n14068), .ZN(
        n14069) );
  OAI21_X1 U17416 ( .B1(n20191), .B2(n14070), .A(n14069), .ZN(n14073) );
  NOR2_X1 U17417 ( .A1(n20216), .A2(n14071), .ZN(n14072) );
  AOI211_X1 U17418 ( .C1(n20213), .C2(n20815), .A(n14073), .B(n14072), .ZN(
        n14074) );
  OAI21_X1 U17419 ( .B1(n14091), .B2(n14075), .A(n14074), .ZN(P1_U2837) );
  INV_X1 U17420 ( .A(n20213), .ZN(n14084) );
  NAND2_X1 U17421 ( .A1(n20206), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n14077) );
  INV_X1 U17422 ( .A(n14112), .ZN(n14550) );
  AOI22_X1 U17423 ( .A1(n20193), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n14550), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n14076) );
  OAI211_X1 U17424 ( .C1(n14084), .C2(n20518), .A(n14077), .B(n14076), .ZN(
        n14080) );
  OAI22_X1 U17425 ( .A1(n20191), .A2(n14078), .B1(n20203), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n14079) );
  AOI211_X1 U17426 ( .C1(n20162), .C2(n14081), .A(n14080), .B(n14079), .ZN(
        n14082) );
  OAI21_X1 U17427 ( .B1(n14091), .B2(n14083), .A(n14082), .ZN(P1_U2839) );
  NAND2_X1 U17428 ( .A1(n20203), .A2(n14112), .ZN(n20189) );
  OAI22_X1 U17429 ( .A1(n20393), .A2(n14084), .B1(n20194), .B2(n13002), .ZN(
        n14087) );
  NOR2_X1 U17430 ( .A1(n20191), .A2(n14085), .ZN(n14086) );
  AOI211_X1 U17431 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(n20189), .A(n14087), .B(
        n14086), .ZN(n14089) );
  OAI21_X1 U17432 ( .B1(n20162), .B2(n20193), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14088) );
  OAI211_X1 U17433 ( .C1(n14091), .C2(n14090), .A(n14089), .B(n14088), .ZN(
        P1_U2840) );
  AOI21_X1 U17434 ( .B1(n14092), .B2(n13933), .A(n14024), .ZN(n19096) );
  INV_X1 U17435 ( .A(n19096), .ZN(n15776) );
  AOI21_X1 U17436 ( .B1(n13931), .B2(n14094), .A(n14093), .ZN(n14095) );
  OR3_X1 U17437 ( .A1(n14023), .A2(n14095), .A3(n15337), .ZN(n14097) );
  NAND2_X1 U17438 ( .A1(n15344), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14096) );
  OAI211_X1 U17439 ( .C1(n15776), .C2(n15344), .A(n14097), .B(n14096), .ZN(
        P2_U2875) );
  AND2_X1 U17440 ( .A1(n14023), .A2(n14098), .ZN(n14101) );
  OAI211_X1 U17441 ( .C1(n14101), .C2(n14100), .A(n15341), .B(n14099), .ZN(
        n14106) );
  NAND2_X1 U17442 ( .A1(n14102), .A2(n14025), .ZN(n14104) );
  INV_X1 U17443 ( .A(n14155), .ZN(n14103) );
  NAND2_X1 U17444 ( .A1(n15319), .A2(n19078), .ZN(n14105) );
  OAI211_X1 U17445 ( .C1(n15319), .C2(n14107), .A(n14106), .B(n14105), .ZN(
        P2_U2873) );
  INV_X1 U17446 ( .A(n14109), .ZN(n14111) );
  INV_X1 U17447 ( .A(n14108), .ZN(n14110) );
  OAI21_X1 U17448 ( .B1(n14111), .B2(n14110), .A(n14230), .ZN(n14271) );
  NAND4_X1 U17449 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n14548)
         );
  INV_X1 U17450 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20750) );
  NAND3_X1 U17451 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n20202) );
  NOR2_X1 U17452 ( .A1(n20750), .A2(n20202), .ZN(n14549) );
  NAND2_X1 U17453 ( .A1(n14549), .A2(n14112), .ZN(n20188) );
  NOR2_X1 U17454 ( .A1(n14548), .A2(n20188), .ZN(n14253) );
  NOR2_X1 U17455 ( .A1(n16031), .A2(n14253), .ZN(n20159) );
  NAND2_X1 U17456 ( .A1(n14114), .A2(n14113), .ZN(n14115) );
  AND2_X1 U17457 ( .A1(n14233), .A2(n14115), .ZN(n16195) );
  INV_X1 U17458 ( .A(n16195), .ZN(n14122) );
  INV_X1 U17459 ( .A(n14267), .ZN(n14116) );
  NAND2_X1 U17460 ( .A1(n20162), .A2(n14116), .ZN(n14121) );
  INV_X1 U17461 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14118) );
  NAND2_X1 U17462 ( .A1(n20193), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14117) );
  OAI211_X1 U17463 ( .C1(n20194), .C2(n14118), .A(n14117), .B(n20207), .ZN(
        n14119) );
  INV_X1 U17464 ( .A(n14119), .ZN(n14120) );
  OAI211_X1 U17465 ( .C1(n14122), .C2(n20191), .A(n14121), .B(n14120), .ZN(
        n14126) );
  NAND3_X1 U17466 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n14124) );
  INV_X1 U17467 ( .A(n14549), .ZN(n14123) );
  NOR3_X1 U17468 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14124), .A3(n20196), .ZN(
        n14125) );
  OR2_X1 U17469 ( .A1(n14126), .A2(n14125), .ZN(n14127) );
  AOI21_X1 U17470 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n20159), .A(n14127), .ZN(
        n14128) );
  OAI21_X1 U17471 ( .B1(n14271), .B2(n16117), .A(n14128), .ZN(P1_U2832) );
  AOI22_X1 U17472 ( .A1(n20222), .A2(n16195), .B1(n14716), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n14129) );
  OAI21_X1 U17473 ( .B1(n14271), .B2(n14701), .A(n14129), .ZN(P1_U2864) );
  NAND2_X1 U17474 ( .A1(n20425), .A2(n20385), .ZN(n14130) );
  NAND2_X1 U17475 ( .A1(n14130), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14131) );
  NAND2_X1 U17476 ( .A1(n14131), .A2(n20809), .ZN(n14135) );
  NAND2_X1 U17477 ( .A1(n9847), .A2(n20437), .ZN(n14133) );
  INV_X1 U17478 ( .A(n20332), .ZN(n14132) );
  NAND2_X1 U17479 ( .A1(n14132), .A2(n20825), .ZN(n14164) );
  OAI22_X1 U17480 ( .A1(n14135), .A2(n14133), .B1(n20520), .B2(n14164), .ZN(
        n20387) );
  INV_X1 U17481 ( .A(n20387), .ZN(n14154) );
  NOR2_X2 U17482 ( .A1(n14798), .A2(n15174), .ZN(n20681) );
  INV_X1 U17483 ( .A(n20681), .ZN(n14188) );
  INV_X1 U17484 ( .A(n14133), .ZN(n14134) );
  NAND3_X1 U17485 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20825), .A3(
        n12111), .ZN(n20397) );
  NOR2_X1 U17486 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20397), .ZN(
        n14139) );
  OAI22_X1 U17487 ( .A1(n14135), .A2(n14134), .B1(n14139), .B2(n20526), .ZN(
        n14136) );
  INV_X1 U17488 ( .A(n14136), .ZN(n14137) );
  OAI21_X1 U17489 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20332), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14168) );
  NAND3_X1 U17490 ( .A1(n20525), .A2(n14137), .A3(n14168), .ZN(n20388) );
  NAND2_X1 U17491 ( .A1(n20388), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n14142) );
  INV_X1 U17492 ( .A(n20425), .ZN(n14150) );
  AOI22_X1 U17493 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n15176), .B1(DATAI_17_), 
        .B2(n15177), .ZN(n20650) );
  INV_X1 U17494 ( .A(n20650), .ZN(n20682) );
  AOI22_X1 U17495 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n15176), .B1(DATAI_25_), 
        .B2(n15177), .ZN(n20685) );
  NOR2_X2 U17496 ( .A1(n15178), .A2(n14138), .ZN(n20680) );
  INV_X1 U17497 ( .A(n20680), .ZN(n20402) );
  INV_X1 U17498 ( .A(n14139), .ZN(n20384) );
  OAI22_X1 U17499 ( .A1(n20385), .A2(n20685), .B1(n20402), .B2(n20384), .ZN(
        n14140) );
  AOI21_X1 U17500 ( .B1(n14150), .B2(n20682), .A(n14140), .ZN(n14141) );
  OAI211_X1 U17501 ( .C1(n14154), .C2(n14188), .A(n14142), .B(n14141), .ZN(
        P1_U3050) );
  INV_X1 U17502 ( .A(n20705), .ZN(n14182) );
  NAND2_X1 U17503 ( .A1(n20388), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n14145) );
  INV_X1 U17504 ( .A(n20617), .ZN(n20706) );
  INV_X1 U17505 ( .A(n20704), .ZN(n14178) );
  OAI22_X1 U17506 ( .A1(n20385), .A2(n20709), .B1(n14178), .B2(n20384), .ZN(
        n14143) );
  AOI21_X1 U17507 ( .B1(n14150), .B2(n20706), .A(n14143), .ZN(n14144) );
  OAI211_X1 U17508 ( .C1(n14154), .C2(n14182), .A(n14145), .B(n14144), .ZN(
        P1_U3054) );
  INV_X1 U17509 ( .A(n20693), .ZN(n14177) );
  NAND2_X1 U17510 ( .A1(n20388), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n14148) );
  INV_X1 U17511 ( .A(n20611), .ZN(n20694) );
  OAI22_X1 U17512 ( .A1(n20385), .A2(n20697), .B1(n20384), .B2(n20410), .ZN(
        n14146) );
  AOI21_X1 U17513 ( .B1(n14150), .B2(n20694), .A(n14146), .ZN(n14147) );
  OAI211_X1 U17514 ( .C1(n14154), .C2(n14177), .A(n14148), .B(n14147), .ZN(
        P1_U3052) );
  INV_X1 U17515 ( .A(n20719), .ZN(n14153) );
  NAND2_X1 U17516 ( .A1(n20388), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n14152) );
  INV_X1 U17517 ( .A(n20593), .ZN(n20720) );
  INV_X1 U17518 ( .A(n20716), .ZN(n20424) );
  OAI22_X1 U17519 ( .A1(n20385), .A2(n20726), .B1(n20424), .B2(n20384), .ZN(
        n14149) );
  AOI21_X1 U17520 ( .B1(n14150), .B2(n20720), .A(n14149), .ZN(n14151) );
  OAI211_X1 U17521 ( .C1(n14154), .C2(n14153), .A(n14152), .B(n14151), .ZN(
        P1_U3056) );
  XNOR2_X1 U17522 ( .A(n14099), .B(n15297), .ZN(n14160) );
  OR2_X1 U17523 ( .A1(n14156), .A2(n14155), .ZN(n14158) );
  INV_X1 U17524 ( .A(n14462), .ZN(n14157) );
  NAND2_X1 U17525 ( .A1(n14158), .A2(n14157), .ZN(n16334) );
  MUX2_X1 U17526 ( .A(n16334), .B(n11585), .S(n9778), .Z(n14159) );
  OAI21_X1 U17527 ( .B1(n14160), .B2(n15337), .A(n14159), .ZN(P2_U2872) );
  OAI21_X1 U17528 ( .B1(n20511), .B2(n20481), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14163) );
  NAND2_X1 U17529 ( .A1(n14163), .A2(n20809), .ZN(n14165) );
  NAND2_X1 U17530 ( .A1(n20487), .A2(n20437), .ZN(n14166) );
  OAI22_X1 U17531 ( .A1(n14165), .A2(n14166), .B1(n20432), .B2(n14164), .ZN(
        n20482) );
  INV_X1 U17532 ( .A(n20482), .ZN(n14189) );
  INV_X1 U17533 ( .A(n20711), .ZN(n14173) );
  INV_X1 U17534 ( .A(n14165), .ZN(n14167) );
  INV_X1 U17535 ( .A(n20492), .ZN(n20488) );
  NOR2_X1 U17536 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20488), .ZN(
        n20480) );
  INV_X1 U17537 ( .A(n20480), .ZN(n14183) );
  AOI22_X1 U17538 ( .A1(n14167), .A2(n14166), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n14183), .ZN(n14169) );
  NAND3_X1 U17539 ( .A1(n20438), .A2(n14169), .A3(n14168), .ZN(n20483) );
  NAND2_X1 U17540 ( .A1(n20483), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n14172) );
  INV_X1 U17541 ( .A(n20662), .ZN(n20712) );
  INV_X1 U17542 ( .A(n20710), .ZN(n20419) );
  OAI22_X1 U17543 ( .A1(n14184), .A2(n20715), .B1(n14183), .B2(n20419), .ZN(
        n14170) );
  AOI21_X1 U17544 ( .B1(n20511), .B2(n20712), .A(n14170), .ZN(n14171) );
  OAI211_X1 U17545 ( .C1(n14189), .C2(n14173), .A(n14172), .B(n14171), .ZN(
        P1_U3087) );
  NAND2_X1 U17546 ( .A1(n20483), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n14176) );
  OAI22_X1 U17547 ( .A1(n14184), .A2(n20697), .B1(n14183), .B2(n20410), .ZN(
        n14174) );
  AOI21_X1 U17548 ( .B1(n20511), .B2(n20694), .A(n14174), .ZN(n14175) );
  OAI211_X1 U17549 ( .C1(n14189), .C2(n14177), .A(n14176), .B(n14175), .ZN(
        P1_U3084) );
  NAND2_X1 U17550 ( .A1(n20483), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n14181) );
  OAI22_X1 U17551 ( .A1(n14184), .A2(n20709), .B1(n14183), .B2(n14178), .ZN(
        n14179) );
  AOI21_X1 U17552 ( .B1(n20511), .B2(n20706), .A(n14179), .ZN(n14180) );
  OAI211_X1 U17553 ( .C1(n14189), .C2(n14182), .A(n14181), .B(n14180), .ZN(
        P1_U3086) );
  NAND2_X1 U17554 ( .A1(n20483), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n14187) );
  OAI22_X1 U17555 ( .A1(n14184), .A2(n20685), .B1(n14183), .B2(n20402), .ZN(
        n14185) );
  AOI21_X1 U17556 ( .B1(n20511), .B2(n20682), .A(n14185), .ZN(n14186) );
  OAI211_X1 U17557 ( .C1(n14189), .C2(n14188), .A(n14187), .B(n14186), .ZN(
        P1_U3082) );
  INV_X1 U17558 ( .A(DATAI_8_), .ZN(n14191) );
  INV_X1 U17559 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n14190) );
  MUX2_X1 U17560 ( .A(n14191), .B(n14190), .S(n14327), .Z(n20251) );
  OAI222_X1 U17561 ( .A1(n14805), .A2(n14271), .B1(n14337), .B2(n20251), .C1(
        n14192), .C2(n14762), .ZN(P1_U2896) );
  AOI22_X1 U17562 ( .A1(n20281), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20284), .ZN(n14194) );
  INV_X1 U17563 ( .A(n15175), .ZN(n14193) );
  NAND2_X1 U17564 ( .A1(n20269), .A2(n14193), .ZN(n14203) );
  NAND2_X1 U17565 ( .A1(n14194), .A2(n14203), .ZN(P1_U2952) );
  AOI22_X1 U17566 ( .A1(n20281), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20284), .ZN(n14196) );
  INV_X1 U17567 ( .A(n14195), .ZN(n14790) );
  NAND2_X1 U17568 ( .A1(n20269), .A2(n14790), .ZN(n14201) );
  NAND2_X1 U17569 ( .A1(n14196), .A2(n14201), .ZN(P1_U2939) );
  AOI22_X1 U17570 ( .A1(n20281), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20284), .ZN(n14198) );
  INV_X1 U17571 ( .A(n14783), .ZN(n14197) );
  NAND2_X1 U17572 ( .A1(n20269), .A2(n14197), .ZN(n14215) );
  NAND2_X1 U17573 ( .A1(n14198), .A2(n14215), .ZN(P1_U2940) );
  AOI22_X1 U17574 ( .A1(n20281), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20284), .ZN(n14200) );
  INV_X1 U17575 ( .A(n14798), .ZN(n14199) );
  NAND2_X1 U17576 ( .A1(n20269), .A2(n14199), .ZN(n14219) );
  NAND2_X1 U17577 ( .A1(n14200), .A2(n14219), .ZN(P1_U2938) );
  AOI22_X1 U17578 ( .A1(n20281), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20284), .ZN(n14202) );
  NAND2_X1 U17579 ( .A1(n14202), .A2(n14201), .ZN(P1_U2954) );
  AOI22_X1 U17580 ( .A1(n20281), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20284), .ZN(n14204) );
  NAND2_X1 U17581 ( .A1(n14204), .A2(n14203), .ZN(P1_U2937) );
  AOI22_X1 U17582 ( .A1(n20281), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20284), .ZN(n14206) );
  NAND2_X1 U17583 ( .A1(n14206), .A2(n14205), .ZN(P1_U2944) );
  AOI22_X1 U17584 ( .A1(n20281), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20284), .ZN(n14210) );
  INV_X1 U17585 ( .A(DATAI_9_), .ZN(n14208) );
  MUX2_X1 U17586 ( .A(n14208), .B(n14207), .S(n14327), .Z(n14753) );
  INV_X1 U17587 ( .A(n14753), .ZN(n14209) );
  NAND2_X1 U17588 ( .A1(n20269), .A2(n14209), .ZN(n20273) );
  NAND2_X1 U17589 ( .A1(n14210), .A2(n20273), .ZN(P1_U2946) );
  AOI22_X1 U17590 ( .A1(n20281), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20284), .ZN(n14212) );
  NAND2_X1 U17591 ( .A1(n14212), .A2(n14211), .ZN(P1_U2943) );
  AOI22_X1 U17592 ( .A1(n20281), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20284), .ZN(n14214) );
  NAND2_X1 U17593 ( .A1(n14214), .A2(n14213), .ZN(P1_U2942) );
  AOI22_X1 U17594 ( .A1(n20281), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20284), .ZN(n14216) );
  NAND2_X1 U17595 ( .A1(n14216), .A2(n14215), .ZN(P1_U2955) );
  AOI22_X1 U17596 ( .A1(n20281), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20284), .ZN(n14218) );
  NAND2_X1 U17597 ( .A1(n14218), .A2(n14217), .ZN(P1_U2941) );
  AOI22_X1 U17598 ( .A1(n20281), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20284), .ZN(n14220) );
  NAND2_X1 U17599 ( .A1(n14220), .A2(n14219), .ZN(P1_U2953) );
  NOR2_X1 U17600 ( .A1(n14234), .A2(n14221), .ZN(n14222) );
  OR2_X1 U17601 ( .A1(n14303), .A2(n14222), .ZN(n16183) );
  INV_X1 U17602 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14226) );
  OAI21_X1 U17603 ( .B1(n14223), .B2(n14225), .A(n14272), .ZN(n16118) );
  OAI222_X1 U17604 ( .A1(n16183), .A2(n14725), .B1(n14226), .B2(n20227), .C1(
        n16118), .C2(n14730), .ZN(P1_U2862) );
  INV_X1 U17605 ( .A(DATAI_10_), .ZN(n21062) );
  MUX2_X1 U17606 ( .A(n21062), .B(n16603), .S(n14327), .Z(n20254) );
  INV_X1 U17607 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14227) );
  OAI222_X1 U17608 ( .A1(n14805), .A2(n16118), .B1(n14337), .B2(n20254), .C1(
        n14227), .C2(n14762), .ZN(P1_U2894) );
  INV_X1 U17609 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20244) );
  OAI222_X1 U17610 ( .A1(n14337), .A2(n14777), .B1(n14805), .B2(n14228), .C1(
        n20244), .C2(n14762), .ZN(P1_U2900) );
  AND2_X1 U17611 ( .A1(n14230), .A2(n14229), .ZN(n14231) );
  OR2_X1 U17612 ( .A1(n14231), .A2(n14223), .ZN(n20160) );
  INV_X1 U17613 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n14236) );
  AND2_X1 U17614 ( .A1(n14233), .A2(n14232), .ZN(n14235) );
  OR2_X1 U17615 ( .A1(n14235), .A2(n14234), .ZN(n20156) );
  OAI222_X1 U17616 ( .A1(n20160), .A2(n14701), .B1(n14236), .B2(n20227), .C1(
        n20156), .C2(n14725), .ZN(P1_U2863) );
  INV_X1 U17617 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n14237) );
  OAI222_X1 U17618 ( .A1(n14805), .A2(n20160), .B1(n14337), .B2(n14753), .C1(
        n14237), .C2(n14762), .ZN(P1_U2895) );
  NOR2_X1 U17619 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14238), .ZN(
        n16222) );
  NAND2_X1 U17620 ( .A1(n15129), .A2(n14239), .ZN(n16220) );
  INV_X1 U17621 ( .A(n16220), .ZN(n14240) );
  NOR2_X1 U17622 ( .A1(n15073), .A2(n14240), .ZN(n14308) );
  OAI21_X1 U17623 ( .B1(n15124), .B2(n14241), .A(n14308), .ZN(n16215) );
  INV_X1 U17624 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16205) );
  NOR3_X1 U17625 ( .A1(n16222), .A2(n16215), .A3(n16205), .ZN(n16214) );
  NOR2_X1 U17626 ( .A1(n14313), .A2(n16214), .ZN(n16196) );
  INV_X1 U17627 ( .A(n16196), .ZN(n14249) );
  NAND2_X1 U17628 ( .A1(n14244), .A2(n14243), .ZN(n14245) );
  XNOR2_X1 U17629 ( .A(n14242), .B(n14245), .ZN(n16150) );
  NAND2_X1 U17630 ( .A1(n16150), .A2(n20318), .ZN(n14248) );
  NOR2_X1 U17631 ( .A1(n16204), .A2(n16205), .ZN(n16198) );
  INV_X1 U17632 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20756) );
  OAI22_X1 U17633 ( .A1(n16218), .A2(n20167), .B1(n20756), .B2(n20207), .ZN(
        n14246) );
  AOI21_X1 U17634 ( .B1(n16198), .B2(n16199), .A(n14246), .ZN(n14247) );
  OAI211_X1 U17635 ( .C1(n14249), .C2(n16199), .A(n14248), .B(n14247), .ZN(
        P1_U3024) );
  OAI21_X1 U17636 ( .B1(n14276), .B2(n14251), .A(n14250), .ZN(n14931) );
  NAND3_X1 U17637 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(P1_REIP_REG_11__SCAN_IN), .ZN(n14252) );
  NAND3_X1 U17638 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(n20158), .ZN(n16093) );
  NOR2_X1 U17639 ( .A1(n14252), .A2(n16093), .ZN(n14353) );
  NAND4_X1 U17640 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(P1_REIP_REG_11__SCAN_IN), .ZN(n14547) );
  NAND3_X1 U17641 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(n14253), .ZN(n16102) );
  NOR2_X1 U17642 ( .A1(n14547), .A2(n16102), .ZN(n14254) );
  OR2_X1 U17643 ( .A1(n14254), .A2(n16031), .ZN(n16087) );
  INV_X1 U17644 ( .A(n16087), .ZN(n14354) );
  OAI21_X1 U17645 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n14353), .A(n14354), 
        .ZN(n14262) );
  INV_X1 U17646 ( .A(n14255), .ZN(n14928) );
  INV_X1 U17647 ( .A(n14279), .ZN(n14323) );
  AOI21_X1 U17648 ( .B1(n14323), .B2(n14278), .A(n14256), .ZN(n14257) );
  OR2_X1 U17649 ( .A1(n14257), .A2(n14348), .ZN(n16166) );
  OAI22_X1 U17650 ( .A1(n16166), .A2(n20191), .B1(n20194), .B2(n20876), .ZN(
        n14258) );
  INV_X1 U17651 ( .A(n14258), .ZN(n14259) );
  OAI211_X1 U17652 ( .C1(n20210), .C2(n14926), .A(n14259), .B(n20207), .ZN(
        n14260) );
  AOI21_X1 U17653 ( .B1(n20162), .B2(n14928), .A(n14260), .ZN(n14261) );
  OAI211_X1 U17654 ( .C1(n14931), .C2(n16117), .A(n14262), .B(n14261), .ZN(
        P1_U2826) );
  XNOR2_X1 U17655 ( .A(n14264), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14265) );
  XNOR2_X1 U17656 ( .A(n14263), .B(n14265), .ZN(n16197) );
  NAND2_X1 U17657 ( .A1(n16197), .A2(n20294), .ZN(n14270) );
  INV_X1 U17658 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n14266) );
  NOR2_X1 U17659 ( .A1(n20207), .A2(n14266), .ZN(n16194) );
  NOR2_X1 U17660 ( .A1(n20298), .A2(n14267), .ZN(n14268) );
  AOI211_X1 U17661 ( .C1(n20287), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16194), .B(n14268), .ZN(n14269) );
  OAI211_X1 U17662 ( .C1(n14954), .C2(n14271), .A(n14270), .B(n14269), .ZN(
        P1_U2991) );
  INV_X1 U17663 ( .A(n14272), .ZN(n14274) );
  OAI21_X1 U17664 ( .B1(n14274), .B2(n14273), .A(n14275), .ZN(n14298) );
  OAI21_X1 U17665 ( .B1(n14298), .B2(n14299), .A(n14275), .ZN(n14318) );
  XNOR2_X1 U17666 ( .A(n14279), .B(n14278), .ZN(n16173) );
  AOI22_X1 U17667 ( .A1(n16173), .A2(n20222), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14716), .ZN(n14280) );
  OAI21_X1 U17668 ( .B1(n14944), .B2(n14730), .A(n14280), .ZN(P1_U2859) );
  AOI22_X1 U17669 ( .A1(n16173), .A2(n20205), .B1(n20206), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14281) );
  OAI211_X1 U17670 ( .C1(n20210), .C2(n14282), .A(n14281), .B(n20207), .ZN(
        n14287) );
  NAND2_X1 U17671 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14283) );
  NOR2_X1 U17672 ( .A1(n14283), .A2(n16093), .ZN(n14285) );
  OAI21_X1 U17673 ( .B1(n14283), .B2(n16102), .A(n20189), .ZN(n16101) );
  INV_X1 U17674 ( .A(n16101), .ZN(n14284) );
  MUX2_X1 U17675 ( .A(n14285), .B(n14284), .S(P1_REIP_REG_13__SCAN_IN), .Z(
        n14286) );
  AOI211_X1 U17676 ( .C1(n20162), .C2(n14941), .A(n14287), .B(n14286), .ZN(
        n14288) );
  OAI21_X1 U17677 ( .B1(n14944), .B2(n16117), .A(n14288), .ZN(P1_U2827) );
  INV_X1 U17678 ( .A(DATAI_14_), .ZN(n14290) );
  INV_X1 U17679 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14289) );
  MUX2_X1 U17680 ( .A(n14290), .B(n14289), .S(n14327), .Z(n20267) );
  OAI222_X1 U17681 ( .A1(n14805), .A2(n14931), .B1(n14337), .B2(n20267), .C1(
        n14291), .C2(n14762), .ZN(P1_U2890) );
  OAI222_X1 U17682 ( .A1(n14730), .A2(n14931), .B1(n20876), .B2(n20227), .C1(
        n16166), .C2(n14725), .ZN(P1_U2858) );
  XNOR2_X1 U17683 ( .A(n15138), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14293) );
  XNOR2_X1 U17684 ( .A(n14292), .B(n14293), .ZN(n14316) );
  INV_X1 U17685 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n14294) );
  OAI22_X1 U17686 ( .A1(n14950), .A2(n12244), .B1(n20207), .B2(n14294), .ZN(
        n14296) );
  NOR2_X1 U17687 ( .A1(n20160), .A2(n14954), .ZN(n14295) );
  AOI211_X1 U17688 ( .C1(n16141), .C2(n20161), .A(n14296), .B(n14295), .ZN(
        n14297) );
  OAI21_X1 U17689 ( .B1(n14316), .B2(n20139), .A(n14297), .ZN(P1_U2990) );
  XOR2_X1 U17690 ( .A(n14299), .B(n14298), .Z(n16145) );
  INV_X1 U17691 ( .A(n16145), .ZN(n14306) );
  INV_X1 U17692 ( .A(DATAI_11_), .ZN(n14300) );
  MUX2_X1 U17693 ( .A(n14300), .B(n21125), .S(n14327), .Z(n20258) );
  OAI222_X1 U17694 ( .A1(n14306), .A2(n14805), .B1(n14301), .B2(n14762), .C1(
        n14337), .C2(n20258), .ZN(P1_U2893) );
  INV_X1 U17695 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14305) );
  OR2_X1 U17696 ( .A1(n14303), .A2(n14302), .ZN(n14304) );
  NAND2_X1 U17697 ( .A1(n14324), .A2(n14304), .ZN(n16103) );
  OAI222_X1 U17698 ( .A1(n14306), .A2(n14701), .B1(n14305), .B2(n20227), .C1(
        n16103), .C2(n14725), .ZN(P1_U2861) );
  NOR2_X1 U17699 ( .A1(n16204), .A2(n14309), .ZN(n16188) );
  OAI22_X1 U17700 ( .A1(n16218), .A2(n20156), .B1(n14294), .B2(n20207), .ZN(
        n14307) );
  AOI21_X1 U17701 ( .B1(n16188), .B2(n16189), .A(n14307), .ZN(n14315) );
  INV_X1 U17702 ( .A(n14308), .ZN(n15127) );
  AOI211_X1 U17703 ( .C1(n14311), .C2(n14310), .A(n14309), .B(n15127), .ZN(
        n14312) );
  NOR2_X1 U17704 ( .A1(n14313), .A2(n14312), .ZN(n16186) );
  NAND2_X1 U17705 ( .A1(n16186), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14314) );
  OAI211_X1 U17706 ( .C1(n14316), .C2(n15137), .A(n14315), .B(n14314), .ZN(
        P1_U3022) );
  INV_X1 U17707 ( .A(DATAI_13_), .ZN(n21074) );
  INV_X1 U17708 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16599) );
  MUX2_X1 U17709 ( .A(n21074), .B(n16599), .S(n14327), .Z(n20264) );
  INV_X1 U17710 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14317) );
  OAI222_X1 U17711 ( .A1(n14805), .A2(n14944), .B1(n14337), .B2(n20264), .C1(
        n14317), .C2(n14762), .ZN(P1_U2891) );
  INV_X1 U17712 ( .A(n14318), .ZN(n14322) );
  INV_X1 U17713 ( .A(n14319), .ZN(n14321) );
  INV_X1 U17714 ( .A(n16139), .ZN(n14331) );
  AOI21_X1 U17715 ( .B1(n14325), .B2(n14324), .A(n14323), .ZN(n16097) );
  AOI22_X1 U17716 ( .A1(n16097), .A2(n20222), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n14716), .ZN(n14326) );
  OAI21_X1 U17717 ( .B1(n14331), .B2(n14701), .A(n14326), .ZN(P1_U2860) );
  INV_X1 U17718 ( .A(DATAI_12_), .ZN(n14329) );
  MUX2_X1 U17719 ( .A(n14329), .B(n14328), .S(n14327), .Z(n20261) );
  OAI222_X1 U17720 ( .A1(n14331), .A2(n14805), .B1(n14330), .B2(n14762), .C1(
        n14337), .C2(n20261), .ZN(P1_U2892) );
  NAND2_X1 U17721 ( .A1(n14250), .A2(n14333), .ZN(n14334) );
  AND2_X1 U17722 ( .A1(n14341), .A2(n14334), .ZN(n16135) );
  XNOR2_X1 U17723 ( .A(n14348), .B(n14344), .ZN(n16082) );
  AOI22_X1 U17724 ( .A1(n16082), .A2(n20222), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n14716), .ZN(n14335) );
  OAI21_X1 U17725 ( .B1(n14339), .B2(n14730), .A(n14335), .ZN(P1_U2857) );
  OAI222_X1 U17726 ( .A1(n14805), .A2(n14339), .B1(n14762), .B2(n14338), .C1(
        n14337), .C2(n14336), .ZN(P1_U2889) );
  AOI21_X1 U17727 ( .B1(n14342), .B2(n14341), .A(n14340), .ZN(n14343) );
  INV_X1 U17728 ( .A(n14343), .ZN(n14916) );
  INV_X1 U17729 ( .A(n14344), .ZN(n14347) );
  INV_X1 U17730 ( .A(n14345), .ZN(n14346) );
  AOI21_X1 U17731 ( .B1(n14348), .B2(n14347), .A(n14346), .ZN(n14349) );
  OR2_X1 U17732 ( .A1(n14678), .A2(n14349), .ZN(n15103) );
  INV_X1 U17733 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14364) );
  OAI22_X1 U17734 ( .A1(n15103), .A2(n20191), .B1(n20194), .B2(n14364), .ZN(
        n14350) );
  INV_X1 U17735 ( .A(n14350), .ZN(n14351) );
  OAI211_X1 U17736 ( .C1(n20210), .C2(n14911), .A(n14351), .B(n20207), .ZN(
        n14352) );
  INV_X1 U17737 ( .A(n14352), .ZN(n14356) );
  NAND2_X1 U17738 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n14353), .ZN(n16068) );
  NOR2_X1 U17739 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n16068), .ZN(n16089) );
  OAI21_X1 U17740 ( .B1(n14354), .B2(n16089), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n14355) );
  NAND2_X1 U17741 ( .A1(n14356), .A2(n14355), .ZN(n14358) );
  INV_X1 U17742 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20764) );
  NOR3_X1 U17743 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n20764), .A3(n16068), 
        .ZN(n14357) );
  AOI211_X1 U17744 ( .C1(n20162), .C2(n14913), .A(n14358), .B(n14357), .ZN(
        n14359) );
  OAI21_X1 U17745 ( .B1(n14916), .B2(n16117), .A(n14359), .ZN(P1_U2824) );
  NAND3_X1 U17746 ( .A1(n14762), .A2(n12083), .A3(n14360), .ZN(n14799) );
  OAI22_X1 U17747 ( .A1(n14799), .A2(n15175), .B1(n14762), .B2(n13663), .ZN(
        n14361) );
  AOI21_X1 U17748 ( .B1(n14801), .B2(BUF1_REG_16__SCAN_IN), .A(n14361), .ZN(
        n14363) );
  NAND2_X1 U17749 ( .A1(n14802), .A2(DATAI_16_), .ZN(n14362) );
  OAI211_X1 U17750 ( .C1(n14916), .C2(n14805), .A(n14363), .B(n14362), .ZN(
        P1_U2888) );
  OAI222_X1 U17751 ( .A1(n14730), .A2(n14916), .B1(n14364), .B2(n20227), .C1(
        n15103), .C2(n14725), .ZN(P1_U2856) );
  AOI22_X1 U17752 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14368) );
  AOI22_X1 U17753 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17295), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14367) );
  AOI22_X1 U17754 ( .A1(n17303), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14366) );
  AOI22_X1 U17755 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14365) );
  NAND4_X1 U17756 ( .A1(n14368), .A2(n14367), .A3(n14366), .A4(n14365), .ZN(
        n14374) );
  AOI22_X1 U17757 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14372) );
  AOI22_X1 U17758 ( .A1(n17305), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14371) );
  AOI22_X1 U17759 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14370) );
  AOI22_X1 U17760 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14369) );
  NAND4_X1 U17761 ( .A1(n14372), .A2(n14371), .A3(n14370), .A4(n14369), .ZN(
        n14373) );
  NOR2_X1 U17762 ( .A1(n14374), .A2(n14373), .ZN(n17450) );
  INV_X1 U17763 ( .A(n17450), .ZN(n14380) );
  NOR2_X1 U17764 ( .A1(n14375), .A2(n17318), .ZN(n17325) );
  INV_X1 U17765 ( .A(n17325), .ZN(n14377) );
  NOR2_X1 U17766 ( .A1(n14376), .A2(n14377), .ZN(n17259) );
  INV_X1 U17767 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16954) );
  INV_X1 U17768 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17291) );
  NOR2_X1 U17769 ( .A1(n17317), .A2(n14377), .ZN(n17316) );
  NAND2_X1 U17770 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17316), .ZN(n17312) );
  NOR3_X1 U17771 ( .A1(n16954), .A2(n17291), .A3(n17312), .ZN(n17275) );
  AOI21_X1 U17772 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17275), .A(
        P3_EBX_REG_11__SCAN_IN), .ZN(n14378) );
  NOR2_X1 U17773 ( .A1(n17259), .A2(n14378), .ZN(n14379) );
  MUX2_X1 U17774 ( .A(n14380), .B(n14379), .S(n17338), .Z(P3_U2692) );
  NAND2_X1 U17775 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17172), .ZN(n17132) );
  NOR3_X1 U17776 ( .A1(n13541), .A2(n14381), .A3(n17132), .ZN(n17084) );
  NAND2_X1 U17777 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17084), .ZN(n14382) );
  NOR2_X1 U17778 ( .A1(n17431), .A2(n14382), .ZN(n14384) );
  NAND2_X1 U17779 ( .A1(n17338), .A2(n14382), .ZN(n17085) );
  INV_X1 U17780 ( .A(n17085), .ZN(n14383) );
  MUX2_X1 U17781 ( .A(n14384), .B(n14383), .S(P3_EBX_REG_31__SCAN_IN), .Z(
        P3_U2672) );
  NAND2_X1 U17782 ( .A1(n14385), .A2(n14513), .ZN(n14394) );
  INV_X1 U17783 ( .A(n16342), .ZN(n14386) );
  INV_X1 U17784 ( .A(n16330), .ZN(n14387) );
  OAI21_X2 U17785 ( .B1(n16332), .B2(n14387), .A(n16331), .ZN(n14468) );
  INV_X1 U17786 ( .A(n14388), .ZN(n14389) );
  INV_X1 U17787 ( .A(n14445), .ZN(n14390) );
  INV_X1 U17788 ( .A(n14391), .ZN(n15532) );
  INV_X1 U17789 ( .A(n14392), .ZN(n15533) );
  XOR2_X1 U17790 ( .A(n14394), .B(n14393), .Z(n14416) );
  INV_X1 U17791 ( .A(n14401), .ZN(n14395) );
  INV_X1 U17792 ( .A(n15798), .ZN(n16407) );
  OAI21_X1 U17793 ( .B1(n14395), .B2(n19396), .A(n16407), .ZN(n15752) );
  AND2_X1 U17794 ( .A1(n15432), .A2(n14396), .ZN(n14397) );
  NOR2_X1 U17795 ( .A1(n15415), .A2(n14397), .ZN(n19020) );
  INV_X1 U17796 ( .A(n19020), .ZN(n15425) );
  OR2_X1 U17797 ( .A1(n15329), .A2(n14399), .ZN(n14400) );
  NAND2_X1 U17798 ( .A1(n14398), .A2(n14400), .ZN(n19022) );
  INV_X1 U17799 ( .A(n19022), .ZN(n14414) );
  OR2_X1 U17800 ( .A1(n14401), .A2(n15800), .ZN(n15736) );
  NAND2_X1 U17801 ( .A1(n19365), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n14409) );
  OAI21_X1 U17802 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15736), .A(
        n14409), .ZN(n14402) );
  AOI21_X1 U17803 ( .B1(n19402), .B2(n14414), .A(n14402), .ZN(n14403) );
  OAI21_X1 U17804 ( .B1(n16433), .B2(n15425), .A(n14403), .ZN(n14408) );
  OR2_X1 U17805 ( .A1(n14404), .A2(n15554), .ZN(n14407) );
  INV_X1 U17806 ( .A(n14407), .ZN(n14405) );
  AND2_X1 U17807 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n14405), .ZN(
        n14522) );
  AND2_X1 U17808 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14406) );
  NAND2_X2 U17809 ( .A1(n14425), .A2(n14406), .ZN(n15555) );
  NOR2_X1 U17810 ( .A1(n15555), .A2(n14407), .ZN(n15537) );
  NAND2_X1 U17811 ( .A1(n19012), .A2(n16370), .ZN(n14410) );
  OAI211_X1 U17812 ( .C1(n16382), .C2(n14411), .A(n14410), .B(n14409), .ZN(
        n14413) );
  OAI21_X1 U17813 ( .B1(n14416), .B2(n9780), .A(n14415), .ZN(P2_U2995) );
  AOI21_X1 U17814 ( .B1(n20287), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14420), .ZN(n14421) );
  OAI21_X1 U17815 ( .B1(n14582), .B2(n20298), .A(n14421), .ZN(n14422) );
  AOI21_X1 U17816 ( .B1(n14689), .B2(n20293), .A(n14422), .ZN(n14423) );
  OAI21_X1 U17817 ( .B1(n14424), .B2(n20139), .A(n14423), .ZN(P1_U2970) );
  OR2_X1 U17818 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n19396), .ZN(
        n14432) );
  NAND2_X1 U17819 ( .A1(n14425), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15564) );
  NAND2_X1 U17820 ( .A1(n19406), .A2(n14426), .ZN(n14431) );
  OAI21_X1 U17821 ( .B1(n14436), .B2(n19396), .A(n16407), .ZN(n16389) );
  INV_X1 U17822 ( .A(n14427), .ZN(n14428) );
  OR2_X1 U17823 ( .A1(n16389), .A2(n14429), .ZN(n14430) );
  NAND2_X1 U17824 ( .A1(n14432), .A2(n14473), .ZN(n14443) );
  INV_X1 U17825 ( .A(n14433), .ZN(n14435) );
  XNOR2_X1 U17826 ( .A(n14435), .B(n14434), .ZN(n15553) );
  INV_X1 U17827 ( .A(n15553), .ZN(n19046) );
  INV_X1 U17828 ( .A(n15800), .ZN(n15724) );
  NAND2_X1 U17829 ( .A1(n15724), .A2(n14436), .ZN(n16386) );
  OAI22_X1 U17830 ( .A1(n15555), .A2(n19406), .B1(n16329), .B2(n16386), .ZN(
        n14471) );
  NAND3_X1 U17831 ( .A1(n14471), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15749), .ZN(n14441) );
  NAND2_X1 U17832 ( .A1(n14437), .A2(n14438), .ZN(n14439) );
  AND2_X1 U17833 ( .A1(n15430), .A2(n14439), .ZN(n19044) );
  AND2_X1 U17834 ( .A1(n19185), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15548) );
  AOI21_X1 U17835 ( .B1(n19391), .B2(n19044), .A(n15548), .ZN(n14440) );
  OAI211_X1 U17836 ( .C1(n19046), .C2(n16411), .A(n14441), .B(n14440), .ZN(
        n14442) );
  AOI21_X1 U17837 ( .B1(n14443), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n14442), .ZN(n14449) );
  NAND2_X1 U17838 ( .A1(n14445), .A2(n14444), .ZN(n14446) );
  OR2_X1 U17839 ( .A1(n15551), .A2(n19395), .ZN(n14448) );
  NAND2_X1 U17840 ( .A1(n14449), .A2(n14448), .ZN(P2_U3029) );
  NOR2_X1 U17841 ( .A1(n14450), .A2(n14529), .ZN(n14455) );
  INV_X1 U17842 ( .A(n16382), .ZN(n19376) );
  NAND2_X1 U17843 ( .A1(n19376), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14452) );
  OAI211_X1 U17844 ( .C1(n19374), .C2(n14451), .A(n14453), .B(n14452), .ZN(
        n14454) );
  OAI21_X1 U17845 ( .B1(n14458), .B2(n9780), .A(n14457), .ZN(P2_U2983) );
  OR2_X1 U17846 ( .A1(n14460), .A2(n14459), .ZN(n14461) );
  NAND2_X1 U17847 ( .A1(n14437), .A2(n14461), .ZN(n19052) );
  OR2_X1 U17848 ( .A1(n14463), .A2(n14462), .ZN(n14464) );
  NAND2_X1 U17849 ( .A1(n14434), .A2(n14464), .ZN(n15345) );
  INV_X1 U17850 ( .A(n15345), .ZN(n19056) );
  NAND2_X1 U17851 ( .A1(n19402), .A2(n19056), .ZN(n14465) );
  NAND2_X1 U17852 ( .A1(n19365), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15557) );
  OAI211_X1 U17853 ( .C1(n16433), .C2(n19052), .A(n14465), .B(n15557), .ZN(
        n14470) );
  AND2_X1 U17854 ( .A1(n14468), .A2(n14467), .ZN(n15559) );
  NOR3_X1 U17855 ( .A1(n14466), .A2(n15559), .A3(n19395), .ZN(n14469) );
  AOI211_X1 U17856 ( .C1(n15554), .C2(n14471), .A(n14470), .B(n14469), .ZN(
        n14472) );
  OAI21_X1 U17857 ( .B1(n14473), .B2(n15554), .A(n14472), .ZN(P2_U3030) );
  NAND2_X1 U17858 ( .A1(n14478), .A2(n14476), .ZN(n14475) );
  NAND3_X1 U17859 ( .A1(n14475), .A2(n14477), .A3(n14474), .ZN(n15476) );
  NOR2_X1 U17860 ( .A1(n15476), .A2(n15655), .ZN(n15475) );
  AOI21_X1 U17861 ( .B1(n14478), .B2(n14477), .A(n14476), .ZN(n14479) );
  NOR2_X1 U17862 ( .A1(n15475), .A2(n14479), .ZN(n14482) );
  XNOR2_X1 U17863 ( .A(n14480), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14481) );
  XNOR2_X1 U17864 ( .A(n14482), .B(n14481), .ZN(n14498) );
  INV_X1 U17865 ( .A(n15258), .ZN(n14491) );
  NOR2_X1 U17866 ( .A1(n13196), .A2(n20041), .ZN(n14490) );
  AOI21_X1 U17867 ( .B1(n19376), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14490), .ZN(n14483) );
  OAI21_X1 U17868 ( .B1(n19374), .B2(n14484), .A(n14483), .ZN(n14486) );
  OAI21_X1 U17869 ( .B1(n15473), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15467), .ZN(n14488) );
  NOR2_X1 U17870 ( .A1(n14488), .A2(n19385), .ZN(n14485) );
  OAI21_X1 U17871 ( .B1(n14498), .B2(n9780), .A(n14487), .ZN(P2_U2986) );
  INV_X1 U17872 ( .A(n14488), .ZN(n14496) );
  INV_X1 U17873 ( .A(n15643), .ZN(n15650) );
  INV_X1 U17874 ( .A(n15637), .ZN(n15656) );
  NAND3_X1 U17875 ( .A1(n15656), .A2(n15640), .A3(n14489), .ZN(n14493) );
  OAI211_X1 U17876 ( .C1(n15650), .C2(n14494), .A(n14493), .B(n14492), .ZN(
        n14495) );
  AOI21_X1 U17877 ( .B1(n14496), .B2(n16450), .A(n14495), .ZN(n14497) );
  OAI21_X1 U17878 ( .B1(n14498), .B2(n19395), .A(n14497), .ZN(P2_U3018) );
  AOI21_X1 U17879 ( .B1(n20804), .B2(n15150), .A(n14502), .ZN(n14504) );
  OAI22_X1 U17880 ( .A1(n20393), .A2(n14499), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15153), .ZN(n15964) );
  OAI22_X1 U17881 ( .A1(n14500), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n20727), .ZN(n14501) );
  AOI21_X1 U17882 ( .B1(n20804), .B2(n15964), .A(n14501), .ZN(n14503) );
  OAI22_X1 U17883 ( .A1(n14504), .A2(n11802), .B1(n14503), .B2(n14502), .ZN(
        P1_U3474) );
  XOR2_X1 U17884 ( .A(n14505), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n14510)
         );
  OR2_X1 U17885 ( .A1(n14506), .A2(n14006), .ZN(n14508) );
  NAND2_X1 U17886 ( .A1(n14508), .A2(n14507), .ZN(n19179) );
  MUX2_X1 U17887 ( .A(n19179), .B(n11545), .S(n9778), .Z(n14509) );
  OAI21_X1 U17888 ( .B1(n14510), .B2(n15337), .A(n14509), .ZN(P2_U2882) );
  INV_X1 U17889 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n19183) );
  NOR2_X1 U17890 ( .A1(n15319), .A2(n19183), .ZN(n14511) );
  AOI21_X1 U17891 ( .B1(n19370), .B2(n15319), .A(n14511), .ZN(n14512) );
  OAI21_X1 U17892 ( .B1(n19186), .B2(n15337), .A(n14512), .ZN(P2_U2883) );
  NAND2_X1 U17893 ( .A1(n14514), .A2(n14513), .ZN(n15520) );
  INV_X1 U17894 ( .A(n15522), .ZN(n14515) );
  INV_X1 U17895 ( .A(n14517), .ZN(n14519) );
  NAND2_X1 U17896 ( .A1(n14519), .A2(n14518), .ZN(n14520) );
  XNOR2_X1 U17897 ( .A(n14521), .B(n14520), .ZN(n15735) );
  NAND2_X1 U17898 ( .A1(n15513), .A2(n14523), .ZN(n15722) );
  INV_X1 U17899 ( .A(n19382), .ZN(n14529) );
  NAND2_X1 U17900 ( .A1(n16370), .A2(n14524), .ZN(n14525) );
  NAND2_X1 U17901 ( .A1(n19365), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15725) );
  OAI211_X1 U17902 ( .C1(n16382), .C2(n14526), .A(n14525), .B(n15725), .ZN(
        n14527) );
  INV_X1 U17903 ( .A(n14527), .ZN(n14528) );
  INV_X1 U17904 ( .A(n14532), .ZN(n14533) );
  OAI21_X1 U17905 ( .B1(n15735), .B2(n9780), .A(n14533), .ZN(P2_U2993) );
  OAI21_X1 U17906 ( .B1(n14534), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n20120), 
        .ZN(n14535) );
  OAI21_X1 U17907 ( .B1(n14536), .B2(n20120), .A(n14535), .ZN(P2_U3612) );
  NAND2_X1 U17908 ( .A1(n15344), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14537) );
  OAI21_X1 U17909 ( .B1(n14450), .B2(n15344), .A(n14537), .ZN(P2_U2856) );
  AND2_X1 U17910 ( .A1(n14540), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14538) );
  AOI21_X1 U17911 ( .B1(n9773), .B2(P1_EBX_REG_31__SCAN_IN), .A(n14538), .ZN(
        n14542) );
  INV_X1 U17912 ( .A(n14542), .ZN(n14539) );
  NAND2_X1 U17913 ( .A1(n14539), .A2(n13064), .ZN(n14544) );
  AND2_X1 U17914 ( .A1(n14540), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14541) );
  AOI21_X1 U17915 ( .B1(n9773), .B2(P1_EBX_REG_30__SCAN_IN), .A(n14541), .ZN(
        n14571) );
  XNOR2_X1 U17916 ( .A(n14542), .B(n14571), .ZN(n14543) );
  MUX2_X1 U17917 ( .A(n14544), .B(n14543), .S(n14570), .Z(n14955) );
  NAND2_X1 U17918 ( .A1(n14545), .A2(n20185), .ZN(n14563) );
  AND2_X1 U17919 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14553) );
  NAND3_X1 U17920 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n16069) );
  NAND4_X1 U17921 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(P1_REIP_REG_9__SCAN_IN), .A4(P1_REIP_REG_10__SCAN_IN), .ZN(n14546)
         );
  NOR4_X1 U17922 ( .A1(n14548), .A2(n14547), .A3(n16069), .A4(n14546), .ZN(
        n16055) );
  NAND3_X1 U17923 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n14549), .A3(n16055), 
        .ZN(n16042) );
  NOR2_X1 U17924 ( .A1(n14550), .A2(n16042), .ZN(n14662) );
  NAND4_X1 U17925 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .A3(P1_REIP_REG_22__SCAN_IN), .A4(n14662), .ZN(n16029) );
  INV_X1 U17926 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20780) );
  NOR2_X1 U17927 ( .A1(n16029), .A2(n20780), .ZN(n14651) );
  AND2_X1 U17928 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14555) );
  NAND2_X1 U17929 ( .A1(n14651), .A2(n14555), .ZN(n14551) );
  NAND2_X1 U17930 ( .A1(n14551), .A2(n20189), .ZN(n14606) );
  NAND2_X1 U17931 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14557) );
  NAND2_X1 U17932 ( .A1(n20189), .A2(n14557), .ZN(n14552) );
  AND2_X1 U17933 ( .A1(n14606), .A2(n14552), .ZN(n14598) );
  OAI21_X1 U17934 ( .B1(n14553), .B2(n16031), .A(n14598), .ZN(n14573) );
  NOR2_X1 U17935 ( .A1(n20203), .A2(n16042), .ZN(n16028) );
  AND3_X1 U17936 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .A3(P1_REIP_REG_22__SCAN_IN), .ZN(n14554) );
  NAND2_X1 U17937 ( .A1(n16028), .A2(n14554), .ZN(n14652) );
  OR2_X1 U17938 ( .A1(n14652), .A2(n20780), .ZN(n14633) );
  INV_X1 U17939 ( .A(n14555), .ZN(n14556) );
  NOR2_X1 U17940 ( .A1(n14633), .A2(n14556), .ZN(n14607) );
  INV_X1 U17941 ( .A(n14557), .ZN(n14558) );
  NAND2_X1 U17942 ( .A1(n14607), .A2(n14558), .ZN(n14581) );
  INV_X1 U17943 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14810) );
  NOR4_X1 U17944 ( .A1(n14581), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14810), 
        .A4(n21141), .ZN(n14561) );
  INV_X1 U17945 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14687) );
  OAI22_X1 U17946 ( .A1(n20194), .A2(n14687), .B1(n14559), .B2(n20210), .ZN(
        n14560) );
  AOI211_X1 U17947 ( .C1(n14573), .C2(P1_REIP_REG_31__SCAN_IN), .A(n14561), 
        .B(n14560), .ZN(n14562) );
  OAI211_X1 U17948 ( .C1(n14955), .C2(n20191), .A(n14563), .B(n14562), .ZN(
        P1_U2809) );
  INV_X1 U17949 ( .A(n14564), .ZN(n20136) );
  NAND2_X1 U17950 ( .A1(n14565), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n14566)
         );
  NAND3_X1 U17951 ( .A1(n14567), .A2(n20136), .A3(n14566), .ZN(P1_U2801) );
  XNOR2_X1 U17952 ( .A(n14572), .B(n14571), .ZN(n14968) );
  INV_X1 U17953 ( .A(n14812), .ZN(n14577) );
  NOR2_X1 U17954 ( .A1(n14581), .A2(n21141), .ZN(n14574) );
  OAI21_X1 U17955 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14574), .A(n14573), 
        .ZN(n14576) );
  AOI22_X1 U17956 ( .A1(n20206), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20193), .ZN(n14575) );
  OAI211_X1 U17957 ( .C1(n14577), .C2(n20216), .A(n14576), .B(n14575), .ZN(
        n14578) );
  AOI21_X1 U17958 ( .B1(n14968), .B2(n20205), .A(n14578), .ZN(n14579) );
  OAI21_X1 U17959 ( .B1(n14815), .B2(n16117), .A(n14579), .ZN(P1_U2810) );
  NAND2_X1 U17960 ( .A1(n14689), .A2(n20185), .ZN(n14587) );
  INV_X1 U17961 ( .A(n14598), .ZN(n14585) );
  AOI22_X1 U17962 ( .A1(n20206), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20193), .ZN(n14580) );
  OAI21_X1 U17963 ( .B1(n14581), .B2(P1_REIP_REG_29__SCAN_IN), .A(n14580), 
        .ZN(n14584) );
  NOR2_X1 U17964 ( .A1(n20216), .A2(n14582), .ZN(n14583) );
  AOI211_X1 U17965 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(n14585), .A(n14584), 
        .B(n14583), .ZN(n14586) );
  OAI211_X1 U17966 ( .C1(n20191), .C2(n14690), .A(n14587), .B(n14586), .ZN(
        P1_U2811) );
  INV_X1 U17967 ( .A(n14417), .ZN(n14590) );
  AOI21_X1 U17968 ( .B1(n9957), .B2(n14605), .A(n14592), .ZN(n14594) );
  OR2_X1 U17969 ( .A1(n14594), .A2(n14593), .ZN(n14976) );
  INV_X1 U17970 ( .A(n14976), .ZN(n14600) );
  AOI21_X1 U17971 ( .B1(n14607), .B2(P1_REIP_REG_27__SCAN_IN), .A(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14597) );
  INV_X1 U17972 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14692) );
  OAI22_X1 U17973 ( .A1(n20194), .A2(n14692), .B1(n14827), .B2(n20210), .ZN(
        n14595) );
  AOI21_X1 U17974 ( .B1(n20162), .B2(n14825), .A(n14595), .ZN(n14596) );
  OAI21_X1 U17975 ( .B1(n14598), .B2(n14597), .A(n14596), .ZN(n14599) );
  AOI21_X1 U17976 ( .B1(n14600), .B2(n20205), .A(n14599), .ZN(n14601) );
  OAI21_X1 U17977 ( .B1(n14743), .B2(n16117), .A(n14601), .ZN(P1_U2812) );
  AOI21_X1 U17978 ( .B1(n14604), .B2(n14602), .A(n14588), .ZN(n14840) );
  INV_X1 U17979 ( .A(n14840), .ZN(n14748) );
  XNOR2_X1 U17980 ( .A(n14622), .B(n14605), .ZN(n14985) );
  INV_X1 U17981 ( .A(n14606), .ZN(n14619) );
  INV_X1 U17982 ( .A(n14607), .ZN(n14609) );
  AOI22_X1 U17983 ( .A1(n20206), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20193), .ZN(n14608) );
  OAI21_X1 U17984 ( .B1(n14609), .B2(P1_REIP_REG_27__SCAN_IN), .A(n14608), 
        .ZN(n14610) );
  AOI21_X1 U17985 ( .B1(n14619), .B2(P1_REIP_REG_27__SCAN_IN), .A(n14610), 
        .ZN(n14611) );
  OAI21_X1 U17986 ( .B1(n14838), .B2(n20216), .A(n14611), .ZN(n14612) );
  AOI21_X1 U17987 ( .B1(n14985), .B2(n20205), .A(n14612), .ZN(n14613) );
  OAI21_X1 U17988 ( .B1(n14748), .B2(n16117), .A(n14613), .ZN(P1_U2813) );
  NAND2_X1 U17989 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14616) );
  INV_X1 U17990 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20782) );
  OAI21_X1 U17991 ( .B1(n14652), .B2(n14616), .A(n20782), .ZN(n14618) );
  INV_X1 U17992 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14694) );
  OAI22_X1 U17993 ( .A1(n20194), .A2(n14694), .B1(n14845), .B2(n20210), .ZN(
        n14617) );
  AOI21_X1 U17994 ( .B1(n14619), .B2(n14618), .A(n14617), .ZN(n14626) );
  NAND2_X1 U17995 ( .A1(n14632), .A2(n14620), .ZN(n14621) );
  NAND2_X1 U17996 ( .A1(n14622), .A2(n14621), .ZN(n14995) );
  INV_X1 U17997 ( .A(n14849), .ZN(n14623) );
  OAI22_X1 U17998 ( .A1(n14995), .A2(n20191), .B1(n14623), .B2(n20216), .ZN(
        n14624) );
  INV_X1 U17999 ( .A(n14624), .ZN(n14625) );
  OAI211_X1 U18000 ( .C1(n14846), .C2(n16117), .A(n14626), .B(n14625), .ZN(
        P1_U2814) );
  AND2_X1 U18001 ( .A1(n14647), .A2(n14628), .ZN(n14629) );
  OR2_X1 U18002 ( .A1(n14629), .A2(n14614), .ZN(n14757) );
  INV_X1 U18003 ( .A(n14757), .ZN(n14858) );
  NAND2_X1 U18004 ( .A1(n14858), .A2(n20185), .ZN(n14643) );
  OR2_X1 U18005 ( .A1(n14649), .A2(n14630), .ZN(n14631) );
  NAND2_X1 U18006 ( .A1(n14632), .A2(n14631), .ZN(n15006) );
  INV_X1 U18007 ( .A(n15006), .ZN(n14641) );
  NAND2_X1 U18008 ( .A1(n20189), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14639) );
  INV_X1 U18009 ( .A(n14633), .ZN(n14637) );
  INV_X1 U18010 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n14636) );
  INV_X1 U18011 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14695) );
  OAI22_X1 U18012 ( .A1(n20194), .A2(n14695), .B1(n14634), .B2(n20210), .ZN(
        n14635) );
  AOI21_X1 U18013 ( .B1(n14637), .B2(n14636), .A(n14635), .ZN(n14638) );
  OAI21_X1 U18014 ( .B1(n14651), .B2(n14639), .A(n14638), .ZN(n14640) );
  AOI21_X1 U18015 ( .B1(n14641), .B2(n20205), .A(n14640), .ZN(n14642) );
  OAI211_X1 U18016 ( .C1(n20216), .C2(n14856), .A(n14643), .B(n14642), .ZN(
        P1_U2815) );
  NAND2_X1 U18017 ( .A1(n14696), .A2(n14645), .ZN(n14646) );
  NAND2_X1 U18018 ( .A1(n14647), .A2(n14646), .ZN(n14864) );
  AOI21_X1 U18019 ( .B1(n9976), .B2(n14698), .A(n14648), .ZN(n14650) );
  OR2_X1 U18020 ( .A1(n14650), .A2(n14649), .ZN(n15013) );
  INV_X1 U18021 ( .A(n14651), .ZN(n14656) );
  AOI21_X1 U18022 ( .B1(n14652), .B2(n20780), .A(n16031), .ZN(n14655) );
  INV_X1 U18023 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14653) );
  INV_X1 U18024 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14863) );
  OAI22_X1 U18025 ( .A1(n20194), .A2(n14653), .B1(n14863), .B2(n20210), .ZN(
        n14654) );
  AOI21_X1 U18026 ( .B1(n14656), .B2(n14655), .A(n14654), .ZN(n14657) );
  OAI21_X1 U18027 ( .B1(n15013), .B2(n20191), .A(n14657), .ZN(n14658) );
  AOI21_X1 U18028 ( .B1(n14867), .B2(n20162), .A(n14658), .ZN(n14659) );
  OAI21_X1 U18029 ( .B1(n14864), .B2(n16117), .A(n14659), .ZN(P1_U2816) );
  AOI21_X1 U18030 ( .B1(n14661), .B2(n9812), .A(n14660), .ZN(n14880) );
  INV_X1 U18031 ( .A(n14880), .ZN(n14771) );
  NOR2_X1 U18032 ( .A1(n16031), .A2(n14662), .ZN(n16054) );
  NOR2_X1 U18033 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n20203), .ZN(n16043) );
  OAI21_X1 U18034 ( .B1(n16054), .B2(n16043), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14670) );
  NAND2_X1 U18035 ( .A1(n9827), .A2(n14663), .ZN(n14664) );
  NAND2_X1 U18036 ( .A1(n14700), .A2(n14664), .ZN(n15036) );
  INV_X1 U18037 ( .A(n15036), .ZN(n14668) );
  AOI22_X1 U18038 ( .A1(n20162), .A2(n14876), .B1(n20206), .B2(
        P1_EBX_REG_22__SCAN_IN), .ZN(n14666) );
  INV_X1 U18039 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20776) );
  NAND3_X1 U18040 ( .A1(n16028), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n20776), 
        .ZN(n14665) );
  OAI211_X1 U18041 ( .C1(n20210), .C2(n14878), .A(n14666), .B(n14665), .ZN(
        n14667) );
  AOI21_X1 U18042 ( .B1(n20205), .B2(n14668), .A(n14667), .ZN(n14669) );
  OAI211_X1 U18043 ( .C1(n14771), .C2(n16117), .A(n14670), .B(n14669), .ZN(
        P1_U2818) );
  INV_X1 U18044 ( .A(n14671), .ZN(n14674) );
  INV_X1 U18045 ( .A(n14340), .ZN(n14673) );
  AOI21_X1 U18046 ( .B1(n14674), .B2(n14673), .A(n14672), .ZN(n16129) );
  INV_X1 U18047 ( .A(n16129), .ZN(n14806) );
  NAND2_X1 U18048 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n14675) );
  INV_X1 U18049 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20767) );
  OAI21_X1 U18050 ( .B1(n14675), .B2(n16068), .A(n20767), .ZN(n14685) );
  INV_X1 U18051 ( .A(n16069), .ZN(n14676) );
  OAI21_X1 U18052 ( .B1(n16031), .B2(n14676), .A(n16087), .ZN(n16074) );
  INV_X1 U18053 ( .A(n16128), .ZN(n14683) );
  OR2_X1 U18054 ( .A1(n14678), .A2(n14677), .ZN(n14679) );
  AND2_X1 U18055 ( .A1(n15075), .A2(n14679), .ZN(n15092) );
  NOR2_X1 U18056 ( .A1(n20194), .A2(n14727), .ZN(n14681) );
  OAI21_X1 U18057 ( .B1(n20210), .B2(n12370), .A(n20207), .ZN(n14680) );
  AOI211_X1 U18058 ( .C1(n15092), .C2(n20205), .A(n14681), .B(n14680), .ZN(
        n14682) );
  OAI21_X1 U18059 ( .B1(n20216), .B2(n14683), .A(n14682), .ZN(n14684) );
  AOI21_X1 U18060 ( .B1(n14685), .B2(n16074), .A(n14684), .ZN(n14686) );
  OAI21_X1 U18061 ( .B1(n14806), .B2(n16117), .A(n14686), .ZN(P1_U2823) );
  OAI22_X1 U18062 ( .A1(n14955), .A2(n14725), .B1(n20227), .B2(n14687), .ZN(
        P1_U2841) );
  AOI22_X1 U18063 ( .A1(n14968), .A2(n20222), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n14716), .ZN(n14688) );
  INV_X1 U18064 ( .A(n14689), .ZN(n14738) );
  INV_X1 U18065 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14691) );
  OAI222_X1 U18066 ( .A1(n14730), .A2(n14738), .B1(n14691), .B2(n20227), .C1(
        n14690), .C2(n14725), .ZN(P1_U2843) );
  OAI222_X1 U18067 ( .A1(n14730), .A2(n14743), .B1(n14692), .B2(n20227), .C1(
        n14976), .C2(n14725), .ZN(P1_U2844) );
  AOI22_X1 U18068 ( .A1(n14985), .A2(n20222), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n14716), .ZN(n14693) );
  OAI21_X1 U18069 ( .B1(n14748), .B2(n14730), .A(n14693), .ZN(P1_U2845) );
  OAI222_X1 U18070 ( .A1(n14730), .A2(n14757), .B1(n14695), .B2(n20227), .C1(
        n15006), .C2(n14725), .ZN(P1_U2847) );
  OAI222_X1 U18071 ( .A1(n14730), .A2(n14864), .B1(n20227), .B2(n14653), .C1(
        n15013), .C2(n14725), .ZN(P1_U2848) );
  OAI21_X1 U18072 ( .B1(n14660), .B2(n14697), .A(n14696), .ZN(n16036) );
  INV_X1 U18073 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n16027) );
  INV_X1 U18074 ( .A(n14698), .ZN(n14699) );
  XNOR2_X1 U18075 ( .A(n14700), .B(n14699), .ZN(n16037) );
  OAI222_X1 U18076 ( .A1(n16036), .A2(n14701), .B1(n16027), .B2(n20227), .C1(
        n14725), .C2(n16037), .ZN(P1_U2849) );
  INV_X1 U18077 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14702) );
  OAI222_X1 U18078 ( .A1(n14730), .A2(n14771), .B1(n14702), .B2(n20227), .C1(
        n15036), .C2(n14725), .ZN(P1_U2850) );
  OAI21_X1 U18079 ( .B1(n14703), .B2(n14711), .A(n14704), .ZN(n14705) );
  AND2_X1 U18080 ( .A1(n14705), .A2(n9812), .ZN(n16049) );
  INV_X1 U18081 ( .A(n16049), .ZN(n14776) );
  OR2_X1 U18082 ( .A1(n14715), .A2(n14706), .ZN(n14707) );
  NAND2_X1 U18083 ( .A1(n9827), .A2(n14707), .ZN(n16047) );
  OAI22_X1 U18084 ( .A1(n16047), .A2(n14725), .B1(n14708), .B2(n20227), .ZN(
        n14709) );
  INV_X1 U18085 ( .A(n14709), .ZN(n14710) );
  OAI21_X1 U18086 ( .B1(n14776), .B2(n14730), .A(n14710), .ZN(P1_U2851) );
  INV_X1 U18087 ( .A(n14711), .ZN(n14712) );
  XNOR2_X1 U18088 ( .A(n14703), .B(n14712), .ZN(n16053) );
  INV_X1 U18089 ( .A(n16053), .ZN(n14781) );
  AND2_X1 U18090 ( .A1(n14724), .A2(n14713), .ZN(n14714) );
  NOR2_X1 U18091 ( .A1(n14715), .A2(n14714), .ZN(n16052) );
  AOI22_X1 U18092 ( .A1(n16052), .A2(n20222), .B1(P1_EBX_REG_20__SCAN_IN), 
        .B2(n14716), .ZN(n14717) );
  OAI21_X1 U18093 ( .B1(n14781), .B2(n14730), .A(n14717), .ZN(P1_U2852) );
  INV_X1 U18094 ( .A(n14788), .ZN(n14718) );
  NAND2_X1 U18095 ( .A1(n14672), .A2(n14718), .ZN(n14720) );
  NAND2_X1 U18096 ( .A1(n14720), .A2(n14719), .ZN(n14721) );
  AND2_X1 U18097 ( .A1(n14721), .A2(n14703), .ZN(n16067) );
  INV_X1 U18098 ( .A(n16067), .ZN(n14787) );
  INV_X1 U18099 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14726) );
  NAND2_X1 U18100 ( .A1(n9785), .A2(n14722), .ZN(n14723) );
  NAND2_X1 U18101 ( .A1(n14724), .A2(n14723), .ZN(n16072) );
  OAI222_X1 U18102 ( .A1(n14730), .A2(n14787), .B1(n20227), .B2(n14726), .C1(
        n16072), .C2(n14725), .ZN(P1_U2853) );
  NOR2_X1 U18103 ( .A1(n20227), .A2(n14727), .ZN(n14728) );
  AOI21_X1 U18104 ( .B1(n15092), .B2(n20222), .A(n14728), .ZN(n14729) );
  OAI21_X1 U18105 ( .B1(n14806), .B2(n14730), .A(n14729), .ZN(P1_U2855) );
  OAI22_X1 U18106 ( .A1(n14799), .A2(n20267), .B1(n14762), .B2(n14731), .ZN(
        n14732) );
  AOI21_X1 U18107 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n14801), .A(n14732), .ZN(
        n14734) );
  NAND2_X1 U18108 ( .A1(n14802), .A2(DATAI_30_), .ZN(n14733) );
  OAI211_X1 U18109 ( .C1(n14815), .C2(n14805), .A(n14734), .B(n14733), .ZN(
        P1_U2874) );
  OAI22_X1 U18110 ( .A1(n14799), .A2(n20264), .B1(n14762), .B2(n13556), .ZN(
        n14735) );
  AOI21_X1 U18111 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n14801), .A(n14735), .ZN(
        n14737) );
  NAND2_X1 U18112 ( .A1(n14802), .A2(DATAI_29_), .ZN(n14736) );
  OAI211_X1 U18113 ( .C1(n14738), .C2(n14805), .A(n14737), .B(n14736), .ZN(
        P1_U2875) );
  OAI22_X1 U18114 ( .A1(n14799), .A2(n20261), .B1(n14762), .B2(n14739), .ZN(
        n14740) );
  AOI21_X1 U18115 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n14801), .A(n14740), .ZN(
        n14742) );
  NAND2_X1 U18116 ( .A1(n14802), .A2(DATAI_28_), .ZN(n14741) );
  OAI211_X1 U18117 ( .C1(n14743), .C2(n14805), .A(n14742), .B(n14741), .ZN(
        P1_U2876) );
  OAI22_X1 U18118 ( .A1(n14799), .A2(n20258), .B1(n14762), .B2(n14744), .ZN(
        n14745) );
  AOI21_X1 U18119 ( .B1(BUF1_REG_27__SCAN_IN), .B2(n14801), .A(n14745), .ZN(
        n14747) );
  NAND2_X1 U18120 ( .A1(n14802), .A2(DATAI_27_), .ZN(n14746) );
  OAI211_X1 U18121 ( .C1(n14748), .C2(n14805), .A(n14747), .B(n14746), .ZN(
        P1_U2877) );
  OAI22_X1 U18122 ( .A1(n14799), .A2(n20254), .B1(n14762), .B2(n14749), .ZN(
        n14750) );
  AOI21_X1 U18123 ( .B1(BUF1_REG_26__SCAN_IN), .B2(n14801), .A(n14750), .ZN(
        n14752) );
  NAND2_X1 U18124 ( .A1(n14802), .A2(DATAI_26_), .ZN(n14751) );
  OAI211_X1 U18125 ( .C1(n14846), .C2(n14805), .A(n14752), .B(n14751), .ZN(
        P1_U2878) );
  OAI22_X1 U18126 ( .A1(n14799), .A2(n14753), .B1(n14762), .B2(n20882), .ZN(
        n14754) );
  AOI21_X1 U18127 ( .B1(BUF1_REG_25__SCAN_IN), .B2(n14801), .A(n14754), .ZN(
        n14756) );
  NAND2_X1 U18128 ( .A1(n14802), .A2(DATAI_25_), .ZN(n14755) );
  OAI211_X1 U18129 ( .C1(n14757), .C2(n14805), .A(n14756), .B(n14755), .ZN(
        P1_U2879) );
  OAI22_X1 U18130 ( .A1(n14799), .A2(n20251), .B1(n14762), .B2(n13550), .ZN(
        n14758) );
  AOI21_X1 U18131 ( .B1(BUF1_REG_24__SCAN_IN), .B2(n14801), .A(n14758), .ZN(
        n14760) );
  NAND2_X1 U18132 ( .A1(n14802), .A2(DATAI_24_), .ZN(n14759) );
  OAI211_X1 U18133 ( .C1(n14864), .C2(n14805), .A(n14760), .B(n14759), .ZN(
        P1_U2880) );
  OAI22_X1 U18134 ( .A1(n14799), .A2(n14763), .B1(n14762), .B2(n14761), .ZN(
        n14764) );
  AOI21_X1 U18135 ( .B1(n14801), .B2(BUF1_REG_23__SCAN_IN), .A(n14764), .ZN(
        n14766) );
  NAND2_X1 U18136 ( .A1(n14802), .A2(DATAI_23_), .ZN(n14765) );
  OAI211_X1 U18137 ( .C1(n16036), .C2(n14805), .A(n14766), .B(n14765), .ZN(
        P1_U2881) );
  OAI22_X1 U18138 ( .A1(n14799), .A2(n14767), .B1(n14762), .B2(n13672), .ZN(
        n14768) );
  AOI21_X1 U18139 ( .B1(n14801), .B2(BUF1_REG_22__SCAN_IN), .A(n14768), .ZN(
        n14770) );
  NAND2_X1 U18140 ( .A1(n14802), .A2(DATAI_22_), .ZN(n14769) );
  OAI211_X1 U18141 ( .C1(n14771), .C2(n14805), .A(n14770), .B(n14769), .ZN(
        P1_U2882) );
  OAI22_X1 U18142 ( .A1(n14799), .A2(n14772), .B1(n14762), .B2(n13667), .ZN(
        n14773) );
  AOI21_X1 U18143 ( .B1(n14801), .B2(BUF1_REG_21__SCAN_IN), .A(n14773), .ZN(
        n14775) );
  NAND2_X1 U18144 ( .A1(n14802), .A2(DATAI_21_), .ZN(n14774) );
  OAI211_X1 U18145 ( .C1(n14776), .C2(n14805), .A(n14775), .B(n14774), .ZN(
        P1_U2883) );
  OAI22_X1 U18146 ( .A1(n14799), .A2(n14777), .B1(n14762), .B2(n13665), .ZN(
        n14778) );
  AOI21_X1 U18147 ( .B1(n14801), .B2(BUF1_REG_20__SCAN_IN), .A(n14778), .ZN(
        n14780) );
  NAND2_X1 U18148 ( .A1(n14802), .A2(DATAI_20_), .ZN(n14779) );
  OAI211_X1 U18149 ( .C1(n14781), .C2(n14805), .A(n14780), .B(n14779), .ZN(
        P1_U2884) );
  OAI22_X1 U18150 ( .A1(n14799), .A2(n14783), .B1(n14762), .B2(n14782), .ZN(
        n14784) );
  AOI21_X1 U18151 ( .B1(n14801), .B2(BUF1_REG_19__SCAN_IN), .A(n14784), .ZN(
        n14786) );
  NAND2_X1 U18152 ( .A1(n14802), .A2(DATAI_19_), .ZN(n14785) );
  OAI211_X1 U18153 ( .C1(n14787), .C2(n14805), .A(n14786), .B(n14785), .ZN(
        P1_U2885) );
  XNOR2_X1 U18154 ( .A(n14672), .B(n14788), .ZN(n16125) );
  INV_X1 U18155 ( .A(n16125), .ZN(n14796) );
  INV_X1 U18156 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n19426) );
  INV_X1 U18157 ( .A(n14799), .ZN(n14791) );
  AOI22_X1 U18158 ( .A1(n14791), .A2(n14790), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n14789), .ZN(n14792) );
  OAI21_X1 U18159 ( .B1(n19426), .B2(n14793), .A(n14792), .ZN(n14794) );
  AOI21_X1 U18160 ( .B1(n14802), .B2(DATAI_18_), .A(n14794), .ZN(n14795) );
  OAI21_X1 U18161 ( .B1(n14796), .B2(n14805), .A(n14795), .ZN(P1_U2886) );
  OAI22_X1 U18162 ( .A1(n14799), .A2(n14798), .B1(n14762), .B2(n14797), .ZN(
        n14800) );
  AOI21_X1 U18163 ( .B1(n14801), .B2(BUF1_REG_17__SCAN_IN), .A(n14800), .ZN(
        n14804) );
  NAND2_X1 U18164 ( .A1(n14802), .A2(DATAI_17_), .ZN(n14803) );
  OAI211_X1 U18165 ( .C1(n14806), .C2(n14805), .A(n14804), .B(n14803), .ZN(
        P1_U2887) );
  NAND2_X1 U18166 ( .A1(n14966), .A2(n20294), .ZN(n14814) );
  NOR2_X1 U18167 ( .A1(n20207), .A2(n14810), .ZN(n14967) );
  NOR2_X1 U18168 ( .A1(n14950), .A2(n21154), .ZN(n14811) );
  AOI211_X1 U18169 ( .C1(n14812), .C2(n16141), .A(n14967), .B(n14811), .ZN(
        n14813) );
  OAI211_X1 U18170 ( .C1(n14954), .C2(n14815), .A(n14814), .B(n14813), .ZN(
        P1_U2969) );
  INV_X1 U18171 ( .A(n14820), .ZN(n14819) );
  NOR4_X1 U18172 ( .A1(n14817), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14818) );
  NAND2_X1 U18173 ( .A1(n14819), .A2(n14818), .ZN(n14822) );
  NAND3_X1 U18174 ( .A1(n14820), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14821) );
  NAND2_X1 U18175 ( .A1(n14825), .A2(n16141), .ZN(n14826) );
  NAND2_X1 U18176 ( .A1(n20299), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14975) );
  OAI211_X1 U18177 ( .C1(n14950), .C2(n14827), .A(n14826), .B(n14975), .ZN(
        n14828) );
  AOI21_X1 U18178 ( .B1(n14829), .B2(n20293), .A(n14828), .ZN(n14830) );
  OAI21_X1 U18179 ( .B1(n20139), .B2(n14983), .A(n14830), .ZN(P1_U2971) );
  NOR2_X1 U18180 ( .A1(n14832), .A2(n14831), .ZN(n14835) );
  INV_X1 U18181 ( .A(n14833), .ZN(n14834) );
  MUX2_X1 U18182 ( .A(n14835), .B(n14834), .S(n15089), .Z(n14836) );
  XNOR2_X1 U18183 ( .A(n14836), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14992) );
  INV_X1 U18184 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21163) );
  NOR2_X1 U18185 ( .A1(n20207), .A2(n21163), .ZN(n14984) );
  AOI21_X1 U18186 ( .B1(n20287), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14984), .ZN(n14837) );
  OAI21_X1 U18187 ( .B1(n14838), .B2(n20298), .A(n14837), .ZN(n14839) );
  AOI21_X1 U18188 ( .B1(n14840), .B2(n20293), .A(n14839), .ZN(n14841) );
  OAI21_X1 U18189 ( .B1(n20139), .B2(n14992), .A(n14841), .ZN(P1_U2972) );
  NAND2_X1 U18190 ( .A1(n14843), .A2(n14842), .ZN(n14844) );
  XOR2_X1 U18191 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n14844), .Z(
        n15003) );
  NAND2_X1 U18192 ( .A1(n20299), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14994) );
  OAI21_X1 U18193 ( .B1(n14950), .B2(n14845), .A(n14994), .ZN(n14848) );
  NOR2_X1 U18194 ( .A1(n14846), .A2(n14954), .ZN(n14847) );
  OAI21_X1 U18195 ( .B1(n20139), .B2(n15003), .A(n14850), .ZN(P1_U2973) );
  INV_X1 U18196 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21064) );
  MUX2_X1 U18197 ( .A(n15016), .B(n14852), .S(n15089), .Z(n14853) );
  AOI21_X1 U18198 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14861), .A(
        n14853), .ZN(n14854) );
  XNOR2_X1 U18199 ( .A(n14854), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15011) );
  NAND2_X1 U18200 ( .A1(n20299), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n15005) );
  NAND2_X1 U18201 ( .A1(n20287), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14855) );
  OAI211_X1 U18202 ( .C1(n14856), .C2(n20298), .A(n15005), .B(n14855), .ZN(
        n14857) );
  AOI21_X1 U18203 ( .B1(n14858), .B2(n20293), .A(n14857), .ZN(n14859) );
  OAI21_X1 U18204 ( .B1(n15011), .B2(n20139), .A(n14859), .ZN(P1_U2974) );
  MUX2_X1 U18205 ( .A(n14861), .B(n14860), .S(n15089), .Z(n14862) );
  XNOR2_X1 U18206 ( .A(n14862), .B(n15016), .ZN(n15024) );
  NAND2_X1 U18207 ( .A1(n20299), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15012) );
  OAI21_X1 U18208 ( .B1(n14950), .B2(n14863), .A(n15012), .ZN(n14866) );
  NOR2_X1 U18209 ( .A1(n14864), .A2(n14954), .ZN(n14865) );
  AOI211_X1 U18210 ( .C1(n16141), .C2(n14867), .A(n14866), .B(n14865), .ZN(
        n14868) );
  OAI21_X1 U18211 ( .B1(n20139), .B2(n15024), .A(n14868), .ZN(P1_U2975) );
  XNOR2_X1 U18212 ( .A(n15089), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14869) );
  XNOR2_X1 U18213 ( .A(n14816), .B(n14869), .ZN(n15026) );
  NAND2_X1 U18214 ( .A1(n15026), .A2(n20294), .ZN(n14872) );
  INV_X1 U18215 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20778) );
  NOR2_X1 U18216 ( .A1(n20207), .A2(n20778), .ZN(n15028) );
  NOR2_X1 U18217 ( .A1(n16026), .A2(n20298), .ZN(n14870) );
  AOI211_X1 U18218 ( .C1(n20287), .C2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15028), .B(n14870), .ZN(n14871) );
  OAI211_X1 U18219 ( .C1(n14954), .C2(n16036), .A(n14872), .B(n14871), .ZN(
        P1_U2976) );
  NAND2_X1 U18220 ( .A1(n14874), .A2(n14873), .ZN(n14875) );
  XOR2_X1 U18221 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n14875), .Z(
        n15040) );
  NAND2_X1 U18222 ( .A1(n14876), .A2(n16141), .ZN(n14877) );
  NAND2_X1 U18223 ( .A1(n20299), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15034) );
  OAI211_X1 U18224 ( .C1(n14950), .C2(n14878), .A(n14877), .B(n15034), .ZN(
        n14879) );
  AOI21_X1 U18225 ( .B1(n14880), .B2(n20293), .A(n14879), .ZN(n14881) );
  OAI21_X1 U18226 ( .B1(n15040), .B2(n20139), .A(n14881), .ZN(P1_U2977) );
  NOR3_X1 U18227 ( .A1(n14882), .A2(n15089), .A3(n12067), .ZN(n14885) );
  NOR3_X1 U18228 ( .A1(n10118), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n14896), .ZN(n14884) );
  NOR2_X1 U18229 ( .A1(n14885), .A2(n14884), .ZN(n14891) );
  NOR2_X1 U18230 ( .A1(n14891), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14890) );
  AOI22_X1 U18231 ( .A1(n14890), .A2(n15089), .B1(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n14885), .ZN(n14886) );
  XNOR2_X1 U18232 ( .A(n14886), .B(n15045), .ZN(n15048) );
  NAND2_X1 U18233 ( .A1(n20299), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15042) );
  NAND2_X1 U18234 ( .A1(n20287), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14887) );
  OAI211_X1 U18235 ( .C1(n16051), .C2(n20298), .A(n15042), .B(n14887), .ZN(
        n14888) );
  AOI21_X1 U18236 ( .B1(n16049), .B2(n20293), .A(n14888), .ZN(n14889) );
  OAI21_X1 U18237 ( .B1(n15048), .B2(n20139), .A(n14889), .ZN(P1_U2978) );
  AOI21_X1 U18238 ( .B1(n14891), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14890), .ZN(n15062) );
  NAND2_X1 U18239 ( .A1(n16141), .A2(n16056), .ZN(n14892) );
  NAND2_X1 U18240 ( .A1(n20299), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15049) );
  OAI211_X1 U18241 ( .C1(n14950), .C2(n14893), .A(n14892), .B(n15049), .ZN(
        n14894) );
  AOI21_X1 U18242 ( .B1(n16053), .B2(n20293), .A(n14894), .ZN(n14895) );
  OAI21_X1 U18243 ( .B1(n15062), .B2(n20139), .A(n14895), .ZN(P1_U2979) );
  MUX2_X1 U18244 ( .A(n15089), .B(n14896), .S(n14882), .Z(n14897) );
  XOR2_X1 U18245 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n14897), .Z(
        n15069) );
  AOI22_X1 U18246 ( .A1(n20287), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n20299), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n14898) );
  OAI21_X1 U18247 ( .B1(n20298), .B2(n16065), .A(n14898), .ZN(n14899) );
  AOI21_X1 U18248 ( .B1(n16067), .B2(n20293), .A(n14899), .ZN(n14900) );
  OAI21_X1 U18249 ( .B1(n15069), .B2(n20139), .A(n14900), .ZN(P1_U2980) );
  OAI21_X1 U18250 ( .B1(n10118), .B2(n14901), .A(n14882), .ZN(n15083) );
  NAND2_X1 U18251 ( .A1(n16141), .A2(n16079), .ZN(n14902) );
  NAND2_X1 U18252 ( .A1(n20299), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15078) );
  OAI211_X1 U18253 ( .C1(n14950), .C2(n16076), .A(n14902), .B(n15078), .ZN(
        n14903) );
  AOI21_X1 U18254 ( .B1(n16125), .B2(n20293), .A(n14903), .ZN(n14904) );
  OAI21_X1 U18255 ( .B1(n20139), .B2(n15083), .A(n14904), .ZN(P1_U2981) );
  OAI211_X1 U18256 ( .C1(n14905), .C2(n14907), .A(n14906), .B(n14917), .ZN(
        n15110) );
  NAND2_X1 U18257 ( .A1(n15110), .A2(n15108), .ZN(n15113) );
  NAND2_X1 U18258 ( .A1(n15113), .A2(n15109), .ZN(n14908) );
  XOR2_X1 U18259 ( .A(n14909), .B(n14908), .Z(n15106) );
  NAND2_X1 U18260 ( .A1(n15106), .A2(n20294), .ZN(n14915) );
  INV_X1 U18261 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14910) );
  OR2_X1 U18262 ( .A1(n20207), .A2(n14910), .ZN(n15101) );
  OAI21_X1 U18263 ( .B1(n14950), .B2(n14911), .A(n15101), .ZN(n14912) );
  AOI21_X1 U18264 ( .B1(n14913), .B2(n16141), .A(n14912), .ZN(n14914) );
  OAI211_X1 U18265 ( .C1(n14954), .C2(n14916), .A(n14915), .B(n14914), .ZN(
        P1_U2983) );
  NAND2_X1 U18266 ( .A1(n14905), .A2(n14917), .ZN(n14921) );
  INV_X1 U18267 ( .A(n14918), .ZN(n14919) );
  AOI21_X1 U18268 ( .B1(n14921), .B2(n14920), .A(n14919), .ZN(n14924) );
  MUX2_X1 U18269 ( .A(n14922), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .S(
        n15138), .Z(n14923) );
  XNOR2_X1 U18270 ( .A(n14924), .B(n14923), .ZN(n16168) );
  NAND2_X1 U18271 ( .A1(n16168), .A2(n20294), .ZN(n14930) );
  INV_X1 U18272 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n14925) );
  OAI22_X1 U18273 ( .A1(n14950), .A2(n14926), .B1(n20207), .B2(n14925), .ZN(
        n14927) );
  AOI21_X1 U18274 ( .B1(n14928), .B2(n16141), .A(n14927), .ZN(n14929) );
  OAI211_X1 U18275 ( .C1(n14954), .C2(n14931), .A(n14930), .B(n14929), .ZN(
        P1_U2985) );
  INV_X1 U18276 ( .A(n14905), .ZN(n15139) );
  INV_X1 U18277 ( .A(n14932), .ZN(n14933) );
  AOI21_X1 U18278 ( .B1(n15139), .B2(n14934), .A(n14933), .ZN(n15121) );
  AND2_X1 U18279 ( .A1(n14935), .A2(n14936), .ZN(n15120) );
  NAND2_X1 U18280 ( .A1(n15121), .A2(n15120), .ZN(n15119) );
  NAND2_X1 U18281 ( .A1(n15119), .A2(n14936), .ZN(n14937) );
  XOR2_X1 U18282 ( .A(n14938), .B(n14937), .Z(n16178) );
  NAND2_X1 U18283 ( .A1(n16178), .A2(n20294), .ZN(n14943) );
  INV_X1 U18284 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n14939) );
  NOR2_X1 U18285 ( .A1(n20207), .A2(n14939), .ZN(n16172) );
  AND2_X1 U18286 ( .A1(n20287), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14940) );
  AOI211_X1 U18287 ( .C1(n14941), .C2(n16141), .A(n16172), .B(n14940), .ZN(
        n14942) );
  OAI211_X1 U18288 ( .C1(n14954), .C2(n14944), .A(n14943), .B(n14942), .ZN(
        P1_U2986) );
  NAND2_X1 U18289 ( .A1(n14945), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14947) );
  XNOR2_X1 U18290 ( .A(n15139), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14946) );
  MUX2_X1 U18291 ( .A(n14947), .B(n14946), .S(n15138), .Z(n14948) );
  OR3_X1 U18292 ( .A1(n14945), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15138), .ZN(n15140) );
  NAND2_X1 U18293 ( .A1(n14948), .A2(n15140), .ZN(n16187) );
  NAND2_X1 U18294 ( .A1(n16187), .A2(n20294), .ZN(n14953) );
  INV_X1 U18295 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14949) );
  NOR2_X1 U18296 ( .A1(n20207), .A2(n14949), .ZN(n16184) );
  NOR2_X1 U18297 ( .A1(n14950), .A2(n16113), .ZN(n14951) );
  AOI211_X1 U18298 ( .C1(n16141), .C2(n16120), .A(n16184), .B(n14951), .ZN(
        n14952) );
  OAI211_X1 U18299 ( .C1(n14954), .C2(n16118), .A(n14953), .B(n14952), .ZN(
        P1_U2989) );
  INV_X1 U18300 ( .A(n14955), .ZN(n14960) );
  INV_X1 U18301 ( .A(n14956), .ZN(n14959) );
  NAND3_X1 U18302 ( .A1(n14990), .A2(n14957), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14969) );
  NOR3_X1 U18303 ( .A1(n14969), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12075), .ZN(n14958) );
  AOI211_X1 U18304 ( .C1(n14960), .C2(n20312), .A(n14959), .B(n14958), .ZN(
        n14964) );
  OAI211_X1 U18305 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15100), .A(
        n14961), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14970) );
  NAND3_X1 U18306 ( .A1(n14970), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14962), .ZN(n14963) );
  OAI211_X1 U18307 ( .C1(n14965), .C2(n15137), .A(n14964), .B(n14963), .ZN(
        P1_U3000) );
  INV_X1 U18308 ( .A(n14966), .ZN(n14974) );
  AOI21_X1 U18309 ( .B1(n14968), .B2(n20312), .A(n14967), .ZN(n14973) );
  INV_X1 U18310 ( .A(n14969), .ZN(n14971) );
  OAI21_X1 U18311 ( .B1(n14971), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n14970), .ZN(n14972) );
  OAI211_X1 U18312 ( .C1(n14974), .C2(n15137), .A(n14973), .B(n14972), .ZN(
        P1_U3001) );
  INV_X1 U18313 ( .A(n14987), .ZN(n14978) );
  OAI21_X1 U18314 ( .B1(n14976), .B2(n16218), .A(n14975), .ZN(n14977) );
  AOI21_X1 U18315 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n14978), .A(
        n14977), .ZN(n14982) );
  NAND3_X1 U18316 ( .A1(n14990), .A2(n14980), .A3(n14979), .ZN(n14981) );
  OAI211_X1 U18317 ( .C1(n14983), .C2(n15137), .A(n14982), .B(n14981), .ZN(
        P1_U3003) );
  AOI21_X1 U18318 ( .B1(n14985), .B2(n20312), .A(n14984), .ZN(n14986) );
  OAI21_X1 U18319 ( .B1(n14987), .B2(n14989), .A(n14986), .ZN(n14988) );
  AOI21_X1 U18320 ( .B1(n14990), .B2(n14989), .A(n14988), .ZN(n14991) );
  OAI21_X1 U18321 ( .B1(n14992), .B2(n15137), .A(n14991), .ZN(P1_U3004) );
  NOR2_X1 U18322 ( .A1(n14993), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15001) );
  OAI21_X1 U18323 ( .B1(n14995), .B2(n16218), .A(n14994), .ZN(n15000) );
  NAND3_X1 U18324 ( .A1(n15025), .A2(n14997), .A3(n14996), .ZN(n15009) );
  AOI21_X1 U18325 ( .B1(n15009), .B2(n15004), .A(n14998), .ZN(n14999) );
  AOI211_X1 U18326 ( .C1(n15025), .C2(n15001), .A(n15000), .B(n14999), .ZN(
        n15002) );
  OAI21_X1 U18327 ( .B1(n15003), .B2(n15137), .A(n15002), .ZN(P1_U3005) );
  INV_X1 U18328 ( .A(n15004), .ZN(n15008) );
  OAI21_X1 U18329 ( .B1(n15006), .B2(n16218), .A(n15005), .ZN(n15007) );
  AOI21_X1 U18330 ( .B1(n15008), .B2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15007), .ZN(n15010) );
  OAI211_X1 U18331 ( .C1(n15011), .C2(n15137), .A(n15010), .B(n15009), .ZN(
        P1_U3006) );
  OAI21_X1 U18332 ( .B1(n15013), .B2(n16218), .A(n15012), .ZN(n15014) );
  AOI21_X1 U18333 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15015), .A(
        n15014), .ZN(n15023) );
  INV_X1 U18334 ( .A(n15046), .ZN(n15017) );
  OAI21_X1 U18335 ( .B1(n15017), .B2(n21064), .A(n15016), .ZN(n15021) );
  OAI21_X1 U18336 ( .B1(n15018), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15019) );
  NAND3_X1 U18337 ( .A1(n15021), .A2(n15020), .A3(n15019), .ZN(n15022) );
  OAI211_X1 U18338 ( .C1(n15024), .C2(n15137), .A(n15023), .B(n15022), .ZN(
        P1_U3007) );
  INV_X1 U18339 ( .A(n15025), .ZN(n15032) );
  NAND2_X1 U18340 ( .A1(n15026), .A2(n20318), .ZN(n15031) );
  NOR2_X1 U18341 ( .A1(n16037), .A2(n16218), .ZN(n15027) );
  AOI211_X1 U18342 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n15029), .A(
        n15028), .B(n15027), .ZN(n15030) );
  OAI211_X1 U18343 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n15032), .A(
        n15031), .B(n15030), .ZN(P1_U3008) );
  XNOR2_X1 U18344 ( .A(n15045), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15038) );
  INV_X1 U18345 ( .A(n15041), .ZN(n15033) );
  NAND2_X1 U18346 ( .A1(n15033), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15035) );
  OAI211_X1 U18347 ( .C1(n16218), .C2(n15036), .A(n15035), .B(n15034), .ZN(
        n15037) );
  AOI21_X1 U18348 ( .B1(n15046), .B2(n15038), .A(n15037), .ZN(n15039) );
  OAI21_X1 U18349 ( .B1(n15040), .B2(n15137), .A(n15039), .ZN(P1_U3009) );
  NOR2_X1 U18350 ( .A1(n15041), .A2(n15045), .ZN(n15044) );
  OAI21_X1 U18351 ( .B1(n16047), .B2(n16218), .A(n15042), .ZN(n15043) );
  AOI211_X1 U18352 ( .C1(n15046), .C2(n15045), .A(n15044), .B(n15043), .ZN(
        n15047) );
  OAI21_X1 U18353 ( .B1(n15048), .B2(n15137), .A(n15047), .ZN(P1_U3010) );
  INV_X1 U18354 ( .A(n15049), .ZN(n15058) );
  NOR2_X1 U18355 ( .A1(n15050), .A2(n16176), .ZN(n15053) );
  AOI22_X1 U18356 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15053), .B1(
        n15052), .B2(n15051), .ZN(n16174) );
  INV_X1 U18357 ( .A(n16174), .ZN(n15055) );
  INV_X1 U18358 ( .A(n16175), .ZN(n15054) );
  OAI21_X1 U18359 ( .B1(n15055), .B2(n15054), .A(n12067), .ZN(n15056) );
  AOI21_X1 U18360 ( .B1(n15056), .B2(n15063), .A(n15059), .ZN(n15057) );
  AOI211_X1 U18361 ( .C1(n20312), .C2(n16052), .A(n15058), .B(n15057), .ZN(
        n15061) );
  NAND3_X1 U18362 ( .A1(n15067), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n15059), .ZN(n15060) );
  OAI211_X1 U18363 ( .C1(n15062), .C2(n15137), .A(n15061), .B(n15060), .ZN(
        P1_U3011) );
  NOR2_X1 U18364 ( .A1(n15063), .A2(n12067), .ZN(n15066) );
  NAND2_X1 U18365 ( .A1(n20299), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n15064) );
  OAI21_X1 U18366 ( .B1(n16072), .B2(n16218), .A(n15064), .ZN(n15065) );
  AOI211_X1 U18367 ( .C1(n15067), .C2(n12067), .A(n15066), .B(n15065), .ZN(
        n15068) );
  OAI21_X1 U18368 ( .B1(n15069), .B2(n15137), .A(n15068), .ZN(P1_U3012) );
  OAI22_X1 U18369 ( .A1(n15124), .A2(n15071), .B1(n15070), .B2(n20314), .ZN(
        n15072) );
  NOR2_X1 U18370 ( .A1(n15073), .A2(n15072), .ZN(n16182) );
  OAI21_X1 U18371 ( .B1(n15100), .B2(n15074), .A(n16182), .ZN(n15095) );
  INV_X1 U18372 ( .A(n15076), .ZN(n15077) );
  OAI21_X1 U18373 ( .B1(n9969), .B2(n15077), .A(n9785), .ZN(n16073) );
  OAI21_X1 U18374 ( .B1(n16073), .B2(n16218), .A(n15078), .ZN(n15081) );
  INV_X1 U18375 ( .A(n15093), .ZN(n16171) );
  NOR3_X1 U18376 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15079), .A3(
        n16171), .ZN(n15080) );
  AOI211_X1 U18377 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n15095), .A(
        n15081), .B(n15080), .ZN(n15082) );
  OAI21_X1 U18378 ( .B1(n15083), .B2(n15137), .A(n15082), .ZN(P1_U3013) );
  NAND2_X1 U18379 ( .A1(n15089), .A2(n15084), .ZN(n15088) );
  OAI21_X1 U18380 ( .B1(n15139), .B2(n15086), .A(n15085), .ZN(n15087) );
  MUX2_X1 U18381 ( .A(n15089), .B(n15088), .S(n15087), .Z(n15091) );
  XNOR2_X1 U18382 ( .A(n15091), .B(n15090), .ZN(n16132) );
  AOI22_X1 U18383 ( .A1(n15092), .A2(n20312), .B1(n20299), .B2(
        P1_REIP_REG_17__SCAN_IN), .ZN(n15098) );
  NAND2_X1 U18384 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15094) );
  NAND2_X1 U18385 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15093), .ZN(
        n15099) );
  OAI21_X1 U18386 ( .B1(n15094), .B2(n15099), .A(n15090), .ZN(n15096) );
  NAND2_X1 U18387 ( .A1(n15096), .A2(n15095), .ZN(n15097) );
  OAI211_X1 U18388 ( .C1(n16132), .C2(n15137), .A(n15098), .B(n15097), .ZN(
        P1_U3014) );
  NOR3_X1 U18389 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n12058), .A3(
        n15099), .ZN(n15105) );
  NOR2_X1 U18390 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15099), .ZN(
        n15116) );
  OAI21_X1 U18391 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15100), .A(
        n16182), .ZN(n15114) );
  OAI21_X1 U18392 ( .B1(n15116), .B2(n15114), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15102) );
  OAI211_X1 U18393 ( .C1(n15103), .C2(n16218), .A(n15102), .B(n15101), .ZN(
        n15104) );
  AOI211_X1 U18394 ( .C1(n15106), .C2(n20318), .A(n15105), .B(n15104), .ZN(
        n15107) );
  INV_X1 U18395 ( .A(n15107), .ZN(P1_U3015) );
  INV_X1 U18396 ( .A(n15109), .ZN(n15112) );
  AND2_X1 U18397 ( .A1(n15109), .A2(n15108), .ZN(n15111) );
  OAI22_X1 U18398 ( .A1(n15113), .A2(n15112), .B1(n15111), .B2(n15110), .ZN(
        n16138) );
  AOI22_X1 U18399 ( .A1(n20299), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15114), .ZN(n15115) );
  INV_X1 U18400 ( .A(n15115), .ZN(n15117) );
  AOI211_X1 U18401 ( .C1(n20312), .C2(n16082), .A(n15117), .B(n15116), .ZN(
        n15118) );
  OAI21_X1 U18402 ( .B1(n16138), .B2(n15137), .A(n15118), .ZN(P1_U3016) );
  OAI21_X1 U18403 ( .B1(n15121), .B2(n15120), .A(n15119), .ZN(n15122) );
  INV_X1 U18404 ( .A(n15122), .ZN(n16144) );
  INV_X1 U18405 ( .A(n15123), .ZN(n15130) );
  INV_X1 U18406 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15143) );
  NAND2_X1 U18407 ( .A1(n15125), .A2(n15143), .ZN(n15145) );
  AOI21_X1 U18408 ( .B1(n15126), .B2(n15125), .A(n15124), .ZN(n15128) );
  AOI211_X1 U18409 ( .C1(n15129), .C2(n15131), .A(n15128), .B(n15127), .ZN(
        n15144) );
  OAI21_X1 U18410 ( .B1(n15130), .B2(n15145), .A(n15144), .ZN(n15133) );
  OAI21_X1 U18411 ( .B1(n15131), .B2(n16204), .A(n15134), .ZN(n15132) );
  OAI21_X1 U18412 ( .B1(n15134), .B2(n15133), .A(n15132), .ZN(n15136) );
  AOI22_X1 U18413 ( .A1(n16097), .A2(n20312), .B1(n20299), .B2(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15135) );
  OAI211_X1 U18414 ( .C1(n16144), .C2(n15137), .A(n15136), .B(n15135), .ZN(
        P1_U3019) );
  NAND3_X1 U18415 ( .A1(n15139), .A2(n15138), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15141) );
  NAND2_X1 U18416 ( .A1(n15141), .A2(n15140), .ZN(n15142) );
  XNOR2_X1 U18417 ( .A(n15142), .B(n15143), .ZN(n16146) );
  OAI22_X1 U18418 ( .A1(n16204), .A2(n15145), .B1(n15144), .B2(n15143), .ZN(
        n15148) );
  INV_X1 U18419 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15146) );
  OAI22_X1 U18420 ( .A1(n16103), .A2(n16218), .B1(n20207), .B2(n15146), .ZN(
        n15147) );
  AOI211_X1 U18421 ( .C1(n16146), .C2(n20318), .A(n15148), .B(n15147), .ZN(
        n15149) );
  INV_X1 U18422 ( .A(n15149), .ZN(P1_U3020) );
  INV_X1 U18423 ( .A(n15150), .ZN(n15966) );
  NAND2_X1 U18424 ( .A1(n15152), .A2(n15151), .ZN(n15156) );
  OAI22_X1 U18425 ( .A1(n15966), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n15156), .B2(n15153), .ZN(n15154) );
  AOI21_X1 U18426 ( .B1(n20437), .B2(n15155), .A(n15154), .ZN(n15967) );
  INV_X1 U18427 ( .A(n20804), .ZN(n15162) );
  INV_X1 U18428 ( .A(n15156), .ZN(n15160) );
  INV_X1 U18429 ( .A(n15157), .ZN(n15158) );
  AOI22_X1 U18430 ( .A1(n20803), .A2(n15160), .B1(n15159), .B2(n15158), .ZN(
        n15161) );
  OAI21_X1 U18431 ( .B1(n15967), .B2(n15162), .A(n15161), .ZN(n15163) );
  MUX2_X1 U18432 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15163), .S(
        n20807), .Z(P1_U3473) );
  INV_X1 U18433 ( .A(n20331), .ZN(n15164) );
  NAND2_X1 U18434 ( .A1(n15164), .A2(n20332), .ZN(n20519) );
  OAI21_X1 U18435 ( .B1(n20623), .B2(n20639), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15168) );
  NAND2_X1 U18436 ( .A1(n15168), .A2(n20809), .ZN(n15173) );
  NAND2_X1 U18437 ( .A1(n20665), .A2(n20518), .ZN(n15172) );
  INV_X1 U18438 ( .A(n15172), .ZN(n15169) );
  NAND3_X1 U18439 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20517), .ZN(n15208) );
  NOR2_X1 U18440 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15208), .ZN(
        n20631) );
  OAI22_X1 U18441 ( .A1(n15173), .A2(n15169), .B1(n20631), .B2(n20526), .ZN(
        n15170) );
  AOI211_X2 U18442 ( .C1(n20519), .C2(P1_STATE2_REG_2__SCAN_IN), .A(n15171), 
        .B(n15170), .ZN(n20628) );
  INV_X1 U18443 ( .A(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15182) );
  OAI22_X1 U18444 ( .A1(n15173), .A2(n15172), .B1(n20519), .B2(n20432), .ZN(
        n20632) );
  NOR2_X2 U18445 ( .A1(n15175), .A2(n15174), .ZN(n20670) );
  AOI22_X1 U18446 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n15176), .B1(DATAI_24_), 
        .B2(n15177), .ZN(n20679) );
  AOI22_X1 U18447 ( .A1(DATAI_16_), .A2(n15177), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n15176), .ZN(n20646) );
  INV_X1 U18448 ( .A(n20646), .ZN(n20676) );
  NOR2_X2 U18449 ( .A1(n15178), .A2(n11788), .ZN(n20669) );
  AOI22_X1 U18450 ( .A1(n20639), .A2(n20676), .B1(n20631), .B2(n20669), .ZN(
        n15179) );
  OAI21_X1 U18451 ( .B1(n20679), .B2(n20636), .A(n15179), .ZN(n15180) );
  AOI21_X1 U18452 ( .B1(n20632), .B2(n20670), .A(n15180), .ZN(n15181) );
  OAI21_X1 U18453 ( .B1(n20628), .B2(n15182), .A(n15181), .ZN(P1_U3129) );
  INV_X1 U18454 ( .A(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15186) );
  AOI22_X1 U18455 ( .A1(n20639), .A2(n20682), .B1(n20631), .B2(n20680), .ZN(
        n15183) );
  OAI21_X1 U18456 ( .B1(n20685), .B2(n20636), .A(n15183), .ZN(n15184) );
  AOI21_X1 U18457 ( .B1(n20632), .B2(n20681), .A(n15184), .ZN(n15185) );
  OAI21_X1 U18458 ( .B1(n20628), .B2(n15186), .A(n15185), .ZN(P1_U3130) );
  INV_X1 U18459 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15190) );
  INV_X1 U18460 ( .A(n20654), .ZN(n20688) );
  AOI22_X1 U18461 ( .A1(n20639), .A2(n20688), .B1(n20631), .B2(n20686), .ZN(
        n15187) );
  OAI21_X1 U18462 ( .B1(n20691), .B2(n20636), .A(n15187), .ZN(n15188) );
  AOI21_X1 U18463 ( .B1(n20632), .B2(n20687), .A(n15188), .ZN(n15189) );
  OAI21_X1 U18464 ( .B1(n20628), .B2(n15190), .A(n15189), .ZN(P1_U3131) );
  INV_X1 U18465 ( .A(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15194) );
  AOI22_X1 U18466 ( .A1(n20639), .A2(n20706), .B1(n20631), .B2(n20704), .ZN(
        n15191) );
  OAI21_X1 U18467 ( .B1(n20709), .B2(n20636), .A(n15191), .ZN(n15192) );
  AOI21_X1 U18468 ( .B1(n20632), .B2(n20705), .A(n15192), .ZN(n15193) );
  OAI21_X1 U18469 ( .B1(n20628), .B2(n15194), .A(n15193), .ZN(P1_U3134) );
  INV_X1 U18470 ( .A(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15198) );
  AOI22_X1 U18471 ( .A1(n20639), .A2(n20712), .B1(n20631), .B2(n20710), .ZN(
        n15195) );
  OAI21_X1 U18472 ( .B1(n20715), .B2(n20636), .A(n15195), .ZN(n15196) );
  AOI21_X1 U18473 ( .B1(n20632), .B2(n20711), .A(n15196), .ZN(n15197) );
  OAI21_X1 U18474 ( .B1(n20628), .B2(n15198), .A(n15197), .ZN(P1_U3135) );
  INV_X1 U18475 ( .A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15202) );
  AOI22_X1 U18476 ( .A1(n20639), .A2(n20720), .B1(n20631), .B2(n20716), .ZN(
        n15199) );
  OAI21_X1 U18477 ( .B1(n20726), .B2(n20636), .A(n15199), .ZN(n15200) );
  AOI21_X1 U18478 ( .B1(n20632), .B2(n20719), .A(n15200), .ZN(n15201) );
  OAI21_X1 U18479 ( .B1(n20628), .B2(n15202), .A(n15201), .ZN(P1_U3136) );
  NAND2_X1 U18480 ( .A1(n20811), .A2(n20810), .ZN(n15204) );
  INV_X1 U18481 ( .A(n20673), .ZN(n15203) );
  AOI21_X1 U18482 ( .B1(n15204), .B2(n15208), .A(n15203), .ZN(n20642) );
  NAND2_X1 U18483 ( .A1(n15236), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n15215) );
  NAND2_X1 U18484 ( .A1(n20665), .A2(n20548), .ZN(n15206) );
  NOR2_X1 U18485 ( .A1(n20547), .A2(n15208), .ZN(n20637) );
  INV_X1 U18486 ( .A(n20637), .ZN(n15205) );
  NAND2_X1 U18487 ( .A1(n15206), .A2(n15205), .ZN(n15207) );
  NAND2_X1 U18488 ( .A1(n15207), .A2(n20809), .ZN(n15211) );
  INV_X1 U18489 ( .A(n15208), .ZN(n15209) );
  NAND2_X1 U18490 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15209), .ZN(n15210) );
  NAND2_X1 U18491 ( .A1(n15211), .A2(n15210), .ZN(n20638) );
  AOI22_X1 U18492 ( .A1(n20681), .A2(n20638), .B1(n20680), .B2(n20637), .ZN(
        n15214) );
  NAND2_X1 U18493 ( .A1(n20658), .A2(n20682), .ZN(n15213) );
  INV_X1 U18494 ( .A(n20685), .ZN(n20647) );
  NAND2_X1 U18495 ( .A1(n20639), .A2(n20647), .ZN(n15212) );
  NAND4_X1 U18496 ( .A1(n15215), .A2(n15214), .A3(n15213), .A4(n15212), .ZN(
        P1_U3138) );
  NAND2_X1 U18497 ( .A1(n15236), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n15219) );
  AOI22_X1 U18498 ( .A1(n20687), .A2(n20638), .B1(n20686), .B2(n20637), .ZN(
        n15218) );
  NAND2_X1 U18499 ( .A1(n20658), .A2(n20688), .ZN(n15217) );
  NAND2_X1 U18500 ( .A1(n20639), .A2(n20651), .ZN(n15216) );
  NAND4_X1 U18501 ( .A1(n15219), .A2(n15218), .A3(n15217), .A4(n15216), .ZN(
        P1_U3139) );
  NAND2_X1 U18502 ( .A1(n15236), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n15223) );
  AOI22_X1 U18503 ( .A1(n20693), .A2(n20638), .B1(n20692), .B2(n20637), .ZN(
        n15222) );
  NAND2_X1 U18504 ( .A1(n20658), .A2(n20694), .ZN(n15221) );
  NAND2_X1 U18505 ( .A1(n20639), .A2(n20608), .ZN(n15220) );
  NAND4_X1 U18506 ( .A1(n15223), .A2(n15222), .A3(n15221), .A4(n15220), .ZN(
        P1_U3140) );
  NAND2_X1 U18507 ( .A1(n15236), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n15227) );
  AOI22_X1 U18508 ( .A1(n20699), .A2(n20638), .B1(n20698), .B2(n20637), .ZN(
        n15226) );
  INV_X1 U18509 ( .A(n20581), .ZN(n20700) );
  NAND2_X1 U18510 ( .A1(n20658), .A2(n20700), .ZN(n15225) );
  NAND2_X1 U18511 ( .A1(n20639), .A2(n20578), .ZN(n15224) );
  NAND4_X1 U18512 ( .A1(n15227), .A2(n15226), .A3(n15225), .A4(n15224), .ZN(
        P1_U3141) );
  NAND2_X1 U18513 ( .A1(n15236), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n15231) );
  AOI22_X1 U18514 ( .A1(n20705), .A2(n20638), .B1(n20704), .B2(n20637), .ZN(
        n15230) );
  NAND2_X1 U18515 ( .A1(n20658), .A2(n20706), .ZN(n15229) );
  NAND2_X1 U18516 ( .A1(n20639), .A2(n20614), .ZN(n15228) );
  NAND4_X1 U18517 ( .A1(n15231), .A2(n15230), .A3(n15229), .A4(n15228), .ZN(
        P1_U3142) );
  NAND2_X1 U18518 ( .A1(n15236), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n15235) );
  AOI22_X1 U18519 ( .A1(n20711), .A2(n20638), .B1(n20710), .B2(n20637), .ZN(
        n15234) );
  NAND2_X1 U18520 ( .A1(n20658), .A2(n20712), .ZN(n15233) );
  NAND2_X1 U18521 ( .A1(n20639), .A2(n20657), .ZN(n15232) );
  NAND4_X1 U18522 ( .A1(n15235), .A2(n15234), .A3(n15233), .A4(n15232), .ZN(
        P1_U3143) );
  NAND2_X1 U18523 ( .A1(n15236), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n15240) );
  AOI22_X1 U18524 ( .A1(n20719), .A2(n20638), .B1(n20716), .B2(n20637), .ZN(
        n15239) );
  NAND2_X1 U18525 ( .A1(n20658), .A2(n20720), .ZN(n15238) );
  NAND2_X1 U18526 ( .A1(n20639), .A2(n20587), .ZN(n15237) );
  NAND4_X1 U18527 ( .A1(n15240), .A2(n15239), .A3(n15238), .A4(n15237), .ZN(
        P1_U3144) );
  INV_X1 U18528 ( .A(n15241), .ZN(n15244) );
  INV_X1 U18529 ( .A(n15242), .ZN(n15243) );
  OR2_X1 U18530 ( .A1(n15248), .A2(n15247), .ZN(n15346) );
  NAND3_X1 U18531 ( .A1(n15346), .A2(n15341), .A3(n15249), .ZN(n15251) );
  NAND2_X1 U18532 ( .A1(n15344), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15250) );
  OAI211_X1 U18533 ( .C1(n15344), .C2(n10229), .A(n15251), .B(n15250), .ZN(
        P2_U2858) );
  NOR2_X1 U18534 ( .A1(n15253), .A2(n15252), .ZN(n15255) );
  XNOR2_X1 U18535 ( .A(n15255), .B(n15254), .ZN(n15361) );
  NAND2_X1 U18536 ( .A1(n15361), .A2(n15341), .ZN(n15257) );
  NAND2_X1 U18537 ( .A1(n15344), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15256) );
  OAI211_X1 U18538 ( .C1(n15344), .C2(n15258), .A(n15257), .B(n15256), .ZN(
        P2_U2859) );
  OAI21_X1 U18539 ( .B1(n15261), .B2(n15260), .A(n15259), .ZN(n15363) );
  OAI21_X1 U18540 ( .B1(n15262), .B2(n15263), .A(n13288), .ZN(n16266) );
  NOR2_X1 U18541 ( .A1(n16266), .A2(n15344), .ZN(n15264) );
  AOI21_X1 U18542 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n9778), .A(n15264), .ZN(
        n15265) );
  OAI21_X1 U18543 ( .B1(n15363), .B2(n15337), .A(n15265), .ZN(P2_U2860) );
  OAI21_X1 U18544 ( .B1(n15268), .B2(n15267), .A(n15266), .ZN(n15379) );
  NOR2_X1 U18545 ( .A1(n15269), .A2(n15270), .ZN(n15271) );
  OR2_X1 U18546 ( .A1(n15262), .A2(n15271), .ZN(n15660) );
  NOR2_X1 U18547 ( .A1(n15660), .A2(n15344), .ZN(n15272) );
  AOI21_X1 U18548 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n15344), .A(n15272), .ZN(
        n15273) );
  OAI21_X1 U18549 ( .B1(n15379), .B2(n15337), .A(n15273), .ZN(P2_U2861) );
  OAI21_X1 U18550 ( .B1(n15276), .B2(n15275), .A(n15274), .ZN(n15389) );
  AND2_X1 U18551 ( .A1(n10230), .A2(n15277), .ZN(n15278) );
  OR2_X1 U18552 ( .A1(n15278), .A2(n15269), .ZN(n15671) );
  MUX2_X1 U18553 ( .A(n15671), .B(n20930), .S(n15344), .Z(n15279) );
  OAI21_X1 U18554 ( .B1(n15389), .B2(n15337), .A(n15279), .ZN(P2_U2862) );
  AOI21_X1 U18555 ( .B1(n15282), .B2(n15281), .A(n15280), .ZN(n15283) );
  XOR2_X1 U18556 ( .A(n15284), .B(n15283), .Z(n15397) );
  NAND2_X1 U18557 ( .A1(n15344), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n15289) );
  NAND2_X1 U18558 ( .A1(n15285), .A2(n15286), .ZN(n15287) );
  NAND2_X1 U18559 ( .A1(n16324), .A2(n15319), .ZN(n15288) );
  OAI211_X1 U18560 ( .C1(n15397), .C2(n15337), .A(n15289), .B(n15288), .ZN(
        P2_U2863) );
  AND2_X1 U18561 ( .A1(n15301), .A2(n15300), .ZN(n15303) );
  OR2_X1 U18562 ( .A1(n15303), .A2(n15290), .ZN(n15291) );
  NAND2_X1 U18563 ( .A1(n15285), .A2(n15291), .ZN(n16311) );
  AOI21_X1 U18564 ( .B1(n15294), .B2(n15293), .A(n15292), .ZN(n16317) );
  NAND2_X1 U18565 ( .A1(n16317), .A2(n15341), .ZN(n15296) );
  NAND2_X1 U18566 ( .A1(n15344), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15295) );
  OAI211_X1 U18567 ( .C1(n16311), .C2(n15344), .A(n15296), .B(n15295), .ZN(
        P2_U2864) );
  NAND2_X1 U18568 ( .A1(n15332), .A2(n15298), .ZN(n15307) );
  AOI21_X1 U18569 ( .B1(n15299), .B2(n15307), .A(n9811), .ZN(n15398) );
  NAND2_X1 U18570 ( .A1(n15398), .A2(n15341), .ZN(n15305) );
  NOR2_X1 U18571 ( .A1(n15301), .A2(n15300), .ZN(n15302) );
  NAND2_X1 U18572 ( .A1(n15962), .A2(n15319), .ZN(n15304) );
  OAI211_X1 U18573 ( .C1(n15319), .C2(n15954), .A(n15305), .B(n15304), .ZN(
        P2_U2865) );
  NAND2_X1 U18574 ( .A1(n15332), .A2(n15326), .ZN(n15325) );
  INV_X1 U18575 ( .A(n15325), .ZN(n15322) );
  OAI21_X1 U18576 ( .B1(n15313), .B2(n15308), .A(n15307), .ZN(n15413) );
  NAND2_X1 U18577 ( .A1(n15344), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n15311) );
  NAND2_X1 U18578 ( .A1(n15727), .A2(n15319), .ZN(n15310) );
  OAI211_X1 U18579 ( .C1(n15413), .C2(n15337), .A(n15311), .B(n15310), .ZN(
        P2_U2866) );
  OR2_X1 U18580 ( .A1(n15325), .A2(n15312), .ZN(n15320) );
  AOI21_X1 U18581 ( .B1(n15314), .B2(n15320), .A(n15313), .ZN(n15420) );
  NAND2_X1 U18582 ( .A1(n15420), .A2(n15341), .ZN(n15318) );
  AOI21_X1 U18583 ( .B1(n15316), .B2(n14398), .A(n11607), .ZN(n19008) );
  NAND2_X1 U18584 ( .A1(n19008), .A2(n15319), .ZN(n15317) );
  OAI211_X1 U18585 ( .C1(n15319), .C2(n11605), .A(n15318), .B(n15317), .ZN(
        P2_U2867) );
  OAI21_X1 U18586 ( .B1(n15322), .B2(n15321), .A(n15320), .ZN(n15428) );
  MUX2_X1 U18587 ( .A(n19022), .B(n15323), .S(n15344), .Z(n15324) );
  OAI21_X1 U18588 ( .B1(n15428), .B2(n15337), .A(n15324), .ZN(P2_U2868) );
  OAI21_X1 U18589 ( .B1(n15332), .B2(n15326), .A(n15325), .ZN(n15438) );
  AND2_X1 U18590 ( .A1(n15328), .A2(n15327), .ZN(n15330) );
  OR2_X1 U18591 ( .A1(n15330), .A2(n15329), .ZN(n15541) );
  MUX2_X1 U18592 ( .A(n15541), .B(n11598), .S(n15344), .Z(n15331) );
  OAI21_X1 U18593 ( .B1(n15438), .B2(n15337), .A(n15331), .ZN(P2_U2869) );
  INV_X1 U18594 ( .A(n15332), .ZN(n15333) );
  OAI21_X1 U18595 ( .B1(n15338), .B2(n15334), .A(n15333), .ZN(n15445) );
  NOR2_X1 U18596 ( .A1(n19046), .A2(n15344), .ZN(n15335) );
  AOI21_X1 U18597 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n15344), .A(n15335), .ZN(
        n15336) );
  OAI21_X1 U18598 ( .B1(n15445), .B2(n15337), .A(n15336), .ZN(P2_U2870) );
  AOI21_X1 U18599 ( .B1(n15340), .B2(n15339), .A(n15338), .ZN(n15449) );
  NAND2_X1 U18600 ( .A1(n15449), .A2(n15341), .ZN(n15343) );
  NAND2_X1 U18601 ( .A1(n15344), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n15342) );
  OAI211_X1 U18602 ( .C1(n15345), .C2(n15344), .A(n15343), .B(n15342), .ZN(
        P2_U2871) );
  NAND3_X1 U18603 ( .A1(n15346), .A2(n15249), .A3(n10867), .ZN(n15355) );
  MUX2_X1 U18604 ( .A(BUF1_REG_13__SCAN_IN), .B(BUF2_REG_13__SCAN_IN), .S(
        n15878), .Z(n19354) );
  AOI22_X1 U18605 ( .A1(n16315), .A2(n19354), .B1(n19262), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n15354) );
  AOI22_X1 U18606 ( .A1(n19215), .A2(BUF2_REG_29__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n15353) );
  INV_X1 U18607 ( .A(n15347), .ZN(n15351) );
  INV_X1 U18608 ( .A(n15348), .ZN(n15350) );
  NAND2_X1 U18609 ( .A1(n16255), .A2(n19263), .ZN(n15352) );
  NAND4_X1 U18610 ( .A1(n15355), .A2(n15354), .A3(n15353), .A4(n15352), .ZN(
        P2_U2890) );
  AOI22_X1 U18611 ( .A1(n16315), .A2(n15356), .B1(n19262), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n15358) );
  AOI22_X1 U18612 ( .A1(n19215), .A2(BUF2_REG_28__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15357) );
  OAI211_X1 U18613 ( .C1(n15359), .C2(n19272), .A(n15358), .B(n15357), .ZN(
        n15360) );
  AOI21_X1 U18614 ( .B1(n15361), .B2(n10867), .A(n15360), .ZN(n15362) );
  INV_X1 U18615 ( .A(n15362), .ZN(P2_U2891) );
  OR2_X1 U18616 ( .A1(n15363), .A2(n19275), .ZN(n15370) );
  AOI22_X1 U18617 ( .A1(n16315), .A2(n19229), .B1(n19262), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n15369) );
  AOI22_X1 U18618 ( .A1(n19215), .A2(BUF2_REG_27__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15368) );
  AND2_X1 U18619 ( .A1(n15373), .A2(n15364), .ZN(n15365) );
  NOR2_X1 U18620 ( .A1(n15366), .A2(n15365), .ZN(n16269) );
  NAND2_X1 U18621 ( .A1(n16269), .A2(n19263), .ZN(n15367) );
  NAND4_X1 U18622 ( .A1(n15370), .A2(n15369), .A3(n15368), .A4(n15367), .ZN(
        P2_U2892) );
  NAND2_X1 U18623 ( .A1(n15383), .A2(n15371), .ZN(n15372) );
  NAND2_X1 U18624 ( .A1(n15373), .A2(n15372), .ZN(n16277) );
  AOI22_X1 U18625 ( .A1(n16315), .A2(n15374), .B1(n19262), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15376) );
  AOI22_X1 U18626 ( .A1(n19215), .A2(BUF2_REG_26__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15375) );
  OAI211_X1 U18627 ( .C1(n16277), .C2(n19272), .A(n15376), .B(n15375), .ZN(
        n15377) );
  INV_X1 U18628 ( .A(n15377), .ZN(n15378) );
  OAI21_X1 U18629 ( .B1(n15379), .B2(n19275), .A(n15378), .ZN(P2_U2893) );
  NAND2_X1 U18630 ( .A1(n15380), .A2(n15381), .ZN(n15382) );
  NAND2_X1 U18631 ( .A1(n15383), .A2(n15382), .ZN(n16292) );
  AOI22_X1 U18632 ( .A1(n16315), .A2(n15384), .B1(n19262), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n15386) );
  AOI22_X1 U18633 ( .A1(n19215), .A2(BUF2_REG_25__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15385) );
  OAI211_X1 U18634 ( .C1(n16292), .C2(n19272), .A(n15386), .B(n15385), .ZN(
        n15387) );
  INV_X1 U18635 ( .A(n15387), .ZN(n15388) );
  OAI21_X1 U18636 ( .B1(n15389), .B2(n19275), .A(n15388), .ZN(P2_U2894) );
  OR2_X1 U18637 ( .A1(n9782), .A2(n15390), .ZN(n15391) );
  NAND2_X1 U18638 ( .A1(n15380), .A2(n15391), .ZN(n16304) );
  AOI22_X1 U18639 ( .A1(n19215), .A2(BUF2_REG_24__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15394) );
  AOI22_X1 U18640 ( .A1(n16315), .A2(n15392), .B1(n19262), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n15393) );
  OAI211_X1 U18641 ( .C1(n19272), .C2(n16304), .A(n15394), .B(n15393), .ZN(
        n15395) );
  INV_X1 U18642 ( .A(n15395), .ZN(n15396) );
  OAI21_X1 U18643 ( .B1(n15397), .B2(n19275), .A(n15396), .ZN(P2_U2895) );
  INV_X1 U18644 ( .A(n15398), .ZN(n15407) );
  AND2_X1 U18645 ( .A1(n15400), .A2(n15399), .ZN(n15401) );
  OR2_X1 U18646 ( .A1(n15401), .A2(n9781), .ZN(n15959) );
  INV_X1 U18647 ( .A(n15959), .ZN(n15404) );
  INV_X1 U18648 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n19307) );
  OAI22_X1 U18649 ( .A1(n15402), .A2(n19443), .B1(n19270), .B2(n19307), .ZN(
        n15403) );
  AOI21_X1 U18650 ( .B1(n19263), .B2(n15404), .A(n15403), .ZN(n15406) );
  AOI22_X1 U18651 ( .A1(n19215), .A2(BUF2_REG_22__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n15405) );
  OAI211_X1 U18652 ( .C1(n15407), .C2(n19275), .A(n15406), .B(n15405), .ZN(
        P2_U2897) );
  AOI22_X1 U18653 ( .A1(n19215), .A2(BUF2_REG_21__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n15410) );
  AOI22_X1 U18654 ( .A1(n16315), .A2(n15408), .B1(n19262), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15409) );
  OAI211_X1 U18655 ( .C1(n19272), .C2(n9821), .A(n15410), .B(n15409), .ZN(
        n15411) );
  INV_X1 U18656 ( .A(n15411), .ZN(n15412) );
  OAI21_X1 U18657 ( .B1(n15413), .B2(n19275), .A(n15412), .ZN(P2_U2898) );
  OR2_X1 U18658 ( .A1(n15415), .A2(n15414), .ZN(n15416) );
  NAND2_X1 U18659 ( .A1(n13244), .A2(n15416), .ZN(n19005) );
  AOI22_X1 U18660 ( .A1(n19215), .A2(BUF2_REG_20__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n15418) );
  AOI22_X1 U18661 ( .A1(n16315), .A2(n19436), .B1(n19262), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n15417) );
  OAI211_X1 U18662 ( .C1(n19272), .C2(n19005), .A(n15418), .B(n15417), .ZN(
        n15419) );
  AOI21_X1 U18663 ( .B1(n15420), .B2(n10867), .A(n15419), .ZN(n15421) );
  INV_X1 U18664 ( .A(n15421), .ZN(P2_U2899) );
  AOI22_X1 U18665 ( .A1(n19215), .A2(BUF2_REG_19__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n15424) );
  AOI22_X1 U18666 ( .A1(n16315), .A2(n15422), .B1(n19262), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n15423) );
  OAI211_X1 U18667 ( .C1(n19272), .C2(n15425), .A(n15424), .B(n15423), .ZN(
        n15426) );
  INV_X1 U18668 ( .A(n15426), .ZN(n15427) );
  OAI21_X1 U18669 ( .B1(n15428), .B2(n19275), .A(n15427), .ZN(P2_U2900) );
  NAND2_X1 U18670 ( .A1(n15430), .A2(n15429), .ZN(n15431) );
  NAND2_X1 U18671 ( .A1(n15432), .A2(n15431), .ZN(n19033) );
  AOI22_X1 U18672 ( .A1(n19215), .A2(BUF2_REG_18__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n15435) );
  AOI22_X1 U18673 ( .A1(n16315), .A2(n15433), .B1(n19262), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n15434) );
  OAI211_X1 U18674 ( .C1(n19272), .C2(n19033), .A(n15435), .B(n15434), .ZN(
        n15436) );
  INV_X1 U18675 ( .A(n15436), .ZN(n15437) );
  OAI21_X1 U18676 ( .B1(n15438), .B2(n19275), .A(n15437), .ZN(P2_U2901) );
  INV_X1 U18677 ( .A(n19044), .ZN(n15442) );
  AOI22_X1 U18678 ( .A1(n19215), .A2(BUF2_REG_17__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n15441) );
  AOI22_X1 U18679 ( .A1(n16315), .A2(n15439), .B1(n19262), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n15440) );
  OAI211_X1 U18680 ( .C1(n19272), .C2(n15442), .A(n15441), .B(n15440), .ZN(
        n15443) );
  INV_X1 U18681 ( .A(n15443), .ZN(n15444) );
  OAI21_X1 U18682 ( .B1(n15445), .B2(n19275), .A(n15444), .ZN(P2_U2902) );
  AOI22_X1 U18683 ( .A1(n19215), .A2(BUF2_REG_16__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n15447) );
  AOI22_X1 U18684 ( .A1(n16315), .A2(n19281), .B1(n19262), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n15446) );
  OAI211_X1 U18685 ( .C1(n19272), .C2(n19052), .A(n15447), .B(n15446), .ZN(
        n15448) );
  AOI21_X1 U18686 ( .B1(n15449), .B2(n10867), .A(n15448), .ZN(n15450) );
  INV_X1 U18687 ( .A(n15450), .ZN(P2_U2903) );
  NAND2_X1 U18688 ( .A1(n15451), .A2(n15463), .ZN(n15456) );
  INV_X1 U18689 ( .A(n15452), .ZN(n15453) );
  NOR2_X1 U18690 ( .A1(n15454), .A2(n15453), .ZN(n15455) );
  XNOR2_X1 U18691 ( .A(n15456), .B(n15455), .ZN(n15634) );
  INV_X1 U18692 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n15458) );
  NOR2_X1 U18693 ( .A1(n13196), .A2(n15458), .ZN(n15626) );
  NOR2_X1 U18694 ( .A1(n19374), .A2(n16246), .ZN(n15459) );
  AOI211_X1 U18695 ( .C1(n19376), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15626), .B(n15459), .ZN(n15460) );
  OAI21_X1 U18696 ( .B1(n15630), .B2(n14529), .A(n15460), .ZN(n15461) );
  AOI21_X1 U18697 ( .B1(n15632), .B2(n16378), .A(n15461), .ZN(n15462) );
  OAI21_X1 U18698 ( .B1(n15634), .B2(n9780), .A(n15462), .ZN(P2_U2984) );
  NAND2_X1 U18699 ( .A1(n15464), .A2(n15463), .ZN(n15466) );
  XOR2_X1 U18700 ( .A(n15466), .B(n15465), .Z(n15647) );
  AOI21_X1 U18701 ( .B1(n15639), .B2(n15467), .A(n15457), .ZN(n15644) );
  NAND2_X1 U18702 ( .A1(n19365), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15636) );
  OAI21_X1 U18703 ( .B1(n16382), .B2(n15468), .A(n15636), .ZN(n15469) );
  AOI21_X1 U18704 ( .B1(n16370), .B2(n16253), .A(n15469), .ZN(n15470) );
  OAI21_X1 U18705 ( .B1(n10229), .B2(n14529), .A(n15470), .ZN(n15471) );
  AOI21_X1 U18706 ( .B1(n15644), .B2(n16378), .A(n15471), .ZN(n15472) );
  OAI21_X1 U18707 ( .B1(n15647), .B2(n9780), .A(n15472), .ZN(P2_U2985) );
  INV_X1 U18708 ( .A(n15473), .ZN(n15474) );
  OAI21_X1 U18709 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n9798), .A(
        n15474), .ZN(n15659) );
  INV_X1 U18710 ( .A(n15475), .ZN(n15649) );
  NAND2_X1 U18711 ( .A1(n15476), .A2(n15655), .ZN(n15648) );
  NAND3_X1 U18712 ( .A1(n15649), .A2(n16379), .A3(n15648), .ZN(n15480) );
  NAND2_X1 U18713 ( .A1(n19365), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15652) );
  OAI21_X1 U18714 ( .B1(n16382), .B2(n16261), .A(n15652), .ZN(n15478) );
  NOR2_X1 U18715 ( .A1(n16266), .A2(n14529), .ZN(n15477) );
  AOI211_X1 U18716 ( .C1(n16370), .C2(n16260), .A(n15478), .B(n15477), .ZN(
        n15479) );
  OAI211_X1 U18717 ( .C1(n19385), .C2(n15659), .A(n15480), .B(n15479), .ZN(
        P2_U2987) );
  OAI21_X1 U18718 ( .B1(n9894), .B2(n15488), .A(n15489), .ZN(n15481) );
  XOR2_X1 U18719 ( .A(n15482), .B(n15481), .Z(n15670) );
  AOI21_X1 U18720 ( .B1(n15662), .B2(n15493), .A(n9798), .ZN(n15668) );
  NOR2_X1 U18721 ( .A1(n15660), .A2(n14529), .ZN(n15486) );
  NAND2_X1 U18722 ( .A1(n19365), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15661) );
  NAND2_X1 U18723 ( .A1(n19376), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15483) );
  OAI211_X1 U18724 ( .C1(n19374), .C2(n15484), .A(n15661), .B(n15483), .ZN(
        n15485) );
  AOI211_X1 U18725 ( .C1(n15668), .C2(n16378), .A(n15486), .B(n15485), .ZN(
        n15487) );
  OAI21_X1 U18726 ( .B1(n15670), .B2(n9780), .A(n15487), .ZN(P2_U2988) );
  INV_X1 U18727 ( .A(n15488), .ZN(n15490) );
  NAND2_X1 U18728 ( .A1(n15490), .A2(n15489), .ZN(n15491) );
  XNOR2_X1 U18729 ( .A(n15492), .B(n15491), .ZN(n15681) );
  INV_X1 U18730 ( .A(n15493), .ZN(n15494) );
  AOI21_X1 U18731 ( .B1(n20936), .B2(n15695), .A(n15494), .ZN(n15679) );
  NAND2_X1 U18732 ( .A1(n19185), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15672) );
  OAI21_X1 U18733 ( .B1(n16382), .B2(n15495), .A(n15672), .ZN(n15496) );
  AOI21_X1 U18734 ( .B1(n16370), .B2(n16284), .A(n15496), .ZN(n15497) );
  OAI21_X1 U18735 ( .B1(n15671), .B2(n14529), .A(n15497), .ZN(n15498) );
  AOI21_X1 U18736 ( .B1(n15679), .B2(n16378), .A(n15498), .ZN(n15499) );
  OAI21_X1 U18737 ( .B1(n15681), .B2(n9780), .A(n15499), .ZN(P2_U2989) );
  OAI21_X1 U18738 ( .B1(n15512), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15693), .ZN(n15711) );
  INV_X1 U18739 ( .A(n16311), .ZN(n15702) );
  NAND2_X1 U18740 ( .A1(n16370), .A2(n16307), .ZN(n15500) );
  NAND2_X1 U18741 ( .A1(n19365), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15700) );
  OAI211_X1 U18742 ( .C1(n16382), .C2(n15501), .A(n15500), .B(n15700), .ZN(
        n15507) );
  NAND2_X1 U18743 ( .A1(n15502), .A2(n15509), .ZN(n15503) );
  NAND2_X1 U18744 ( .A1(n15503), .A2(n15510), .ZN(n15505) );
  NOR2_X1 U18745 ( .A1(n15505), .A2(n15504), .ZN(n15706) );
  AND2_X1 U18746 ( .A1(n15505), .A2(n15504), .ZN(n15705) );
  NOR3_X1 U18747 ( .A1(n15706), .A2(n15705), .A3(n19379), .ZN(n15506) );
  AOI211_X1 U18748 ( .C1(n19382), .C2(n15702), .A(n15507), .B(n15506), .ZN(
        n15508) );
  OAI21_X1 U18749 ( .B1(n15711), .B2(n19385), .A(n15508), .ZN(P2_U2991) );
  NAND2_X1 U18750 ( .A1(n15510), .A2(n15509), .ZN(n15511) );
  XOR2_X1 U18751 ( .A(n15511), .B(n15502), .Z(n15721) );
  AOI21_X1 U18752 ( .B1(n15717), .B2(n15513), .A(n15512), .ZN(n15712) );
  NAND2_X1 U18753 ( .A1(n15712), .A2(n16378), .ZN(n15518) );
  INV_X1 U18754 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20029) );
  NOR2_X1 U18755 ( .A1(n13196), .A2(n20029), .ZN(n15714) );
  AOI21_X1 U18756 ( .B1(n19376), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15714), .ZN(n15514) );
  OAI21_X1 U18757 ( .B1(n19374), .B2(n15515), .A(n15514), .ZN(n15516) );
  AOI21_X1 U18758 ( .B1(n15962), .B2(n19382), .A(n15516), .ZN(n15517) );
  OAI211_X1 U18759 ( .C1(n15721), .C2(n9780), .A(n15518), .B(n15517), .ZN(
        P2_U2992) );
  NAND2_X1 U18760 ( .A1(n15520), .A2(n15519), .ZN(n15524) );
  NAND2_X1 U18761 ( .A1(n15522), .A2(n15521), .ZN(n15523) );
  XNOR2_X1 U18762 ( .A(n15524), .B(n15523), .ZN(n15745) );
  AOI21_X1 U18763 ( .B1(n15526), .B2(n9789), .A(n15525), .ZN(n15743) );
  NAND2_X1 U18764 ( .A1(n19008), .A2(n19382), .ZN(n15528) );
  NOR2_X1 U18765 ( .A1(n13196), .A2(n20025), .ZN(n15739) );
  AOI21_X1 U18766 ( .B1(n19376), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15739), .ZN(n15527) );
  OAI211_X1 U18767 ( .C1(n19374), .C2(n15529), .A(n15528), .B(n15527), .ZN(
        n15530) );
  AOI21_X1 U18768 ( .B1(n15743), .B2(n16378), .A(n15530), .ZN(n15531) );
  OAI21_X1 U18769 ( .B1(n15745), .B2(n9780), .A(n15531), .ZN(P2_U2994) );
  NOR2_X1 U18770 ( .A1(n15533), .A2(n15532), .ZN(n15534) );
  XNOR2_X1 U18771 ( .A(n15535), .B(n15534), .ZN(n15756) );
  INV_X1 U18772 ( .A(n15547), .ZN(n15536) );
  AOI21_X1 U18773 ( .B1(n15536), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15538) );
  INV_X1 U18774 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15539) );
  NAND2_X1 U18775 ( .A1(n19365), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n15746) );
  OAI21_X1 U18776 ( .B1(n16382), .B2(n15539), .A(n15746), .ZN(n15540) );
  INV_X1 U18777 ( .A(n15540), .ZN(n15543) );
  NAND2_X1 U18778 ( .A1(n19382), .A2(n19031), .ZN(n15542) );
  OAI211_X1 U18779 ( .C1(n19374), .C2(n15544), .A(n15543), .B(n15542), .ZN(
        n15545) );
  AOI21_X1 U18780 ( .B1(n15753), .B2(n16378), .A(n15545), .ZN(n15546) );
  OAI21_X1 U18781 ( .B1(n15756), .B2(n9780), .A(n15546), .ZN(P2_U2996) );
  INV_X1 U18782 ( .A(n19036), .ZN(n15550) );
  AOI21_X1 U18783 ( .B1(n19376), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15548), .ZN(n15549) );
  OAI21_X1 U18784 ( .B1(n15550), .B2(n19374), .A(n15549), .ZN(n15552) );
  XNOR2_X1 U18785 ( .A(n15555), .B(n15554), .ZN(n15563) );
  INV_X1 U18786 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n19059) );
  INV_X1 U18787 ( .A(n19051), .ZN(n15556) );
  NAND2_X1 U18788 ( .A1(n16370), .A2(n15556), .ZN(n15558) );
  OAI211_X1 U18789 ( .C1(n19059), .C2(n16382), .A(n15558), .B(n15557), .ZN(
        n15561) );
  NOR3_X1 U18790 ( .A1(n14466), .A2(n15559), .A3(n19379), .ZN(n15560) );
  AOI211_X1 U18791 ( .C1(n19382), .C2(n19056), .A(n15561), .B(n15560), .ZN(
        n15562) );
  OAI21_X1 U18792 ( .B1(n19385), .B2(n15563), .A(n15562), .ZN(P2_U2998) );
  OAI21_X1 U18793 ( .B1(n14425), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15564), .ZN(n15772) );
  INV_X1 U18794 ( .A(n15566), .ZN(n15569) );
  AND2_X1 U18795 ( .A1(n15566), .A2(n15565), .ZN(n15567) );
  OAI22_X1 U18796 ( .A1(n15570), .A2(n15569), .B1(n15568), .B2(n15567), .ZN(
        n15769) );
  AOI22_X1 U18797 ( .A1(n19382), .A2(n19078), .B1(n19376), .B2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15573) );
  INV_X1 U18798 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20017) );
  OAI22_X1 U18799 ( .A1(n20017), .A2(n13196), .B1(n19374), .B2(n19075), .ZN(
        n15571) );
  INV_X1 U18800 ( .A(n15571), .ZN(n15572) );
  OAI211_X1 U18801 ( .C1(n15769), .C2(n9780), .A(n15573), .B(n15572), .ZN(
        n15574) );
  INV_X1 U18802 ( .A(n15574), .ZN(n15575) );
  OAI21_X1 U18803 ( .B1(n15772), .B2(n19385), .A(n15575), .ZN(P2_U3000) );
  NOR2_X1 U18804 ( .A1(n15577), .A2(n9992), .ZN(n15578) );
  XNOR2_X1 U18805 ( .A(n15579), .B(n15578), .ZN(n15783) );
  NAND2_X1 U18806 ( .A1(n16353), .A2(n20867), .ZN(n15773) );
  NAND3_X1 U18807 ( .A1(n15580), .A2(n16378), .A3(n15773), .ZN(n15585) );
  NOR2_X1 U18808 ( .A1(n14529), .A2(n15776), .ZN(n15583) );
  INV_X1 U18809 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20014) );
  OAI22_X1 U18810 ( .A1(n20014), .A2(n13196), .B1(n19374), .B2(n19092), .ZN(
        n15582) );
  AOI211_X1 U18811 ( .C1(n19376), .C2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15583), .B(n15582), .ZN(n15584) );
  OAI211_X1 U18812 ( .C1(n15783), .C2(n9780), .A(n15585), .B(n15584), .ZN(
        P2_U3002) );
  INV_X1 U18813 ( .A(n15587), .ZN(n15588) );
  AOI21_X1 U18814 ( .B1(n16423), .B2(n15586), .A(n15588), .ZN(n16426) );
  INV_X1 U18815 ( .A(n15589), .ZN(n15789) );
  OR2_X1 U18816 ( .A1(n15590), .A2(n15789), .ZN(n15594) );
  AND2_X1 U18817 ( .A1(n15592), .A2(n15591), .ZN(n15593) );
  XNOR2_X1 U18818 ( .A(n15594), .B(n15593), .ZN(n16429) );
  AOI22_X1 U18819 ( .A1(n19382), .A2(n9846), .B1(n19376), .B2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15597) );
  INV_X1 U18820 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20011) );
  OAI22_X1 U18821 ( .A1(n20011), .A2(n13196), .B1(n19374), .B2(n19116), .ZN(
        n15595) );
  INV_X1 U18822 ( .A(n15595), .ZN(n15596) );
  OAI211_X1 U18823 ( .C1(n16429), .C2(n9780), .A(n15597), .B(n15596), .ZN(
        n15598) );
  AOI21_X1 U18824 ( .B1(n16426), .B2(n16378), .A(n15598), .ZN(n15599) );
  INV_X1 U18825 ( .A(n15599), .ZN(P2_U3004) );
  OAI21_X1 U18826 ( .B1(n15602), .B2(n15601), .A(n15600), .ZN(n15603) );
  INV_X1 U18827 ( .A(n15603), .ZN(n16438) );
  NAND2_X1 U18828 ( .A1(n15604), .A2(n15804), .ZN(n15605) );
  NAND2_X1 U18829 ( .A1(n15605), .A2(n15805), .ZN(n15609) );
  AND2_X1 U18830 ( .A1(n15607), .A2(n15606), .ZN(n15608) );
  XNOR2_X1 U18831 ( .A(n15609), .B(n15608), .ZN(n16441) );
  AOI22_X1 U18832 ( .A1(n19382), .A2(n19139), .B1(n19185), .B2(
        P2_REIP_REG_8__SCAN_IN), .ZN(n15612) );
  INV_X1 U18833 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n21066) );
  OAI22_X1 U18834 ( .A1(n21066), .A2(n16382), .B1(n19374), .B2(n19136), .ZN(
        n15610) );
  INV_X1 U18835 ( .A(n15610), .ZN(n15611) );
  OAI211_X1 U18836 ( .C1(n16441), .C2(n9780), .A(n15612), .B(n15611), .ZN(
        n15613) );
  AOI21_X1 U18837 ( .B1(n16438), .B2(n16378), .A(n15613), .ZN(n15614) );
  INV_X1 U18838 ( .A(n15614), .ZN(P2_U3006) );
  OAI21_X1 U18839 ( .B1(n15616), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15615), .ZN(n15834) );
  XOR2_X1 U18840 ( .A(n15618), .B(n15617), .Z(n15832) );
  INV_X1 U18841 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20003) );
  OAI22_X1 U18842 ( .A1(n20003), .A2(n13196), .B1(n19374), .B2(n19160), .ZN(
        n15621) );
  INV_X1 U18843 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n15619) );
  OAI22_X1 U18844 ( .A1(n14529), .A2(n19165), .B1(n16382), .B2(n15619), .ZN(
        n15620) );
  AOI211_X1 U18845 ( .C1(n15832), .C2(n16379), .A(n15621), .B(n15620), .ZN(
        n15622) );
  OAI21_X1 U18846 ( .B1(n19385), .B2(n15834), .A(n15622), .ZN(P2_U3008) );
  NOR2_X1 U18847 ( .A1(n15637), .A2(n15623), .ZN(n15625) );
  OAI21_X1 U18848 ( .B1(n15625), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n15624), .ZN(n15629) );
  AOI21_X1 U18849 ( .B1(n15627), .B2(n19391), .A(n15626), .ZN(n15628) );
  OAI211_X1 U18850 ( .C1(n15630), .C2(n16411), .A(n15629), .B(n15628), .ZN(
        n15631) );
  AOI21_X1 U18851 ( .B1(n15632), .B2(n16450), .A(n15631), .ZN(n15633) );
  OAI21_X1 U18852 ( .B1(n15634), .B2(n19395), .A(n15633), .ZN(P2_U3016) );
  NAND2_X1 U18853 ( .A1(n16255), .A2(n19391), .ZN(n15635) );
  OAI211_X1 U18854 ( .C1(n10229), .C2(n16411), .A(n15636), .B(n15635), .ZN(
        n15642) );
  AOI211_X1 U18855 ( .C1(n15640), .C2(n15639), .A(n15638), .B(n15637), .ZN(
        n15641) );
  NAND2_X1 U18856 ( .A1(n15644), .A2(n16450), .ZN(n15645) );
  OAI211_X1 U18857 ( .C1(n15647), .C2(n19395), .A(n15646), .B(n15645), .ZN(
        P2_U3017) );
  NAND3_X1 U18858 ( .A1(n15649), .A2(n16451), .A3(n15648), .ZN(n15658) );
  NOR2_X1 U18859 ( .A1(n15650), .A2(n15655), .ZN(n15654) );
  NAND2_X1 U18860 ( .A1(n16269), .A2(n19391), .ZN(n15651) );
  OAI211_X1 U18861 ( .C1(n16266), .C2(n16411), .A(n15652), .B(n15651), .ZN(
        n15653) );
  AOI211_X1 U18862 ( .C1(n15656), .C2(n15655), .A(n15654), .B(n15653), .ZN(
        n15657) );
  OAI211_X1 U18863 ( .C1(n15659), .C2(n19406), .A(n15658), .B(n15657), .ZN(
        P2_U3019) );
  XNOR2_X1 U18864 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15666) );
  INV_X1 U18865 ( .A(n15660), .ZN(n16280) );
  OAI21_X1 U18866 ( .B1(n16277), .B2(n16433), .A(n15661), .ZN(n15664) );
  NOR2_X1 U18867 ( .A1(n15673), .A2(n15662), .ZN(n15663) );
  AOI211_X1 U18868 ( .C1(n16280), .C2(n19402), .A(n15664), .B(n15663), .ZN(
        n15665) );
  OAI21_X1 U18869 ( .B1(n15677), .B2(n15666), .A(n15665), .ZN(n15667) );
  AOI21_X1 U18870 ( .B1(n15668), .B2(n16450), .A(n15667), .ZN(n15669) );
  OAI21_X1 U18871 ( .B1(n15670), .B2(n19395), .A(n15669), .ZN(P2_U3020) );
  INV_X1 U18872 ( .A(n15671), .ZN(n16290) );
  OAI21_X1 U18873 ( .B1(n16292), .B2(n16433), .A(n15672), .ZN(n15675) );
  NOR2_X1 U18874 ( .A1(n15673), .A2(n20936), .ZN(n15674) );
  AOI211_X1 U18875 ( .C1(n16290), .C2(n19402), .A(n15675), .B(n15674), .ZN(
        n15676) );
  OAI21_X1 U18876 ( .B1(n15677), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15676), .ZN(n15678) );
  AOI21_X1 U18877 ( .B1(n15679), .B2(n16450), .A(n15678), .ZN(n15680) );
  OAI21_X1 U18878 ( .B1(n15681), .B2(n19395), .A(n15680), .ZN(P2_U3021) );
  INV_X1 U18879 ( .A(n15682), .ZN(n15683) );
  NOR2_X1 U18880 ( .A1(n15684), .A2(n15683), .ZN(n15685) );
  XNOR2_X1 U18881 ( .A(n15686), .B(n15685), .ZN(n16322) );
  AOI21_X1 U18882 ( .B1(n15692), .B2(n15688), .A(n15687), .ZN(n15689) );
  AOI21_X1 U18883 ( .B1(n19185), .B2(P2_REIP_REG_24__SCAN_IN), .A(n15689), 
        .ZN(n15690) );
  OAI21_X1 U18884 ( .B1(n16433), .B2(n16304), .A(n15690), .ZN(n15691) );
  AOI21_X1 U18885 ( .B1(n16324), .B2(n19402), .A(n15691), .ZN(n15697) );
  NAND2_X1 U18886 ( .A1(n15693), .A2(n15692), .ZN(n15694) );
  NAND2_X1 U18887 ( .A1(n15695), .A2(n15694), .ZN(n16321) );
  OR2_X1 U18888 ( .A1(n16321), .A2(n19406), .ZN(n15696) );
  OAI211_X1 U18889 ( .C1(n16322), .C2(n19395), .A(n15697), .B(n15696), .ZN(
        P2_U3022) );
  XNOR2_X1 U18890 ( .A(n15717), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15709) );
  NOR2_X1 U18891 ( .A1(n9781), .A2(n15698), .ZN(n15699) );
  OR2_X1 U18892 ( .A1(n9782), .A2(n15699), .ZN(n16305) );
  OAI21_X1 U18893 ( .B1(n16433), .B2(n16305), .A(n15700), .ZN(n15701) );
  AOI21_X1 U18894 ( .B1(n15702), .B2(n19402), .A(n15701), .ZN(n15703) );
  OAI21_X1 U18895 ( .B1(n15731), .B2(n15704), .A(n15703), .ZN(n15708) );
  NOR3_X1 U18896 ( .A1(n15706), .A2(n15705), .A3(n19395), .ZN(n15707) );
  AOI211_X1 U18897 ( .C1(n15718), .C2(n15709), .A(n15708), .B(n15707), .ZN(
        n15710) );
  OAI21_X1 U18898 ( .B1(n15711), .B2(n19406), .A(n15710), .ZN(P2_U3023) );
  NAND2_X1 U18899 ( .A1(n15712), .A2(n16450), .ZN(n15720) );
  NOR2_X1 U18900 ( .A1(n16433), .A2(n15959), .ZN(n15713) );
  AOI211_X1 U18901 ( .C1(n15962), .C2(n19402), .A(n15714), .B(n15713), .ZN(
        n15715) );
  OAI21_X1 U18902 ( .B1(n15731), .B2(n15717), .A(n15715), .ZN(n15716) );
  AOI21_X1 U18903 ( .B1(n15718), .B2(n15717), .A(n15716), .ZN(n15719) );
  OAI211_X1 U18904 ( .C1(n15721), .C2(n19395), .A(n15720), .B(n15719), .ZN(
        P2_U3024) );
  INV_X1 U18905 ( .A(n15722), .ZN(n15733) );
  NAND3_X1 U18906 ( .A1(n15724), .A2(n15723), .A3(n15730), .ZN(n15729) );
  OAI21_X1 U18907 ( .B1(n16433), .B2(n9821), .A(n15725), .ZN(n15726) );
  AOI21_X1 U18908 ( .B1(n15727), .B2(n19402), .A(n15726), .ZN(n15728) );
  OAI211_X1 U18909 ( .C1(n15731), .C2(n15730), .A(n15729), .B(n15728), .ZN(
        n15732) );
  AOI21_X1 U18910 ( .B1(n15733), .B2(n16450), .A(n15732), .ZN(n15734) );
  OAI21_X1 U18911 ( .B1(n15735), .B2(n19395), .A(n15734), .ZN(P2_U3025) );
  NAND2_X1 U18912 ( .A1(n15752), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15741) );
  XNOR2_X1 U18913 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15737) );
  NOR2_X1 U18914 ( .A1(n15737), .A2(n15736), .ZN(n15738) );
  AOI211_X1 U18915 ( .C1(n19008), .C2(n19402), .A(n15739), .B(n15738), .ZN(
        n15740) );
  OAI211_X1 U18916 ( .C1(n16433), .C2(n19005), .A(n15741), .B(n15740), .ZN(
        n15742) );
  AOI21_X1 U18917 ( .B1(n15743), .B2(n16450), .A(n15742), .ZN(n15744) );
  OAI21_X1 U18918 ( .B1(n15745), .B2(n19395), .A(n15744), .ZN(P2_U3026) );
  NAND2_X1 U18919 ( .A1(n19402), .A2(n19031), .ZN(n15747) );
  OAI211_X1 U18920 ( .C1(n16433), .C2(n19033), .A(n15747), .B(n15746), .ZN(
        n15751) );
  NOR4_X1 U18921 ( .A1(n16386), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15749), .A4(n15748), .ZN(n15750) );
  AOI211_X1 U18922 ( .C1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n15752), .A(
        n15751), .B(n15750), .ZN(n15755) );
  NAND2_X1 U18923 ( .A1(n15753), .A2(n16450), .ZN(n15754) );
  OAI211_X1 U18924 ( .C1(n15756), .C2(n19395), .A(n15755), .B(n15754), .ZN(
        P2_U3028) );
  NOR2_X1 U18925 ( .A1(n15786), .A2(n15800), .ZN(n16424) );
  NAND2_X1 U18926 ( .A1(n16415), .A2(n16424), .ZN(n16395) );
  NAND2_X1 U18927 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16415), .ZN(
        n15757) );
  AOI21_X1 U18928 ( .B1(n15757), .B2(n15815), .A(n15798), .ZN(n15778) );
  OAI21_X1 U18929 ( .B1(n16395), .B2(n15758), .A(n15778), .ZN(n16399) );
  NAND3_X1 U18930 ( .A1(n15760), .A2(n16415), .A3(n15759), .ZN(n15767) );
  OR2_X1 U18931 ( .A1(n15762), .A2(n15761), .ZN(n15763) );
  NAND2_X1 U18932 ( .A1(n15763), .A2(n16384), .ZN(n19223) );
  OAI22_X1 U18933 ( .A1(n16433), .A2(n19223), .B1(n20017), .B2(n13196), .ZN(
        n15764) );
  INV_X1 U18934 ( .A(n15764), .ZN(n15766) );
  NAND2_X1 U18935 ( .A1(n19402), .A2(n19078), .ZN(n15765) );
  OAI211_X1 U18936 ( .C1(n15800), .C2(n15767), .A(n15766), .B(n15765), .ZN(
        n15768) );
  AOI21_X1 U18937 ( .B1(n16399), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15768), .ZN(n15771) );
  OR2_X1 U18938 ( .A1(n15769), .A2(n19395), .ZN(n15770) );
  OAI211_X1 U18939 ( .C1(n15772), .C2(n19406), .A(n15771), .B(n15770), .ZN(
        P2_U3032) );
  NAND3_X1 U18940 ( .A1(n15580), .A2(n16450), .A3(n15773), .ZN(n15782) );
  XOR2_X1 U18941 ( .A(n15774), .B(n15775), .Z(n19226) );
  NOR2_X1 U18942 ( .A1(n16411), .A2(n15776), .ZN(n15780) );
  NAND2_X1 U18943 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19365), .ZN(n15777) );
  OAI221_X1 U18944 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16395), 
        .C1(n20867), .C2(n15778), .A(n15777), .ZN(n15779) );
  AOI211_X1 U18945 ( .C1(n19391), .C2(n19226), .A(n15780), .B(n15779), .ZN(
        n15781) );
  OAI211_X1 U18946 ( .C1(n15783), .C2(n19395), .A(n15782), .B(n15781), .ZN(
        P2_U3034) );
  INV_X1 U18947 ( .A(n15784), .ZN(n15787) );
  INV_X1 U18948 ( .A(n15586), .ZN(n15785) );
  AOI21_X1 U18949 ( .B1(n15787), .B2(n15786), .A(n15785), .ZN(n16361) );
  INV_X1 U18950 ( .A(n16361), .ZN(n15803) );
  NOR2_X1 U18951 ( .A1(n15789), .A2(n15788), .ZN(n15790) );
  XNOR2_X1 U18952 ( .A(n15791), .B(n15790), .ZN(n16360) );
  NAND2_X1 U18953 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19365), .ZN(n15796) );
  AOI21_X1 U18954 ( .B1(n15794), .B2(n15792), .A(n15793), .ZN(n19234) );
  NAND2_X1 U18955 ( .A1(n19391), .A2(n19234), .ZN(n15795) );
  OAI211_X1 U18956 ( .C1(n16411), .C2(n19131), .A(n15796), .B(n15795), .ZN(
        n15797) );
  AOI21_X1 U18957 ( .B1(n15798), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15797), .ZN(n15799) );
  OAI21_X1 U18958 ( .B1(n15800), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15799), .ZN(n15801) );
  AOI21_X1 U18959 ( .B1(n16360), .B2(n16451), .A(n15801), .ZN(n15802) );
  OAI21_X1 U18960 ( .B1(n15803), .B2(n19406), .A(n15802), .ZN(P2_U3037) );
  NAND2_X1 U18961 ( .A1(n15805), .A2(n15804), .ZN(n15806) );
  XOR2_X1 U18962 ( .A(n15806), .B(n15604), .Z(n16365) );
  NOR2_X1 U18963 ( .A1(n15808), .A2(n15807), .ZN(n16364) );
  INV_X1 U18964 ( .A(n16364), .ZN(n15810) );
  NAND3_X1 U18965 ( .A1(n15810), .A2(n16450), .A3(n15809), .ZN(n15821) );
  AOI21_X1 U18966 ( .B1(n15813), .B2(n15812), .A(n15811), .ZN(n19241) );
  NOR2_X1 U18967 ( .A1(n16411), .A2(n19153), .ZN(n15819) );
  INV_X1 U18968 ( .A(n15814), .ZN(n15816) );
  AOI21_X1 U18969 ( .B1(n15816), .B2(n15815), .A(n16447), .ZN(n16435) );
  NAND2_X1 U18970 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19365), .ZN(n15817) );
  OAI221_X1 U18971 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16430), .C1(
        n20950), .C2(n16435), .A(n15817), .ZN(n15818) );
  AOI211_X1 U18972 ( .C1(n19391), .C2(n19241), .A(n15819), .B(n15818), .ZN(
        n15820) );
  OAI211_X1 U18973 ( .C1(n16365), .C2(n19395), .A(n15821), .B(n15820), .ZN(
        P2_U3039) );
  INV_X1 U18974 ( .A(n16454), .ZN(n15822) );
  NOR2_X1 U18975 ( .A1(n16453), .A2(n15822), .ZN(n15824) );
  INV_X1 U18976 ( .A(n16435), .ZN(n15823) );
  MUX2_X1 U18977 ( .A(n15824), .B(n15823), .S(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(n15831) );
  NOR2_X1 U18978 ( .A1(n15826), .A2(n15825), .ZN(n15827) );
  AOI22_X1 U18979 ( .A1(n19391), .A2(n9848), .B1(n19185), .B2(
        P2_REIP_REG_6__SCAN_IN), .ZN(n15829) );
  OAI21_X1 U18980 ( .B1(n16411), .B2(n19165), .A(n15829), .ZN(n15830) );
  AOI211_X1 U18981 ( .C1(n15832), .C2(n16451), .A(n15831), .B(n15830), .ZN(
        n15833) );
  OAI21_X1 U18982 ( .B1(n19406), .B2(n15834), .A(n15833), .ZN(P2_U3040) );
  INV_X1 U18983 ( .A(n15836), .ZN(n15848) );
  INV_X1 U18984 ( .A(n11403), .ZN(n15838) );
  NAND2_X1 U18985 ( .A1(n10381), .A2(n15838), .ZN(n15856) );
  NOR2_X1 U18986 ( .A1(n13834), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15852) );
  NAND2_X1 U18987 ( .A1(n15840), .A2(n15839), .ZN(n15841) );
  NAND2_X1 U18988 ( .A1(n15841), .A2(n15842), .ZN(n15854) );
  AND2_X1 U18989 ( .A1(n16477), .A2(n16472), .ZN(n15853) );
  OAI21_X1 U18990 ( .B1(n15852), .B2(n15854), .A(n15853), .ZN(n15844) );
  INV_X1 U18991 ( .A(n15852), .ZN(n15855) );
  NAND3_X1 U18992 ( .A1(n15854), .A2(n15842), .A3(n15855), .ZN(n15843) );
  NAND2_X1 U18993 ( .A1(n15844), .A2(n15843), .ZN(n15845) );
  OAI21_X1 U18994 ( .B1(n15837), .B2(n15856), .A(n15845), .ZN(n15846) );
  AOI21_X1 U18995 ( .B1(n15847), .B2(n15860), .A(n15846), .ZN(n16468) );
  OAI222_X1 U18996 ( .A1(n16494), .A2(n20072), .B1(n15849), .B2(n15848), .C1(
        n16468), .C2(n20061), .ZN(n15850) );
  MUX2_X1 U18997 ( .A(n15850), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15862), .Z(P2_U3599) );
  AOI21_X1 U18998 ( .B1(n10381), .B2(n11403), .A(n10636), .ZN(n15851) );
  OAI21_X1 U18999 ( .B1(n15853), .B2(n15852), .A(n15851), .ZN(n15858) );
  NAND3_X1 U19000 ( .A1(n15856), .A2(n15855), .A3(n15854), .ZN(n15857) );
  MUX2_X1 U19001 ( .A(n15858), .B(n15857), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15859) );
  AOI21_X1 U19002 ( .B1(n15861), .B2(n15860), .A(n15859), .ZN(n16489) );
  OAI22_X1 U19003 ( .A1(n15893), .A2(n16494), .B1(n16489), .B2(n20061), .ZN(
        n15863) );
  MUX2_X1 U19004 ( .A(n15863), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15862), .Z(P2_U3596) );
  NAND2_X1 U19005 ( .A1(n15893), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19581) );
  NOR2_X1 U19006 ( .A1(n19581), .A2(n15894), .ZN(n20063) );
  NOR2_X1 U19007 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15886), .ZN(
        n15870) );
  AOI21_X1 U19008 ( .B1(n20113), .B2(n13298), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n20115) );
  INV_X1 U19009 ( .A(n20115), .ZN(n15864) );
  OAI21_X1 U19010 ( .B1(n20063), .B2(n15870), .A(n19883), .ZN(n15869) );
  INV_X1 U19011 ( .A(n19517), .ZN(n19756) );
  NOR2_X1 U19012 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20076), .ZN(
        n19611) );
  NAND2_X1 U19013 ( .A1(n19756), .A2(n19611), .ZN(n19664) );
  AND2_X1 U19014 ( .A1(n19664), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n15865) );
  NAND2_X1 U19015 ( .A1(n15866), .A2(n15865), .ZN(n15872) );
  NAND2_X1 U19016 ( .A1(n19664), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15867) );
  NAND2_X1 U19017 ( .A1(n15872), .A2(n15867), .ZN(n15868) );
  INV_X1 U19018 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15884) );
  INV_X1 U19019 ( .A(n15870), .ZN(n15874) );
  INV_X1 U19020 ( .A(n15871), .ZN(n19615) );
  INV_X1 U19021 ( .A(n15872), .ZN(n15873) );
  AOI211_X2 U19022 ( .C1(n15874), .C2(n20113), .A(n19615), .B(n15873), .ZN(
        n19657) );
  NAND2_X1 U19023 ( .A1(n19281), .A2(n19883), .ZN(n19889) );
  INV_X1 U19024 ( .A(n19453), .ZN(n15877) );
  NAND2_X1 U19025 ( .A1(n15877), .A2(n15876), .ZN(n19408) );
  AOI22_X1 U19026 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19451), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19450), .ZN(n19803) );
  INV_X1 U19027 ( .A(n19803), .ZN(n19877) );
  NAND2_X1 U19028 ( .A1(n15885), .A2(n19549), .ZN(n19645) );
  INV_X1 U19029 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16583) );
  INV_X1 U19030 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18309) );
  OAI22_X2 U19031 ( .A1(n16583), .A2(n19446), .B1(n18309), .B2(n19448), .ZN(
        n19886) );
  AOI22_X1 U19032 ( .A1(n19683), .A2(n19877), .B1(n19658), .B2(n19886), .ZN(
        n15881) );
  OAI21_X1 U19033 ( .B1(n19408), .B2(n19664), .A(n15881), .ZN(n15882) );
  AOI21_X1 U19034 ( .B1(n19657), .B2(n19833), .A(n15882), .ZN(n15883) );
  OAI21_X1 U19035 ( .B1(n19656), .B2(n15884), .A(n15883), .ZN(P2_U3104) );
  NOR2_X1 U19036 ( .A1(n15893), .A2(n20107), .ZN(n19835) );
  NAND2_X1 U19037 ( .A1(n19835), .A2(n15885), .ZN(n15890) );
  OR2_X1 U19038 ( .A1(n20069), .A2(n15886), .ZN(n19873) );
  INV_X1 U19039 ( .A(n19412), .ZN(n19954) );
  AND2_X1 U19040 ( .A1(n19412), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n15887) );
  NAND2_X1 U19041 ( .A1(n15888), .A2(n15887), .ZN(n15892) );
  OAI211_X1 U19042 ( .C1(n19954), .C2(n19879), .A(n15892), .B(n19883), .ZN(
        n15889) );
  INV_X1 U19043 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15898) );
  OAI21_X1 U19044 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19873), .A(n20113), 
        .ZN(n15891) );
  AND2_X1 U19045 ( .A1(n15892), .A2(n15891), .ZN(n19956) );
  AOI22_X1 U19046 ( .A1(n19958), .A2(n19886), .B1(n19960), .B2(n19877), .ZN(
        n15895) );
  OAI21_X1 U19047 ( .B1(n19408), .B2(n19412), .A(n15895), .ZN(n15896) );
  AOI21_X1 U19048 ( .B1(n19833), .B2(n19956), .A(n15896), .ZN(n15897) );
  OAI21_X1 U19049 ( .B1(n19964), .B2(n15898), .A(n15897), .ZN(P2_U3168) );
  NAND2_X1 U19050 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17259), .ZN(n17260) );
  NOR2_X1 U19051 ( .A1(n16914), .A2(n17260), .ZN(n17244) );
  INV_X1 U19052 ( .A(n17260), .ZN(n15899) );
  AOI22_X1 U19053 ( .A1(n18348), .A2(n15899), .B1(P3_EBX_REG_13__SCAN_IN), 
        .B2(n17338), .ZN(n15912) );
  AOI22_X1 U19054 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15905) );
  AOI22_X1 U19055 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15904) );
  AOI22_X1 U19056 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15903) );
  AOI22_X1 U19057 ( .A1(n15901), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13466), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15902) );
  NAND4_X1 U19058 ( .A1(n15905), .A2(n15904), .A3(n15903), .A4(n15902), .ZN(
        n15911) );
  AOI22_X1 U19059 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17277), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15909) );
  AOI22_X1 U19060 ( .A1(n12749), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9754), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15908) );
  AOI22_X1 U19061 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15907) );
  AOI22_X1 U19062 ( .A1(n17303), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12838), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15906) );
  NAND4_X1 U19063 ( .A1(n15909), .A2(n15908), .A3(n15907), .A4(n15906), .ZN(
        n15910) );
  NOR2_X1 U19064 ( .A1(n15911), .A2(n15910), .ZN(n17441) );
  OAI22_X1 U19065 ( .A1(n17244), .A2(n15912), .B1(n17441), .B2(n17338), .ZN(
        P3_U2690) );
  NOR2_X1 U19066 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18935), .ZN(
        n18295) );
  INV_X1 U19067 ( .A(n18295), .ZN(n18355) );
  INV_X1 U19068 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18294) );
  NAND3_X1 U19069 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(P3_STATE2_REG_0__SCAN_IN), .ZN(n18913)
         );
  INV_X1 U19070 ( .A(n18758), .ZN(n18765) );
  AOI211_X1 U19071 ( .C1(n18765), .C2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n17302), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18292) );
  OAI221_X1 U19072 ( .B1(n18294), .B2(n18913), .C1(n18292), .C2(n18913), .A(
        n18612), .ZN(n18304) );
  NAND2_X1 U19073 ( .A1(n18355), .A2(n18304), .ZN(n18298) );
  INV_X1 U19074 ( .A(n18298), .ZN(n15914) );
  INV_X1 U19075 ( .A(n18663), .ZN(n18611) );
  INV_X1 U19076 ( .A(n17922), .ZN(n18297) );
  INV_X1 U19077 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18607) );
  OAI22_X1 U19078 ( .A1(n18956), .A2(n18297), .B1(n18607), .B2(n18935), .ZN(
        n18300) );
  NAND3_X1 U19079 ( .A1(n18793), .A2(n18304), .A3(n18300), .ZN(n15913) );
  OAI221_X1 U19080 ( .B1(n18793), .B2(n15914), .C1(n18793), .C2(n18611), .A(
        n15913), .ZN(P3_U2864) );
  NOR2_X1 U19081 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18935), .ZN(n18307) );
  INV_X1 U19082 ( .A(n15915), .ZN(n15918) );
  AOI221_X1 U19083 ( .B1(n15919), .B2(n15918), .C1(n15917), .C2(n15918), .A(
        n15916), .ZN(n15937) );
  NAND2_X1 U19084 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n20932), .ZN(n18969) );
  NAND2_X1 U19085 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n18950), .ZN(n18900) );
  NOR2_X1 U19086 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n18828) );
  INV_X1 U19087 ( .A(n18828), .ZN(n15920) );
  NAND3_X1 U19088 ( .A1(n20932), .A2(n18893), .A3(n15920), .ZN(n18834) );
  NOR2_X1 U19089 ( .A1(n16682), .A2(n18834), .ZN(n17499) );
  NAND2_X1 U19090 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18953) );
  OAI211_X1 U19091 ( .C1(n17499), .C2(n16683), .A(n18748), .B(n18953), .ZN(
        n15922) );
  OAI211_X1 U19092 ( .C1(n15924), .C2(n15923), .A(n15937), .B(n15922), .ZN(
        n18786) );
  INV_X1 U19093 ( .A(n18786), .ZN(n18796) );
  OAI22_X1 U19094 ( .A1(n18796), .A2(n18817), .B1(n18294), .B2(n18913), .ZN(
        n15925) );
  NOR2_X1 U19095 ( .A1(n18307), .A2(n15925), .ZN(n21190) );
  INV_X1 U19096 ( .A(n21190), .ZN(n21187) );
  AOI21_X1 U19097 ( .B1(n18765), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15926) );
  NOR2_X1 U19098 ( .A1(n15926), .A2(n18772), .ZN(n18807) );
  NAND3_X1 U19099 ( .A1(n21187), .A2(n21185), .A3(n18807), .ZN(n15927) );
  OAI21_X1 U19100 ( .B1(n21187), .B2(n18754), .A(n15927), .ZN(P3_U3284) );
  OAI21_X1 U19101 ( .B1(n15929), .B2(n15928), .A(n18328), .ZN(n15935) );
  AND4_X1 U19102 ( .A1(n18959), .A2(n17349), .A3(n18318), .A4(n18749), .ZN(
        n15934) );
  INV_X1 U19103 ( .A(n18834), .ZN(n18958) );
  AOI22_X1 U19104 ( .A1(n18313), .A2(n18318), .B1(n15929), .B2(n18959), .ZN(
        n15930) );
  OAI21_X1 U19105 ( .B1(n18958), .B2(n15930), .A(n18953), .ZN(n16667) );
  NOR3_X1 U19106 ( .A1(n15932), .A2(n15931), .A3(n16667), .ZN(n15933) );
  AOI211_X1 U19107 ( .C1(n18745), .C2(n15935), .A(n15934), .B(n15933), .ZN(
        n15936) );
  AOI21_X2 U19108 ( .B1(n15937), .B2(n15936), .A(n18817), .ZN(n18271) );
  NOR2_X1 U19109 ( .A1(n18125), .A2(n18286), .ZN(n18237) );
  INV_X1 U19110 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21067) );
  NAND2_X1 U19111 ( .A1(n18789), .A2(n18757), .ZN(n18167) );
  NOR3_X1 U19112 ( .A1(n18243), .A2(n18246), .A3(n18231), .ZN(n18077) );
  NAND3_X1 U19113 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n18077), .ZN(n18192) );
  NAND3_X1 U19114 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18076) );
  NOR2_X1 U19115 ( .A1(n18192), .A2(n18076), .ZN(n18122) );
  NAND2_X1 U19116 ( .A1(n16508), .A2(n18122), .ZN(n18031) );
  INV_X1 U19117 ( .A(n18031), .ZN(n18069) );
  NAND2_X1 U19118 ( .A1(n16509), .A2(n18069), .ZN(n15945) );
  INV_X1 U19119 ( .A(n15945), .ZN(n15940) );
  NAND2_X1 U19120 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15940), .ZN(
        n15938) );
  INV_X1 U19121 ( .A(n17682), .ZN(n17970) );
  INV_X1 U19122 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18924) );
  OAI21_X1 U19123 ( .B1(n18924), .B2(n18925), .A(n18261), .ZN(n18233) );
  NAND2_X1 U19124 ( .A1(n18077), .A2(n18233), .ZN(n18193) );
  NOR2_X1 U19125 ( .A1(n18076), .A2(n18193), .ZN(n18091) );
  NAND2_X1 U19126 ( .A1(n16508), .A2(n18091), .ZN(n18070) );
  NOR2_X1 U19127 ( .A1(n17970), .A2(n18070), .ZN(n17992) );
  AOI21_X1 U19128 ( .B1(n17973), .B2(n17992), .A(n18757), .ZN(n17969) );
  AOI221_X1 U19129 ( .B1(n21067), .B2(n18787), .C1(n15938), .C2(n18787), .A(
        n17969), .ZN(n15939) );
  OAI211_X1 U19130 ( .C1(n18789), .C2(n15940), .A(n18271), .B(n15939), .ZN(
        n16010) );
  AOI21_X1 U19131 ( .B1(n21067), .B2(n18167), .A(n16010), .ZN(n16555) );
  NAND2_X1 U19132 ( .A1(n18744), .A2(n18271), .ZN(n18216) );
  NAND2_X1 U19133 ( .A1(n16539), .A2(n17967), .ZN(n16514) );
  NAND2_X1 U19134 ( .A1(n16553), .A2(n18271), .ZN(n18279) );
  NOR2_X1 U19135 ( .A1(n16552), .A2(n18279), .ZN(n18135) );
  INV_X1 U19136 ( .A(n16515), .ZN(n16523) );
  AOI22_X1 U19137 ( .A1(n18282), .A2(n16514), .B1(n18135), .B2(n16523), .ZN(
        n16013) );
  OAI21_X1 U19138 ( .B1(n18285), .B2(n16555), .A(n16013), .ZN(n15941) );
  AOI21_X1 U19139 ( .B1(n18237), .B2(n17606), .A(n15941), .ZN(n15950) );
  NAND2_X1 U19140 ( .A1(n17872), .A2(n17606), .ZN(n16559) );
  INV_X1 U19141 ( .A(n16559), .ZN(n15942) );
  AOI21_X1 U19142 ( .B1(n16551), .B2(n15943), .A(n15942), .ZN(n15944) );
  XNOR2_X1 U19143 ( .A(n15944), .B(n16536), .ZN(n16534) );
  INV_X1 U19144 ( .A(n18135), .ZN(n18206) );
  AOI221_X1 U19145 ( .B1(n18755), .B2(n18789), .C1(n18925), .C2(n18789), .A(
        n15945), .ZN(n15946) );
  NOR2_X1 U19146 ( .A1(n18757), .A2(n18070), .ZN(n16561) );
  OAI211_X1 U19147 ( .C1(n15946), .C2(n16561), .A(n16509), .B(n18271), .ZN(
        n16540) );
  OAI21_X1 U19148 ( .B1(n18206), .B2(n17605), .A(n16540), .ZN(n15947) );
  AOI21_X1 U19149 ( .B1(n17967), .B2(n18282), .A(n15947), .ZN(n16016) );
  NOR3_X1 U19150 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16016), .A3(
        n16522), .ZN(n15948) );
  AOI21_X1 U19151 ( .B1(n16534), .B2(n9863), .A(n15948), .ZN(n15949) );
  NAND2_X1 U19152 ( .A1(n18285), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16532) );
  OAI211_X1 U19153 ( .C1(n15950), .C2(n16536), .A(n15949), .B(n16532), .ZN(
        P3_U2833) );
  AOI211_X1 U19154 ( .C1(n15953), .C2(n15951), .A(n15952), .B(n19972), .ZN(
        n15961) );
  AOI22_X1 U19155 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19166), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19204), .ZN(n15958) );
  OAI22_X1 U19156 ( .A1(n15955), .A2(n19169), .B1(n19207), .B2(n15954), .ZN(
        n15956) );
  INV_X1 U19157 ( .A(n15956), .ZN(n15957) );
  OAI211_X1 U19158 ( .C1(n15959), .C2(n19182), .A(n15958), .B(n15957), .ZN(
        n15960) );
  AOI211_X1 U19159 ( .C1(n19187), .C2(n15962), .A(n15961), .B(n15960), .ZN(
        n15963) );
  INV_X1 U19160 ( .A(n15963), .ZN(P2_U2833) );
  INV_X1 U19161 ( .A(n15979), .ZN(n15983) );
  INV_X1 U19162 ( .A(n15964), .ZN(n15965) );
  OAI211_X1 U19163 ( .C1(n11802), .C2(n15966), .A(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n15965), .ZN(n15969) );
  INV_X1 U19164 ( .A(n15967), .ZN(n15968) );
  OAI21_X1 U19165 ( .B1(n20517), .B2(n15969), .A(n15968), .ZN(n15971) );
  NAND2_X1 U19166 ( .A1(n20517), .A2(n15969), .ZN(n15970) );
  OAI21_X1 U19167 ( .B1(n15972), .B2(n15971), .A(n15970), .ZN(n15975) );
  AND2_X1 U19168 ( .A1(n12111), .A2(n15975), .ZN(n15973) );
  OR2_X1 U19169 ( .A1(n15974), .A2(n15973), .ZN(n15978) );
  INV_X1 U19170 ( .A(n15975), .ZN(n15976) );
  NAND2_X1 U19171 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n15976), .ZN(
        n15977) );
  NAND2_X1 U19172 ( .A1(n15978), .A2(n15977), .ZN(n15982) );
  INV_X1 U19173 ( .A(n15982), .ZN(n15980) );
  OAI21_X1 U19174 ( .B1(n15980), .B2(n15979), .A(n20825), .ZN(n15981) );
  OAI21_X1 U19175 ( .B1(n15983), .B2(n15982), .A(n15981), .ZN(n15990) );
  NOR2_X1 U19176 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n15986) );
  OAI211_X1 U19177 ( .C1(n15987), .C2(n15986), .A(n15985), .B(n15984), .ZN(
        n15988) );
  AOI211_X1 U19178 ( .C1(n15990), .C2(n20326), .A(n15989), .B(n15988), .ZN(
        n15991) );
  NAND2_X1 U19179 ( .A1(n15992), .A2(n15991), .ZN(n16000) );
  INV_X1 U19180 ( .A(n15993), .ZN(n15997) );
  OAI21_X1 U19181 ( .B1(n20846), .B2(n15995), .A(n15994), .ZN(n15996) );
  OAI21_X1 U19182 ( .B1(n15998), .B2(n15997), .A(n15996), .ZN(n16232) );
  AOI221_X1 U19183 ( .B1(n9918), .B2(n20727), .C1(n16000), .C2(n20727), .A(
        n16232), .ZN(n16236) );
  AOI21_X1 U19184 ( .B1(n16001), .B2(n16000), .A(n15999), .ZN(n16003) );
  OAI211_X1 U19185 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20846), .A(n16003), 
        .B(n16002), .ZN(n16004) );
  NOR2_X1 U19186 ( .A1(n16236), .A2(n16004), .ZN(n16007) );
  NAND2_X1 U19187 ( .A1(n16229), .A2(n20803), .ZN(n16005) );
  NAND2_X1 U19188 ( .A1(n9918), .A2(n16005), .ZN(n16006) );
  OAI22_X1 U19189 ( .A1(n16007), .A2(n9918), .B1(n16236), .B2(n16006), .ZN(
        P1_U3161) );
  NAND2_X1 U19190 ( .A1(n16539), .A2(n16012), .ZN(n16520) );
  AOI21_X1 U19191 ( .B1(n16009), .B2(n16012), .A(n16008), .ZN(n16516) );
  AOI22_X1 U19192 ( .A1(n18237), .A2(n16011), .B1(n16866), .B2(n16010), .ZN(
        n16542) );
  AOI21_X1 U19193 ( .B1(n16542), .B2(n16013), .A(n16012), .ZN(n16014) );
  AOI21_X1 U19194 ( .B1(n9863), .B2(n16516), .A(n16014), .ZN(n16015) );
  INV_X1 U19195 ( .A(n16866), .ZN(n18245) );
  NAND2_X1 U19196 ( .A1(n18245), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16510) );
  OAI211_X1 U19197 ( .C1(n16016), .C2(n16520), .A(n16015), .B(n16510), .ZN(
        P3_U2832) );
  INV_X1 U19198 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20130) );
  INV_X1 U19199 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20739) );
  NOR2_X1 U19200 ( .A1(n20738), .A2(n20739), .ZN(n20736) );
  INV_X1 U19201 ( .A(HOLD), .ZN(n20743) );
  OAI222_X1 U19202 ( .A1(n20736), .A2(P1_STATE_REG_1__SCAN_IN), .B1(n20736), 
        .B2(HOLD), .C1(n20743), .C2(n11789), .ZN(n16018) );
  OAI211_X1 U19203 ( .C1(n20846), .C2(n20130), .A(n16018), .B(n16017), .ZN(
        P1_U3195) );
  AND2_X1 U19204 ( .A1(n20239), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NAND2_X1 U19205 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20118), .ZN(n19966) );
  AOI21_X1 U19206 ( .B1(n20078), .B2(n20119), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16019) );
  INV_X1 U19207 ( .A(n16500), .ZN(n16505) );
  AOI221_X1 U19208 ( .B1(n19966), .B2(n16019), .C1(n13298), .C2(n16019), .A(
        n16505), .ZN(P2_U3178) );
  INV_X1 U19209 ( .A(n16020), .ZN(n20102) );
  AOI221_X1 U19210 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16505), .C1(n20102), .C2(
        n16505), .A(n19883), .ZN(n20093) );
  INV_X1 U19211 ( .A(n20093), .ZN(n20090) );
  NOR2_X1 U19212 ( .A1(n16493), .A2(n20090), .ZN(P2_U3047) );
  NAND3_X1 U19213 ( .A1(n18308), .A2(n18313), .A3(n16021), .ZN(n16022) );
  NAND2_X1 U19214 ( .A1(n18348), .A2(n17498), .ZN(n17484) );
  INV_X1 U19215 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17571) );
  NAND2_X2 U19216 ( .A1(n17498), .A2(n17431), .ZN(n17486) );
  NAND2_X1 U19217 ( .A1(n16024), .A2(n17375), .ZN(n17490) );
  INV_X1 U19218 ( .A(n17490), .ZN(n17493) );
  NAND2_X1 U19219 ( .A1(n18788), .A2(n17498), .ZN(n17487) );
  OAI221_X1 U19220 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17484), .C1(n17571), 
        .C2(n17498), .A(n16025), .ZN(P3_U2735) );
  INV_X1 U19221 ( .A(n16026), .ZN(n16035) );
  OAI22_X1 U19222 ( .A1(n20194), .A2(n16027), .B1(n12467), .B2(n20210), .ZN(
        n16034) );
  NAND3_X1 U19223 ( .A1(n16028), .A2(P1_REIP_REG_21__SCAN_IN), .A3(
        P1_REIP_REG_22__SCAN_IN), .ZN(n16032) );
  INV_X1 U19224 ( .A(n16029), .ZN(n16030) );
  AOI211_X1 U19225 ( .C1(n20778), .C2(n16032), .A(n16031), .B(n16030), .ZN(
        n16033) );
  AOI211_X1 U19226 ( .C1(n20162), .C2(n16035), .A(n16034), .B(n16033), .ZN(
        n16041) );
  INV_X1 U19227 ( .A(n16036), .ZN(n16039) );
  INV_X1 U19228 ( .A(n16037), .ZN(n16038) );
  AOI22_X1 U19229 ( .A1(n16039), .A2(n20185), .B1(n20205), .B2(n16038), .ZN(
        n16040) );
  NAND2_X1 U19230 ( .A1(n16041), .A2(n16040), .ZN(P1_U2817) );
  INV_X1 U19231 ( .A(n16042), .ZN(n16044) );
  AOI22_X1 U19232 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n16054), .B1(n16044), 
        .B2(n16043), .ZN(n16046) );
  AOI22_X1 U19233 ( .A1(n20206), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20193), .ZN(n16045) );
  OAI211_X1 U19234 ( .C1(n16047), .C2(n20191), .A(n16046), .B(n16045), .ZN(
        n16048) );
  AOI21_X1 U19235 ( .B1(n16049), .B2(n20185), .A(n16048), .ZN(n16050) );
  OAI21_X1 U19236 ( .B1(n16051), .B2(n20216), .A(n16050), .ZN(P1_U2819) );
  AOI22_X1 U19237 ( .A1(n20206), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20193), .ZN(n16060) );
  AOI22_X1 U19238 ( .A1(n16053), .A2(n20185), .B1(n16052), .B2(n20205), .ZN(
        n16059) );
  INV_X1 U19239 ( .A(n20196), .ZN(n20179) );
  OAI221_X1 U19240 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(n16055), .C1(
        P1_REIP_REG_20__SCAN_IN), .C2(n20179), .A(n16054), .ZN(n16058) );
  NAND2_X1 U19241 ( .A1(n16056), .A2(n20162), .ZN(n16057) );
  NAND4_X1 U19242 ( .A1(n16060), .A2(n16059), .A3(n16058), .A4(n16057), .ZN(
        P1_U2820) );
  NOR2_X1 U19243 ( .A1(n16069), .A2(n16068), .ZN(n16061) );
  INV_X1 U19244 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20771) );
  NAND3_X1 U19245 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n16061), .A3(n20771), 
        .ZN(n16064) );
  OAI21_X1 U19246 ( .B1(n20210), .B2(n12377), .A(n20207), .ZN(n16062) );
  AOI21_X1 U19247 ( .B1(n20206), .B2(P1_EBX_REG_19__SCAN_IN), .A(n16062), .ZN(
        n16063) );
  OAI211_X1 U19248 ( .C1(n16065), .C2(n20216), .A(n16064), .B(n16063), .ZN(
        n16066) );
  AOI21_X1 U19249 ( .B1(n16067), .B2(n20185), .A(n16066), .ZN(n16071) );
  NOR3_X1 U19250 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n16069), .A3(n16068), 
        .ZN(n16078) );
  OAI21_X1 U19251 ( .B1(n16074), .B2(n16078), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n16070) );
  OAI211_X1 U19252 ( .C1(n16072), .C2(n20191), .A(n16071), .B(n16070), .ZN(
        P1_U2821) );
  INV_X1 U19253 ( .A(n16073), .ZN(n16124) );
  AOI22_X1 U19254 ( .A1(n16125), .A2(n20185), .B1(n20205), .B2(n16124), .ZN(
        n16081) );
  AOI22_X1 U19255 ( .A1(n16074), .A2(P1_REIP_REG_18__SCAN_IN), .B1(n20206), 
        .B2(P1_EBX_REG_18__SCAN_IN), .ZN(n16075) );
  OAI211_X1 U19256 ( .C1(n20210), .C2(n16076), .A(n16075), .B(n20207), .ZN(
        n16077) );
  AOI211_X1 U19257 ( .C1(n20162), .C2(n16079), .A(n16078), .B(n16077), .ZN(
        n16080) );
  NAND2_X1 U19258 ( .A1(n16081), .A2(n16080), .ZN(P1_U2822) );
  AOI22_X1 U19259 ( .A1(n16083), .A2(n20162), .B1(n20205), .B2(n16082), .ZN(
        n16092) );
  NAND2_X1 U19260 ( .A1(n20193), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16084) );
  NAND2_X1 U19261 ( .A1(n16084), .A2(n20207), .ZN(n16085) );
  AOI21_X1 U19262 ( .B1(n20206), .B2(P1_EBX_REG_15__SCAN_IN), .A(n16085), .ZN(
        n16086) );
  OAI21_X1 U19263 ( .B1(n16087), .B2(n20764), .A(n16086), .ZN(n16088) );
  OR2_X1 U19264 ( .A1(n16089), .A2(n16088), .ZN(n16090) );
  AOI21_X1 U19265 ( .B1(n16135), .B2(n20185), .A(n16090), .ZN(n16091) );
  NAND2_X1 U19266 ( .A1(n16092), .A2(n16091), .ZN(P1_U2825) );
  INV_X1 U19267 ( .A(n16093), .ZN(n16110) );
  AOI21_X1 U19268 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n16110), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n16100) );
  NAND2_X1 U19269 ( .A1(n20206), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n16094) );
  OAI211_X1 U19270 ( .C1(n16095), .C2(n20210), .A(n16094), .B(n20207), .ZN(
        n16096) );
  AOI21_X1 U19271 ( .B1(n16097), .B2(n20205), .A(n16096), .ZN(n16099) );
  AOI22_X1 U19272 ( .A1(n16140), .A2(n20162), .B1(n20185), .B2(n16139), .ZN(
        n16098) );
  OAI211_X1 U19273 ( .C1(n16101), .C2(n16100), .A(n16099), .B(n16098), .ZN(
        P1_U2828) );
  NAND2_X1 U19274 ( .A1(n20189), .A2(n16102), .ZN(n16122) );
  INV_X1 U19275 ( .A(n16122), .ZN(n16109) );
  INV_X1 U19276 ( .A(n16103), .ZN(n16104) );
  NAND2_X1 U19277 ( .A1(n16104), .A2(n20205), .ZN(n16107) );
  NAND2_X1 U19278 ( .A1(n20206), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n16106) );
  NAND2_X1 U19279 ( .A1(n20193), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16105) );
  NAND4_X1 U19280 ( .A1(n16107), .A2(n16106), .A3(n20207), .A4(n16105), .ZN(
        n16108) );
  AOI21_X1 U19281 ( .B1(n16109), .B2(P1_REIP_REG_11__SCAN_IN), .A(n16108), 
        .ZN(n16112) );
  AOI22_X1 U19282 ( .A1(n16145), .A2(n20185), .B1(n16110), .B2(n15146), .ZN(
        n16111) );
  OAI211_X1 U19283 ( .C1(n16149), .C2(n20216), .A(n16112), .B(n16111), .ZN(
        P1_U2829) );
  NAND2_X1 U19284 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n20158), .ZN(n16123) );
  OAI21_X1 U19285 ( .B1(n20210), .B2(n16113), .A(n20207), .ZN(n16115) );
  NOR2_X1 U19286 ( .A1(n20191), .A2(n16183), .ZN(n16114) );
  AOI211_X1 U19287 ( .C1(n20206), .C2(P1_EBX_REG_10__SCAN_IN), .A(n16115), .B(
        n16114), .ZN(n16116) );
  OAI21_X1 U19288 ( .B1(n16118), .B2(n16117), .A(n16116), .ZN(n16119) );
  AOI21_X1 U19289 ( .B1(n16120), .B2(n20162), .A(n16119), .ZN(n16121) );
  OAI221_X1 U19290 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n16123), .C1(n14949), 
        .C2(n16122), .A(n16121), .ZN(P1_U2830) );
  INV_X1 U19291 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n16127) );
  AOI22_X1 U19292 ( .A1(n16125), .A2(n20223), .B1(n20222), .B2(n16124), .ZN(
        n16126) );
  OAI21_X1 U19293 ( .B1(n20227), .B2(n16127), .A(n16126), .ZN(P1_U2854) );
  AOI22_X1 U19294 ( .A1(n20287), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20299), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16131) );
  AOI22_X1 U19295 ( .A1(n16129), .A2(n20293), .B1(n16141), .B2(n16128), .ZN(
        n16130) );
  OAI211_X1 U19296 ( .C1(n20139), .C2(n16132), .A(n16131), .B(n16130), .ZN(
        P1_U2982) );
  AOI22_X1 U19297 ( .A1(n20287), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20299), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16137) );
  NOR2_X1 U19298 ( .A1(n20298), .A2(n16133), .ZN(n16134) );
  AOI21_X1 U19299 ( .B1(n16135), .B2(n20293), .A(n16134), .ZN(n16136) );
  OAI211_X1 U19300 ( .C1(n16138), .C2(n20139), .A(n16137), .B(n16136), .ZN(
        P1_U2984) );
  AOI22_X1 U19301 ( .A1(n20287), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20299), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16143) );
  AOI22_X1 U19302 ( .A1(n16141), .A2(n16140), .B1(n20293), .B2(n16139), .ZN(
        n16142) );
  OAI211_X1 U19303 ( .C1(n16144), .C2(n20139), .A(n16143), .B(n16142), .ZN(
        P1_U2987) );
  AOI22_X1 U19304 ( .A1(n20287), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20299), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16148) );
  AOI22_X1 U19305 ( .A1(n20294), .A2(n16146), .B1(n20293), .B2(n16145), .ZN(
        n16147) );
  OAI211_X1 U19306 ( .C1(n20298), .C2(n16149), .A(n16148), .B(n16147), .ZN(
        P1_U2988) );
  AOI22_X1 U19307 ( .A1(n20287), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20299), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16152) );
  AOI22_X1 U19308 ( .A1(n16150), .A2(n20294), .B1(n20293), .B2(n20174), .ZN(
        n16151) );
  OAI211_X1 U19309 ( .C1(n20298), .C2(n20178), .A(n16152), .B(n16151), .ZN(
        P1_U2992) );
  AOI22_X1 U19310 ( .A1(n20287), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20299), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16157) );
  XNOR2_X1 U19311 ( .A(n16154), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16155) );
  XNOR2_X1 U19312 ( .A(n16153), .B(n16155), .ZN(n16210) );
  AOI22_X1 U19313 ( .A1(n16210), .A2(n20294), .B1(n20293), .B2(n20224), .ZN(
        n16156) );
  OAI211_X1 U19314 ( .C1(n20298), .C2(n20187), .A(n16157), .B(n16156), .ZN(
        P1_U2993) );
  AOI22_X1 U19315 ( .A1(n20287), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20299), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16164) );
  OAI21_X1 U19316 ( .B1(n16160), .B2(n16159), .A(n16158), .ZN(n16161) );
  INV_X1 U19317 ( .A(n16161), .ZN(n16216) );
  INV_X1 U19318 ( .A(n16162), .ZN(n20198) );
  AOI22_X1 U19319 ( .A1(n16216), .A2(n20294), .B1(n20293), .B2(n20198), .ZN(
        n16163) );
  OAI211_X1 U19320 ( .C1(n20298), .C2(n20201), .A(n16164), .B(n16163), .ZN(
        P1_U2994) );
  INV_X1 U19321 ( .A(n16182), .ZN(n16165) );
  AOI22_X1 U19322 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16165), .B1(
        n20299), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16170) );
  INV_X1 U19323 ( .A(n16166), .ZN(n16167) );
  AOI22_X1 U19324 ( .A1(n16168), .A2(n20318), .B1(n20312), .B2(n16167), .ZN(
        n16169) );
  OAI211_X1 U19325 ( .C1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n16171), .A(
        n16170), .B(n16169), .ZN(P1_U3017) );
  AOI21_X1 U19326 ( .B1(n16173), .B2(n20312), .A(n16172), .ZN(n16180) );
  OAI21_X1 U19327 ( .B1(n16176), .B2(n16175), .A(n16174), .ZN(n16177) );
  AOI22_X1 U19328 ( .A1(n16178), .A2(n20318), .B1(n16181), .B2(n16177), .ZN(
        n16179) );
  OAI211_X1 U19329 ( .C1(n16182), .C2(n16181), .A(n16180), .B(n16179), .ZN(
        P1_U3018) );
  INV_X1 U19330 ( .A(n16183), .ZN(n16185) );
  AOI21_X1 U19331 ( .B1(n16185), .B2(n20312), .A(n16184), .ZN(n16193) );
  AOI22_X1 U19332 ( .A1(n16187), .A2(n20318), .B1(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16186), .ZN(n16192) );
  OAI221_X1 U19333 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n16190), .C2(n16189), .A(
        n16188), .ZN(n16191) );
  NAND3_X1 U19334 ( .A1(n16193), .A2(n16192), .A3(n16191), .ZN(P1_U3021) );
  AOI21_X1 U19335 ( .B1(n20312), .B2(n16195), .A(n16194), .ZN(n16203) );
  AOI22_X1 U19336 ( .A1(n16197), .A2(n20318), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16196), .ZN(n16202) );
  INV_X1 U19337 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16200) );
  OAI221_X1 U19338 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16200), .C2(n16199), .A(
        n16198), .ZN(n16201) );
  NAND3_X1 U19339 ( .A1(n16203), .A2(n16202), .A3(n16201), .ZN(P1_U3023) );
  AND2_X1 U19340 ( .A1(n16205), .A2(n16204), .ZN(n16213) );
  AND2_X1 U19341 ( .A1(n16207), .A2(n16206), .ZN(n16208) );
  NOR2_X1 U19342 ( .A1(n16209), .A2(n16208), .ZN(n20221) );
  AOI22_X1 U19343 ( .A1(n16210), .A2(n20318), .B1(n20312), .B2(n20221), .ZN(
        n16212) );
  NAND2_X1 U19344 ( .A1(n20299), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n16211) );
  OAI211_X1 U19345 ( .C1(n16214), .C2(n16213), .A(n16212), .B(n16211), .ZN(
        P1_U3025) );
  AOI22_X1 U19346 ( .A1(n16216), .A2(n20318), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16215), .ZN(n16224) );
  INV_X1 U19347 ( .A(n16217), .ZN(n16219) );
  OAI22_X1 U19348 ( .A1(n16220), .A2(n16219), .B1(n16218), .B2(n20190), .ZN(
        n16221) );
  AOI211_X1 U19349 ( .C1(P1_REIP_REG_5__SCAN_IN), .C2(n20299), .A(n16222), .B(
        n16221), .ZN(n16223) );
  NAND2_X1 U19350 ( .A1(n16224), .A2(n16223), .ZN(P1_U3026) );
  NAND2_X1 U19351 ( .A1(n16225), .A2(n20804), .ZN(n16227) );
  OAI22_X1 U19352 ( .A1(n16228), .A2(n16227), .B1(n16226), .B2(n20807), .ZN(
        P1_U3468) );
  INV_X1 U19353 ( .A(n16229), .ZN(n20843) );
  NAND4_X1 U19354 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20839), .A4(n20846), .ZN(n16230) );
  OAI21_X1 U19355 ( .B1(n16231), .B2(n20840), .A(n16230), .ZN(n20728) );
  OAI21_X1 U19356 ( .B1(n16233), .B2(n20728), .A(n16232), .ZN(n16234) );
  OAI221_X1 U19357 ( .B1(n20843), .B2(n20526), .C1(n20843), .C2(n20846), .A(
        n16234), .ZN(n16235) );
  AOI221_X1 U19358 ( .B1(n16236), .B2(n20727), .C1(n9918), .C2(n20727), .A(
        n16235), .ZN(P1_U3162) );
  NOR2_X1 U19359 ( .A1(n16236), .A2(n9918), .ZN(n16238) );
  OAI22_X1 U19360 ( .A1(n20526), .A2(n16238), .B1(n16237), .B2(n9918), .ZN(
        P1_U3466) );
  INV_X1 U19361 ( .A(n19169), .ZN(n19202) );
  NAND2_X1 U19362 ( .A1(n19202), .A2(n16239), .ZN(n16240) );
  INV_X1 U19363 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20048) );
  OAI22_X1 U19364 ( .A1(n16241), .A2(n16240), .B1(n20048), .B2(n19154), .ZN(
        n16245) );
  INV_X1 U19365 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16243) );
  OAI22_X1 U19366 ( .A1(n21126), .A2(n19144), .B1(n16243), .B2(n16242), .ZN(
        n16244) );
  AOI211_X1 U19367 ( .C1(n19203), .C2(n19216), .A(n16245), .B(n16244), .ZN(
        n16248) );
  NAND4_X1 U19368 ( .A1(n19198), .A2(n16252), .A3(n16246), .A4(n19173), .ZN(
        n16247) );
  OAI211_X1 U19369 ( .C1(n14450), .C2(n19199), .A(n16248), .B(n16247), .ZN(
        P2_U2824) );
  AOI22_X1 U19370 ( .A1(n16249), .A2(n19202), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19211), .ZN(n16250) );
  OAI21_X1 U19371 ( .B1(n20043), .B2(n19154), .A(n16250), .ZN(n16251) );
  AOI21_X1 U19372 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n19167), .A(n16251), .ZN(
        n16256) );
  INV_X1 U19373 ( .A(n16257), .ZN(n16258) );
  AOI211_X1 U19374 ( .C1(n16260), .C2(n16259), .A(n16258), .B(n19972), .ZN(
        n16268) );
  OAI22_X1 U19375 ( .A1(n16262), .A2(n19169), .B1(n16261), .B2(n19144), .ZN(
        n16263) );
  INV_X1 U19376 ( .A(n16263), .ZN(n16265) );
  AOI22_X1 U19377 ( .A1(P2_EBX_REG_27__SCAN_IN), .A2(n19167), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19204), .ZN(n16264) );
  OAI211_X1 U19378 ( .C1(n16266), .C2(n19199), .A(n16265), .B(n16264), .ZN(
        n16267) );
  AOI211_X1 U19379 ( .C1(n19203), .C2(n16269), .A(n16268), .B(n16267), .ZN(
        n16270) );
  INV_X1 U19380 ( .A(n16270), .ZN(P2_U2828) );
  AOI211_X1 U19381 ( .C1(n16273), .C2(n16272), .A(n16271), .B(n19972), .ZN(
        n16279) );
  AOI22_X1 U19382 ( .A1(n16274), .A2(n19202), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19166), .ZN(n16276) );
  AOI22_X1 U19383 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n19167), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19204), .ZN(n16275) );
  OAI211_X1 U19384 ( .C1(n16277), .C2(n19182), .A(n16276), .B(n16275), .ZN(
        n16278) );
  AOI211_X1 U19385 ( .C1(n19187), .C2(n16280), .A(n16279), .B(n16278), .ZN(
        n16281) );
  INV_X1 U19386 ( .A(n16281), .ZN(P2_U2829) );
  AOI211_X1 U19387 ( .C1(n16284), .C2(n16283), .A(n16282), .B(n19972), .ZN(
        n16289) );
  AOI22_X1 U19388 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19211), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19204), .ZN(n16287) );
  OAI211_X1 U19389 ( .C1(n16293), .C2(n20930), .A(n19202), .B(n16285), .ZN(
        n16286) );
  OAI211_X1 U19390 ( .C1(n19207), .C2(n20930), .A(n16287), .B(n16286), .ZN(
        n16288) );
  AOI211_X1 U19391 ( .C1(n19187), .C2(n16290), .A(n16289), .B(n16288), .ZN(
        n16291) );
  OAI21_X1 U19392 ( .B1(n16292), .B2(n19182), .A(n16291), .ZN(P2_U2830) );
  AOI211_X1 U19393 ( .C1(P2_EBX_REG_24__SCAN_IN), .C2(n16294), .A(n19169), .B(
        n16293), .ZN(n16297) );
  INV_X1 U19394 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16295) );
  OAI22_X1 U19395 ( .A1(n16295), .A2(n19144), .B1(n20033), .B2(n19154), .ZN(
        n16296) );
  AOI211_X1 U19396 ( .C1(P2_EBX_REG_24__SCAN_IN), .C2(n19167), .A(n16297), .B(
        n16296), .ZN(n16303) );
  AOI211_X1 U19397 ( .C1(n16300), .C2(n16298), .A(n16299), .B(n19972), .ZN(
        n16301) );
  AOI21_X1 U19398 ( .B1(n19187), .B2(n16324), .A(n16301), .ZN(n16302) );
  OAI211_X1 U19399 ( .C1(n16304), .C2(n19182), .A(n16303), .B(n16302), .ZN(
        P2_U2831) );
  INV_X1 U19400 ( .A(n16305), .ZN(n16316) );
  AOI211_X1 U19401 ( .C1(n16307), .C2(n16306), .A(n9838), .B(n19972), .ZN(
        n16313) );
  AOI22_X1 U19402 ( .A1(n16308), .A2(n19202), .B1(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19211), .ZN(n16310) );
  AOI22_X1 U19403 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(n19167), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19204), .ZN(n16309) );
  OAI211_X1 U19404 ( .C1(n16311), .C2(n19199), .A(n16310), .B(n16309), .ZN(
        n16312) );
  AOI211_X1 U19405 ( .C1(n19203), .C2(n16316), .A(n16313), .B(n16312), .ZN(
        n16314) );
  INV_X1 U19406 ( .A(n16314), .ZN(P2_U2832) );
  AOI22_X1 U19407 ( .A1(n16315), .A2(n19240), .B1(n19262), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16320) );
  AOI22_X1 U19408 ( .A1(n19215), .A2(BUF2_REG_23__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n16319) );
  AOI22_X1 U19409 ( .A1(n16317), .A2(n10867), .B1(n19263), .B2(n16316), .ZN(
        n16318) );
  NAND3_X1 U19410 ( .A1(n16320), .A2(n16319), .A3(n16318), .ZN(P2_U2896) );
  AOI22_X1 U19411 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19376), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19365), .ZN(n16326) );
  OAI22_X1 U19412 ( .A1(n16322), .A2(n9780), .B1(n19385), .B2(n16321), .ZN(
        n16323) );
  AOI21_X1 U19413 ( .B1(n19382), .B2(n16324), .A(n16323), .ZN(n16325) );
  OAI211_X1 U19414 ( .C1(n19374), .C2(n16327), .A(n16326), .B(n16325), .ZN(
        P2_U2990) );
  AOI22_X1 U19415 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19365), .B1(n16370), 
        .B2(n19065), .ZN(n16339) );
  AOI21_X1 U19416 ( .B1(n15564), .B2(n16329), .A(n16328), .ZN(n16390) );
  NAND2_X1 U19417 ( .A1(n16331), .A2(n16330), .ZN(n16333) );
  XOR2_X1 U19418 ( .A(n16333), .B(n16332), .Z(n16393) );
  INV_X1 U19419 ( .A(n16393), .ZN(n16335) );
  INV_X1 U19420 ( .A(n16334), .ZN(n19067) );
  INV_X1 U19421 ( .A(n16336), .ZN(n16337) );
  AOI21_X1 U19422 ( .B1(n16390), .B2(n16378), .A(n16337), .ZN(n16338) );
  OAI211_X1 U19423 ( .C1(n16340), .C2(n16382), .A(n16339), .B(n16338), .ZN(
        P2_U2999) );
  AOI22_X1 U19424 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19365), .B1(n16370), 
        .B2(n19086), .ZN(n16346) );
  AOI21_X1 U19425 ( .B1(n16394), .B2(n15580), .A(n14425), .ZN(n16402) );
  NAND2_X1 U19426 ( .A1(n16342), .A2(n16341), .ZN(n16344) );
  XOR2_X1 U19427 ( .A(n16344), .B(n16343), .Z(n16401) );
  INV_X1 U19428 ( .A(n19090), .ZN(n16400) );
  AOI222_X1 U19429 ( .A1(n16402), .A2(n16378), .B1(n16379), .B2(n16401), .C1(
        n19382), .C2(n16400), .ZN(n16345) );
  OAI211_X1 U19430 ( .C1(n16347), .C2(n16382), .A(n16346), .B(n16345), .ZN(
        P2_U3001) );
  AOI22_X1 U19431 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19185), .B1(n16370), 
        .B2(n19108), .ZN(n16357) );
  NOR2_X1 U19432 ( .A1(n9804), .A2(n16348), .ZN(n16352) );
  NOR2_X1 U19433 ( .A1(n16350), .A2(n16349), .ZN(n16351) );
  XNOR2_X1 U19434 ( .A(n16352), .B(n16351), .ZN(n16414) );
  INV_X1 U19435 ( .A(n19111), .ZN(n16355) );
  AOI21_X1 U19436 ( .B1(n16354), .B2(n15587), .A(n15581), .ZN(n16410) );
  AOI222_X1 U19437 ( .A1(n16414), .A2(n16379), .B1(n19382), .B2(n16355), .C1(
        n16378), .C2(n16410), .ZN(n16356) );
  OAI211_X1 U19438 ( .C1(n16358), .C2(n16382), .A(n16357), .B(n16356), .ZN(
        P2_U3003) );
  AOI22_X1 U19439 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19365), .B1(n16370), 
        .B2(n19127), .ZN(n16363) );
  INV_X1 U19440 ( .A(n19131), .ZN(n16359) );
  AOI222_X1 U19441 ( .A1(n16361), .A2(n16378), .B1(n16379), .B2(n16360), .C1(
        n19382), .C2(n16359), .ZN(n16362) );
  OAI211_X1 U19442 ( .C1(n19123), .C2(n16382), .A(n16363), .B(n16362), .ZN(
        P2_U3005) );
  AOI22_X1 U19443 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19365), .B1(n16370), 
        .B2(n19149), .ZN(n16369) );
  NOR2_X1 U19444 ( .A1(n16364), .A2(n19385), .ZN(n16367) );
  OAI22_X1 U19445 ( .A1(n16365), .A2(n9780), .B1(n14529), .B2(n19153), .ZN(
        n16366) );
  AOI21_X1 U19446 ( .B1(n16367), .B2(n15809), .A(n16366), .ZN(n16368) );
  OAI211_X1 U19447 ( .C1(n19145), .C2(n16382), .A(n16369), .B(n16368), .ZN(
        P2_U3007) );
  AOI22_X1 U19448 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19185), .B1(n16370), 
        .B2(n19175), .ZN(n16381) );
  XOR2_X1 U19449 ( .A(n16371), .B(n16372), .Z(n16452) );
  INV_X1 U19450 ( .A(n16373), .ZN(n16375) );
  NOR2_X1 U19451 ( .A1(n16375), .A2(n16374), .ZN(n16376) );
  XNOR2_X1 U19452 ( .A(n16377), .B(n16376), .ZN(n16449) );
  INV_X1 U19453 ( .A(n19179), .ZN(n16448) );
  AOI222_X1 U19454 ( .A1(n16452), .A2(n16379), .B1(n16378), .B2(n16449), .C1(
        n19382), .C2(n16448), .ZN(n16380) );
  OAI211_X1 U19455 ( .C1(n16383), .C2(n16382), .A(n16381), .B(n16380), .ZN(
        P2_U3009) );
  NOR2_X1 U19456 ( .A1(n11032), .A2(n13196), .ZN(n16388) );
  XNOR2_X1 U19457 ( .A(n16385), .B(n16384), .ZN(n19221) );
  OAI22_X1 U19458 ( .A1(n16386), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n19221), .B2(n16433), .ZN(n16387) );
  AOI211_X1 U19459 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16389), .A(
        n16388), .B(n16387), .ZN(n16392) );
  AOI22_X1 U19460 ( .A1(n16390), .A2(n16450), .B1(n19402), .B2(n19067), .ZN(
        n16391) );
  OAI211_X1 U19461 ( .C1(n16393), .C2(n19395), .A(n16392), .B(n16391), .ZN(
        P2_U3031) );
  OAI21_X1 U19462 ( .B1(n20867), .B2(n16395), .A(n16394), .ZN(n16398) );
  AOI21_X1 U19463 ( .B1(n16397), .B2(n16396), .A(n15761), .ZN(n19224) );
  AOI22_X1 U19464 ( .A1(n16399), .A2(n16398), .B1(n19391), .B2(n19224), .ZN(
        n16404) );
  AOI222_X1 U19465 ( .A1(n16402), .A2(n16450), .B1(n16451), .B2(n16401), .C1(
        n19402), .C2(n16400), .ZN(n16403) );
  OAI211_X1 U19466 ( .C1(n11025), .C2(n13196), .A(n16404), .B(n16403), .ZN(
        P2_U3033) );
  INV_X1 U19467 ( .A(n16405), .ZN(n16406) );
  AOI21_X1 U19468 ( .B1(n16407), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16406), .ZN(n16425) );
  AOI21_X1 U19469 ( .B1(n16409), .B2(n16408), .A(n15774), .ZN(n19230) );
  AOI22_X1 U19470 ( .A1(n16425), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n19391), .B2(n19230), .ZN(n16420) );
  INV_X1 U19471 ( .A(n16410), .ZN(n16412) );
  OAI22_X1 U19472 ( .A1(n16412), .A2(n19406), .B1(n16411), .B2(n19111), .ZN(
        n16413) );
  AOI21_X1 U19473 ( .B1(n16451), .B2(n16414), .A(n16413), .ZN(n16419) );
  NAND2_X1 U19474 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19365), .ZN(n16418) );
  INV_X1 U19475 ( .A(n16415), .ZN(n16416) );
  OAI211_X1 U19476 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n16424), .B(n16416), .ZN(
        n16417) );
  NAND4_X1 U19477 ( .A1(n16420), .A2(n16419), .A3(n16418), .A4(n16417), .ZN(
        P2_U3035) );
  OAI21_X1 U19478 ( .B1(n16421), .B2(n15793), .A(n16408), .ZN(n19233) );
  OAI22_X1 U19479 ( .A1(n16433), .A2(n19233), .B1(n20011), .B2(n13196), .ZN(
        n16422) );
  AOI221_X1 U19480 ( .B1(n16425), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), 
        .C1(n16424), .C2(n16423), .A(n16422), .ZN(n16428) );
  AOI22_X1 U19481 ( .A1(n16426), .A2(n16450), .B1(n19402), .B2(n9846), .ZN(
        n16427) );
  OAI211_X1 U19482 ( .C1(n16429), .C2(n19395), .A(n16428), .B(n16427), .ZN(
        P2_U3036) );
  AOI211_X1 U19483 ( .C1(n20950), .C2(n16434), .A(n16431), .B(n16430), .ZN(
        n16437) );
  OAI21_X1 U19484 ( .B1(n16432), .B2(n15811), .A(n15792), .ZN(n19239) );
  OAI22_X1 U19485 ( .A1(n16435), .A2(n16434), .B1(n16433), .B2(n19239), .ZN(
        n16436) );
  AOI211_X1 U19486 ( .C1(n19365), .C2(P2_REIP_REG_8__SCAN_IN), .A(n16437), .B(
        n16436), .ZN(n16440) );
  AOI22_X1 U19487 ( .A1(n16438), .A2(n16450), .B1(n19402), .B2(n19139), .ZN(
        n16439) );
  OAI211_X1 U19488 ( .C1(n16441), .C2(n19395), .A(n16440), .B(n16439), .ZN(
        P2_U3038) );
  INV_X1 U19489 ( .A(n16442), .ZN(n16446) );
  INV_X1 U19490 ( .A(n16443), .ZN(n16444) );
  AOI21_X1 U19491 ( .B1(n16446), .B2(n16445), .A(n16444), .ZN(n19245) );
  AOI22_X1 U19492 ( .A1(n16447), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n19391), .B2(n19245), .ZN(n16458) );
  AOI222_X1 U19493 ( .A1(n16452), .A2(n16451), .B1(n16450), .B2(n16449), .C1(
        n19402), .C2(n16448), .ZN(n16457) );
  NAND2_X1 U19494 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19185), .ZN(n16456) );
  OAI211_X1 U19495 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n16454), .B(n16453), .ZN(n16455) );
  NAND4_X1 U19496 ( .A1(n16458), .A2(n16457), .A3(n16456), .A4(n16455), .ZN(
        P2_U3041) );
  NAND2_X1 U19497 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20113), .ZN(n19968) );
  INV_X1 U19498 ( .A(n19968), .ZN(n16460) );
  AOI21_X1 U19499 ( .B1(n20114), .B2(n16460), .A(n16459), .ZN(n16499) );
  NAND2_X1 U19500 ( .A1(n16465), .A2(n20085), .ZN(n16463) );
  NOR2_X1 U19501 ( .A1(n16461), .A2(n20092), .ZN(n16462) );
  NAND2_X1 U19502 ( .A1(n16463), .A2(n16462), .ZN(n16464) );
  OAI211_X1 U19503 ( .C1(n16465), .C2(n20085), .A(n16464), .B(n16488), .ZN(
        n16466) );
  AOI21_X1 U19504 ( .B1(n16489), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n16466), .ZN(n16469) );
  NOR2_X1 U19505 ( .A1(n16488), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16467) );
  AOI21_X1 U19506 ( .B1(n16468), .B2(n16488), .A(n16467), .ZN(n16485) );
  OAI211_X1 U19507 ( .C1(n16469), .C2(n20076), .A(n16485), .B(n20069), .ZN(
        n16471) );
  NAND2_X1 U19508 ( .A1(n16469), .A2(n20076), .ZN(n16470) );
  NAND2_X1 U19509 ( .A1(n16471), .A2(n16470), .ZN(n16492) );
  INV_X1 U19510 ( .A(n16472), .ZN(n16475) );
  INV_X1 U19511 ( .A(n10859), .ZN(n16474) );
  AOI22_X1 U19512 ( .A1(n16478), .A2(n16475), .B1(n16474), .B2(n16473), .ZN(
        n16476) );
  OAI21_X1 U19513 ( .B1(n16478), .B2(n16477), .A(n16476), .ZN(n20099) );
  OAI21_X1 U19514 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n16479), .ZN(n16481) );
  OAI211_X1 U19515 ( .C1(n20109), .C2(n11408), .A(n16481), .B(n16480), .ZN(
        n16482) );
  AOI211_X1 U19516 ( .C1(n16483), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n20099), .B(n16482), .ZN(n16484) );
  INV_X1 U19517 ( .A(n16484), .ZN(n16491) );
  NOR2_X1 U19518 ( .A1(n16488), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16487) );
  AOI21_X1 U19519 ( .B1(n16493), .B2(n20069), .A(n16485), .ZN(n16486) );
  AOI211_X1 U19520 ( .C1(n16489), .C2(n16488), .A(n16487), .B(n16486), .ZN(
        n16490) );
  AOI211_X1 U19521 ( .C1(n16493), .C2(n16492), .A(n16491), .B(n16490), .ZN(
        n16504) );
  NAND4_X1 U19522 ( .A1(n16504), .A2(n16502), .A3(n20106), .A4(n16501), .ZN(
        n16497) );
  NAND2_X1 U19523 ( .A1(n20119), .A2(n20089), .ZN(n19287) );
  AOI21_X1 U19524 ( .B1(n20119), .B2(n16494), .A(n20115), .ZN(n16495) );
  AOI21_X1 U19525 ( .B1(n19350), .B2(n20114), .A(n16495), .ZN(n16496) );
  AOI21_X1 U19526 ( .B1(n16497), .B2(n20123), .A(n16496), .ZN(n16498) );
  OAI211_X1 U19527 ( .C1(n20102), .C2(n16500), .A(n16499), .B(n16498), .ZN(
        P2_U3176) );
  NAND3_X1 U19528 ( .A1(n16502), .A2(n20106), .A3(n16501), .ZN(n16503) );
  AND3_X1 U19529 ( .A1(n16504), .A2(n20123), .A3(n16503), .ZN(n19965) );
  AOI211_X1 U19530 ( .C1(n19965), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n16506), 
        .B(n16505), .ZN(n16507) );
  INV_X1 U19531 ( .A(n16507), .ZN(P2_U3593) );
  INV_X1 U19532 ( .A(n18159), .ZN(n18134) );
  AOI22_X1 U19533 ( .A1(n17801), .A2(n18163), .B1(n17953), .B2(n18134), .ZN(
        n17862) );
  NAND2_X1 U19534 ( .A1(n16509), .A2(n17755), .ZN(n17629) );
  XOR2_X1 U19535 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n16524), .Z(
        n16719) );
  INV_X1 U19536 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16720) );
  OAI221_X1 U19537 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16512), .C1(
        n16720), .C2(n16511), .A(n16510), .ZN(n16513) );
  AOI21_X1 U19538 ( .B1(n17800), .B2(n16719), .A(n16513), .ZN(n16519) );
  NAND2_X1 U19539 ( .A1(n17953), .A2(n16514), .ZN(n16537) );
  OAI21_X1 U19540 ( .B1(n16515), .B2(n17876), .A(n16537), .ZN(n16517) );
  AOI22_X1 U19541 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16517), .B1(
        n17873), .B2(n16516), .ZN(n16518) );
  OAI211_X1 U19542 ( .C1(n16520), .C2(n17629), .A(n16519), .B(n16518), .ZN(
        P3_U2800) );
  INV_X1 U19543 ( .A(n16522), .ZN(n16521) );
  NAND2_X1 U19544 ( .A1(n16521), .A2(n17967), .ZN(n16557) );
  NOR2_X1 U19545 ( .A1(n17605), .A2(n16522), .ZN(n16556) );
  OAI211_X1 U19546 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16556), .A(
        n17801), .B(n16523), .ZN(n16531) );
  AOI21_X1 U19547 ( .B1(n16728), .B2(n9860), .A(n16524), .ZN(n16727) );
  OAI21_X1 U19548 ( .B1(n16525), .B2(n17800), .A(n16727), .ZN(n16530) );
  NOR2_X1 U19549 ( .A1(n16526), .A2(n18340), .ZN(n16528) );
  OAI21_X1 U19550 ( .B1(n16528), .B2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16527), .ZN(n16529) );
  NAND4_X1 U19551 ( .A1(n16532), .A2(n16531), .A3(n16530), .A4(n16529), .ZN(
        n16533) );
  AOI21_X1 U19552 ( .B1(n17873), .B2(n16534), .A(n16533), .ZN(n16535) );
  OAI221_X1 U19553 ( .B1(n16537), .B2(n16536), .C1(n16537), .C2(n16557), .A(
        n16535), .ZN(P3_U2801) );
  NAND2_X1 U19554 ( .A1(n16539), .A2(n16538), .ZN(n16541) );
  OAI22_X1 U19555 ( .A1(n16542), .A2(n18923), .B1(n16541), .B2(n16540), .ZN(
        n16543) );
  AOI211_X1 U19556 ( .C1(n16545), .C2(n18237), .A(n16544), .B(n16543), .ZN(
        n16549) );
  AOI22_X1 U19557 ( .A1(n9863), .A2(n16547), .B1(n18135), .B2(n16546), .ZN(
        n16548) );
  OAI211_X1 U19558 ( .C1(n16550), .C2(n18216), .A(n16549), .B(n16548), .ZN(
        P3_U2831) );
  NAND2_X1 U19559 ( .A1(n17468), .A2(n16553), .ZN(n18162) );
  INV_X1 U19560 ( .A(n17624), .ZN(n16564) );
  OAI21_X1 U19561 ( .B1(n17625), .B2(n17802), .A(n16564), .ZN(n17620) );
  AOI22_X1 U19562 ( .A1(n17872), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n17606), .B2(n17802), .ZN(n17619) );
  NAND2_X1 U19563 ( .A1(n17620), .A2(n17619), .ZN(n17618) );
  NAND4_X1 U19564 ( .A1(n16553), .A2(n16552), .A3(n16551), .A4(n17618), .ZN(
        n16554) );
  OAI211_X1 U19565 ( .C1(n16556), .C2(n18162), .A(n16555), .B(n16554), .ZN(
        n16558) );
  OAI221_X1 U19566 ( .B1(n16558), .B2(n18744), .C1(n16558), .C2(n16557), .A(
        n16866), .ZN(n16567) );
  NOR3_X1 U19567 ( .A1(n18279), .A2(n16559), .A3(n17620), .ZN(n16563) );
  INV_X1 U19568 ( .A(n16560), .ZN(n18035) );
  NOR2_X1 U19569 ( .A1(n18029), .A2(n18035), .ZN(n18034) );
  INV_X1 U19570 ( .A(n18028), .ZN(n18104) );
  AOI22_X1 U19571 ( .A1(n18744), .A2(n18104), .B1(n18105), .B2(n18140), .ZN(
        n18078) );
  OAI21_X1 U19572 ( .B1(n18755), .B2(n18925), .A(n18789), .ZN(n18262) );
  AOI21_X1 U19573 ( .B1(n18069), .B2(n18262), .A(n16561), .ZN(n17998) );
  NAND2_X1 U19574 ( .A1(n18078), .A2(n17998), .ZN(n17983) );
  NAND2_X1 U19575 ( .A1(n18034), .A2(n17983), .ZN(n18036) );
  NOR2_X1 U19576 ( .A1(n18043), .A2(n18036), .ZN(n18023) );
  NAND2_X1 U19577 ( .A1(n17973), .A2(n18023), .ZN(n17977) );
  NOR4_X1 U19578 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n21067), .A3(
        n18286), .A4(n17977), .ZN(n16562) );
  AOI211_X1 U19579 ( .C1(n18285), .C2(P3_REIP_REG_28__SCAN_IN), .A(n16563), 
        .B(n16562), .ZN(n16566) );
  OR3_X1 U19580 ( .A1(n16564), .A2(n18175), .A3(n17619), .ZN(n16565) );
  OAI211_X1 U19581 ( .C1(n17606), .C2(n16567), .A(n16566), .B(n16565), .ZN(
        P3_U2834) );
  NOR3_X1 U19582 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16569) );
  NOR4_X1 U19583 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16568) );
  NAND4_X1 U19584 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16569), .A3(n16568), .A4(
        U215), .ZN(U213) );
  INV_X1 U19585 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19288) );
  NOR2_X1 U19586 ( .A1(n16621), .A2(n16570), .ZN(n16573) );
  INV_X1 U19587 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16657) );
  OAI222_X1 U19588 ( .A1(U212), .A2(n19288), .B1(n16623), .B2(n16571), .C1(
        U214), .C2(n16657), .ZN(U216) );
  AOI222_X1 U19589 ( .A1(n16621), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16573), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n16620), .C2(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n16572) );
  INV_X1 U19590 ( .A(n16572), .ZN(U217) );
  AOI222_X1 U19591 ( .A1(n16620), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(n16573), 
        .B2(BUF1_REG_29__SCAN_IN), .C1(n16621), .C2(P1_DATAO_REG_29__SCAN_IN), 
        .ZN(n16574) );
  INV_X1 U19592 ( .A(n16574), .ZN(U218) );
  INV_X1 U19593 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16576) );
  AOI22_X1 U19594 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16620), .ZN(n16575) );
  OAI21_X1 U19595 ( .B1(n16576), .B2(n16623), .A(n16575), .ZN(U219) );
  INV_X1 U19596 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n19431) );
  AOI22_X1 U19597 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16620), .ZN(n16577) );
  OAI21_X1 U19598 ( .B1(n19431), .B2(n16623), .A(n16577), .ZN(U220) );
  INV_X1 U19599 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16579) );
  AOI22_X1 U19600 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16620), .ZN(n16578) );
  OAI21_X1 U19601 ( .B1(n16579), .B2(n16623), .A(n16578), .ZN(U221) );
  INV_X1 U19602 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16581) );
  AOI22_X1 U19603 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16620), .ZN(n16580) );
  OAI21_X1 U19604 ( .B1(n16581), .B2(n16623), .A(n16580), .ZN(U222) );
  AOI22_X1 U19605 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16620), .ZN(n16582) );
  OAI21_X1 U19606 ( .B1(n16583), .B2(n16623), .A(n16582), .ZN(U223) );
  INV_X1 U19607 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n19447) );
  AOI22_X1 U19608 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16620), .ZN(n16584) );
  OAI21_X1 U19609 ( .B1(n19447), .B2(n16623), .A(n16584), .ZN(U224) );
  INV_X1 U19610 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16586) );
  AOI22_X1 U19611 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16620), .ZN(n16585) );
  OAI21_X1 U19612 ( .B1(n16586), .B2(n16623), .A(n16585), .ZN(U225) );
  INV_X1 U19613 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16588) );
  AOI22_X1 U19614 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16620), .ZN(n16587) );
  OAI21_X1 U19615 ( .B1(n16588), .B2(n16623), .A(n16587), .ZN(U226) );
  INV_X1 U19616 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n21048) );
  AOI22_X1 U19617 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16620), .ZN(n16589) );
  OAI21_X1 U19618 ( .B1(n21048), .B2(n16623), .A(n16589), .ZN(U227) );
  INV_X1 U19619 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16591) );
  AOI22_X1 U19620 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16620), .ZN(n16590) );
  OAI21_X1 U19621 ( .B1(n16591), .B2(n16623), .A(n16590), .ZN(U228) );
  AOI22_X1 U19622 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16620), .ZN(n16592) );
  OAI21_X1 U19623 ( .B1(n19426), .B2(n16623), .A(n16592), .ZN(U229) );
  INV_X1 U19624 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n19421) );
  AOI22_X1 U19625 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16620), .ZN(n16593) );
  OAI21_X1 U19626 ( .B1(n19421), .B2(n16623), .A(n16593), .ZN(U230) );
  INV_X1 U19627 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16595) );
  AOI22_X1 U19628 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16620), .ZN(n16594) );
  OAI21_X1 U19629 ( .B1(n16595), .B2(n16623), .A(n16594), .ZN(U231) );
  AOI22_X1 U19630 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16620), .ZN(n16596) );
  OAI21_X1 U19631 ( .B1(n13606), .B2(n16623), .A(n16596), .ZN(U232) );
  AOI22_X1 U19632 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16620), .ZN(n16597) );
  OAI21_X1 U19633 ( .B1(n14289), .B2(n16623), .A(n16597), .ZN(U233) );
  AOI22_X1 U19634 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16620), .ZN(n16598) );
  OAI21_X1 U19635 ( .B1(n16599), .B2(n16623), .A(n16598), .ZN(U234) );
  AOI22_X1 U19636 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16620), .ZN(n16600) );
  OAI21_X1 U19637 ( .B1(n14328), .B2(n16623), .A(n16600), .ZN(U235) );
  AOI22_X1 U19638 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16620), .ZN(n16601) );
  OAI21_X1 U19639 ( .B1(n21125), .B2(n16623), .A(n16601), .ZN(U236) );
  AOI22_X1 U19640 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16620), .ZN(n16602) );
  OAI21_X1 U19641 ( .B1(n16603), .B2(n16623), .A(n16602), .ZN(U237) );
  AOI22_X1 U19642 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16620), .ZN(n16604) );
  OAI21_X1 U19643 ( .B1(n14207), .B2(n16623), .A(n16604), .ZN(U238) );
  AOI22_X1 U19644 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16620), .ZN(n16605) );
  OAI21_X1 U19645 ( .B1(n14190), .B2(n16623), .A(n16605), .ZN(U239) );
  AOI22_X1 U19646 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16620), .ZN(n16606) );
  OAI21_X1 U19647 ( .B1(n16607), .B2(n16623), .A(n16606), .ZN(U240) );
  INV_X1 U19648 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16609) );
  AOI22_X1 U19649 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16620), .ZN(n16608) );
  OAI21_X1 U19650 ( .B1(n16609), .B2(n16623), .A(n16608), .ZN(U241) );
  INV_X1 U19651 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16611) );
  AOI22_X1 U19652 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16620), .ZN(n16610) );
  OAI21_X1 U19653 ( .B1(n16611), .B2(n16623), .A(n16610), .ZN(U242) );
  AOI22_X1 U19654 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16620), .ZN(n16612) );
  OAI21_X1 U19655 ( .B1(n16613), .B2(n16623), .A(n16612), .ZN(U243) );
  INV_X1 U19656 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16615) );
  AOI22_X1 U19657 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16620), .ZN(n16614) );
  OAI21_X1 U19658 ( .B1(n16615), .B2(n16623), .A(n16614), .ZN(U244) );
  INV_X1 U19659 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16617) );
  AOI22_X1 U19660 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16620), .ZN(n16616) );
  OAI21_X1 U19661 ( .B1(n16617), .B2(n16623), .A(n16616), .ZN(U245) );
  INV_X1 U19662 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16619) );
  AOI22_X1 U19663 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16620), .ZN(n16618) );
  OAI21_X1 U19664 ( .B1(n16619), .B2(n16623), .A(n16618), .ZN(U246) );
  INV_X1 U19665 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16624) );
  AOI22_X1 U19666 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16621), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16620), .ZN(n16622) );
  OAI21_X1 U19667 ( .B1(n16624), .B2(n16623), .A(n16622), .ZN(U247) );
  OAI22_X1 U19668 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16654), .ZN(n16625) );
  INV_X1 U19669 ( .A(n16625), .ZN(U251) );
  OAI22_X1 U19670 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16654), .ZN(n16626) );
  INV_X1 U19671 ( .A(n16626), .ZN(U252) );
  INV_X1 U19672 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16627) );
  INV_X1 U19673 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18317) );
  AOI22_X1 U19674 ( .A1(n16654), .A2(n16627), .B1(n18317), .B2(U215), .ZN(U253) );
  INV_X1 U19675 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16628) );
  INV_X1 U19676 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18322) );
  AOI22_X1 U19677 ( .A1(n16654), .A2(n16628), .B1(n18322), .B2(U215), .ZN(U254) );
  INV_X1 U19678 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16629) );
  AOI22_X1 U19679 ( .A1(n16654), .A2(n16629), .B1(n18327), .B2(U215), .ZN(U255) );
  INV_X1 U19680 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16630) );
  INV_X1 U19681 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18333) );
  AOI22_X1 U19682 ( .A1(n16654), .A2(n16630), .B1(n18333), .B2(U215), .ZN(U256) );
  INV_X1 U19683 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16631) );
  INV_X1 U19684 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18338) );
  AOI22_X1 U19685 ( .A1(n16655), .A2(n16631), .B1(n18338), .B2(U215), .ZN(U257) );
  INV_X1 U19686 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16632) );
  AOI22_X1 U19687 ( .A1(n16654), .A2(n16632), .B1(n18345), .B2(U215), .ZN(U258) );
  OAI22_X1 U19688 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16655), .ZN(n16633) );
  INV_X1 U19689 ( .A(n16633), .ZN(U259) );
  INV_X1 U19690 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16634) );
  INV_X1 U19691 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n21044) );
  AOI22_X1 U19692 ( .A1(n16655), .A2(n16634), .B1(n21044), .B2(U215), .ZN(U260) );
  OAI22_X1 U19693 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16654), .ZN(n16635) );
  INV_X1 U19694 ( .A(n16635), .ZN(U261) );
  INV_X1 U19695 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16636) );
  INV_X1 U19696 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17453) );
  AOI22_X1 U19697 ( .A1(n16654), .A2(n16636), .B1(n17453), .B2(U215), .ZN(U262) );
  INV_X1 U19698 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16637) );
  INV_X1 U19699 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17449) );
  AOI22_X1 U19700 ( .A1(n16654), .A2(n16637), .B1(n17449), .B2(U215), .ZN(U263) );
  INV_X1 U19701 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16638) );
  INV_X1 U19702 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17444) );
  AOI22_X1 U19703 ( .A1(n16654), .A2(n16638), .B1(n17444), .B2(U215), .ZN(U264) );
  OAI22_X1 U19704 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16654), .ZN(n16639) );
  INV_X1 U19705 ( .A(n16639), .ZN(U265) );
  OAI22_X1 U19706 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16655), .ZN(n16640) );
  INV_X1 U19707 ( .A(n16640), .ZN(U266) );
  OAI22_X1 U19708 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16654), .ZN(n16641) );
  INV_X1 U19709 ( .A(n16641), .ZN(U267) );
  INV_X1 U19710 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n16642) );
  INV_X1 U19711 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n19420) );
  AOI22_X1 U19712 ( .A1(n16655), .A2(n16642), .B1(n19420), .B2(U215), .ZN(U268) );
  INV_X1 U19713 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n16643) );
  INV_X1 U19714 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n20927) );
  AOI22_X1 U19715 ( .A1(n16654), .A2(n16643), .B1(n20927), .B2(U215), .ZN(U269) );
  INV_X1 U19716 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n16644) );
  INV_X1 U19717 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n21059) );
  AOI22_X1 U19718 ( .A1(n16655), .A2(n16644), .B1(n21059), .B2(U215), .ZN(U270) );
  INV_X1 U19719 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16645) );
  INV_X1 U19720 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n20915) );
  AOI22_X1 U19721 ( .A1(n16654), .A2(n16645), .B1(n20915), .B2(U215), .ZN(U271) );
  OAI22_X1 U19722 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16654), .ZN(n16646) );
  INV_X1 U19723 ( .A(n16646), .ZN(U272) );
  OAI22_X1 U19724 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16655), .ZN(n16647) );
  INV_X1 U19725 ( .A(n16647), .ZN(U273) );
  INV_X1 U19726 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n16648) );
  INV_X1 U19727 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n19449) );
  AOI22_X1 U19728 ( .A1(n16655), .A2(n16648), .B1(n19449), .B2(U215), .ZN(U274) );
  INV_X1 U19729 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n16649) );
  AOI22_X1 U19730 ( .A1(n16655), .A2(n16649), .B1(n18309), .B2(U215), .ZN(U275) );
  OAI22_X1 U19731 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16654), .ZN(n16650) );
  INV_X1 U19732 ( .A(n16650), .ZN(U276) );
  OAI22_X1 U19733 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16654), .ZN(n16651) );
  INV_X1 U19734 ( .A(n16651), .ZN(U277) );
  INV_X1 U19735 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n16652) );
  INV_X1 U19736 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n19430) );
  AOI22_X1 U19737 ( .A1(n16654), .A2(n16652), .B1(n19430), .B2(U215), .ZN(U278) );
  INV_X1 U19738 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16653) );
  INV_X1 U19739 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n21060) );
  AOI22_X1 U19740 ( .A1(n16654), .A2(n16653), .B1(n21060), .B2(U215), .ZN(U279) );
  INV_X1 U19741 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n19292) );
  INV_X1 U19742 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18332) );
  AOI22_X1 U19743 ( .A1(n16654), .A2(n19292), .B1(n18332), .B2(U215), .ZN(U280) );
  INV_X1 U19744 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n20891) );
  AOI22_X1 U19745 ( .A1(n16654), .A2(n20891), .B1(n11079), .B2(U215), .ZN(U281) );
  INV_X1 U19746 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18344) );
  AOI22_X1 U19747 ( .A1(n16655), .A2(n19288), .B1(n18344), .B2(U215), .ZN(U282) );
  INV_X1 U19748 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16656) );
  AOI222_X1 U19749 ( .A1(n19288), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16657), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n16656), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16658) );
  INV_X1 U19750 ( .A(n16660), .ZN(n16659) );
  INV_X1 U19751 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18859) );
  INV_X1 U19752 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20012) );
  AOI22_X1 U19753 ( .A1(n16659), .A2(n18859), .B1(n20012), .B2(n16660), .ZN(
        U347) );
  INV_X1 U19754 ( .A(n16660), .ZN(n16661) );
  INV_X1 U19755 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18857) );
  INV_X1 U19756 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20010) );
  AOI22_X1 U19757 ( .A1(n16661), .A2(n18857), .B1(n20010), .B2(n16660), .ZN(
        U348) );
  INV_X1 U19758 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18854) );
  INV_X1 U19759 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20008) );
  AOI22_X1 U19760 ( .A1(n16659), .A2(n18854), .B1(n20008), .B2(n16660), .ZN(
        U349) );
  INV_X1 U19761 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18853) );
  INV_X1 U19762 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20006) );
  AOI22_X1 U19763 ( .A1(n16659), .A2(n18853), .B1(n20006), .B2(n16660), .ZN(
        U350) );
  INV_X1 U19764 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18851) );
  INV_X1 U19765 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20004) );
  AOI22_X1 U19766 ( .A1(n16659), .A2(n18851), .B1(n20004), .B2(n16660), .ZN(
        U351) );
  INV_X1 U19767 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18848) );
  INV_X1 U19768 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20002) );
  AOI22_X1 U19769 ( .A1(n16659), .A2(n18848), .B1(n20002), .B2(n16660), .ZN(
        U352) );
  INV_X1 U19770 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18847) );
  INV_X1 U19771 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20000) );
  AOI22_X1 U19772 ( .A1(n16661), .A2(n18847), .B1(n20000), .B2(n16660), .ZN(
        U353) );
  INV_X1 U19773 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18845) );
  AOI22_X1 U19774 ( .A1(n16659), .A2(n18845), .B1(n19997), .B2(n16660), .ZN(
        U354) );
  INV_X1 U19775 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18898) );
  INV_X1 U19776 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20047) );
  AOI22_X1 U19777 ( .A1(n16659), .A2(n18898), .B1(n20047), .B2(n16660), .ZN(
        U355) );
  INV_X1 U19778 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18895) );
  INV_X1 U19779 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20044) );
  AOI22_X1 U19780 ( .A1(n16659), .A2(n18895), .B1(n20044), .B2(n16660), .ZN(
        U356) );
  INV_X1 U19781 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18891) );
  INV_X1 U19782 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20042) );
  AOI22_X1 U19783 ( .A1(n16659), .A2(n18891), .B1(n20042), .B2(n16660), .ZN(
        U357) );
  INV_X1 U19784 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18890) );
  INV_X1 U19785 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20039) );
  AOI22_X1 U19786 ( .A1(n16659), .A2(n18890), .B1(n20039), .B2(n16660), .ZN(
        U358) );
  INV_X1 U19787 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18888) );
  INV_X1 U19788 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20038) );
  AOI22_X1 U19789 ( .A1(n16659), .A2(n18888), .B1(n20038), .B2(n16660), .ZN(
        U359) );
  INV_X1 U19790 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18886) );
  INV_X1 U19791 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20036) );
  AOI22_X1 U19792 ( .A1(n16659), .A2(n18886), .B1(n20036), .B2(n16660), .ZN(
        U360) );
  INV_X1 U19793 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18884) );
  INV_X1 U19794 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20034) );
  AOI22_X1 U19795 ( .A1(n16659), .A2(n18884), .B1(n20034), .B2(n16660), .ZN(
        U361) );
  INV_X1 U19796 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18882) );
  INV_X1 U19797 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20032) );
  AOI22_X1 U19798 ( .A1(n16659), .A2(n18882), .B1(n20032), .B2(n16660), .ZN(
        U362) );
  INV_X1 U19799 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18880) );
  INV_X1 U19800 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20030) );
  AOI22_X1 U19801 ( .A1(n16659), .A2(n18880), .B1(n20030), .B2(n16660), .ZN(
        U363) );
  INV_X1 U19802 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18878) );
  INV_X1 U19803 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20028) );
  AOI22_X1 U19804 ( .A1(n16659), .A2(n18878), .B1(n20028), .B2(n16660), .ZN(
        U364) );
  INV_X1 U19805 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18844) );
  INV_X1 U19806 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19995) );
  AOI22_X1 U19807 ( .A1(n16659), .A2(n18844), .B1(n19995), .B2(n16660), .ZN(
        U365) );
  INV_X1 U19808 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18876) );
  INV_X1 U19809 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20026) );
  AOI22_X1 U19810 ( .A1(n16659), .A2(n18876), .B1(n20026), .B2(n16660), .ZN(
        U366) );
  INV_X1 U19811 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18874) );
  INV_X1 U19812 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20024) );
  AOI22_X1 U19813 ( .A1(n16659), .A2(n18874), .B1(n20024), .B2(n16660), .ZN(
        U367) );
  INV_X1 U19814 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18872) );
  INV_X1 U19815 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20023) );
  AOI22_X1 U19816 ( .A1(n16659), .A2(n18872), .B1(n20023), .B2(n16660), .ZN(
        U368) );
  INV_X1 U19817 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18870) );
  INV_X1 U19818 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20021) );
  AOI22_X1 U19819 ( .A1(n16659), .A2(n18870), .B1(n20021), .B2(n16660), .ZN(
        U369) );
  INV_X1 U19820 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18869) );
  INV_X1 U19821 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20888) );
  AOI22_X1 U19822 ( .A1(n16659), .A2(n18869), .B1(n20888), .B2(n16660), .ZN(
        U370) );
  INV_X1 U19823 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18867) );
  INV_X1 U19824 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20019) );
  AOI22_X1 U19825 ( .A1(n16661), .A2(n18867), .B1(n20019), .B2(n16660), .ZN(
        U371) );
  INV_X1 U19826 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18865) );
  INV_X1 U19827 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20018) );
  AOI22_X1 U19828 ( .A1(n16661), .A2(n18865), .B1(n20018), .B2(n16660), .ZN(
        U372) );
  INV_X1 U19829 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18864) );
  INV_X1 U19830 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20016) );
  AOI22_X1 U19831 ( .A1(n16661), .A2(n18864), .B1(n20016), .B2(n16660), .ZN(
        U373) );
  INV_X1 U19832 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18862) );
  INV_X1 U19833 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20015) );
  AOI22_X1 U19834 ( .A1(n16661), .A2(n18862), .B1(n20015), .B2(n16660), .ZN(
        U374) );
  INV_X1 U19835 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18861) );
  INV_X1 U19836 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20013) );
  AOI22_X1 U19837 ( .A1(n16661), .A2(n18861), .B1(n20013), .B2(n16660), .ZN(
        U375) );
  INV_X1 U19838 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18842) );
  INV_X1 U19839 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19994) );
  AOI22_X1 U19840 ( .A1(n16661), .A2(n18842), .B1(n19994), .B2(n16660), .ZN(
        U376) );
  INV_X1 U19841 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16662) );
  INV_X1 U19842 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n21159) );
  NAND2_X1 U19843 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n21159), .ZN(n18832) );
  AOI21_X1 U19844 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(n18832), .A(n18950), 
        .ZN(n18912) );
  INV_X1 U19845 ( .A(n18912), .ZN(n18908) );
  OAI21_X1 U19846 ( .B1(n16662), .B2(n20932), .A(n18908), .ZN(P3_U2633) );
  NAND2_X1 U19847 ( .A1(n18957), .A2(n18748), .ZN(n17538) );
  OAI21_X1 U19848 ( .B1(n16663), .B2(n17538), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16664) );
  OAI21_X1 U19849 ( .B1(n16665), .B2(n18821), .A(n16664), .ZN(P3_U2634) );
  AOI22_X1 U19850 ( .A1(P3_D_C_N_REG_SCAN_IN), .A2(n18969), .B1(n18828), .B2(
        n20932), .ZN(n16666) );
  OAI21_X1 U19851 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n18969), .A(n16666), 
        .ZN(P3_U2635) );
  OAI21_X1 U19852 ( .B1(n18828), .B2(BS16), .A(n18912), .ZN(n18910) );
  OAI21_X1 U19853 ( .B1(n18912), .B2(n16685), .A(n18910), .ZN(P3_U2636) );
  AND3_X1 U19854 ( .A1(n18748), .A2(n16668), .A3(n16667), .ZN(n18751) );
  NOR2_X1 U19855 ( .A1(n18751), .A2(n18817), .ZN(n18951) );
  OAI21_X1 U19856 ( .B1(n18951), .B2(n18294), .A(n9796), .ZN(P3_U2637) );
  NOR4_X1 U19857 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16672) );
  NOR4_X1 U19858 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16671) );
  NOR4_X1 U19859 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16670) );
  NOR4_X1 U19860 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16669) );
  NAND4_X1 U19861 ( .A1(n16672), .A2(n16671), .A3(n16670), .A4(n16669), .ZN(
        n16678) );
  NOR4_X1 U19862 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16676) );
  AOI211_X1 U19863 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_20__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16675) );
  NOR4_X1 U19864 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16674) );
  NOR4_X1 U19865 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16673) );
  NAND4_X1 U19866 ( .A1(n16676), .A2(n16675), .A3(n16674), .A4(n16673), .ZN(
        n16677) );
  NOR2_X1 U19867 ( .A1(n16678), .A2(n16677), .ZN(n18948) );
  INV_X1 U19868 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18905) );
  NOR3_X1 U19869 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16680) );
  OAI21_X1 U19870 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16680), .A(n18948), .ZN(
        n16679) );
  OAI21_X1 U19871 ( .B1(n18948), .B2(n18905), .A(n16679), .ZN(P3_U2638) );
  INV_X1 U19872 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18941) );
  INV_X1 U19873 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18911) );
  AOI21_X1 U19874 ( .B1(n18941), .B2(n18911), .A(n16680), .ZN(n16681) );
  INV_X1 U19875 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18902) );
  INV_X1 U19876 ( .A(n18948), .ZN(n18943) );
  AOI22_X1 U19877 ( .A1(n18948), .A2(n16681), .B1(n18902), .B2(n18943), .ZN(
        P3_U2639) );
  INV_X1 U19878 ( .A(n16682), .ZN(n16684) );
  NAND3_X1 U19879 ( .A1(n18971), .A2(n18962), .A3(n16685), .ZN(n18826) );
  NOR2_X2 U19880 ( .A1(n18926), .A2(n18826), .ZN(n17056) );
  INV_X1 U19881 ( .A(n18819), .ZN(n18686) );
  NOR2_X1 U19882 ( .A1(n18821), .A2(n18686), .ZN(n18814) );
  NOR4_X2 U19883 ( .A1(n18285), .A2(n18973), .A3(n17056), .A4(n18814), .ZN(
        n17060) );
  INV_X1 U19884 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n16700) );
  OAI211_X1 U19885 ( .C1(n18959), .C2(n18958), .A(n18953), .B(n16685), .ZN(
        n18810) );
  OAI211_X2 U19886 ( .C1(n16700), .C2(n18313), .A(n18810), .B(n16702), .ZN(
        n17065) );
  INV_X1 U19887 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18899) );
  INV_X1 U19888 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18885) );
  INV_X1 U19889 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18881) );
  INV_X1 U19890 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n21089) );
  INV_X1 U19891 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n21045) );
  NAND3_X1 U19892 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n17010) );
  NAND2_X1 U19893 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .ZN(n16928) );
  NOR2_X1 U19894 ( .A1(n17010), .A2(n16928), .ZN(n16943) );
  INV_X1 U19895 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18855) );
  NAND2_X1 U19896 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n16984) );
  NOR2_X1 U19897 ( .A1(n18855), .A2(n16984), .ZN(n16927) );
  INV_X1 U19898 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18858) );
  INV_X1 U19899 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18856) );
  NOR2_X1 U19900 ( .A1(n18858), .A2(n18856), .ZN(n16929) );
  NAND4_X1 U19901 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16943), .A3(n16927), 
        .A4(n16929), .ZN(n16921) );
  NOR2_X1 U19902 ( .A1(n21045), .A2(n16921), .ZN(n16911) );
  NAND2_X1 U19903 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16911), .ZN(n16893) );
  NOR2_X1 U19904 ( .A1(n21089), .A2(n16893), .ZN(n16803) );
  INV_X1 U19905 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n21129) );
  NAND2_X1 U19906 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16856) );
  NOR2_X1 U19907 ( .A1(n21129), .A2(n16856), .ZN(n16806) );
  INV_X1 U19908 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18877) );
  NAND3_X1 U19909 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .ZN(n16817) );
  NOR2_X1 U19910 ( .A1(n18877), .A2(n16817), .ZN(n16805) );
  NAND4_X1 U19911 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16803), .A3(n16806), 
        .A4(n16805), .ZN(n16793) );
  NOR2_X1 U19912 ( .A1(n18881), .A2(n16793), .ZN(n16791) );
  NAND2_X1 U19913 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16791), .ZN(n16771) );
  NOR2_X1 U19914 ( .A1(n18885), .A2(n16771), .ZN(n16758) );
  NAND2_X1 U19915 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16758), .ZN(n16704) );
  NOR2_X1 U19916 ( .A1(n17057), .A2(n16704), .ZN(n16752) );
  NAND4_X1 U19917 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16752), .ZN(n16706) );
  NOR3_X1 U19918 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18899), .A3(n16706), 
        .ZN(n16687) );
  AOI21_X1 U19919 ( .B1(n17048), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16687), .ZN(
        n16715) );
  OAI21_X1 U19920 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16688), .A(
        n9860), .ZN(n17615) );
  INV_X1 U19921 ( .A(n17615), .ZN(n16740) );
  NOR3_X1 U19922 ( .A1(n17954), .A2(n17673), .A3(n17672), .ZN(n17647) );
  NAND3_X1 U19923 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(n17647), .ZN(n17612) );
  INV_X1 U19924 ( .A(n17612), .ZN(n16698) );
  NAND2_X1 U19925 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16698), .ZN(
        n16697) );
  AOI21_X1 U19926 ( .B1(n16749), .B2(n16697), .A(n16688), .ZN(n17627) );
  INV_X1 U19927 ( .A(n17647), .ZN(n16690) );
  NOR2_X1 U19928 ( .A1(n10046), .A2(n16690), .ZN(n16689) );
  OAI21_X1 U19929 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16689), .A(
        n17612), .ZN(n17648) );
  INV_X1 U19930 ( .A(n17648), .ZN(n16770) );
  AOI21_X1 U19931 ( .B1(n10046), .B2(n16690), .A(n16689), .ZN(n17664) );
  NOR2_X1 U19932 ( .A1(n17954), .A2(n17673), .ZN(n16691) );
  NOR2_X1 U19933 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n16691), .ZN(
        n17671) );
  NOR2_X1 U19934 ( .A1(n17647), .A2(n17671), .ZN(n17677) );
  INV_X1 U19935 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17690) );
  NAND3_X1 U19936 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17687), .A3(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16692) );
  AOI21_X1 U19937 ( .B1(n17690), .B2(n16692), .A(n16691), .ZN(n17693) );
  NAND2_X1 U19938 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17687), .ZN(
        n16693) );
  XNOR2_X1 U19939 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n16693), .ZN(
        n17708) );
  INV_X1 U19940 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17777) );
  NAND2_X1 U19941 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16694) );
  NAND2_X1 U19942 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17854), .ZN(
        n16976) );
  NOR2_X1 U19943 ( .A1(n16694), .A2(n16976), .ZN(n16930) );
  NAND2_X1 U19944 ( .A1(n16903), .A2(n16930), .ZN(n17796) );
  NOR2_X1 U19945 ( .A1(n17810), .A2(n17796), .ZN(n16902) );
  NAND2_X1 U19946 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16902), .ZN(
        n17761) );
  NOR2_X1 U19947 ( .A1(n17777), .A2(n17761), .ZN(n16881) );
  NAND2_X1 U19948 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16881), .ZN(
        n16857) );
  NOR2_X1 U19949 ( .A1(n17752), .A2(n16857), .ZN(n17724) );
  NAND3_X1 U19950 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A3(n17724), .ZN(n17685) );
  AOI22_X1 U19951 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17687), .B1(
        n17688), .B2(n17685), .ZN(n17718) );
  INV_X1 U19952 ( .A(n16695), .ZN(n17717) );
  NOR2_X1 U19953 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17954), .ZN(
        n17042) );
  AOI21_X1 U19954 ( .B1(n17717), .B2(n17042), .A(n16696), .ZN(n16826) );
  NOR2_X1 U19955 ( .A1(n17718), .A2(n16826), .ZN(n16825) );
  NOR2_X1 U19956 ( .A1(n16825), .A2(n17029), .ZN(n16814) );
  NOR2_X1 U19957 ( .A1(n17677), .A2(n16790), .ZN(n16789) );
  NOR2_X1 U19958 ( .A1(n16789), .A2(n17029), .ZN(n16783) );
  NOR2_X1 U19959 ( .A1(n17664), .A2(n16783), .ZN(n16782) );
  NOR2_X1 U19960 ( .A1(n16782), .A2(n17029), .ZN(n16769) );
  NOR2_X1 U19961 ( .A1(n16770), .A2(n16769), .ZN(n16768) );
  OAI21_X1 U19962 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n16698), .A(
        n16697), .ZN(n17640) );
  INV_X1 U19963 ( .A(n17640), .ZN(n16762) );
  NOR2_X1 U19964 ( .A1(n16760), .A2(n17029), .ZN(n16748) );
  NOR2_X1 U19965 ( .A1(n17627), .A2(n16748), .ZN(n16747) );
  NOR2_X1 U19966 ( .A1(n16747), .A2(n17029), .ZN(n16739) );
  NOR2_X1 U19967 ( .A1(n16740), .A2(n16739), .ZN(n16738) );
  NOR2_X1 U19968 ( .A1(n16738), .A2(n17029), .ZN(n16726) );
  NOR2_X1 U19969 ( .A1(n16727), .A2(n16726), .ZN(n16725) );
  INV_X1 U19970 ( .A(n16718), .ZN(n16713) );
  INV_X1 U19971 ( .A(n17056), .ZN(n18824) );
  OR2_X1 U19972 ( .A1(n16719), .A2(n18824), .ZN(n16699) );
  INV_X1 U19973 ( .A(n18953), .ZN(n18960) );
  NOR2_X1 U19974 ( .A1(n16700), .A2(n18313), .ZN(n16701) );
  OAI211_X2 U19975 ( .C1(P3_STATEBS16_REG_SCAN_IN), .C2(n18960), .A(n16702), 
        .B(n16701), .ZN(n17064) );
  NOR3_X1 U19976 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n17038) );
  INV_X1 U19977 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17328) );
  NAND2_X1 U19978 ( .A1(n17038), .A2(n17328), .ZN(n17034) );
  NOR2_X1 U19979 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17034), .ZN(n17018) );
  INV_X1 U19980 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17006) );
  NAND2_X1 U19981 ( .A1(n17018), .A2(n17006), .ZN(n17005) );
  NOR2_X1 U19982 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17005), .ZN(n16990) );
  NAND2_X1 U19983 ( .A1(n16990), .A2(n17319), .ZN(n16980) );
  NOR2_X1 U19984 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16980), .ZN(n16960) );
  NAND2_X1 U19985 ( .A1(n16960), .A2(n16954), .ZN(n16946) );
  NOR2_X1 U19986 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16946), .ZN(n16945) );
  NAND2_X1 U19987 ( .A1(n16945), .A2(n16937), .ZN(n16936) );
  NOR2_X1 U19988 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16936), .ZN(n16919) );
  NAND2_X1 U19989 ( .A1(n16919), .A2(n16914), .ZN(n16905) );
  NOR2_X1 U19990 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16905), .ZN(n16892) );
  INV_X1 U19991 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16886) );
  NAND2_X1 U19992 ( .A1(n16892), .A2(n16886), .ZN(n16884) );
  NOR2_X1 U19993 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16884), .ZN(n16869) );
  NAND2_X1 U19994 ( .A1(n16869), .A2(n17200), .ZN(n16864) );
  NOR2_X1 U19995 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16864), .ZN(n16846) );
  NAND2_X1 U19996 ( .A1(n16846), .A2(n16838), .ZN(n16836) );
  NOR2_X1 U19997 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16836), .ZN(n16823) );
  INV_X1 U19998 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17145) );
  NAND2_X1 U19999 ( .A1(n16823), .A2(n17145), .ZN(n16820) );
  NOR2_X1 U20000 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16820), .ZN(n16801) );
  INV_X1 U20001 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16797) );
  NAND2_X1 U20002 ( .A1(n16801), .A2(n16797), .ZN(n16796) );
  NOR2_X1 U20003 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16796), .ZN(n16781) );
  INV_X1 U20004 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16776) );
  NAND2_X1 U20005 ( .A1(n16781), .A2(n16776), .ZN(n16775) );
  NOR2_X1 U20006 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16775), .ZN(n16759) );
  NAND2_X1 U20007 ( .A1(n16759), .A2(n17096), .ZN(n16753) );
  NOR2_X1 U20008 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16753), .ZN(n16737) );
  NAND2_X1 U20009 ( .A1(n16737), .A2(n13541), .ZN(n16717) );
  NOR2_X1 U20010 ( .A1(n17064), .A2(n16717), .ZN(n16723) );
  INV_X1 U20011 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16703) );
  NAND2_X1 U20012 ( .A1(n16723), .A2(n16703), .ZN(n16710) );
  NAND3_X1 U20013 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16705) );
  AND2_X1 U20014 ( .A1(n17050), .A2(n16704), .ZN(n16757) );
  NOR2_X1 U20015 ( .A1(n17060), .A2(n16757), .ZN(n16756) );
  INV_X1 U20016 ( .A(n16756), .ZN(n16765) );
  AOI21_X1 U20017 ( .B1(n17050), .B2(n16705), .A(n16765), .ZN(n16736) );
  NOR2_X1 U20018 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16706), .ZN(n16722) );
  INV_X1 U20019 ( .A(n16722), .ZN(n16707) );
  AOI21_X1 U20020 ( .B1(n16736), .B2(n16707), .A(n18897), .ZN(n16708) );
  INV_X1 U20021 ( .A(n16708), .ZN(n16709) );
  OAI211_X1 U20022 ( .C1(n16716), .C2(n17053), .A(n16715), .B(n16714), .ZN(
        P3_U2640) );
  NAND2_X1 U20023 ( .A1(n17035), .A2(n16717), .ZN(n16732) );
  OAI22_X1 U20024 ( .A1(n16736), .A2(n18899), .B1(n16720), .B2(n17053), .ZN(
        n16721) );
  OAI21_X1 U20025 ( .B1(n17048), .B2(n16723), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16724) );
  INV_X1 U20026 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18894) );
  AOI211_X1 U20027 ( .C1(n16727), .C2(n16726), .A(n16725), .B(n18824), .ZN(
        n16731) );
  NAND3_X1 U20028 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16752), .ZN(n16729) );
  OAI22_X1 U20029 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16729), .B1(n16728), 
        .B2(n17053), .ZN(n16730) );
  AOI211_X1 U20030 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n17048), .A(n16731), .B(
        n16730), .ZN(n16735) );
  INV_X1 U20031 ( .A(n16732), .ZN(n16733) );
  OAI21_X1 U20032 ( .B1(n16737), .B2(n13541), .A(n16733), .ZN(n16734) );
  OAI211_X1 U20033 ( .C1(n16736), .C2(n18894), .A(n16735), .B(n16734), .ZN(
        P3_U2642) );
  AOI22_X1 U20034 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17054), .B1(
        n17048), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16746) );
  AOI211_X1 U20035 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16753), .A(n16737), .B(
        n17064), .ZN(n16742) );
  AOI211_X1 U20036 ( .C1(n16740), .C2(n16739), .A(n16738), .B(n18824), .ZN(
        n16741) );
  AOI211_X1 U20037 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16765), .A(n16742), 
        .B(n16741), .ZN(n16745) );
  NAND2_X1 U20038 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16743) );
  OAI211_X1 U20039 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16752), .B(n16743), .ZN(n16744) );
  NAND3_X1 U20040 ( .A1(n16746), .A2(n16745), .A3(n16744), .ZN(P3_U2643) );
  INV_X1 U20041 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18889) );
  AOI211_X1 U20042 ( .C1(n17627), .C2(n16748), .A(n16747), .B(n18824), .ZN(
        n16751) );
  OAI22_X1 U20043 ( .A1(n16749), .A2(n17053), .B1(n17065), .B2(n17096), .ZN(
        n16750) );
  AOI211_X1 U20044 ( .C1(n16752), .C2(n18889), .A(n16751), .B(n16750), .ZN(
        n16755) );
  OAI211_X1 U20045 ( .C1(n16759), .C2(n17096), .A(n17035), .B(n16753), .ZN(
        n16754) );
  OAI211_X1 U20046 ( .C1(n16756), .C2(n18889), .A(n16755), .B(n16754), .ZN(
        P3_U2644) );
  AOI22_X1 U20047 ( .A1(n17048), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n16758), 
        .B2(n16757), .ZN(n16767) );
  AOI211_X1 U20048 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16775), .A(n16759), .B(
        n17064), .ZN(n16764) );
  AOI211_X1 U20049 ( .C1(n16762), .C2(n16761), .A(n16760), .B(n18824), .ZN(
        n16763) );
  AOI211_X1 U20050 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16765), .A(n16764), 
        .B(n16763), .ZN(n16766) );
  OAI211_X1 U20051 ( .C1(n17639), .C2(n17053), .A(n16767), .B(n16766), .ZN(
        P3_U2645) );
  INV_X1 U20052 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18883) );
  OAI21_X1 U20053 ( .B1(n16791), .B2(n17057), .A(n17068), .ZN(n16788) );
  AOI21_X1 U20054 ( .B1(n17050), .B2(n18883), .A(n16788), .ZN(n16779) );
  AOI211_X1 U20055 ( .C1(n16770), .C2(n16769), .A(n16768), .B(n18824), .ZN(
        n16774) );
  NOR3_X1 U20056 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n17057), .A3(n16771), 
        .ZN(n16773) );
  OAI22_X1 U20057 ( .A1(n10047), .A2(n17053), .B1(n17065), .B2(n16776), .ZN(
        n16772) );
  NOR3_X1 U20058 ( .A1(n16774), .A2(n16773), .A3(n16772), .ZN(n16778) );
  OAI211_X1 U20059 ( .C1(n16781), .C2(n16776), .A(n17035), .B(n16775), .ZN(
        n16777) );
  OAI211_X1 U20060 ( .C1(n16779), .C2(n18885), .A(n16778), .B(n16777), .ZN(
        P3_U2646) );
  NOR2_X1 U20061 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17057), .ZN(n16780) );
  AOI22_X1 U20062 ( .A1(n17048), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16791), 
        .B2(n16780), .ZN(n16787) );
  AOI211_X1 U20063 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16796), .A(n16781), .B(
        n17064), .ZN(n16785) );
  AOI211_X1 U20064 ( .C1(n17664), .C2(n16783), .A(n16782), .B(n18824), .ZN(
        n16784) );
  AOI211_X1 U20065 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16788), .A(n16785), 
        .B(n16784), .ZN(n16786) );
  OAI211_X1 U20066 ( .C1(n10046), .C2(n17053), .A(n16787), .B(n16786), .ZN(
        P3_U2647) );
  INV_X1 U20067 ( .A(n16788), .ZN(n16800) );
  AOI211_X1 U20068 ( .C1(n17677), .C2(n16790), .A(n16789), .B(n18824), .ZN(
        n16795) );
  OR2_X1 U20069 ( .A1(n17057), .A2(n16791), .ZN(n16792) );
  OAI22_X1 U20070 ( .A1(n17065), .A2(n16797), .B1(n16793), .B2(n16792), .ZN(
        n16794) );
  AOI211_X1 U20071 ( .C1(n17054), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16795), .B(n16794), .ZN(n16799) );
  OAI211_X1 U20072 ( .C1(n16801), .C2(n16797), .A(n17035), .B(n16796), .ZN(
        n16798) );
  OAI211_X1 U20073 ( .C1(n16800), .C2(n18881), .A(n16799), .B(n16798), .ZN(
        P3_U2648) );
  AOI211_X1 U20074 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16820), .A(n16801), .B(
        n17064), .ZN(n16802) );
  AOI21_X1 U20075 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17048), .A(n16802), .ZN(
        n16812) );
  INV_X1 U20076 ( .A(n16806), .ZN(n16804) );
  NAND2_X1 U20077 ( .A1(n16803), .A2(n17068), .ZN(n16894) );
  NOR2_X1 U20078 ( .A1(n16804), .A2(n16894), .ZN(n16841) );
  NOR2_X1 U20079 ( .A1(n17060), .A2(n17050), .ZN(n16873) );
  AOI21_X1 U20080 ( .B1(n16805), .B2(n16841), .A(n16873), .ZN(n16815) );
  NOR3_X1 U20081 ( .A1(n17057), .A2(n21089), .A3(n16893), .ZN(n16874) );
  NAND2_X1 U20082 ( .A1(n16806), .A2(n16874), .ZN(n16842) );
  NOR4_X1 U20083 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n18877), .A3(n16817), 
        .A4(n16842), .ZN(n16810) );
  AOI211_X1 U20084 ( .C1(n17693), .C2(n16808), .A(n16807), .B(n18824), .ZN(
        n16809) );
  AOI211_X1 U20085 ( .C1(n16815), .C2(P3_REIP_REG_22__SCAN_IN), .A(n16810), 
        .B(n16809), .ZN(n16811) );
  OAI211_X1 U20086 ( .C1(n17690), .C2(n17053), .A(n16812), .B(n16811), .ZN(
        P3_U2649) );
  INV_X1 U20087 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17705) );
  AOI211_X1 U20088 ( .C1(n17708), .C2(n16814), .A(n16813), .B(n18824), .ZN(
        n16819) );
  INV_X1 U20089 ( .A(n16815), .ZN(n16816) );
  AOI221_X1 U20090 ( .B1(n16817), .B2(n18877), .C1(n16842), .C2(n18877), .A(
        n16816), .ZN(n16818) );
  AOI211_X1 U20091 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n17048), .A(n16819), .B(
        n16818), .ZN(n16822) );
  OAI211_X1 U20092 ( .C1(n16823), .C2(n17145), .A(n17035), .B(n16820), .ZN(
        n16821) );
  OAI211_X1 U20093 ( .C1(n17053), .C2(n17705), .A(n16822), .B(n16821), .ZN(
        P3_U2650) );
  AOI211_X1 U20094 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16836), .A(n16823), .B(
        n17064), .ZN(n16824) );
  AOI21_X1 U20095 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17048), .A(n16824), .ZN(
        n16833) );
  INV_X1 U20096 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18873) );
  INV_X1 U20097 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18871) );
  NOR2_X1 U20098 ( .A1(n18873), .A2(n18871), .ZN(n16827) );
  AOI21_X1 U20099 ( .B1(n16827), .B2(n16841), .A(n16873), .ZN(n16831) );
  AOI211_X1 U20100 ( .C1(n17718), .C2(n16826), .A(n16825), .B(n18824), .ZN(
        n16830) );
  INV_X1 U20101 ( .A(n16827), .ZN(n16828) );
  NOR3_X1 U20102 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16828), .A3(n16842), 
        .ZN(n16829) );
  AOI211_X1 U20103 ( .C1(P3_REIP_REG_20__SCAN_IN), .C2(n16831), .A(n16830), 
        .B(n16829), .ZN(n16832) );
  OAI211_X1 U20104 ( .C1(n17688), .C2(n17053), .A(n16833), .B(n16832), .ZN(
        P3_U2651) );
  NAND2_X1 U20105 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17724), .ZN(
        n16849) );
  INV_X1 U20106 ( .A(n16849), .ZN(n16834) );
  OAI21_X1 U20107 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16834), .A(
        n17685), .ZN(n17728) );
  INV_X1 U20108 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16991) );
  NAND2_X1 U20109 ( .A1(n16881), .A2(n16991), .ZN(n16871) );
  OAI21_X1 U20110 ( .B1(n16849), .B2(n16871), .A(n10031), .ZN(n16835) );
  XNOR2_X1 U20111 ( .A(n17728), .B(n16835), .ZN(n16845) );
  NOR3_X1 U20112 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n18871), .A3(n16842), 
        .ZN(n16840) );
  OAI211_X1 U20113 ( .C1(n16846), .C2(n16838), .A(n17035), .B(n16836), .ZN(
        n16837) );
  OAI211_X1 U20114 ( .C1(n17065), .C2(n16838), .A(n16866), .B(n16837), .ZN(
        n16839) );
  AOI211_X1 U20115 ( .C1(n17054), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16840), .B(n16839), .ZN(n16844) );
  NOR2_X1 U20116 ( .A1(n16873), .A2(n16841), .ZN(n16863) );
  NOR2_X1 U20117 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16842), .ZN(n16853) );
  OAI21_X1 U20118 ( .B1(n16863), .B2(n16853), .A(P3_REIP_REG_19__SCAN_IN), 
        .ZN(n16843) );
  OAI211_X1 U20119 ( .C1(n18824), .C2(n16845), .A(n16844), .B(n16843), .ZN(
        P3_U2652) );
  INV_X1 U20120 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17742) );
  AOI211_X1 U20121 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16864), .A(n16846), .B(
        n17064), .ZN(n16847) );
  AOI211_X1 U20122 ( .C1(n17048), .C2(P3_EBX_REG_18__SCAN_IN), .A(n18285), .B(
        n16847), .ZN(n16855) );
  AOI21_X1 U20123 ( .B1(n16991), .B2(n17724), .A(n17029), .ZN(n16848) );
  INV_X1 U20124 ( .A(n16848), .ZN(n16851) );
  OAI21_X1 U20125 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17724), .A(
        n16849), .ZN(n17739) );
  OAI21_X1 U20126 ( .B1(n16851), .B2(n17739), .A(n17056), .ZN(n16850) );
  AOI21_X1 U20127 ( .B1(n16851), .B2(n17739), .A(n16850), .ZN(n16852) );
  AOI211_X1 U20128 ( .C1(n16863), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16853), 
        .B(n16852), .ZN(n16854) );
  OAI211_X1 U20129 ( .C1(n17742), .C2(n17053), .A(n16855), .B(n16854), .ZN(
        P3_U2653) );
  AOI22_X1 U20130 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17054), .B1(
        n17048), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16868) );
  INV_X1 U20131 ( .A(n16874), .ZN(n16875) );
  NOR2_X1 U20132 ( .A1(n16856), .A2(n16875), .ZN(n16862) );
  AOI21_X1 U20133 ( .B1(n17752), .B2(n16857), .A(n17724), .ZN(n17754) );
  INV_X1 U20134 ( .A(n16871), .ZN(n16858) );
  OAI21_X1 U20135 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16881), .A(
        n16857), .ZN(n17762) );
  AOI21_X1 U20136 ( .B1(n16858), .B2(n17762), .A(n17029), .ZN(n16860) );
  OAI21_X1 U20137 ( .B1(n17754), .B2(n16860), .A(n17056), .ZN(n16859) );
  AOI21_X1 U20138 ( .B1(n17754), .B2(n16860), .A(n16859), .ZN(n16861) );
  AOI221_X1 U20139 ( .B1(n16863), .B2(P3_REIP_REG_17__SCAN_IN), .C1(n16862), 
        .C2(n21129), .A(n16861), .ZN(n16867) );
  OAI211_X1 U20140 ( .C1(n16869), .C2(n17200), .A(n17035), .B(n16864), .ZN(
        n16865) );
  NAND4_X1 U20141 ( .A1(n16868), .A2(n16867), .A3(n16866), .A4(n16865), .ZN(
        P3_U2654) );
  INV_X1 U20142 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17763) );
  AOI211_X1 U20143 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16884), .A(n16869), .B(
        n17064), .ZN(n16870) );
  AOI211_X1 U20144 ( .C1(n17048), .C2(P3_EBX_REG_16__SCAN_IN), .A(n18285), .B(
        n16870), .ZN(n16880) );
  NAND2_X1 U20145 ( .A1(n10031), .A2(n16871), .ZN(n16872) );
  XOR2_X1 U20146 ( .A(n17762), .B(n16872), .Z(n16878) );
  INV_X1 U20147 ( .A(n16873), .ZN(n17066) );
  NAND2_X1 U20148 ( .A1(n17066), .A2(n16894), .ZN(n16897) );
  INV_X1 U20149 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18866) );
  NAND2_X1 U20150 ( .A1(n16874), .A2(n18866), .ZN(n16889) );
  INV_X1 U20151 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18868) );
  AOI21_X1 U20152 ( .B1(n16897), .B2(n16889), .A(n18868), .ZN(n16877) );
  NOR3_X1 U20153 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n18866), .A3(n16875), 
        .ZN(n16876) );
  AOI211_X1 U20154 ( .C1(n16878), .C2(n17056), .A(n16877), .B(n16876), .ZN(
        n16879) );
  OAI211_X1 U20155 ( .C1(n17763), .C2(n17053), .A(n16880), .B(n16879), .ZN(
        P3_U2655) );
  AOI21_X1 U20156 ( .B1(n17777), .B2(n17761), .A(n16881), .ZN(n17781) );
  AOI21_X1 U20157 ( .B1(n17775), .B2(n17042), .A(n17029), .ZN(n16883) );
  OAI21_X1 U20158 ( .B1(n17781), .B2(n16883), .A(n17056), .ZN(n16882) );
  AOI21_X1 U20159 ( .B1(n17781), .B2(n16883), .A(n16882), .ZN(n16888) );
  OAI211_X1 U20160 ( .C1(n16892), .C2(n16886), .A(n17035), .B(n16884), .ZN(
        n16885) );
  OAI211_X1 U20161 ( .C1(n17065), .C2(n16886), .A(n16866), .B(n16885), .ZN(
        n16887) );
  AOI211_X1 U20162 ( .C1(n17054), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16888), .B(n16887), .ZN(n16890) );
  OAI211_X1 U20163 ( .C1(n16897), .C2(n18866), .A(n16890), .B(n16889), .ZN(
        P3_U2656) );
  OAI21_X1 U20164 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16902), .A(
        n17761), .ZN(n17787) );
  AOI21_X1 U20165 ( .B1(n16902), .B2(n16991), .A(n17029), .ZN(n16891) );
  XOR2_X1 U20166 ( .A(n17787), .B(n16891), .Z(n16901) );
  AOI211_X1 U20167 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16905), .A(n16892), .B(
        n17064), .ZN(n16899) );
  NOR2_X1 U20168 ( .A1(n17057), .A2(n16893), .ZN(n16895) );
  AOI22_X1 U20169 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n17054), .B1(
        n16895), .B2(n16894), .ZN(n16896) );
  OAI211_X1 U20170 ( .C1(n21089), .C2(n16897), .A(n16896), .B(n16866), .ZN(
        n16898) );
  AOI211_X1 U20171 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17048), .A(n16899), .B(
        n16898), .ZN(n16900) );
  OAI21_X1 U20172 ( .B1(n18824), .B2(n16901), .A(n16900), .ZN(P3_U2657) );
  INV_X1 U20173 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16907) );
  INV_X1 U20174 ( .A(n17796), .ZN(n16916) );
  NAND2_X1 U20175 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16916), .ZN(
        n16915) );
  AOI21_X1 U20176 ( .B1(n16907), .B2(n16915), .A(n16902), .ZN(n17799) );
  INV_X1 U20177 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17818) );
  INV_X1 U20178 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n21050) );
  INV_X1 U20179 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n21122) );
  NAND2_X1 U20180 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17890), .ZN(
        n16999) );
  NOR2_X1 U20181 ( .A1(n21122), .A2(n16999), .ZN(n16988) );
  NAND2_X1 U20182 ( .A1(n16988), .A2(n16991), .ZN(n16977) );
  NOR2_X1 U20183 ( .A1(n17879), .A2(n16977), .ZN(n16967) );
  NAND2_X1 U20184 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16967), .ZN(
        n16956) );
  NOR2_X1 U20185 ( .A1(n21050), .A2(n16956), .ZN(n16942) );
  NAND2_X1 U20186 ( .A1(n16903), .A2(n16942), .ZN(n16917) );
  OAI21_X1 U20187 ( .B1(n17818), .B2(n16917), .A(n10031), .ZN(n16904) );
  XNOR2_X1 U20188 ( .A(n17799), .B(n16904), .ZN(n16910) );
  AOI21_X1 U20189 ( .B1(n17050), .B2(n16921), .A(n17060), .ZN(n16933) );
  NAND2_X1 U20190 ( .A1(n17050), .A2(n21045), .ZN(n16920) );
  INV_X1 U20191 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18863) );
  AOI21_X1 U20192 ( .B1(n16933), .B2(n16920), .A(n18863), .ZN(n16909) );
  OAI211_X1 U20193 ( .C1(n16919), .C2(n16914), .A(n17035), .B(n16905), .ZN(
        n16906) );
  OAI211_X1 U20194 ( .C1(n16907), .C2(n17053), .A(n16866), .B(n16906), .ZN(
        n16908) );
  AOI211_X1 U20195 ( .C1(n16910), .C2(n17056), .A(n16909), .B(n16908), .ZN(
        n16913) );
  NAND3_X1 U20196 ( .A1(n17050), .A2(n16911), .A3(n18863), .ZN(n16912) );
  OAI211_X1 U20197 ( .C1(n16914), .C2(n17065), .A(n16913), .B(n16912), .ZN(
        P3_U2658) );
  AOI22_X1 U20198 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17054), .B1(
        n17048), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n16926) );
  OAI21_X1 U20199 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n16916), .A(
        n16915), .ZN(n17822) );
  NAND2_X1 U20200 ( .A1(n10031), .A2(n16917), .ZN(n16918) );
  XOR2_X1 U20201 ( .A(n17822), .B(n16918), .Z(n16924) );
  AOI211_X1 U20202 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16936), .A(n16919), .B(
        n17064), .ZN(n16923) );
  OAI21_X1 U20203 ( .B1(n16921), .B2(n16920), .A(n16866), .ZN(n16922) );
  AOI211_X1 U20204 ( .C1(n16924), .C2(n17056), .A(n16923), .B(n16922), .ZN(
        n16925) );
  OAI211_X1 U20205 ( .C1(n16933), .C2(n21045), .A(n16926), .B(n16925), .ZN(
        P3_U2659) );
  INV_X1 U20206 ( .A(n16927), .ZN(n16944) );
  NOR3_X1 U20207 ( .A1(n17057), .A2(n17010), .A3(n16928), .ZN(n16985) );
  INV_X1 U20208 ( .A(n16985), .ZN(n16998) );
  NOR2_X1 U20209 ( .A1(n16944), .A2(n16998), .ZN(n16950) );
  AOI21_X1 U20210 ( .B1(n16929), .B2(n16950), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16934) );
  INV_X1 U20211 ( .A(n16930), .ZN(n16955) );
  NOR2_X1 U20212 ( .A1(n17841), .A2(n16955), .ZN(n16941) );
  OAI21_X1 U20213 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16941), .A(
        n17796), .ZN(n17830) );
  AOI21_X1 U20214 ( .B1(n16941), .B2(n16991), .A(n17029), .ZN(n16931) );
  XOR2_X1 U20215 ( .A(n17830), .B(n16931), .Z(n16932) );
  OAI22_X1 U20216 ( .A1(n16934), .A2(n16933), .B1(n18824), .B2(n16932), .ZN(
        n16935) );
  AOI211_X1 U20217 ( .C1(n17048), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18285), .B(
        n16935), .ZN(n16939) );
  OAI211_X1 U20218 ( .C1(n16945), .C2(n16937), .A(n17035), .B(n16936), .ZN(
        n16938) );
  OAI211_X1 U20219 ( .C1(n17053), .C2(n16940), .A(n16939), .B(n16938), .ZN(
        P3_U2660) );
  AOI21_X1 U20220 ( .B1(n17841), .B2(n16955), .A(n16941), .ZN(n17844) );
  NOR2_X1 U20221 ( .A1(n16942), .A2(n17029), .ZN(n16958) );
  XNOR2_X1 U20222 ( .A(n17844), .B(n16958), .ZN(n16953) );
  NAND2_X1 U20223 ( .A1(n16943), .A2(n17068), .ZN(n16975) );
  OAI21_X1 U20224 ( .B1(n16944), .B2(n16975), .A(n17066), .ZN(n16970) );
  NAND2_X1 U20225 ( .A1(n16950), .A2(n18856), .ZN(n16964) );
  AOI21_X1 U20226 ( .B1(n16970), .B2(n16964), .A(n18858), .ZN(n16949) );
  AOI211_X1 U20227 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16946), .A(n16945), .B(
        n17064), .ZN(n16948) );
  OAI22_X1 U20228 ( .A1(n17841), .A2(n17053), .B1(n17065), .B2(n17274), .ZN(
        n16947) );
  NOR4_X1 U20229 ( .A1(n18285), .A2(n16949), .A3(n16948), .A4(n16947), .ZN(
        n16952) );
  NAND3_X1 U20230 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16950), .A3(n18858), 
        .ZN(n16951) );
  OAI211_X1 U20231 ( .C1(n18824), .C2(n16953), .A(n16952), .B(n16951), .ZN(
        P3_U2661) );
  NOR2_X1 U20232 ( .A1(n16960), .A2(n17064), .ZN(n16969) );
  AOI22_X1 U20233 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17054), .B1(
        n16969), .B2(n16954), .ZN(n16963) );
  INV_X1 U20234 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17863) );
  NOR2_X1 U20235 ( .A1(n17863), .A2(n16976), .ZN(n16966) );
  OAI21_X1 U20236 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16966), .A(
        n16955), .ZN(n17856) );
  INV_X1 U20237 ( .A(n17856), .ZN(n16959) );
  NOR2_X1 U20238 ( .A1(n10031), .A2(n18824), .ZN(n17017) );
  AOI21_X1 U20239 ( .B1(n16959), .B2(n16956), .A(n18824), .ZN(n16957) );
  OAI22_X1 U20240 ( .A1(n16959), .A2(n16958), .B1(n17017), .B2(n16957), .ZN(
        n16962) );
  OAI221_X1 U20241 ( .B1(n17048), .B2(n17035), .C1(n17048), .C2(n16960), .A(
        P3_EBX_REG_9__SCAN_IN), .ZN(n16961) );
  AND4_X1 U20242 ( .A1(n16963), .A2(n16866), .A3(n16962), .A4(n16961), .ZN(
        n16965) );
  OAI211_X1 U20243 ( .C1(n16970), .C2(n18856), .A(n16965), .B(n16964), .ZN(
        P3_U2662) );
  AOI21_X1 U20244 ( .B1(n17863), .B2(n16976), .A(n16966), .ZN(n17867) );
  OR2_X1 U20245 ( .A1(n16967), .A2(n17029), .ZN(n16979) );
  XOR2_X1 U20246 ( .A(n17867), .B(n16979), .Z(n16974) );
  NAND2_X1 U20247 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16980), .ZN(n16968) );
  AOI22_X1 U20248 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17048), .B1(n16969), .B2(
        n16968), .ZN(n16973) );
  AOI221_X1 U20249 ( .B1(n16984), .B2(n18855), .C1(n16998), .C2(n18855), .A(
        n16970), .ZN(n16971) );
  AOI211_X1 U20250 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17054), .A(
        n18285), .B(n16971), .ZN(n16972) );
  OAI211_X1 U20251 ( .C1(n18824), .C2(n16974), .A(n16973), .B(n16972), .ZN(
        P3_U2663) );
  NAND2_X1 U20252 ( .A1(n17066), .A2(n16975), .ZN(n17002) );
  INV_X1 U20253 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18852) );
  OAI21_X1 U20254 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16988), .A(
        n16976), .ZN(n17889) );
  INV_X1 U20255 ( .A(n17017), .ZN(n17045) );
  INV_X1 U20256 ( .A(n16977), .ZN(n16989) );
  OAI21_X1 U20257 ( .B1(n16989), .B2(n17889), .A(n17056), .ZN(n16978) );
  AOI22_X1 U20258 ( .A1(n17889), .A2(n16979), .B1(n17045), .B2(n16978), .ZN(
        n16983) );
  OAI211_X1 U20259 ( .C1(n16990), .C2(n17319), .A(n17035), .B(n16980), .ZN(
        n16981) );
  OAI211_X1 U20260 ( .C1(n17065), .C2(n17319), .A(n16866), .B(n16981), .ZN(
        n16982) );
  AOI211_X1 U20261 ( .C1(n17054), .C2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n16983), .B(n16982), .ZN(n16987) );
  OAI211_X1 U20262 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(P3_REIP_REG_6__SCAN_IN), 
        .A(n16985), .B(n16984), .ZN(n16986) );
  OAI211_X1 U20263 ( .C1(n17002), .C2(n18852), .A(n16987), .B(n16986), .ZN(
        P3_U2664) );
  INV_X1 U20264 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18850) );
  AOI21_X1 U20265 ( .B1(n21122), .B2(n16999), .A(n16988), .ZN(n17898) );
  NOR4_X1 U20266 ( .A1(n17898), .A2(n16989), .A3(n18824), .A4(n17029), .ZN(
        n16996) );
  AOI211_X1 U20267 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17005), .A(n16990), .B(
        n17064), .ZN(n16995) );
  NOR2_X1 U20268 ( .A1(n17029), .A2(n16991), .ZN(n17055) );
  AOI211_X1 U20269 ( .C1(n10031), .C2(n16999), .A(n17055), .B(n18824), .ZN(
        n16992) );
  AOI22_X1 U20270 ( .A1(n17048), .A2(P3_EBX_REG_6__SCAN_IN), .B1(n17898), .B2(
        n16992), .ZN(n16993) );
  OAI21_X1 U20271 ( .B1(n21122), .B2(n17053), .A(n16993), .ZN(n16994) );
  NOR4_X1 U20272 ( .A1(n18285), .A2(n16996), .A3(n16995), .A4(n16994), .ZN(
        n16997) );
  OAI221_X1 U20273 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16998), .C1(n18850), 
        .C2(n17002), .A(n16997), .ZN(P3_U2665) );
  INV_X1 U20274 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17009) );
  NOR2_X1 U20275 ( .A1(n17057), .A2(n17010), .ZN(n17015) );
  AOI21_X1 U20276 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n17015), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17003) );
  NAND2_X1 U20277 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17901), .ZN(
        n17012) );
  INV_X1 U20278 ( .A(n16999), .ZN(n17000) );
  AOI21_X1 U20279 ( .B1(n17009), .B2(n17012), .A(n17000), .ZN(n17909) );
  OAI21_X1 U20280 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17012), .A(
        n10031), .ZN(n17014) );
  XOR2_X1 U20281 ( .A(n17909), .B(n17014), .Z(n17001) );
  OAI22_X1 U20282 ( .A1(n17003), .A2(n17002), .B1(n18824), .B2(n17001), .ZN(
        n17004) );
  AOI211_X1 U20283 ( .C1(n17048), .C2(P3_EBX_REG_5__SCAN_IN), .A(n18285), .B(
        n17004), .ZN(n17008) );
  OAI211_X1 U20284 ( .C1(n17018), .C2(n17006), .A(n17035), .B(n17005), .ZN(
        n17007) );
  OAI211_X1 U20285 ( .C1(n17053), .C2(n17009), .A(n17008), .B(n17007), .ZN(
        P3_U2666) );
  INV_X1 U20286 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18846) );
  AOI21_X1 U20287 ( .B1(n17050), .B2(n17010), .A(n17060), .ZN(n17030) );
  NOR2_X1 U20288 ( .A1(n17954), .A2(n17011), .ZN(n17028) );
  OAI21_X1 U20289 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17028), .A(
        n17012), .ZN(n17926) );
  INV_X1 U20290 ( .A(n17926), .ZN(n17016) );
  INV_X1 U20291 ( .A(n17042), .ZN(n17013) );
  NAND2_X1 U20292 ( .A1(n17923), .A2(n17024), .ZN(n17918) );
  OAI22_X1 U20293 ( .A1(n17016), .A2(n17014), .B1(n17013), .B2(n17918), .ZN(
        n17026) );
  AOI22_X1 U20294 ( .A1(n17017), .A2(n17016), .B1(n17015), .B2(n18846), .ZN(
        n17023) );
  AOI211_X1 U20295 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17034), .A(n17018), .B(
        n17064), .ZN(n17021) );
  NAND2_X1 U20296 ( .A1(n18308), .A2(n18973), .ZN(n17071) );
  AOI21_X1 U20297 ( .B1(n17019), .B2(n18754), .A(n17071), .ZN(n17020) );
  AOI211_X1 U20298 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17048), .A(n17021), .B(
        n17020), .ZN(n17022) );
  OAI211_X1 U20299 ( .C1(n17024), .C2(n17053), .A(n17023), .B(n17022), .ZN(
        n17025) );
  AOI211_X1 U20300 ( .C1(n17056), .C2(n17026), .A(n18245), .B(n17025), .ZN(
        n17027) );
  OAI21_X1 U20301 ( .B1(n18846), .B2(n17030), .A(n17027), .ZN(P3_U2667) );
  NAND2_X1 U20302 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17040) );
  AOI21_X1 U20303 ( .B1(n17932), .B2(n17040), .A(n17028), .ZN(n17936) );
  AOI21_X1 U20304 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17042), .A(
        n17029), .ZN(n17041) );
  XOR2_X1 U20305 ( .A(n17936), .B(n17041), .Z(n17033) );
  INV_X1 U20306 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n21047) );
  NAND2_X1 U20307 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17049) );
  AOI221_X1 U20308 ( .B1(n17057), .B2(n21047), .C1(n17049), .C2(n21047), .A(
        n17030), .ZN(n17032) );
  NAND2_X1 U20309 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18765), .ZN(
        n18770) );
  AOI21_X1 U20310 ( .B1(n18770), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n17279), .ZN(n18915) );
  OAI22_X1 U20311 ( .A1(n18915), .A2(n17071), .B1(n17065), .B2(n17328), .ZN(
        n17031) );
  AOI211_X1 U20312 ( .C1(n17056), .C2(n17033), .A(n17032), .B(n17031), .ZN(
        n17037) );
  OAI211_X1 U20313 ( .C1(n17038), .C2(n17328), .A(n17035), .B(n17034), .ZN(
        n17036) );
  OAI211_X1 U20314 ( .C1(n17053), .C2(n17932), .A(n17037), .B(n17036), .ZN(
        P3_U2668) );
  INV_X1 U20315 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17345) );
  INV_X1 U20316 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17339) );
  NAND2_X1 U20317 ( .A1(n17345), .A2(n17339), .ZN(n17039) );
  AOI211_X1 U20318 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17039), .A(n17038), .B(
        n17064), .ZN(n17047) );
  OAI21_X1 U20319 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17040), .ZN(n17945) );
  NOR2_X1 U20320 ( .A1(n21189), .A2(n18940), .ZN(n18781) );
  NOR2_X1 U20321 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18781), .ZN(
        n18768) );
  AOI21_X1 U20322 ( .B1(n18765), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n18768), .ZN(n18931) );
  INV_X1 U20323 ( .A(n17071), .ZN(n18975) );
  AOI22_X1 U20324 ( .A1(n17060), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n18931), 
        .B2(n18975), .ZN(n17044) );
  OAI211_X1 U20325 ( .C1(n17042), .C2(n17945), .A(n17056), .B(n17041), .ZN(
        n17043) );
  OAI211_X1 U20326 ( .C1(n17045), .C2(n17945), .A(n17044), .B(n17043), .ZN(
        n17046) );
  AOI211_X1 U20327 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17048), .A(n17047), .B(
        n17046), .ZN(n17052) );
  OAI211_X1 U20328 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17050), .B(n17049), .ZN(n17051) );
  OAI211_X1 U20329 ( .C1(n17053), .C2(n17949), .A(n17052), .B(n17051), .ZN(
        P3_U2669) );
  OR2_X1 U20330 ( .A1(n18824), .A2(n17055), .ZN(n17063) );
  AOI21_X1 U20331 ( .B1(n17056), .B2(n17055), .A(n17054), .ZN(n17062) );
  OAI22_X1 U20332 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17057), .B1(n17065), 
        .B2(n17339), .ZN(n17059) );
  OAI21_X1 U20333 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17334), .ZN(n17340) );
  OAI22_X1 U20334 ( .A1(n17064), .A2(n17340), .B1(n21180), .B2(n17071), .ZN(
        n17058) );
  AOI211_X1 U20335 ( .C1(n17060), .C2(P3_REIP_REG_1__SCAN_IN), .A(n17059), .B(
        n17058), .ZN(n17061) );
  OAI221_X1 U20336 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17063), .C1(
        n17954), .C2(n17062), .A(n17061), .ZN(P3_U2670) );
  NAND2_X1 U20337 ( .A1(n17065), .A2(n17064), .ZN(n17067) );
  AOI22_X1 U20338 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17067), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n17066), .ZN(n17070) );
  NAND3_X1 U20339 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18928), .A3(
        n17068), .ZN(n17069) );
  OAI211_X1 U20340 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n17071), .A(
        n17070), .B(n17069), .ZN(P3_U2671) );
  AOI22_X1 U20341 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17248), .ZN(n17075) );
  AOI22_X1 U20342 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n17267), .ZN(n17074) );
  AOI22_X1 U20343 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17247), .B1(
        n17294), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17073) );
  AOI22_X1 U20344 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n9758), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n17304), .ZN(n17072) );
  NAND4_X1 U20345 ( .A1(n17075), .A2(n17074), .A3(n17073), .A4(n17072), .ZN(
        n17081) );
  AOI22_X1 U20346 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n17284), .ZN(n17079) );
  AOI22_X1 U20347 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17278), .B1(
        n17305), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17078) );
  AOI22_X1 U20348 ( .A1(n12749), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17295), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17077) );
  AOI22_X1 U20349 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17262), .B1(
        n17277), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17076) );
  NAND4_X1 U20350 ( .A1(n17079), .A2(n17078), .A3(n17077), .A4(n17076), .ZN(
        n17080) );
  NOR2_X1 U20351 ( .A1(n17081), .A2(n17080), .ZN(n17082) );
  XOR2_X1 U20352 ( .A(n17083), .B(n17082), .Z(n17353) );
  NOR2_X1 U20353 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17084), .ZN(n17086) );
  OAI22_X1 U20354 ( .A1(n17353), .A2(n17338), .B1(n17086), .B2(n17085), .ZN(
        P3_U2673) );
  OAI21_X1 U20355 ( .B1(n17092), .B2(n17088), .A(n17087), .ZN(n17365) );
  OAI21_X1 U20356 ( .B1(n17096), .B2(n17097), .A(n20963), .ZN(n17090) );
  NAND2_X1 U20357 ( .A1(n17090), .A2(n17089), .ZN(n17091) );
  OAI21_X1 U20358 ( .B1(n17365), .B2(n17338), .A(n17091), .ZN(P3_U2675) );
  AOI21_X1 U20359 ( .B1(n17093), .B2(n17098), .A(n17092), .ZN(n17366) );
  NAND2_X1 U20360 ( .A1(n17366), .A2(n17343), .ZN(n17094) );
  OAI221_X1 U20361 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17097), .C1(n17096), 
        .C2(n17095), .A(n17094), .ZN(P3_U2676) );
  INV_X1 U20362 ( .A(n17097), .ZN(n17101) );
  AOI21_X1 U20363 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17338), .A(n17106), .ZN(
        n17100) );
  OAI21_X1 U20364 ( .B1(n17102), .B2(n17099), .A(n17098), .ZN(n17374) );
  OAI22_X1 U20365 ( .A1(n17101), .A2(n17100), .B1(n17374), .B2(n17338), .ZN(
        P3_U2677) );
  INV_X1 U20366 ( .A(n17131), .ZN(n17111) );
  AND3_X1 U20367 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n17111), .ZN(n17117) );
  AND2_X1 U20368 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17117), .ZN(n17110) );
  AOI21_X1 U20369 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17338), .A(n17110), .ZN(
        n17105) );
  AOI21_X1 U20370 ( .B1(n17103), .B2(n17107), .A(n17102), .ZN(n17377) );
  INV_X1 U20371 ( .A(n17377), .ZN(n17104) );
  OAI22_X1 U20372 ( .A1(n17106), .A2(n17105), .B1(n17104), .B2(n17338), .ZN(
        P3_U2678) );
  AOI21_X1 U20373 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17338), .A(n17117), .ZN(
        n17109) );
  OAI21_X1 U20374 ( .B1(n17112), .B2(n17108), .A(n17107), .ZN(n17386) );
  OAI22_X1 U20375 ( .A1(n17110), .A2(n17109), .B1(n17386), .B2(n17338), .ZN(
        P3_U2679) );
  AOI22_X1 U20376 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17338), .B1(
        P3_EBX_REG_22__SCAN_IN), .B2(n17111), .ZN(n17116) );
  AOI21_X1 U20377 ( .B1(n17114), .B2(n17113), .A(n17112), .ZN(n17387) );
  INV_X1 U20378 ( .A(n17387), .ZN(n17115) );
  OAI22_X1 U20379 ( .A1(n17117), .A2(n17116), .B1(n17115), .B2(n17338), .ZN(
        P3_U2680) );
  AOI22_X1 U20380 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17128) );
  AOI22_X1 U20381 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17305), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20382 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9754), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17118) );
  OAI21_X1 U20383 ( .B1(n17119), .B2(n20962), .A(n17118), .ZN(n17125) );
  AOI22_X1 U20384 ( .A1(n17248), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17123) );
  AOI22_X1 U20385 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17122) );
  AOI22_X1 U20386 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17121) );
  AOI22_X1 U20387 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17120) );
  NAND4_X1 U20388 ( .A1(n17123), .A2(n17122), .A3(n17121), .A4(n17120), .ZN(
        n17124) );
  AOI211_X1 U20389 ( .C1(n17296), .C2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n17125), .B(n17124), .ZN(n17126) );
  NAND3_X1 U20390 ( .A1(n17128), .A2(n17127), .A3(n17126), .ZN(n17393) );
  INV_X1 U20391 ( .A(n17393), .ZN(n17130) );
  NAND3_X1 U20392 ( .A1(n17131), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17338), 
        .ZN(n17129) );
  OAI221_X1 U20393 ( .B1(n17131), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17338), 
        .C2(n17130), .A(n17129), .ZN(P3_U2681) );
  NAND2_X1 U20394 ( .A1(n17338), .A2(n17132), .ZN(n17159) );
  AOI22_X1 U20395 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13466), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17142) );
  AOI22_X1 U20396 ( .A1(n17248), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17305), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U20397 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17133) );
  OAI21_X1 U20398 ( .B1(n17218), .B2(n18337), .A(n17133), .ZN(n17139) );
  AOI22_X1 U20399 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17137) );
  AOI22_X1 U20400 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17136) );
  AOI22_X1 U20401 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17135) );
  AOI22_X1 U20402 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17134) );
  NAND4_X1 U20403 ( .A1(n17137), .A2(n17136), .A3(n17135), .A4(n17134), .ZN(
        n17138) );
  AOI211_X1 U20404 ( .C1(n17294), .C2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n17139), .B(n17138), .ZN(n17140) );
  NAND3_X1 U20405 ( .A1(n17142), .A2(n17141), .A3(n17140), .ZN(n17399) );
  AOI22_X1 U20406 ( .A1(n17343), .A2(n17399), .B1(n17143), .B2(n17145), .ZN(
        n17144) );
  OAI21_X1 U20407 ( .B1(n17145), .B2(n17159), .A(n17144), .ZN(P3_U2682) );
  AOI22_X1 U20408 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U20409 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17277), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17154) );
  INV_X1 U20410 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18331) );
  AOI22_X1 U20411 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13466), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17146) );
  OAI21_X1 U20412 ( .B1(n17218), .B2(n18331), .A(n17146), .ZN(n17152) );
  AOI22_X1 U20413 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17305), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17150) );
  AOI22_X1 U20414 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17149) );
  AOI22_X1 U20415 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17148) );
  AOI22_X1 U20416 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17147) );
  NAND4_X1 U20417 ( .A1(n17150), .A2(n17149), .A3(n17148), .A4(n17147), .ZN(
        n17151) );
  AOI211_X1 U20418 ( .C1(n17248), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n17152), .B(n17151), .ZN(n17153) );
  NAND3_X1 U20419 ( .A1(n17155), .A2(n17154), .A3(n17153), .ZN(n17404) );
  NAND2_X1 U20420 ( .A1(n17343), .A2(n17404), .ZN(n17156) );
  OAI221_X1 U20421 ( .B1(n17159), .B2(n17158), .C1(n17159), .C2(n17157), .A(
        n17156), .ZN(P3_U2683) );
  INV_X1 U20422 ( .A(n17173), .ZN(n17160) );
  OAI21_X1 U20423 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17160), .A(n17338), .ZN(
        n17171) );
  AOI22_X1 U20424 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17295), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17164) );
  AOI22_X1 U20425 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17163) );
  AOI22_X1 U20426 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17162) );
  AOI22_X1 U20427 ( .A1(n17248), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17161) );
  NAND4_X1 U20428 ( .A1(n17164), .A2(n17163), .A3(n17162), .A4(n17161), .ZN(
        n17170) );
  AOI22_X1 U20429 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17168) );
  AOI22_X1 U20430 ( .A1(n17305), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13466), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17167) );
  AOI22_X1 U20431 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17166) );
  AOI22_X1 U20432 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9754), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17165) );
  NAND4_X1 U20433 ( .A1(n17168), .A2(n17167), .A3(n17166), .A4(n17165), .ZN(
        n17169) );
  NOR2_X1 U20434 ( .A1(n17170), .A2(n17169), .ZN(n17412) );
  OAI22_X1 U20435 ( .A1(n17172), .A2(n17171), .B1(n17412), .B2(n17338), .ZN(
        P3_U2684) );
  NAND2_X1 U20436 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17173), .ZN(n17187) );
  AOI22_X1 U20437 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17305), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17177) );
  AOI22_X1 U20438 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17176) );
  AOI22_X1 U20439 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17175) );
  AOI22_X1 U20440 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17174) );
  NAND4_X1 U20441 ( .A1(n17177), .A2(n17176), .A3(n17175), .A4(n17174), .ZN(
        n17183) );
  AOI22_X1 U20442 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17181) );
  AOI22_X1 U20443 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U20444 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U20445 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17178) );
  NAND4_X1 U20446 ( .A1(n17181), .A2(n17180), .A3(n17179), .A4(n17178), .ZN(
        n17182) );
  NOR2_X1 U20447 ( .A1(n17183), .A2(n17182), .ZN(n17418) );
  INV_X1 U20448 ( .A(n17341), .ZN(n17342) );
  INV_X1 U20449 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17184) );
  NAND3_X1 U20450 ( .A1(n17185), .A2(n17342), .A3(n17184), .ZN(n17186) );
  OAI221_X1 U20451 ( .B1(n17343), .B2(n17187), .C1(n17338), .C2(n17418), .A(
        n17186), .ZN(P3_U2685) );
  AOI22_X1 U20452 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17191) );
  AOI22_X1 U20453 ( .A1(n17305), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17190) );
  AOI22_X1 U20454 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17189) );
  AOI22_X1 U20455 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17188) );
  NAND4_X1 U20456 ( .A1(n17191), .A2(n17190), .A3(n17189), .A4(n17188), .ZN(
        n17198) );
  AOI22_X1 U20457 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17196) );
  AOI22_X1 U20458 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17195) );
  AOI22_X1 U20459 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17194) );
  AOI22_X1 U20460 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17193) );
  NAND4_X1 U20461 ( .A1(n17196), .A2(n17195), .A3(n17194), .A4(n17193), .ZN(
        n17197) );
  NOR2_X1 U20462 ( .A1(n17198), .A2(n17197), .ZN(n17423) );
  OR3_X1 U20463 ( .A1(n17199), .A2(n17341), .A3(P3_EBX_REG_17__SCAN_IN), .ZN(
        n17203) );
  NAND2_X1 U20464 ( .A1(n18348), .A2(n17199), .ZN(n17216) );
  AOI21_X1 U20465 ( .B1(n17216), .B2(n17346), .A(n17200), .ZN(n17201) );
  INV_X1 U20466 ( .A(n17201), .ZN(n17202) );
  OAI211_X1 U20467 ( .C1(n17423), .C2(n17338), .A(n17203), .B(n17202), .ZN(
        P3_U2686) );
  NAND3_X1 U20468 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(n17244), .ZN(n17215) );
  AOI22_X1 U20469 ( .A1(n17248), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17207) );
  AOI22_X1 U20470 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17206) );
  AOI22_X1 U20471 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17205) );
  AOI22_X1 U20472 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17204) );
  NAND4_X1 U20473 ( .A1(n17207), .A2(n17206), .A3(n17205), .A4(n17204), .ZN(
        n17213) );
  AOI22_X1 U20474 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17294), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17211) );
  AOI22_X1 U20475 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U20476 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17209) );
  AOI22_X1 U20477 ( .A1(n17305), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17208) );
  NAND4_X1 U20478 ( .A1(n17211), .A2(n17210), .A3(n17209), .A4(n17208), .ZN(
        n17212) );
  NOR2_X1 U20479 ( .A1(n17213), .A2(n17212), .ZN(n17430) );
  INV_X1 U20480 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17214) );
  NAND2_X1 U20481 ( .A1(n17338), .A2(n17215), .ZN(n17229) );
  OAI222_X1 U20482 ( .A1(n17216), .A2(n17215), .B1(n17338), .B2(n17430), .C1(
        n17214), .C2(n17229), .ZN(P3_U2687) );
  AOI22_X1 U20483 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17278), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n17247), .ZN(n17228) );
  AOI22_X1 U20484 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17305), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17262), .ZN(n17227) );
  INV_X1 U20485 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n20951) );
  AOI22_X1 U20486 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17267), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17284), .ZN(n17217) );
  OAI21_X1 U20487 ( .B1(n17218), .B2(n20951), .A(n17217), .ZN(n17225) );
  AOI22_X1 U20488 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17223) );
  AOI22_X1 U20489 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9754), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U20490 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17248), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n17219), .ZN(n17221) );
  AOI22_X1 U20491 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n9758), .ZN(n17220) );
  NAND4_X1 U20492 ( .A1(n17223), .A2(n17222), .A3(n17221), .A4(n17220), .ZN(
        n17224) );
  AOI211_X1 U20493 ( .C1(n17277), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n17225), .B(n17224), .ZN(n17226) );
  NAND3_X1 U20494 ( .A1(n17228), .A2(n17227), .A3(n17226), .ZN(n17433) );
  INV_X1 U20495 ( .A(n17433), .ZN(n17231) );
  AOI21_X1 U20496 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17244), .A(
        P3_EBX_REG_15__SCAN_IN), .ZN(n17230) );
  OAI22_X1 U20497 ( .A1(n17231), .A2(n17338), .B1(n17230), .B2(n17229), .ZN(
        P3_U2688) );
  AOI22_X1 U20498 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17242) );
  AOI22_X1 U20499 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17241) );
  AOI22_X1 U20500 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17248), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17232) );
  OAI21_X1 U20501 ( .B1(n17233), .B2(n20962), .A(n17232), .ZN(n17239) );
  AOI22_X1 U20502 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17237) );
  AOI22_X1 U20503 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17236) );
  AOI22_X1 U20504 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17235) );
  AOI22_X1 U20505 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17234) );
  NAND4_X1 U20506 ( .A1(n17237), .A2(n17236), .A3(n17235), .A4(n17234), .ZN(
        n17238) );
  AOI211_X1 U20507 ( .C1(n17279), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n17239), .B(n17238), .ZN(n17240) );
  NAND3_X1 U20508 ( .A1(n17242), .A2(n17241), .A3(n17240), .ZN(n17437) );
  INV_X1 U20509 ( .A(n17437), .ZN(n17246) );
  NAND2_X1 U20510 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17244), .ZN(n17243) );
  OAI21_X1 U20511 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17244), .A(n17243), .ZN(
        n17245) );
  AOI22_X1 U20512 ( .A1(n17343), .A2(n17246), .B1(n17245), .B2(n17338), .ZN(
        P3_U2689) );
  AOI22_X1 U20513 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17252) );
  AOI22_X1 U20514 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17251) );
  AOI22_X1 U20515 ( .A1(n17248), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17250) );
  AOI22_X1 U20516 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17249) );
  NAND4_X1 U20517 ( .A1(n17252), .A2(n17251), .A3(n17250), .A4(n17249), .ZN(
        n17258) );
  AOI22_X1 U20518 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17256) );
  AOI22_X1 U20519 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17255) );
  AOI22_X1 U20520 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17277), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17254) );
  AOI22_X1 U20521 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17305), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17253) );
  NAND4_X1 U20522 ( .A1(n17256), .A2(n17255), .A3(n17254), .A4(n17253), .ZN(
        n17257) );
  NOR2_X1 U20523 ( .A1(n17258), .A2(n17257), .ZN(n17446) );
  AOI221_X1 U20524 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17260), .C1(n17259), 
        .C2(n17260), .A(n17343), .ZN(n17261) );
  AOI21_X1 U20525 ( .B1(n17446), .B2(n17343), .A(n17261), .ZN(P3_U2691) );
  AOI22_X1 U20526 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17266) );
  AOI22_X1 U20527 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17265) );
  AOI22_X1 U20528 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13466), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17264) );
  AOI22_X1 U20529 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17247), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17263) );
  NAND4_X1 U20530 ( .A1(n17266), .A2(n17265), .A3(n17264), .A4(n17263), .ZN(
        n17273) );
  AOI22_X1 U20531 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17271) );
  AOI22_X1 U20532 ( .A1(n17303), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17294), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17270) );
  AOI22_X1 U20533 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17279), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17269) );
  AOI22_X1 U20534 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17305), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17268) );
  NAND4_X1 U20535 ( .A1(n17271), .A2(n17270), .A3(n17269), .A4(n17268), .ZN(
        n17272) );
  NOR2_X1 U20536 ( .A1(n17273), .A2(n17272), .ZN(n17457) );
  NOR2_X1 U20537 ( .A1(n17343), .A2(n17275), .ZN(n17292) );
  OAI222_X1 U20538 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18348), .B1(
        P3_EBX_REG_10__SCAN_IN), .B2(n17275), .C1(n17292), .C2(n17274), .ZN(
        n17276) );
  OAI21_X1 U20539 ( .B1(n17457), .B2(n17338), .A(n17276), .ZN(P3_U2693) );
  AOI22_X1 U20540 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17283) );
  AOI22_X1 U20541 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17305), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17282) );
  AOI22_X1 U20542 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17281) );
  AOI22_X1 U20543 ( .A1(n17279), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17280) );
  NAND4_X1 U20544 ( .A1(n17283), .A2(n17282), .A3(n17281), .A4(n17280), .ZN(
        n17290) );
  AOI22_X1 U20545 ( .A1(n17294), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17288) );
  AOI22_X1 U20546 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17295), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17287) );
  AOI22_X1 U20547 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U20548 ( .A1(n17303), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17285) );
  NAND4_X1 U20549 ( .A1(n17288), .A2(n17287), .A3(n17286), .A4(n17285), .ZN(
        n17289) );
  NOR2_X1 U20550 ( .A1(n17290), .A2(n17289), .ZN(n17460) );
  NOR2_X1 U20551 ( .A1(n17291), .A2(n17312), .ZN(n17315) );
  OAI21_X1 U20552 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17315), .A(n17292), .ZN(
        n17293) );
  OAI21_X1 U20553 ( .B1(n17460), .B2(n17338), .A(n17293), .ZN(P3_U2694) );
  AOI22_X1 U20554 ( .A1(n17295), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17294), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17300) );
  AOI22_X1 U20555 ( .A1(n17296), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17299) );
  AOI22_X1 U20556 ( .A1(n12749), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15900), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17298) );
  AOI22_X1 U20557 ( .A1(n9754), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(n9758), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17297) );
  NAND4_X1 U20558 ( .A1(n17300), .A2(n17299), .A3(n17298), .A4(n17297), .ZN(
        n17311) );
  AOI22_X1 U20559 ( .A1(n17247), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17309) );
  AOI22_X1 U20560 ( .A1(n17303), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17308) );
  AOI22_X1 U20561 ( .A1(n17305), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17307) );
  AOI22_X1 U20562 ( .A1(n17277), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13466), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17306) );
  NAND4_X1 U20563 ( .A1(n17309), .A2(n17308), .A3(n17307), .A4(n17306), .ZN(
        n17310) );
  NOR2_X1 U20564 ( .A1(n17311), .A2(n17310), .ZN(n17467) );
  INV_X1 U20565 ( .A(n17312), .ZN(n17313) );
  OAI21_X1 U20566 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17313), .A(n17338), .ZN(
        n17314) );
  OAI22_X1 U20567 ( .A1(n17467), .A2(n17338), .B1(n17315), .B2(n17314), .ZN(
        P3_U2695) );
  OR2_X1 U20568 ( .A1(n17316), .A2(n17319), .ZN(n17322) );
  INV_X1 U20569 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18353) );
  INV_X1 U20570 ( .A(n17317), .ZN(n17320) );
  NOR2_X1 U20571 ( .A1(n17318), .A2(n17341), .ZN(n17330) );
  NAND3_X1 U20572 ( .A1(n17320), .A2(n17330), .A3(n17319), .ZN(n17321) );
  OAI221_X1 U20573 ( .B1(n17343), .B2(n17322), .C1(n17338), .C2(n18353), .A(
        n17321), .ZN(P3_U2696) );
  NAND2_X1 U20574 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17330), .ZN(n17324) );
  INV_X1 U20575 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18343) );
  NAND3_X1 U20576 ( .A1(n17324), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n17338), .ZN(
        n17323) );
  OAI221_X1 U20577 ( .B1(n17324), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n17338), 
        .C2(n18343), .A(n17323), .ZN(P3_U2697) );
  OAI211_X1 U20578 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n17325), .A(n17324), .B(
        n17338), .ZN(n17326) );
  OAI21_X1 U20579 ( .B1(n17338), .B2(n18337), .A(n17326), .ZN(P3_U2698) );
  NAND2_X1 U20580 ( .A1(n17327), .A2(n17342), .ZN(n17331) );
  NOR2_X1 U20581 ( .A1(n17328), .A2(n17331), .ZN(n17333) );
  AOI21_X1 U20582 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17338), .A(n17333), .ZN(
        n17329) );
  OAI22_X1 U20583 ( .A1(n17330), .A2(n17329), .B1(n18331), .B2(n17338), .ZN(
        P3_U2699) );
  INV_X1 U20584 ( .A(n17331), .ZN(n17336) );
  AOI21_X1 U20585 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17338), .A(n17336), .ZN(
        n17332) );
  INV_X1 U20586 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18326) );
  OAI22_X1 U20587 ( .A1(n17333), .A2(n17332), .B1(n18326), .B2(n17338), .ZN(
        P3_U2700) );
  INV_X1 U20588 ( .A(n17334), .ZN(n17335) );
  AOI221_X1 U20589 ( .B1(n17335), .B2(n17346), .C1(n17431), .C2(n17346), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17337) );
  AOI211_X1 U20590 ( .C1(n17343), .C2(n18321), .A(n17337), .B(n17336), .ZN(
        P3_U2701) );
  INV_X1 U20591 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18316) );
  OAI222_X1 U20592 ( .A1(n17341), .A2(n17340), .B1(n17339), .B2(n17346), .C1(
        n18316), .C2(n17338), .ZN(P3_U2702) );
  AOI22_X1 U20593 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17343), .B1(
        n17342), .B2(n17345), .ZN(n17344) );
  OAI21_X1 U20594 ( .B1(n17346), .B2(n17345), .A(n17344), .ZN(P3_U2703) );
  INV_X1 U20595 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17565) );
  INV_X1 U20596 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17559) );
  INV_X1 U20597 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17553) );
  INV_X1 U20598 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17544) );
  INV_X1 U20599 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17604) );
  NAND2_X1 U20600 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n17494) );
  INV_X1 U20601 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17580) );
  INV_X1 U20602 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17578) );
  NAND4_X1 U20603 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17347) );
  NOR4_X1 U20604 ( .A1(n17494), .A2(n17580), .A3(n17578), .A4(n17347), .ZN(
        n17436) );
  NAND2_X1 U20605 ( .A1(n17498), .A2(n17436), .ZN(n17464) );
  NAND4_X1 U20606 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n17348)
         );
  INV_X1 U20607 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n20860) );
  INV_X1 U20608 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17549) );
  INV_X1 U20609 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17547) );
  NOR3_X1 U20610 ( .A1(n20860), .A2(n17549), .A3(n17547), .ZN(n17408) );
  NAND2_X1 U20611 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17408), .ZN(n17398) );
  NAND2_X1 U20612 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17389), .ZN(n17388) );
  INV_X1 U20613 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17569) );
  OR2_X1 U20614 ( .A1(n17358), .A2(n17569), .ZN(n17351) );
  NAND2_X1 U20615 ( .A1(n17349), .A2(n17375), .ZN(n17392) );
  OAI21_X1 U20616 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17351), .A(n17350), .ZN(
        P3_U2704) );
  NOR2_X2 U20617 ( .A1(n17352), .A2(n17486), .ZN(n17425) );
  OAI22_X1 U20618 ( .A1(n17353), .A2(n17487), .B1(n11079), .B2(n17392), .ZN(
        n17354) );
  AOI21_X1 U20619 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17425), .A(n17354), .ZN(
        n17355) );
  OAI221_X1 U20620 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17358), .C1(n17569), 
        .C2(n17356), .A(n17355), .ZN(P3_U2705) );
  AOI22_X1 U20621 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17425), .B1(n17492), .B2(
        n17357), .ZN(n17360) );
  OAI211_X1 U20622 ( .C1(n17361), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17486), .B(
        n17358), .ZN(n17359) );
  OAI211_X1 U20623 ( .C1(n17392), .C2(n18332), .A(n17360), .B(n17359), .ZN(
        P3_U2706) );
  AOI22_X1 U20624 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17425), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17424), .ZN(n17364) );
  AOI211_X1 U20625 ( .C1(n17565), .C2(n17367), .A(n17361), .B(n17375), .ZN(
        n17362) );
  INV_X1 U20626 ( .A(n17362), .ZN(n17363) );
  OAI211_X1 U20627 ( .C1(n17365), .C2(n17487), .A(n17364), .B(n17363), .ZN(
        P3_U2707) );
  AOI22_X1 U20628 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17425), .B1(n17492), .B2(
        n17366), .ZN(n17370) );
  OAI211_X1 U20629 ( .C1(n17368), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17486), .B(
        n17367), .ZN(n17369) );
  OAI211_X1 U20630 ( .C1(n17392), .C2(n19430), .A(n17370), .B(n17369), .ZN(
        P3_U2708) );
  AOI22_X1 U20631 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17425), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17424), .ZN(n17373) );
  OAI211_X1 U20632 ( .C1(n17381), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17486), .B(
        n17371), .ZN(n17372) );
  OAI211_X1 U20633 ( .C1(n17374), .C2(n17487), .A(n17373), .B(n17372), .ZN(
        P3_U2709) );
  OAI21_X1 U20634 ( .B1(n17559), .B2(n17375), .A(n17382), .ZN(n17376) );
  INV_X1 U20635 ( .A(n17376), .ZN(n17380) );
  AOI22_X1 U20636 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n17424), .B1(n17492), .B2(
        n17377), .ZN(n17379) );
  NAND2_X1 U20637 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17425), .ZN(n17378) );
  OAI211_X1 U20638 ( .C1(n17381), .C2(n17380), .A(n17379), .B(n17378), .ZN(
        P3_U2710) );
  AOI22_X1 U20639 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17425), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17424), .ZN(n17385) );
  OAI211_X1 U20640 ( .C1(n17383), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17486), .B(
        n17382), .ZN(n17384) );
  OAI211_X1 U20641 ( .C1(n17386), .C2(n17487), .A(n17385), .B(n17384), .ZN(
        P3_U2711) );
  AOI22_X1 U20642 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17425), .B1(n17492), .B2(
        n17387), .ZN(n17391) );
  OAI211_X1 U20643 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17389), .A(n17486), .B(
        n17388), .ZN(n17390) );
  OAI211_X1 U20644 ( .C1(n17392), .C2(n19449), .A(n17391), .B(n17390), .ZN(
        P3_U2712) );
  NAND2_X1 U20645 ( .A1(n17415), .A2(n17553), .ZN(n17397) );
  AOI22_X1 U20646 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17424), .B1(n17492), .B2(
        n17393), .ZN(n17396) );
  NAND2_X1 U20647 ( .A1(n17408), .A2(n17415), .ZN(n17403) );
  NAND2_X1 U20648 ( .A1(n17486), .A2(n17403), .ZN(n17400) );
  OAI21_X1 U20649 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17484), .A(n17400), .ZN(
        n17394) );
  AOI22_X1 U20650 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17425), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17394), .ZN(n17395) );
  OAI211_X1 U20651 ( .C1(n17398), .C2(n17397), .A(n17396), .B(n17395), .ZN(
        P3_U2713) );
  AOI22_X1 U20652 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17424), .B1(n17492), .B2(
        n17399), .ZN(n17402) );
  INV_X1 U20653 ( .A(n17400), .ZN(n17405) );
  AOI22_X1 U20654 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17425), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n17405), .ZN(n17401) );
  OAI211_X1 U20655 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n17403), .A(n17402), .B(
        n17401), .ZN(P3_U2714) );
  NAND3_X1 U20656 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(n17415), .ZN(n17409) );
  AOI22_X1 U20657 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17424), .B1(n17492), .B2(
        n17404), .ZN(n17407) );
  AOI22_X1 U20658 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17425), .B1(
        P3_EAX_REG_20__SCAN_IN), .B2(n17405), .ZN(n17406) );
  OAI211_X1 U20659 ( .C1(n17408), .C2(n17409), .A(n17407), .B(n17406), .ZN(
        P3_U2715) );
  AOI22_X1 U20660 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17425), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17424), .ZN(n17411) );
  INV_X1 U20661 ( .A(n17415), .ZN(n17419) );
  NOR2_X1 U20662 ( .A1(n20860), .A2(n17419), .ZN(n17413) );
  OAI211_X1 U20663 ( .C1(n17413), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17486), .B(
        n17409), .ZN(n17410) );
  OAI211_X1 U20664 ( .C1(n17412), .C2(n17487), .A(n17411), .B(n17410), .ZN(
        P3_U2716) );
  AOI22_X1 U20665 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17425), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17424), .ZN(n17417) );
  INV_X1 U20666 ( .A(n17413), .ZN(n17414) );
  OAI211_X1 U20667 ( .C1(n17415), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17486), .B(
        n17414), .ZN(n17416) );
  OAI211_X1 U20668 ( .C1(n17418), .C2(n17487), .A(n17417), .B(n17416), .ZN(
        P3_U2717) );
  AOI22_X1 U20669 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17425), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17424), .ZN(n17422) );
  INV_X1 U20670 ( .A(n17426), .ZN(n17420) );
  OAI211_X1 U20671 ( .C1(n17420), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17486), .B(
        n17419), .ZN(n17421) );
  OAI211_X1 U20672 ( .C1(n17423), .C2(n17487), .A(n17422), .B(n17421), .ZN(
        P3_U2718) );
  AOI22_X1 U20673 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17425), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17424), .ZN(n17429) );
  OAI211_X1 U20674 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17427), .A(n17486), .B(
        n17426), .ZN(n17428) );
  OAI211_X1 U20675 ( .C1(n17430), .C2(n17487), .A(n17429), .B(n17428), .ZN(
        P3_U2719) );
  OR2_X1 U20676 ( .A1(n17431), .A2(n17432), .ZN(n17435) );
  NAND2_X1 U20677 ( .A1(n17486), .A2(n17432), .ZN(n17439) );
  AOI22_X1 U20678 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17493), .B1(n17492), .B2(
        n17433), .ZN(n17434) );
  OAI221_X1 U20679 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n17435), .C1(n17604), 
        .C2(n17439), .A(n17434), .ZN(P3_U2720) );
  INV_X1 U20680 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n21116) );
  INV_X1 U20681 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17590) );
  INV_X1 U20682 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17586) );
  INV_X1 U20683 ( .A(n17484), .ZN(n17495) );
  NAND2_X1 U20684 ( .A1(n17436), .A2(n17495), .ZN(n17463) );
  NOR2_X1 U20685 ( .A1(n17586), .A2(n17463), .ZN(n17459) );
  NAND2_X1 U20686 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17459), .ZN(n17458) );
  NOR2_X1 U20687 ( .A1(n17590), .A2(n17458), .ZN(n17454) );
  NAND2_X1 U20688 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17454), .ZN(n17445) );
  NOR2_X1 U20689 ( .A1(n21116), .A2(n17445), .ZN(n17448) );
  NAND2_X1 U20690 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17448), .ZN(n17440) );
  INV_X1 U20691 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17599) );
  AOI22_X1 U20692 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17493), .B1(n17492), .B2(
        n17437), .ZN(n17438) );
  OAI221_X1 U20693 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17440), .C1(n17599), 
        .C2(n17439), .A(n17438), .ZN(P3_U2721) );
  INV_X1 U20694 ( .A(n17440), .ZN(n17443) );
  AOI21_X1 U20695 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17486), .A(n17448), .ZN(
        n17442) );
  OAI222_X1 U20696 ( .A1(n17490), .A2(n17444), .B1(n17443), .B2(n17442), .C1(
        n17487), .C2(n17441), .ZN(P3_U2722) );
  INV_X1 U20697 ( .A(n17445), .ZN(n17452) );
  AOI21_X1 U20698 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17486), .A(n17452), .ZN(
        n17447) );
  OAI222_X1 U20699 ( .A1(n17490), .A2(n17449), .B1(n17448), .B2(n17447), .C1(
        n17487), .C2(n17446), .ZN(P3_U2723) );
  AOI21_X1 U20700 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17486), .A(n17454), .ZN(
        n17451) );
  OAI222_X1 U20701 ( .A1(n17490), .A2(n17453), .B1(n17452), .B2(n17451), .C1(
        n17487), .C2(n17450), .ZN(P3_U2724) );
  AOI21_X1 U20702 ( .B1(n17590), .B2(n17458), .A(n17454), .ZN(n17455) );
  AOI22_X1 U20703 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17493), .B1(n17455), .B2(
        n17486), .ZN(n17456) );
  OAI21_X1 U20704 ( .B1(n17457), .B2(n17487), .A(n17456), .ZN(P3_U2725) );
  INV_X1 U20705 ( .A(n17458), .ZN(n17462) );
  AOI21_X1 U20706 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17486), .A(n17459), .ZN(
        n17461) );
  OAI222_X1 U20707 ( .A1(n17490), .A2(n21044), .B1(n17462), .B2(n17461), .C1(
        n17487), .C2(n17460), .ZN(P3_U2726) );
  INV_X1 U20708 ( .A(n17463), .ZN(n17470) );
  AOI22_X1 U20709 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17493), .B1(n17470), .B2(
        n17586), .ZN(n17466) );
  NAND3_X1 U20710 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17486), .A3(n17464), .ZN(
        n17465) );
  OAI211_X1 U20711 ( .C1(n17467), .C2(n17487), .A(n17466), .B(n17465), .ZN(
        P3_U2727) );
  INV_X1 U20712 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17582) );
  INV_X1 U20713 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17574) );
  NOR3_X1 U20714 ( .A1(n17494), .A2(n17574), .A3(n17484), .ZN(n17489) );
  NAND2_X1 U20715 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17489), .ZN(n17478) );
  NOR2_X1 U20716 ( .A1(n17578), .A2(n17478), .ZN(n17481) );
  NAND2_X1 U20717 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17481), .ZN(n17471) );
  NOR2_X1 U20718 ( .A1(n17582), .A2(n17471), .ZN(n17474) );
  AOI21_X1 U20719 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17486), .A(n17474), .ZN(
        n17469) );
  OAI222_X1 U20720 ( .A1(n17490), .A2(n18345), .B1(n17470), .B2(n17469), .C1(
        n17487), .C2(n17468), .ZN(P3_U2728) );
  INV_X1 U20721 ( .A(n17471), .ZN(n17477) );
  AOI21_X1 U20722 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17486), .A(n17477), .ZN(
        n17473) );
  OAI222_X1 U20723 ( .A1(n18338), .A2(n17490), .B1(n17474), .B2(n17473), .C1(
        n17487), .C2(n17472), .ZN(P3_U2729) );
  AOI21_X1 U20724 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17486), .A(n17481), .ZN(
        n17476) );
  OAI222_X1 U20725 ( .A1(n18333), .A2(n17490), .B1(n17477), .B2(n17476), .C1(
        n17487), .C2(n17475), .ZN(P3_U2730) );
  INV_X1 U20726 ( .A(n17478), .ZN(n17483) );
  AOI21_X1 U20727 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17486), .A(n17483), .ZN(
        n17480) );
  OAI222_X1 U20728 ( .A1(n18327), .A2(n17490), .B1(n17481), .B2(n17480), .C1(
        n17487), .C2(n17479), .ZN(P3_U2731) );
  AOI21_X1 U20729 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17486), .A(n17489), .ZN(
        n17482) );
  OAI222_X1 U20730 ( .A1(n18322), .A2(n17490), .B1(n17483), .B2(n17482), .C1(
        n17487), .C2(n12762), .ZN(P3_U2732) );
  NOR2_X1 U20731 ( .A1(n17494), .A2(n17484), .ZN(n17485) );
  AOI21_X1 U20732 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17486), .A(n17485), .ZN(
        n17488) );
  OAI222_X1 U20733 ( .A1(n18317), .A2(n17490), .B1(n17489), .B2(n17488), .C1(
        n17487), .C2(n12919), .ZN(P3_U2733) );
  INV_X1 U20734 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n21082) );
  AOI22_X1 U20735 ( .A1(n17493), .A2(BUF2_REG_1__SCAN_IN), .B1(n17492), .B2(
        n17491), .ZN(n17497) );
  OAI211_X1 U20736 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(P3_EAX_REG_0__SCAN_IN), 
        .A(n17495), .B(n17494), .ZN(n17496) );
  OAI211_X1 U20737 ( .C1(n17498), .C2(n21082), .A(n17497), .B(n17496), .ZN(
        P3_U2734) );
  INV_X1 U20738 ( .A(n17797), .ZN(n17962) );
  NOR2_X1 U20739 ( .A1(n18926), .A2(n17962), .ZN(n18954) );
  INV_X1 U20740 ( .A(n17538), .ZN(n17539) );
  AND2_X1 U20741 ( .A1(n17514), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20742 ( .A1(n17501), .A2(n17500), .ZN(n17518) );
  AOI22_X1 U20743 ( .A1(n18954), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17502) );
  OAI21_X1 U20744 ( .B1(n17569), .B2(n17518), .A(n17502), .ZN(P3_U2737) );
  INV_X1 U20745 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17567) );
  AOI22_X1 U20746 ( .A1(n18954), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17514), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17503) );
  OAI21_X1 U20747 ( .B1(n17567), .B2(n17518), .A(n17503), .ZN(P3_U2738) );
  AOI22_X1 U20748 ( .A1(n18954), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17514), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17504) );
  OAI21_X1 U20749 ( .B1(n17565), .B2(n17518), .A(n17504), .ZN(P3_U2739) );
  INV_X1 U20750 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17563) );
  AOI22_X1 U20751 ( .A1(n18954), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17505) );
  OAI21_X1 U20752 ( .B1(n17563), .B2(n17518), .A(n17505), .ZN(P3_U2740) );
  INV_X1 U20753 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17561) );
  AOI22_X1 U20754 ( .A1(n18954), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17514), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17506) );
  OAI21_X1 U20755 ( .B1(n17561), .B2(n17518), .A(n17506), .ZN(P3_U2741) );
  AOI22_X1 U20756 ( .A1(n18954), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17514), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17507) );
  OAI21_X1 U20757 ( .B1(n17559), .B2(n17518), .A(n17507), .ZN(P3_U2742) );
  INV_X1 U20758 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17557) );
  AOI22_X1 U20759 ( .A1(n18954), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17514), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17508) );
  OAI21_X1 U20760 ( .B1(n17557), .B2(n17518), .A(n17508), .ZN(P3_U2743) );
  INV_X1 U20761 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17555) );
  AOI22_X1 U20762 ( .A1(n17535), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(
        P3_DATAO_REG_23__SCAN_IN), .B2(n17534), .ZN(n17509) );
  OAI21_X1 U20763 ( .B1(n17555), .B2(n17518), .A(n17509), .ZN(P3_U2744) );
  AOI22_X1 U20764 ( .A1(n17535), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17514), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17510) );
  OAI21_X1 U20765 ( .B1(n17553), .B2(n17518), .A(n17510), .ZN(P3_U2745) );
  INV_X1 U20766 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17551) );
  AOI22_X1 U20767 ( .A1(n17535), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17514), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17511) );
  OAI21_X1 U20768 ( .B1(n17551), .B2(n17518), .A(n17511), .ZN(P3_U2746) );
  AOI22_X1 U20769 ( .A1(n17535), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17514), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17512) );
  OAI21_X1 U20770 ( .B1(n17549), .B2(n17518), .A(n17512), .ZN(P3_U2747) );
  AOI22_X1 U20771 ( .A1(n17535), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17514), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17513) );
  OAI21_X1 U20772 ( .B1(n17547), .B2(n17518), .A(n17513), .ZN(P3_U2748) );
  AOI22_X1 U20773 ( .A1(n17535), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17514), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17515) );
  OAI21_X1 U20774 ( .B1(n20860), .B2(n17518), .A(n17515), .ZN(P3_U2749) );
  AOI22_X1 U20775 ( .A1(n17535), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17516) );
  OAI21_X1 U20776 ( .B1(n17544), .B2(n17518), .A(n17516), .ZN(P3_U2750) );
  INV_X1 U20777 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17542) );
  AOI22_X1 U20778 ( .A1(n17535), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17517) );
  OAI21_X1 U20779 ( .B1(n17542), .B2(n17518), .A(n17517), .ZN(P3_U2751) );
  AOI22_X1 U20780 ( .A1(n17535), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17519) );
  OAI21_X1 U20781 ( .B1(n17604), .B2(n17537), .A(n17519), .ZN(P3_U2752) );
  AOI22_X1 U20782 ( .A1(n17535), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17520) );
  OAI21_X1 U20783 ( .B1(n17599), .B2(n17537), .A(n17520), .ZN(P3_U2753) );
  INV_X1 U20784 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17596) );
  AOI22_X1 U20785 ( .A1(n17535), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17521) );
  OAI21_X1 U20786 ( .B1(n17596), .B2(n17537), .A(n17521), .ZN(P3_U2754) );
  AOI22_X1 U20787 ( .A1(n17535), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17522) );
  OAI21_X1 U20788 ( .B1(n21116), .B2(n17537), .A(n17522), .ZN(P3_U2755) );
  INV_X1 U20789 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17592) );
  AOI22_X1 U20790 ( .A1(n17535), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17523) );
  OAI21_X1 U20791 ( .B1(n17592), .B2(n17537), .A(n17523), .ZN(P3_U2756) );
  AOI22_X1 U20792 ( .A1(n17535), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17524) );
  OAI21_X1 U20793 ( .B1(n17590), .B2(n17537), .A(n17524), .ZN(P3_U2757) );
  INV_X1 U20794 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17588) );
  AOI22_X1 U20795 ( .A1(n17535), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17525) );
  OAI21_X1 U20796 ( .B1(n17588), .B2(n17537), .A(n17525), .ZN(P3_U2758) );
  AOI22_X1 U20797 ( .A1(n17535), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17526) );
  OAI21_X1 U20798 ( .B1(n17586), .B2(n17537), .A(n17526), .ZN(P3_U2759) );
  INV_X1 U20799 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17584) );
  AOI22_X1 U20800 ( .A1(n17535), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(
        P3_DATAO_REG_7__SCAN_IN), .B2(n17534), .ZN(n17527) );
  OAI21_X1 U20801 ( .B1(n17584), .B2(n17537), .A(n17527), .ZN(P3_U2760) );
  AOI22_X1 U20802 ( .A1(n17535), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17528) );
  OAI21_X1 U20803 ( .B1(n17582), .B2(n17537), .A(n17528), .ZN(P3_U2761) );
  AOI22_X1 U20804 ( .A1(n17535), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17529) );
  OAI21_X1 U20805 ( .B1(n17580), .B2(n17537), .A(n17529), .ZN(P3_U2762) );
  AOI22_X1 U20806 ( .A1(n17535), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17530) );
  OAI21_X1 U20807 ( .B1(n17578), .B2(n17537), .A(n17530), .ZN(P3_U2763) );
  INV_X1 U20808 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17576) );
  AOI22_X1 U20809 ( .A1(n17535), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17531) );
  OAI21_X1 U20810 ( .B1(n17576), .B2(n17537), .A(n17531), .ZN(P3_U2764) );
  AOI22_X1 U20811 ( .A1(n17535), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17532) );
  OAI21_X1 U20812 ( .B1(n17574), .B2(n17537), .A(n17532), .ZN(P3_U2765) );
  AOI22_X1 U20813 ( .A1(n17535), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17533) );
  OAI21_X1 U20814 ( .B1(n21082), .B2(n17537), .A(n17533), .ZN(P3_U2766) );
  AOI22_X1 U20815 ( .A1(n17535), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17534), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17536) );
  OAI21_X1 U20816 ( .B1(n17571), .B2(n17537), .A(n17536), .ZN(P3_U2767) );
  NAND2_X1 U20817 ( .A1(n18313), .A2(n17540), .ZN(n18809) );
  OAI211_X1 U20818 ( .C1(n18313), .C2(n18953), .A(n17540), .B(n17539), .ZN(
        n17597) );
  AOI22_X1 U20819 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17601), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17600), .ZN(n17541) );
  OAI21_X1 U20820 ( .B1(n17542), .B2(n17603), .A(n17541), .ZN(P3_U2768) );
  AOI22_X1 U20821 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17601), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17600), .ZN(n17543) );
  OAI21_X1 U20822 ( .B1(n17544), .B2(n17603), .A(n17543), .ZN(P3_U2769) );
  AOI22_X1 U20823 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17601), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17600), .ZN(n17545) );
  OAI21_X1 U20824 ( .B1(n20860), .B2(n17603), .A(n17545), .ZN(P3_U2770) );
  AOI22_X1 U20825 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17593), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17600), .ZN(n17546) );
  OAI21_X1 U20826 ( .B1(n17547), .B2(n17603), .A(n17546), .ZN(P3_U2771) );
  AOI22_X1 U20827 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17593), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17600), .ZN(n17548) );
  OAI21_X1 U20828 ( .B1(n17549), .B2(n17603), .A(n17548), .ZN(P3_U2772) );
  AOI22_X1 U20829 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17593), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17600), .ZN(n17550) );
  OAI21_X1 U20830 ( .B1(n17551), .B2(n17603), .A(n17550), .ZN(P3_U2773) );
  AOI22_X1 U20831 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17593), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17600), .ZN(n17552) );
  OAI21_X1 U20832 ( .B1(n17553), .B2(n17603), .A(n17552), .ZN(P3_U2774) );
  AOI22_X1 U20833 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17593), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17600), .ZN(n17554) );
  OAI21_X1 U20834 ( .B1(n17555), .B2(n17603), .A(n17554), .ZN(P3_U2775) );
  AOI22_X1 U20835 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17593), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17600), .ZN(n17556) );
  OAI21_X1 U20836 ( .B1(n17557), .B2(n17603), .A(n17556), .ZN(P3_U2776) );
  AOI22_X1 U20837 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17593), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17600), .ZN(n17558) );
  OAI21_X1 U20838 ( .B1(n17559), .B2(n17603), .A(n17558), .ZN(P3_U2777) );
  AOI22_X1 U20839 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17593), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17600), .ZN(n17560) );
  OAI21_X1 U20840 ( .B1(n17561), .B2(n17603), .A(n17560), .ZN(P3_U2778) );
  AOI22_X1 U20841 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17593), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17600), .ZN(n17562) );
  OAI21_X1 U20842 ( .B1(n17563), .B2(n17603), .A(n17562), .ZN(P3_U2779) );
  AOI22_X1 U20843 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17601), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17600), .ZN(n17564) );
  OAI21_X1 U20844 ( .B1(n17565), .B2(n17603), .A(n17564), .ZN(P3_U2780) );
  AOI22_X1 U20845 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17601), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17600), .ZN(n17566) );
  OAI21_X1 U20846 ( .B1(n17567), .B2(n17603), .A(n17566), .ZN(P3_U2781) );
  AOI22_X1 U20847 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17601), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17600), .ZN(n17568) );
  OAI21_X1 U20848 ( .B1(n17569), .B2(n17603), .A(n17568), .ZN(P3_U2782) );
  AOI22_X1 U20849 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17601), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17600), .ZN(n17570) );
  OAI21_X1 U20850 ( .B1(n17571), .B2(n17603), .A(n17570), .ZN(P3_U2783) );
  AOI22_X1 U20851 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17601), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17600), .ZN(n17572) );
  OAI21_X1 U20852 ( .B1(n21082), .B2(n17603), .A(n17572), .ZN(P3_U2784) );
  AOI22_X1 U20853 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17601), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17600), .ZN(n17573) );
  OAI21_X1 U20854 ( .B1(n17574), .B2(n17603), .A(n17573), .ZN(P3_U2785) );
  AOI22_X1 U20855 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17601), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17597), .ZN(n17575) );
  OAI21_X1 U20856 ( .B1(n17576), .B2(n17603), .A(n17575), .ZN(P3_U2786) );
  AOI22_X1 U20857 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17601), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17597), .ZN(n17577) );
  OAI21_X1 U20858 ( .B1(n17578), .B2(n17603), .A(n17577), .ZN(P3_U2787) );
  AOI22_X1 U20859 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17601), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17597), .ZN(n17579) );
  OAI21_X1 U20860 ( .B1(n17580), .B2(n17603), .A(n17579), .ZN(P3_U2788) );
  AOI22_X1 U20861 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17601), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17597), .ZN(n17581) );
  OAI21_X1 U20862 ( .B1(n17582), .B2(n17603), .A(n17581), .ZN(P3_U2789) );
  AOI22_X1 U20863 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17601), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17597), .ZN(n17583) );
  OAI21_X1 U20864 ( .B1(n17584), .B2(n17603), .A(n17583), .ZN(P3_U2790) );
  AOI22_X1 U20865 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17601), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17597), .ZN(n17585) );
  OAI21_X1 U20866 ( .B1(n17586), .B2(n17603), .A(n17585), .ZN(P3_U2791) );
  AOI22_X1 U20867 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17601), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17597), .ZN(n17587) );
  OAI21_X1 U20868 ( .B1(n17588), .B2(n17603), .A(n17587), .ZN(P3_U2792) );
  AOI22_X1 U20869 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17593), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17600), .ZN(n17589) );
  OAI21_X1 U20870 ( .B1(n17590), .B2(n17603), .A(n17589), .ZN(P3_U2793) );
  AOI22_X1 U20871 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17601), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17597), .ZN(n17591) );
  OAI21_X1 U20872 ( .B1(n17592), .B2(n17603), .A(n17591), .ZN(P3_U2794) );
  AOI22_X1 U20873 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17593), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17600), .ZN(n17594) );
  OAI21_X1 U20874 ( .B1(n21116), .B2(n17603), .A(n17594), .ZN(P3_U2795) );
  AOI22_X1 U20875 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17601), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17597), .ZN(n17595) );
  OAI21_X1 U20876 ( .B1(n17596), .B2(n17603), .A(n17595), .ZN(P3_U2796) );
  AOI22_X1 U20877 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17601), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17597), .ZN(n17598) );
  OAI21_X1 U20878 ( .B1(n17599), .B2(n17603), .A(n17598), .ZN(P3_U2797) );
  AOI22_X1 U20879 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17601), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17600), .ZN(n17602) );
  OAI21_X1 U20880 ( .B1(n17604), .B2(n17603), .A(n17602), .ZN(P3_U2798) );
  NAND2_X1 U20881 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17606), .ZN(
        n17623) );
  NOR2_X1 U20882 ( .A1(n17801), .A2(n17953), .ZN(n17714) );
  INV_X1 U20883 ( .A(n17605), .ZN(n17968) );
  OAI22_X1 U20884 ( .A1(n17968), .A2(n17876), .B1(n17967), .B2(n17966), .ZN(
        n17643) );
  NOR2_X1 U20885 ( .A1(n21067), .A2(n17643), .ZN(n17628) );
  NOR3_X1 U20886 ( .A1(n17714), .A2(n17628), .A3(n17606), .ZN(n17617) );
  INV_X1 U20887 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17607) );
  NAND3_X1 U20888 ( .A1(n17608), .A2(n17774), .A3(n17607), .ZN(n17614) );
  INV_X1 U20889 ( .A(n17774), .ZN(n17809) );
  NOR3_X1 U20890 ( .A1(n17809), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        n17609), .ZN(n17631) );
  OAI21_X1 U20891 ( .B1(n17610), .B2(n17922), .A(n17961), .ZN(n17611) );
  AOI21_X1 U20892 ( .B1(n17797), .B2(n17612), .A(n17611), .ZN(n17637) );
  OAI21_X1 U20893 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17749), .A(
        n17637), .ZN(n17632) );
  OAI21_X1 U20894 ( .B1(n17631), .B2(n17632), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17613) );
  OAI211_X1 U20895 ( .C1(n17823), .C2(n17615), .A(n17614), .B(n17613), .ZN(
        n17616) );
  AOI211_X1 U20896 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n18285), .A(n17617), 
        .B(n17616), .ZN(n17622) );
  OAI211_X1 U20897 ( .C1(n17620), .C2(n17619), .A(n17873), .B(n17618), .ZN(
        n17621) );
  OAI211_X1 U20898 ( .C1(n17623), .C2(n17629), .A(n17622), .B(n17621), .ZN(
        P3_U2802) );
  NOR2_X1 U20899 ( .A1(n17625), .A2(n17624), .ZN(n17626) );
  XNOR2_X1 U20900 ( .A(n17626), .B(n17802), .ZN(n17982) );
  AOI22_X1 U20901 ( .A1(n18245), .A2(P3_REIP_REG_27__SCAN_IN), .B1(n17800), 
        .B2(n17627), .ZN(n17634) );
  AOI21_X1 U20902 ( .B1(n21067), .B2(n17629), .A(n17628), .ZN(n17630) );
  AOI211_X1 U20903 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17632), .A(
        n17631), .B(n17630), .ZN(n17633) );
  OAI211_X1 U20904 ( .C1(n17982), .C2(n17837), .A(n17634), .B(n17633), .ZN(
        P3_U2803) );
  AOI21_X1 U20905 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17636), .A(
        n17635), .ZN(n17991) );
  AOI221_X1 U20906 ( .B1(n18349), .B2(n17639), .C1(n17638), .C2(n17639), .A(
        n17637), .ZN(n17642) );
  INV_X1 U20907 ( .A(n17749), .ZN(n17689) );
  NAND2_X1 U20908 ( .A1(n18245), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17989) );
  OAI221_X1 U20909 ( .B1(n17640), .B2(n17823), .C1(n17640), .C2(n17749), .A(
        n17989), .ZN(n17641) );
  AOI211_X1 U20910 ( .C1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n17643), .A(
        n17642), .B(n17641), .ZN(n17645) );
  NOR2_X1 U20911 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17994), .ZN(
        n17988) );
  NAND3_X1 U20912 ( .A1(n17682), .A2(n17755), .A3(n17988), .ZN(n17644) );
  OAI211_X1 U20913 ( .C1(n17991), .C2(n17837), .A(n17645), .B(n17644), .ZN(
        P3_U2804) );
  INV_X1 U20914 ( .A(n18105), .ZN(n18027) );
  NOR2_X1 U20915 ( .A1(n18027), .A2(n17997), .ZN(n18009) );
  NAND2_X1 U20916 ( .A1(n18009), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17646) );
  XNOR2_X1 U20917 ( .A(n17646), .B(n17995), .ZN(n18006) );
  OR2_X1 U20918 ( .A1(n18349), .A2(n9859), .ZN(n17674) );
  OAI211_X1 U20919 ( .C1(n17647), .C2(n17962), .A(n17961), .B(n17674), .ZN(
        n17661) );
  NOR2_X1 U20920 ( .A1(n16866), .A2(n18885), .ZN(n17999) );
  NOR2_X1 U20921 ( .A1(n10046), .A2(n10047), .ZN(n17650) );
  OAI211_X1 U20922 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n9859), .B(n17774), .ZN(n17649)
         );
  OAI22_X1 U20923 ( .A1(n17650), .A2(n17649), .B1(n17648), .B2(n17823), .ZN(
        n17651) );
  AOI211_X1 U20924 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17661), .A(
        n17999), .B(n17651), .ZN(n17657) );
  NOR3_X1 U20925 ( .A1(n17997), .A2(n18028), .A3(n18014), .ZN(n17652) );
  XNOR2_X1 U20926 ( .A(n17995), .B(n17652), .ZN(n18003) );
  OAI21_X1 U20927 ( .B1(n17802), .B2(n17654), .A(n17653), .ZN(n17655) );
  XNOR2_X1 U20928 ( .A(n17655), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18002) );
  AOI22_X1 U20929 ( .A1(n17953), .A2(n18003), .B1(n17873), .B2(n18002), .ZN(
        n17656) );
  OAI211_X1 U20930 ( .C1(n17876), .C2(n18006), .A(n17657), .B(n17656), .ZN(
        P3_U2805) );
  OAI21_X1 U20931 ( .B1(n18014), .B2(n17659), .A(n17658), .ZN(n17660) );
  INV_X1 U20932 ( .A(n17660), .ZN(n18021) );
  NAND2_X1 U20933 ( .A1(n9859), .A2(n17774), .ZN(n17662) );
  INV_X1 U20934 ( .A(n17661), .ZN(n17670) );
  NAND2_X1 U20935 ( .A1(n18245), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18019) );
  OAI221_X1 U20936 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17662), .C1(
        n10046), .C2(n17670), .A(n18019), .ZN(n17663) );
  AOI21_X1 U20937 ( .B1(n17800), .B2(n17664), .A(n17663), .ZN(n17666) );
  NOR2_X1 U20938 ( .A1(n18028), .A2(n17997), .ZN(n18008) );
  OAI22_X1 U20939 ( .A1(n18009), .A2(n17876), .B1(n18008), .B2(n17966), .ZN(
        n17680) );
  NOR2_X1 U20940 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17997), .ZN(
        n18017) );
  AOI22_X1 U20941 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17680), .B1(
        n17755), .B2(n18017), .ZN(n17665) );
  OAI211_X1 U20942 ( .C1(n18021), .C2(n17837), .A(n17666), .B(n17665), .ZN(
        P3_U2806) );
  OAI22_X1 U20943 ( .A1(n17667), .A2(n17695), .B1(n17872), .B2(n18043), .ZN(
        n17668) );
  NOR2_X1 U20944 ( .A1(n17668), .A2(n17712), .ZN(n17669) );
  XNOR2_X1 U20945 ( .A(n17669), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18026) );
  AOI211_X1 U20946 ( .C1(n17749), .C2(n17672), .A(n17671), .B(n17670), .ZN(
        n17676) );
  NAND2_X1 U20947 ( .A1(n18245), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18025) );
  OAI21_X1 U20948 ( .B1(n17674), .B2(n17673), .A(n18025), .ZN(n17675) );
  AOI211_X1 U20949 ( .C1(n17677), .C2(n17800), .A(n17676), .B(n17675), .ZN(
        n17684) );
  OR2_X1 U20950 ( .A1(n17876), .A2(n18009), .ZN(n17679) );
  OR2_X1 U20951 ( .A1(n17966), .A2(n18008), .ZN(n17678) );
  OAI22_X1 U20952 ( .A1(n18027), .A2(n17679), .B1(n18028), .B2(n17678), .ZN(
        n17681) );
  AOI22_X1 U20953 ( .A1(n17682), .A2(n17681), .B1(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17680), .ZN(n17683) );
  OAI211_X1 U20954 ( .C1(n17837), .C2(n18026), .A(n17684), .B(n17683), .ZN(
        P3_U2807) );
  NAND2_X1 U20955 ( .A1(n17687), .A2(n17774), .ZN(n17706) );
  AOI221_X1 U20956 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n17705), .C2(n17690), .A(
        n17706), .ZN(n17692) );
  NAND2_X1 U20957 ( .A1(n17797), .A2(n17685), .ZN(n17686) );
  OAI211_X1 U20958 ( .C1(n17687), .C2(n17922), .A(n17961), .B(n17686), .ZN(
        n17716) );
  AOI21_X1 U20959 ( .B1(n17689), .B2(n17688), .A(n17716), .ZN(n17704) );
  NAND2_X1 U20960 ( .A1(n18245), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18041) );
  OAI21_X1 U20961 ( .B1(n17704), .B2(n17690), .A(n18041), .ZN(n17691) );
  AOI211_X1 U20962 ( .C1(n17693), .C2(n17800), .A(n17692), .B(n17691), .ZN(
        n17699) );
  AOI22_X1 U20963 ( .A1(n17801), .A2(n18027), .B1(n17953), .B2(n18028), .ZN(
        n17768) );
  OAI21_X1 U20964 ( .B1(n18034), .B2(n17714), .A(n17768), .ZN(n17709) );
  OAI221_X1 U20965 ( .B1(n17695), .B2(n17694), .C1(n17695), .C2(n18034), .A(
        n12788), .ZN(n17696) );
  XNOR2_X1 U20966 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17696), .ZN(
        n18039) );
  AOI22_X1 U20967 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17709), .B1(
        n17873), .B2(n18039), .ZN(n17698) );
  NAND3_X1 U20968 ( .A1(n17755), .A2(n18034), .A3(n18043), .ZN(n17697) );
  NAND3_X1 U20969 ( .A1(n17699), .A2(n17698), .A3(n17697), .ZN(P3_U2808) );
  NAND3_X1 U20970 ( .A1(n17872), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17700), .ZN(n17730) );
  INV_X1 U20971 ( .A(n17701), .ZN(n17737) );
  OAI22_X1 U20972 ( .A1(n18049), .A2(n17730), .B1(n17737), .B2(n17702), .ZN(
        n17703) );
  XNOR2_X1 U20973 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17703), .ZN(
        n18056) );
  NAND2_X1 U20974 ( .A1(n18245), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18054) );
  OAI221_X1 U20975 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17706), .C1(
        n17705), .C2(n17704), .A(n18054), .ZN(n17707) );
  AOI21_X1 U20976 ( .B1(n17800), .B2(n17708), .A(n17707), .ZN(n17711) );
  NOR2_X1 U20977 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18049), .ZN(
        n18053) );
  AOI22_X1 U20978 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17709), .B1(
        n18053), .B2(n17732), .ZN(n17710) );
  OAI211_X1 U20979 ( .C1(n18056), .C2(n17837), .A(n17711), .B(n17710), .ZN(
        P3_U2809) );
  INV_X1 U20980 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21131) );
  AOI221_X1 U20981 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17730), 
        .C1(n21131), .C2(n17736), .A(n17712), .ZN(n17713) );
  XNOR2_X1 U20982 ( .A(n17713), .B(n20926), .ZN(n18057) );
  NOR2_X1 U20983 ( .A1(n18029), .A2(n21131), .ZN(n18058) );
  OAI21_X1 U20984 ( .B1(n17714), .B2(n18058), .A(n17768), .ZN(n17715) );
  INV_X1 U20985 ( .A(n17715), .ZN(n17735) );
  NAND2_X1 U20986 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n20926), .ZN(
        n18063) );
  NAND2_X1 U20987 ( .A1(n18285), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17721) );
  OAI221_X1 U20988 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17717), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n18692), .A(n17716), .ZN(
        n17720) );
  OAI21_X1 U20989 ( .B1(n17800), .B2(n17689), .A(n17718), .ZN(n17719) );
  NAND4_X1 U20990 ( .A1(n17722), .A2(n17721), .A3(n17720), .A4(n17719), .ZN(
        P3_U2810) );
  INV_X1 U20991 ( .A(n17961), .ZN(n17933) );
  INV_X1 U20992 ( .A(n17723), .ZN(n17725) );
  OAI21_X1 U20993 ( .B1(n17933), .B2(n17725), .A(n17956), .ZN(n17750) );
  OAI21_X1 U20994 ( .B1(n17724), .B2(n17962), .A(n17750), .ZN(n17741) );
  NOR2_X1 U20995 ( .A1(n17809), .A2(n17725), .ZN(n17743) );
  NAND2_X1 U20996 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17726) );
  OAI211_X1 U20997 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17743), .B(n17726), .ZN(n17727) );
  NAND2_X1 U20998 ( .A1(n18285), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18066) );
  OAI211_X1 U20999 ( .C1(n17823), .C2(n17728), .A(n17727), .B(n18066), .ZN(
        n17729) );
  AOI21_X1 U21000 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17741), .A(
        n17729), .ZN(n17734) );
  OAI21_X1 U21001 ( .B1(n17737), .B2(n17736), .A(n17730), .ZN(n17731) );
  XNOR2_X1 U21002 ( .A(n17731), .B(n21131), .ZN(n18064) );
  AOI22_X1 U21003 ( .A1(n17873), .A2(n18064), .B1(n17732), .B2(n21131), .ZN(
        n17733) );
  OAI211_X1 U21004 ( .C1(n17735), .C2(n21131), .A(n17734), .B(n17733), .ZN(
        P3_U2811) );
  OAI21_X1 U21005 ( .B1(n21092), .B2(n17802), .A(n17736), .ZN(n17738) );
  XNOR2_X1 U21006 ( .A(n17738), .B(n17737), .ZN(n18083) );
  NAND2_X1 U21007 ( .A1(n18245), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18081) );
  OAI21_X1 U21008 ( .B1(n17823), .B2(n17739), .A(n18081), .ZN(n17740) );
  AOI221_X1 U21009 ( .B1(n17743), .B2(n17742), .C1(n17741), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17740), .ZN(n17746) );
  OAI21_X1 U21010 ( .B1(n18072), .B2(n17769), .A(n17768), .ZN(n17756) );
  NOR2_X1 U21011 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17744), .ZN(
        n18079) );
  AOI22_X1 U21012 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17756), .B1(
        n17755), .B2(n18079), .ZN(n17745) );
  OAI211_X1 U21013 ( .C1(n17837), .C2(n18083), .A(n17746), .B(n17745), .ZN(
        P3_U2812) );
  AOI21_X1 U21014 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17748), .A(
        n17747), .ZN(n18090) );
  NOR2_X1 U21015 ( .A1(n16866), .A2(n21129), .ZN(n18086) );
  AOI221_X1 U21016 ( .B1(n18340), .B2(n17752), .C1(n17751), .C2(n17752), .A(
        n17750), .ZN(n17753) );
  AOI211_X1 U21017 ( .C1(n17754), .C2(n17955), .A(n18086), .B(n17753), .ZN(
        n17758) );
  NOR2_X1 U21018 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18097), .ZN(
        n18088) );
  AOI22_X1 U21019 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17756), .B1(
        n17755), .B2(n18088), .ZN(n17757) );
  OAI211_X1 U21020 ( .C1(n18090), .C2(n17837), .A(n17758), .B(n17757), .ZN(
        P3_U2813) );
  OAI21_X1 U21021 ( .B1(n17802), .B2(n17694), .A(n17759), .ZN(n17760) );
  XNOR2_X1 U21022 ( .A(n17760), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n18099) );
  OAI21_X1 U21023 ( .B1(n17775), .B2(n17922), .A(n17961), .ZN(n17790) );
  AOI21_X1 U21024 ( .B1(n17797), .B2(n17761), .A(n17790), .ZN(n17776) );
  OAI22_X1 U21025 ( .A1(n17776), .A2(n17763), .B1(n17823), .B2(n17762), .ZN(
        n17766) );
  OAI211_X1 U21026 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17775), .B(n17774), .ZN(n17764) );
  OAI22_X1 U21027 ( .A1(n10217), .A2(n17764), .B1(n16866), .B2(n18868), .ZN(
        n17765) );
  AOI211_X1 U21028 ( .C1(n17873), .C2(n18099), .A(n17766), .B(n17765), .ZN(
        n17767) );
  OAI221_X1 U21029 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17769), 
        .C1(n18097), .C2(n17768), .A(n17767), .ZN(P3_U2814) );
  AND2_X1 U21030 ( .A1(n17770), .A2(n17802), .ZN(n17815) );
  AOI22_X1 U21031 ( .A1(n17803), .A2(n17771), .B1(n17815), .B2(n21139), .ZN(
        n17772) );
  AOI221_X1 U21032 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18148), 
        .C1(n17802), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17772), .ZN(
        n17773) );
  XNOR2_X1 U21033 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17773), .ZN(
        n18112) );
  AOI211_X1 U21034 ( .C1(n18106), .C2(n18118), .A(n18105), .B(n17876), .ZN(
        n17780) );
  NAND2_X1 U21035 ( .A1(n17775), .A2(n17774), .ZN(n17778) );
  NAND2_X1 U21036 ( .A1(n18245), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18116) );
  OAI221_X1 U21037 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17778), .C1(
        n17777), .C2(n17776), .A(n18116), .ZN(n17779) );
  AOI211_X1 U21038 ( .C1(n17800), .C2(n17781), .A(n17780), .B(n17779), .ZN(
        n17783) );
  OAI211_X1 U21039 ( .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18102), .A(
        n17953), .B(n18028), .ZN(n17782) );
  OAI211_X1 U21040 ( .C1(n18112), .C2(n17837), .A(n17783), .B(n17782), .ZN(
        P3_U2815) );
  NOR2_X1 U21041 ( .A1(n18148), .A2(n17784), .ZN(n18124) );
  OAI221_X1 U21042 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18163), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18124), .A(n18106), .ZN(
        n18133) );
  NOR2_X1 U21043 ( .A1(n18349), .A2(n17808), .ZN(n17831) );
  INV_X1 U21044 ( .A(n17831), .ZN(n17786) );
  OAI21_X1 U21045 ( .B1(n17810), .B2(n17786), .A(n17785), .ZN(n17789) );
  OAI22_X1 U21046 ( .A1(n17946), .A2(n17787), .B1(n16866), .B2(n21089), .ZN(
        n17788) );
  AOI21_X1 U21047 ( .B1(n17790), .B2(n17789), .A(n17788), .ZN(n17795) );
  INV_X1 U21048 ( .A(n18124), .ZN(n18121) );
  AOI221_X1 U21049 ( .B1(n18159), .B2(n20868), .C1(n18121), .C2(n20868), .A(
        n18102), .ZN(n18130) );
  NOR2_X1 U21050 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17792) );
  NAND2_X1 U21051 ( .A1(n17872), .A2(n17791), .ZN(n17850) );
  INV_X1 U21052 ( .A(n17850), .ZN(n17816) );
  AOI22_X1 U21053 ( .A1(n17792), .A2(n17815), .B1(n17816), .B2(n18124), .ZN(
        n17793) );
  XNOR2_X1 U21054 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17793), .ZN(
        n18129) );
  AOI22_X1 U21055 ( .A1(n17953), .A2(n18130), .B1(n17873), .B2(n18129), .ZN(
        n17794) );
  OAI211_X1 U21056 ( .C1(n17876), .C2(n18133), .A(n17795), .B(n17794), .ZN(
        P3_U2816) );
  AOI22_X1 U21057 ( .A1(n17797), .A2(n17796), .B1(n18297), .B2(n17808), .ZN(
        n17798) );
  NAND2_X1 U21058 ( .A1(n17798), .A2(n17961), .ZN(n17820) );
  AOI22_X1 U21059 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17820), .B1(
        n17800), .B2(n17799), .ZN(n17814) );
  INV_X1 U21060 ( .A(n18151), .ZN(n18168) );
  NOR2_X1 U21061 ( .A1(n18148), .A2(n18168), .ZN(n18123) );
  AND2_X1 U21062 ( .A1(n21139), .A2(n18123), .ZN(n18138) );
  NAND2_X1 U21063 ( .A1(n18163), .A2(n18123), .ZN(n18139) );
  NAND2_X1 U21064 ( .A1(n18123), .A2(n18134), .ZN(n18141) );
  AOI22_X1 U21065 ( .A1(n17801), .A2(n18139), .B1(n17953), .B2(n18141), .ZN(
        n17827) );
  AOI22_X1 U21066 ( .A1(n18123), .A2(n17803), .B1(n17802), .B2(n18148), .ZN(
        n17805) );
  NOR2_X1 U21067 ( .A1(n17805), .A2(n17804), .ZN(n17806) );
  XNOR2_X1 U21068 ( .A(n17806), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18147) );
  OAI22_X1 U21069 ( .A1(n17827), .A2(n21139), .B1(n17837), .B2(n18147), .ZN(
        n17807) );
  AOI21_X1 U21070 ( .B1(n18138), .B2(n17834), .A(n17807), .ZN(n17813) );
  NAND2_X1 U21071 ( .A1(n18245), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17812) );
  NOR2_X1 U21072 ( .A1(n17809), .A2(n17808), .ZN(n17819) );
  OAI211_X1 U21073 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17819), .B(n17810), .ZN(n17811) );
  NAND4_X1 U21074 ( .A1(n17814), .A2(n17813), .A3(n17812), .A4(n17811), .ZN(
        P3_U2817) );
  AOI21_X1 U21075 ( .B1(n18151), .B2(n17816), .A(n17815), .ZN(n17817) );
  XNOR2_X1 U21076 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n17817), .ZN(
        n18152) );
  NOR3_X1 U21077 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17862), .A3(
        n18168), .ZN(n17825) );
  AOI22_X1 U21078 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17820), .B1(
        n17819), .B2(n17818), .ZN(n17821) );
  NAND2_X1 U21079 ( .A1(n18245), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18153) );
  OAI211_X1 U21080 ( .C1(n17823), .C2(n17822), .A(n17821), .B(n18153), .ZN(
        n17824) );
  AOI211_X1 U21081 ( .C1(n17873), .C2(n18152), .A(n17825), .B(n17824), .ZN(
        n17826) );
  OAI21_X1 U21082 ( .B1(n17827), .B2(n18148), .A(n17826), .ZN(P3_U2818) );
  NAND2_X1 U21083 ( .A1(n12780), .A2(n12779), .ZN(n17846) );
  NAND2_X1 U21084 ( .A1(n17828), .A2(n18199), .ZN(n17851) );
  OAI22_X1 U21085 ( .A1(n18166), .A2(n17850), .B1(n17846), .B2(n17851), .ZN(
        n17829) );
  XNOR2_X1 U21086 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17829), .ZN(
        n18176) );
  NOR2_X1 U21087 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18166), .ZN(
        n18173) );
  INV_X1 U21088 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18860) );
  NOR2_X1 U21089 ( .A1(n16866), .A2(n18860), .ZN(n18171) );
  NAND4_X1 U21090 ( .A1(n18692), .A2(n17854), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17853) );
  NOR2_X1 U21091 ( .A1(n17841), .A2(n17853), .ZN(n17839) );
  AOI21_X1 U21092 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17956), .A(
        n17839), .ZN(n17832) );
  OAI22_X1 U21093 ( .A1(n17832), .A2(n17831), .B1(n17946), .B2(n17830), .ZN(
        n17833) );
  AOI211_X1 U21094 ( .C1(n18173), .C2(n17834), .A(n18171), .B(n17833), .ZN(
        n17836) );
  AND2_X1 U21095 ( .A1(n18166), .A2(n17834), .ZN(n17847) );
  OAI22_X1 U21096 ( .A1(n18163), .A2(n17876), .B1(n17966), .B2(n18134), .ZN(
        n17838) );
  OAI21_X1 U21097 ( .B1(n17847), .B2(n17838), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17835) );
  OAI211_X1 U21098 ( .C1(n18176), .C2(n17837), .A(n17836), .B(n17835), .ZN(
        P3_U2819) );
  INV_X1 U21099 ( .A(n17838), .ZN(n17861) );
  INV_X1 U21100 ( .A(n17956), .ZN(n17840) );
  AOI211_X1 U21101 ( .C1(n17853), .C2(n17841), .A(n17840), .B(n17839), .ZN(
        n17843) );
  NOR2_X1 U21102 ( .A1(n16866), .A2(n18858), .ZN(n17842) );
  AOI211_X1 U21103 ( .C1(n17844), .C2(n17955), .A(n17843), .B(n17842), .ZN(
        n17849) );
  AOI22_X1 U21104 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17850), .B1(
        n17851), .B2(n12780), .ZN(n17845) );
  XNOR2_X1 U21105 ( .A(n12779), .B(n17845), .ZN(n18179) );
  AOI22_X1 U21106 ( .A1(n17873), .A2(n18179), .B1(n17847), .B2(n17846), .ZN(
        n17848) );
  OAI211_X1 U21107 ( .C1(n17861), .C2(n12779), .A(n17849), .B(n17848), .ZN(
        P3_U2820) );
  NAND2_X1 U21108 ( .A1(n17851), .A2(n17850), .ZN(n17852) );
  XNOR2_X1 U21109 ( .A(n17852), .B(n12780), .ZN(n18187) );
  NOR2_X1 U21110 ( .A1(n16866), .A2(n18856), .ZN(n18186) );
  INV_X1 U21111 ( .A(n17853), .ZN(n17858) );
  NAND2_X1 U21112 ( .A1(n18692), .A2(n17854), .ZN(n17864) );
  NOR2_X1 U21113 ( .A1(n17863), .A2(n17864), .ZN(n17855) );
  AOI21_X1 U21114 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17956), .A(
        n17855), .ZN(n17857) );
  OAI22_X1 U21115 ( .A1(n17858), .A2(n17857), .B1(n17946), .B2(n17856), .ZN(
        n17859) );
  AOI211_X1 U21116 ( .C1(n17873), .C2(n18187), .A(n18186), .B(n17859), .ZN(
        n17860) );
  OAI221_X1 U21117 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17862), .C1(
        n12780), .C2(n17861), .A(n17860), .ZN(P3_U2821) );
  INV_X1 U21118 ( .A(n17871), .ZN(n18207) );
  AOI21_X1 U21119 ( .B1(n18297), .B2(n17878), .A(n17933), .ZN(n17880) );
  NAND2_X1 U21120 ( .A1(n18692), .A2(n17879), .ZN(n17877) );
  AOI21_X1 U21121 ( .B1(n17880), .B2(n17877), .A(n17863), .ZN(n17866) );
  OAI22_X1 U21122 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17864), .B1(
        n16866), .B2(n18855), .ZN(n17865) );
  AOI211_X1 U21123 ( .C1(n17867), .C2(n17955), .A(n17866), .B(n17865), .ZN(
        n17875) );
  AOI21_X1 U21124 ( .B1(n17869), .B2(n18199), .A(n17868), .ZN(n18203) );
  OAI21_X1 U21125 ( .B1(n17872), .B2(n17871), .A(n17870), .ZN(n18201) );
  AOI22_X1 U21126 ( .A1(n17953), .A2(n18203), .B1(n17873), .B2(n18201), .ZN(
        n17874) );
  OAI211_X1 U21127 ( .C1(n17876), .C2(n18207), .A(n17875), .B(n17874), .ZN(
        P3_U2822) );
  OAI22_X1 U21128 ( .A1(n17880), .A2(n17879), .B1(n17878), .B2(n17877), .ZN(
        n17887) );
  OAI21_X1 U21129 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17882), .A(
        n17881), .ZN(n18209) );
  NAND2_X1 U21130 ( .A1(n17884), .A2(n17883), .ZN(n17885) );
  INV_X1 U21131 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18195) );
  XNOR2_X1 U21132 ( .A(n17885), .B(n18195), .ZN(n18215) );
  OAI22_X1 U21133 ( .A1(n17965), .A2(n18209), .B1(n17966), .B2(n18215), .ZN(
        n17886) );
  AOI211_X1 U21134 ( .C1(n18285), .C2(P3_REIP_REG_7__SCAN_IN), .A(n17887), .B(
        n17886), .ZN(n17888) );
  OAI21_X1 U21135 ( .B1(n17946), .B2(n17889), .A(n17888), .ZN(P3_U2823) );
  NAND2_X1 U21136 ( .A1(n18692), .A2(n17890), .ZN(n17894) );
  NAND2_X1 U21137 ( .A1(n17956), .A2(n17894), .ZN(n17913) );
  OAI21_X1 U21138 ( .B1(n17891), .B2(n17893), .A(n17892), .ZN(n18224) );
  OAI22_X1 U21139 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17894), .B1(
        n17965), .B2(n18224), .ZN(n17895) );
  AOI21_X1 U21140 ( .B1(n18285), .B2(P3_REIP_REG_6__SCAN_IN), .A(n17895), .ZN(
        n17900) );
  AOI21_X1 U21141 ( .B1(n18219), .B2(n17897), .A(n17896), .ZN(n18222) );
  AOI22_X1 U21142 ( .A1(n17953), .A2(n18222), .B1(n17898), .B2(n17955), .ZN(
        n17899) );
  OAI211_X1 U21143 ( .C1(n21122), .C2(n17913), .A(n17900), .B(n17899), .ZN(
        P3_U2824) );
  AOI21_X1 U21144 ( .B1(n17901), .B2(n17961), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17914) );
  AOI21_X1 U21145 ( .B1(n17904), .B2(n17903), .A(n17902), .ZN(n18225) );
  AOI22_X1 U21146 ( .A1(n17953), .A2(n18225), .B1(n18285), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17912) );
  AOI21_X1 U21147 ( .B1(n17907), .B2(n17906), .A(n17905), .ZN(n17908) );
  XNOR2_X1 U21148 ( .A(n17908), .B(n18231), .ZN(n18226) );
  AOI22_X1 U21149 ( .A1(n17910), .A2(n18226), .B1(n17909), .B2(n17955), .ZN(
        n17911) );
  OAI211_X1 U21150 ( .C1(n17914), .C2(n17913), .A(n17912), .B(n17911), .ZN(
        P3_U2825) );
  OAI21_X1 U21151 ( .B1(n17917), .B2(n17916), .A(n17915), .ZN(n18238) );
  OAI22_X1 U21152 ( .A1(n17965), .A2(n18238), .B1(n18340), .B2(n17918), .ZN(
        n17919) );
  AOI21_X1 U21153 ( .B1(n18285), .B2(P3_REIP_REG_4__SCAN_IN), .A(n17919), .ZN(
        n17925) );
  AOI21_X1 U21154 ( .B1(n18243), .B2(n17921), .A(n17920), .ZN(n18240) );
  OAI21_X1 U21155 ( .B1(n17923), .B2(n17922), .A(n17961), .ZN(n17935) );
  AOI22_X1 U21156 ( .A1(n17953), .A2(n18240), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17935), .ZN(n17924) );
  OAI211_X1 U21157 ( .C1(n17946), .C2(n17926), .A(n17925), .B(n17924), .ZN(
        P3_U2826) );
  OAI21_X1 U21158 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17928), .A(
        n17927), .ZN(n18253) );
  AOI21_X1 U21159 ( .B1(n17931), .B2(n17930), .A(n17929), .ZN(n18250) );
  AOI22_X1 U21160 ( .A1(n17953), .A2(n18250), .B1(n18285), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17938) );
  OAI21_X1 U21161 ( .B1(n17933), .B2(n17949), .A(n17932), .ZN(n17934) );
  AOI22_X1 U21162 ( .A1(n17936), .A2(n17955), .B1(n17935), .B2(n17934), .ZN(
        n17937) );
  OAI211_X1 U21163 ( .C1(n17965), .C2(n18253), .A(n17938), .B(n17937), .ZN(
        P3_U2827) );
  AOI21_X1 U21164 ( .B1(n17941), .B2(n17940), .A(n17939), .ZN(n18260) );
  INV_X1 U21165 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18843) );
  NOR2_X1 U21166 ( .A1(n16866), .A2(n18843), .ZN(n18266) );
  OAI21_X1 U21167 ( .B1(n17944), .B2(n17943), .A(n17942), .ZN(n18269) );
  OAI22_X1 U21168 ( .A1(n17946), .A2(n17945), .B1(n17965), .B2(n18269), .ZN(
        n17947) );
  AOI211_X1 U21169 ( .C1(n17953), .C2(n18260), .A(n18266), .B(n17947), .ZN(
        n17948) );
  OAI221_X1 U21170 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18349), .C1(
        n17949), .C2(n17961), .A(n17948), .ZN(P3_U2828) );
  OAI21_X1 U21171 ( .B1(n17959), .B2(n17951), .A(n17950), .ZN(n18280) );
  NAND2_X1 U21172 ( .A1(n18925), .A2(n17960), .ZN(n17952) );
  XNOR2_X1 U21173 ( .A(n17952), .B(n17951), .ZN(n18276) );
  AOI22_X1 U21174 ( .A1(n17953), .A2(n18276), .B1(n18245), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17958) );
  AOI22_X1 U21175 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17956), .B1(
        n17955), .B2(n17954), .ZN(n17957) );
  OAI211_X1 U21176 ( .C1(n17965), .C2(n18280), .A(n17958), .B(n17957), .ZN(
        P3_U2829) );
  AOI21_X1 U21177 ( .B1(n17960), .B2(n18925), .A(n17959), .ZN(n18284) );
  INV_X1 U21178 ( .A(n18284), .ZN(n18281) );
  NAND3_X1 U21179 ( .A1(n18926), .A2(n17962), .A3(n17961), .ZN(n17963) );
  AOI22_X1 U21180 ( .A1(n18245), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17963), .ZN(n17964) );
  OAI221_X1 U21181 ( .B1(n18284), .B2(n17966), .C1(n18281), .C2(n17965), .A(
        n17964), .ZN(P3_U2830) );
  AOI21_X1 U21182 ( .B1(n18287), .B2(n17985), .A(n21067), .ZN(n17976) );
  INV_X1 U21183 ( .A(n18744), .ZN(n18007) );
  OAI22_X1 U21184 ( .A1(n17968), .A2(n18162), .B1(n17967), .B2(n18007), .ZN(
        n17975) );
  AOI21_X1 U21185 ( .B1(n18287), .B2(n17994), .A(n17969), .ZN(n17972) );
  NOR2_X1 U21186 ( .A1(n18925), .A2(n18031), .ZN(n18044) );
  INV_X1 U21187 ( .A(n18044), .ZN(n18093) );
  OAI22_X1 U21188 ( .A1(n18787), .A2(n18043), .B1(n17970), .B2(n18093), .ZN(
        n18037) );
  NAND3_X1 U21189 ( .A1(n18034), .A2(n18069), .A3(n18037), .ZN(n17971) );
  NAND2_X1 U21190 ( .A1(n18254), .A2(n17971), .ZN(n17993) );
  OAI211_X1 U21191 ( .C1(n18755), .C2(n17973), .A(n17972), .B(n17993), .ZN(
        n17974) );
  OAI21_X1 U21192 ( .B1(n17975), .B2(n17974), .A(n18271), .ZN(n17986) );
  OAI21_X1 U21193 ( .B1(n17976), .B2(n18286), .A(n17986), .ZN(n17979) );
  NOR2_X1 U21194 ( .A1(n18285), .A2(n18271), .ZN(n18267) );
  INV_X1 U21195 ( .A(n17977), .ZN(n17978) );
  AOI222_X1 U21196 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17979), 
        .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18267), .C1(n17979), 
        .C2(n17978), .ZN(n17981) );
  NAND2_X1 U21197 ( .A1(n18285), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17980) );
  OAI211_X1 U21198 ( .C1(n17982), .C2(n18175), .A(n17981), .B(n17980), .ZN(
        P3_U2835) );
  INV_X1 U21199 ( .A(n18029), .ZN(n18045) );
  NAND3_X1 U21200 ( .A1(n18271), .A2(n18045), .A3(n17983), .ZN(n18068) );
  NOR2_X1 U21201 ( .A1(n17984), .A2(n18068), .ZN(n18018) );
  INV_X1 U21202 ( .A(n18267), .ZN(n18272) );
  AOI21_X1 U21203 ( .B1(n18272), .B2(n17986), .A(n17985), .ZN(n17987) );
  AOI21_X1 U21204 ( .B1(n17988), .B2(n18018), .A(n17987), .ZN(n17990) );
  OAI211_X1 U21205 ( .C1(n17991), .C2(n18175), .A(n17990), .B(n17989), .ZN(
        P3_U2836) );
  NOR2_X1 U21206 ( .A1(n17992), .A2(n18757), .ZN(n18012) );
  INV_X1 U21207 ( .A(n17993), .ZN(n18011) );
  AOI211_X1 U21208 ( .C1(n18196), .C2(n17994), .A(n18012), .B(n18011), .ZN(
        n17996) );
  OAI22_X1 U21209 ( .A1(n17996), .A2(n18286), .B1(n17995), .B2(n18272), .ZN(
        n18001) );
  NOR3_X1 U21210 ( .A1(n17998), .A2(n17997), .A3(n18014), .ZN(n18000) );
  AOI221_X1 U21211 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18001), 
        .C1(n18000), .C2(n18001), .A(n17999), .ZN(n18005) );
  AOI22_X1 U21212 ( .A1(n18282), .A2(n18003), .B1(n9863), .B2(n18002), .ZN(
        n18004) );
  OAI211_X1 U21213 ( .C1(n18206), .C2(n18006), .A(n18005), .B(n18004), .ZN(
        P3_U2837) );
  OAI22_X1 U21214 ( .A1(n18009), .A2(n18162), .B1(n18008), .B2(n18007), .ZN(
        n18010) );
  NOR3_X1 U21215 ( .A1(n18267), .A2(n18011), .A3(n18010), .ZN(n18015) );
  NOR2_X1 U21216 ( .A1(n18012), .A2(n20898), .ZN(n18013) );
  AOI21_X1 U21217 ( .B1(n18015), .B2(n18013), .A(n18285), .ZN(n18022) );
  AOI21_X1 U21218 ( .B1(n18125), .B2(n18015), .A(n18014), .ZN(n18016) );
  AOI22_X1 U21219 ( .A1(n18018), .A2(n18017), .B1(n18022), .B2(n18016), .ZN(
        n18020) );
  OAI211_X1 U21220 ( .C1(n18021), .C2(n18175), .A(n18020), .B(n18019), .ZN(
        P3_U2838) );
  OAI221_X1 U21221 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18023), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n18272), .A(n18022), .ZN(
        n18024) );
  OAI211_X1 U21222 ( .C1(n18026), .C2(n18175), .A(n18025), .B(n18024), .ZN(
        P3_U2839) );
  AOI22_X1 U21223 ( .A1(n18744), .A2(n18028), .B1(n18140), .B2(n18027), .ZN(
        n18073) );
  OAI21_X1 U21224 ( .B1(n18029), .B2(n18070), .A(n18785), .ZN(n18033) );
  INV_X1 U21225 ( .A(n18058), .ZN(n18030) );
  OAI21_X1 U21226 ( .B1(n18031), .B2(n18030), .A(n18287), .ZN(n18032) );
  NAND3_X1 U21227 ( .A1(n18073), .A2(n18033), .A3(n18032), .ZN(n18046) );
  NOR2_X1 U21228 ( .A1(n18744), .A2(n18140), .ZN(n18157) );
  OAI22_X1 U21229 ( .A1(n18789), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n18034), .B2(n18157), .ZN(n18048) );
  AOI211_X1 U21230 ( .C1(n18035), .C2(n18167), .A(n18046), .B(n18048), .ZN(
        n18038) );
  AOI22_X1 U21231 ( .A1(n18038), .A2(n18037), .B1(n18043), .B2(n18036), .ZN(
        n18040) );
  AOI22_X1 U21232 ( .A1(n18271), .A2(n18040), .B1(n9863), .B2(n18039), .ZN(
        n18042) );
  OAI211_X1 U21233 ( .C1(n18272), .C2(n18043), .A(n18042), .B(n18041), .ZN(
        P3_U2840) );
  INV_X1 U21234 ( .A(n18068), .ZN(n18052) );
  AOI21_X1 U21235 ( .B1(n18045), .B2(n18044), .A(n18755), .ZN(n18047) );
  NOR3_X1 U21236 ( .A1(n18047), .A2(n18046), .A3(n18286), .ZN(n18059) );
  AOI21_X1 U21237 ( .B1(n18270), .B2(n18049), .A(n18048), .ZN(n18050) );
  AOI211_X1 U21238 ( .C1(n18059), .C2(n18050), .A(n18245), .B(n21148), .ZN(
        n18051) );
  AOI21_X1 U21239 ( .B1(n18053), .B2(n18052), .A(n18051), .ZN(n18055) );
  OAI211_X1 U21240 ( .C1(n18056), .C2(n18175), .A(n18055), .B(n18054), .ZN(
        P3_U2841) );
  AOI22_X1 U21241 ( .A1(n18245), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n9863), 
        .B2(n18057), .ZN(n18062) );
  AOI221_X1 U21242 ( .B1(n18157), .B2(n18059), .C1(n18058), .C2(n18059), .A(
        n18245), .ZN(n18065) );
  AND3_X1 U21243 ( .A1(n18270), .A2(n21131), .A3(P3_STATE2_REG_2__SCAN_IN), 
        .ZN(n18060) );
  OAI21_X1 U21244 ( .B1(n18065), .B2(n18060), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18061) );
  OAI211_X1 U21245 ( .C1(n18063), .C2(n18068), .A(n18062), .B(n18061), .ZN(
        P3_U2842) );
  AOI22_X1 U21246 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18065), .B1(
        n9863), .B2(n18064), .ZN(n18067) );
  OAI211_X1 U21247 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18068), .A(
        n18067), .B(n18066), .ZN(P3_U2843) );
  NAND2_X1 U21248 ( .A1(n18787), .A2(n18925), .ZN(n18256) );
  NAND3_X1 U21249 ( .A1(n18069), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18256), .ZN(n18075) );
  NAND2_X1 U21250 ( .A1(n18785), .A2(n18070), .ZN(n18071) );
  AOI22_X1 U21251 ( .A1(n18072), .A2(n18071), .B1(n18157), .B2(n18757), .ZN(
        n18074) );
  NAND2_X1 U21252 ( .A1(n18271), .A2(n18073), .ZN(n18096) );
  AOI211_X1 U21253 ( .C1(n18254), .C2(n18075), .A(n18074), .B(n18096), .ZN(
        n18085) );
  AOI221_X1 U21254 ( .B1(n18236), .B2(n18085), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n18085), .A(n18245), .ZN(
        n18080) );
  INV_X1 U21255 ( .A(n18076), .ZN(n18120) );
  NOR2_X1 U21256 ( .A1(n18261), .A2(n18924), .ZN(n18235) );
  AOI22_X1 U21257 ( .A1(n18785), .A2(n18233), .B1(n18235), .B2(n18262), .ZN(
        n18247) );
  INV_X1 U21258 ( .A(n18077), .ZN(n18119) );
  NOR2_X1 U21259 ( .A1(n18247), .A2(n18119), .ZN(n18208) );
  NAND3_X1 U21260 ( .A1(n18095), .A2(n18120), .A3(n18208), .ZN(n18107) );
  AOI211_X1 U21261 ( .C1(n18078), .C2(n18107), .A(n18118), .B(n18286), .ZN(
        n18098) );
  AOI22_X1 U21262 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18080), .B1(
        n18098), .B2(n18079), .ZN(n18082) );
  OAI211_X1 U21263 ( .C1(n18175), .C2(n18083), .A(n18082), .B(n18081), .ZN(
        P3_U2844) );
  NOR3_X1 U21264 ( .A1(n18245), .A2(n18085), .A3(n18084), .ZN(n18087) );
  AOI211_X1 U21265 ( .C1(n18088), .C2(n18098), .A(n18087), .B(n18086), .ZN(
        n18089) );
  OAI21_X1 U21266 ( .B1(n18090), .B2(n18175), .A(n18089), .ZN(P3_U2845) );
  INV_X1 U21267 ( .A(n18167), .ZN(n18177) );
  OAI22_X1 U21268 ( .A1(n18757), .A2(n18091), .B1(n18789), .B2(n18122), .ZN(
        n18092) );
  INV_X1 U21269 ( .A(n18092), .ZN(n18161) );
  OAI21_X1 U21270 ( .B1(n18118), .B2(n18787), .A(n18093), .ZN(n18094) );
  OAI211_X1 U21271 ( .C1(n18095), .C2(n18177), .A(n18161), .B(n18094), .ZN(
        n18109) );
  OAI221_X1 U21272 ( .B1(n18096), .B2(n18196), .C1(n18096), .C2(n18109), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18101) );
  AOI22_X1 U21273 ( .A1(n18099), .A2(n9863), .B1(n18098), .B2(n18097), .ZN(
        n18100) );
  OAI221_X1 U21274 ( .B1(n18285), .B2(n18101), .C1(n16866), .C2(n18868), .A(
        n18100), .ZN(P3_U2846) );
  NOR2_X1 U21275 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18102), .ZN(
        n18103) );
  NOR2_X1 U21276 ( .A1(n18104), .A2(n18103), .ZN(n18115) );
  NOR2_X1 U21277 ( .A1(n18105), .A2(n18162), .ZN(n18111) );
  NAND2_X1 U21278 ( .A1(n18106), .A2(n18118), .ZN(n18110) );
  NAND2_X1 U21279 ( .A1(n18118), .A2(n18107), .ZN(n18108) );
  AOI22_X1 U21280 ( .A1(n18111), .A2(n18110), .B1(n18109), .B2(n18108), .ZN(
        n18113) );
  OAI22_X1 U21281 ( .A1(n18113), .A2(n18286), .B1(n18175), .B2(n18112), .ZN(
        n18114) );
  AOI21_X1 U21282 ( .B1(n18115), .B2(n18282), .A(n18114), .ZN(n18117) );
  OAI211_X1 U21283 ( .C1(n18272), .C2(n18118), .A(n18117), .B(n18116), .ZN(
        P3_U2847) );
  NOR3_X1 U21284 ( .A1(n18247), .A2(n18119), .A3(n18286), .ZN(n18191) );
  NAND2_X1 U21285 ( .A1(n18120), .A2(n18191), .ZN(n18136) );
  OAI22_X1 U21286 ( .A1(n20868), .A2(n18286), .B1(n18136), .B2(n18121), .ZN(
        n18128) );
  NAND2_X1 U21287 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18122), .ZN(
        n18184) );
  INV_X1 U21288 ( .A(n18184), .ZN(n18158) );
  NAND2_X1 U21289 ( .A1(n18123), .A2(n18158), .ZN(n18150) );
  NAND2_X1 U21290 ( .A1(n18787), .A2(n18150), .ZN(n18143) );
  OAI211_X1 U21291 ( .C1(n18125), .C2(n18124), .A(n18161), .B(n18143), .ZN(
        n18127) );
  OAI22_X1 U21292 ( .A1(n20868), .A2(n18272), .B1(n16866), .B2(n21089), .ZN(
        n18126) );
  AOI221_X1 U21293 ( .B1(n20868), .B2(n18128), .C1(n18127), .C2(n18128), .A(
        n18126), .ZN(n18132) );
  AOI22_X1 U21294 ( .A1(n18282), .A2(n18130), .B1(n9863), .B2(n18129), .ZN(
        n18131) );
  OAI211_X1 U21295 ( .C1(n18206), .C2(n18133), .A(n18132), .B(n18131), .ZN(
        P3_U2848) );
  AOI22_X1 U21296 ( .A1(n18163), .A2(n18135), .B1(n18282), .B2(n18134), .ZN(
        n18137) );
  NAND2_X1 U21297 ( .A1(n18137), .A2(n18136), .ZN(n18183) );
  AOI22_X1 U21298 ( .A1(n18245), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18138), 
        .B2(n18183), .ZN(n18146) );
  AOI22_X1 U21299 ( .A1(n18744), .A2(n18141), .B1(n18140), .B2(n18139), .ZN(
        n18142) );
  OAI211_X1 U21300 ( .C1(n18151), .C2(n18177), .A(n18161), .B(n18142), .ZN(
        n18149) );
  OAI211_X1 U21301 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18177), .A(
        n18271), .B(n18143), .ZN(n18144) );
  OAI211_X1 U21302 ( .C1(n18149), .C2(n18144), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n16866), .ZN(n18145) );
  OAI211_X1 U21303 ( .C1(n18175), .C2(n18147), .A(n18146), .B(n18145), .ZN(
        P3_U2849) );
  AOI211_X1 U21304 ( .C1(n18150), .C2(n18787), .A(n18149), .B(n18148), .ZN(
        n18156) );
  AOI22_X1 U21305 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18271), .B1(
        n18151), .B2(n18183), .ZN(n18155) );
  AOI22_X1 U21306 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18267), .B1(
        n9863), .B2(n18152), .ZN(n18154) );
  OAI211_X1 U21307 ( .C1(n18156), .C2(n18155), .A(n18154), .B(n18153), .ZN(
        P3_U2850) );
  INV_X1 U21308 ( .A(n18157), .ZN(n18165) );
  AOI21_X1 U21309 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18158), .A(
        n18755), .ZN(n18164) );
  AOI21_X1 U21310 ( .B1(n18744), .B2(n18159), .A(n18286), .ZN(n18160) );
  OAI211_X1 U21311 ( .C1(n18163), .C2(n18162), .A(n18161), .B(n18160), .ZN(
        n18185) );
  AOI211_X1 U21312 ( .C1(n18166), .C2(n18165), .A(n18164), .B(n18185), .ZN(
        n18178) );
  AOI22_X1 U21313 ( .A1(n18787), .A2(n12779), .B1(n18168), .B2(n18167), .ZN(
        n18170) );
  AOI211_X1 U21314 ( .C1(n18178), .C2(n18170), .A(n18245), .B(n18169), .ZN(
        n18172) );
  AOI211_X1 U21315 ( .C1(n18173), .C2(n18183), .A(n18172), .B(n18171), .ZN(
        n18174) );
  OAI21_X1 U21316 ( .B1(n18176), .B2(n18175), .A(n18174), .ZN(P3_U2851) );
  AOI221_X1 U21317 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18178), .C1(
        n18177), .C2(n18178), .A(n18245), .ZN(n18180) );
  AOI22_X1 U21318 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18180), .B1(
        n9863), .B2(n18179), .ZN(n18182) );
  NAND3_X1 U21319 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n12779), .A3(
        n18183), .ZN(n18181) );
  OAI211_X1 U21320 ( .C1(n18858), .C2(n16866), .A(n18182), .B(n18181), .ZN(
        P3_U2852) );
  INV_X1 U21321 ( .A(n18183), .ZN(n18190) );
  OAI221_X1 U21322 ( .B1(n18185), .B2(n18787), .C1(n18185), .C2(n18184), .A(
        n16866), .ZN(n18189) );
  AOI21_X1 U21323 ( .B1(n9863), .B2(n18187), .A(n18186), .ZN(n18188) );
  OAI221_X1 U21324 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18190), .C1(
        n12780), .C2(n18189), .A(n18188), .ZN(P3_U2853) );
  INV_X1 U21325 ( .A(n18191), .ZN(n18220) );
  NOR3_X1 U21326 ( .A1(n18219), .A2(n18195), .A3(n18220), .ZN(n18200) );
  AOI22_X1 U21327 ( .A1(n18785), .A2(n18193), .B1(n18254), .B2(n18192), .ZN(
        n18194) );
  NAND2_X1 U21328 ( .A1(n18194), .A2(n18256), .ZN(n18217) );
  AOI211_X1 U21329 ( .C1(n18196), .C2(n18219), .A(n18195), .B(n18217), .ZN(
        n18211) );
  INV_X1 U21330 ( .A(n18237), .ZN(n18273) );
  OAI21_X1 U21331 ( .B1(n18211), .B2(n18273), .A(n18272), .ZN(n18198) );
  NOR2_X1 U21332 ( .A1(n16866), .A2(n18855), .ZN(n18197) );
  AOI221_X1 U21333 ( .B1(n18200), .B2(n18199), .C1(n18198), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18197), .ZN(n18205) );
  AOI22_X1 U21334 ( .A1(n18282), .A2(n18203), .B1(n9863), .B2(n18201), .ZN(
        n18204) );
  OAI211_X1 U21335 ( .C1(n18207), .C2(n18206), .A(n18205), .B(n18204), .ZN(
        P3_U2854) );
  NOR2_X1 U21336 ( .A1(n16866), .A2(n18852), .ZN(n18213) );
  OAI221_X1 U21337 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18208), .A(n18271), .ZN(
        n18210) );
  OAI22_X1 U21338 ( .A1(n18211), .A2(n18210), .B1(n18279), .B2(n18209), .ZN(
        n18212) );
  AOI211_X1 U21339 ( .C1(n18267), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18213), .B(n18212), .ZN(n18214) );
  OAI21_X1 U21340 ( .B1(n18216), .B2(n18215), .A(n18214), .ZN(P3_U2855) );
  OAI21_X1 U21341 ( .B1(n18286), .B2(n18217), .A(n16866), .ZN(n18230) );
  NAND2_X1 U21342 ( .A1(n18285), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n18218) );
  OAI221_X1 U21343 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18220), .C1(
        n18219), .C2(n18230), .A(n18218), .ZN(n18221) );
  AOI21_X1 U21344 ( .B1(n18282), .B2(n18222), .A(n18221), .ZN(n18223) );
  OAI21_X1 U21345 ( .B1(n18279), .B2(n18224), .A(n18223), .ZN(P3_U2856) );
  AOI22_X1 U21346 ( .A1(n18245), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18282), 
        .B2(n18225), .ZN(n18229) );
  NOR4_X1 U21347 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18247), .A3(
        n18246), .A4(n18286), .ZN(n18227) );
  INV_X1 U21348 ( .A(n18279), .ZN(n18283) );
  AOI22_X1 U21349 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18227), .B1(
        n18283), .B2(n18226), .ZN(n18228) );
  OAI211_X1 U21350 ( .C1(n18231), .C2(n18230), .A(n18229), .B(n18228), .ZN(
        P3_U2857) );
  NOR2_X1 U21351 ( .A1(n18247), .A2(n18286), .ZN(n18232) );
  NAND2_X1 U21352 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18232), .ZN(
        n18244) );
  NOR2_X1 U21353 ( .A1(n18757), .A2(n18233), .ZN(n18259) );
  NOR2_X1 U21354 ( .A1(n18259), .A2(n18246), .ZN(n18234) );
  OAI211_X1 U21355 ( .C1(n18236), .C2(n18235), .A(n18234), .B(n18256), .ZN(
        n18248) );
  AOI21_X1 U21356 ( .B1(n18237), .B2(n18248), .A(n18267), .ZN(n18242) );
  OAI22_X1 U21357 ( .A1(n16866), .A2(n18846), .B1(n18279), .B2(n18238), .ZN(
        n18239) );
  AOI21_X1 U21358 ( .B1(n18282), .B2(n18240), .A(n18239), .ZN(n18241) );
  OAI221_X1 U21359 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18244), .C1(
        n18243), .C2(n18242), .A(n18241), .ZN(P3_U2858) );
  AOI22_X1 U21360 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18267), .B1(
        n18245), .B2(P3_REIP_REG_3__SCAN_IN), .ZN(n18252) );
  AOI21_X1 U21361 ( .B1(n18247), .B2(n18246), .A(n18286), .ZN(n18249) );
  AOI22_X1 U21362 ( .A1(n18282), .A2(n18250), .B1(n18249), .B2(n18248), .ZN(
        n18251) );
  OAI211_X1 U21363 ( .C1(n18279), .C2(n18253), .A(n18252), .B(n18251), .ZN(
        P3_U2859) );
  NOR2_X1 U21364 ( .A1(n18924), .A2(n18925), .ZN(n18255) );
  AOI22_X1 U21365 ( .A1(n18785), .A2(n18255), .B1(n18254), .B2(n18924), .ZN(
        n18257) );
  AOI21_X1 U21366 ( .B1(n18257), .B2(n18256), .A(n18261), .ZN(n18258) );
  AOI211_X1 U21367 ( .C1(n18260), .C2(n18744), .A(n18259), .B(n18258), .ZN(
        n18264) );
  NAND3_X1 U21368 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18262), .A3(
        n18261), .ZN(n18263) );
  AOI21_X1 U21369 ( .B1(n18264), .B2(n18263), .A(n18286), .ZN(n18265) );
  AOI211_X1 U21370 ( .C1(n18267), .C2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n18266), .B(n18265), .ZN(n18268) );
  OAI21_X1 U21371 ( .B1(n18279), .B2(n18269), .A(n18268), .ZN(P3_U2860) );
  NAND3_X1 U21372 ( .A1(n18271), .A2(n18270), .A3(n18925), .ZN(n18289) );
  AOI21_X1 U21373 ( .B1(n18272), .B2(n18289), .A(n18924), .ZN(n18275) );
  AOI211_X1 U21374 ( .C1(n18789), .C2(n18925), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18273), .ZN(n18274) );
  AOI211_X1 U21375 ( .C1(n18282), .C2(n18276), .A(n18275), .B(n18274), .ZN(
        n18278) );
  NAND2_X1 U21376 ( .A1(n18285), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18277) );
  OAI211_X1 U21377 ( .C1(n18280), .C2(n18279), .A(n18278), .B(n18277), .ZN(
        P3_U2861) );
  AOI22_X1 U21378 ( .A1(n18284), .A2(n18283), .B1(n18282), .B2(n18281), .ZN(
        n18291) );
  NAND2_X1 U21379 ( .A1(n18285), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18290) );
  OAI211_X1 U21380 ( .C1(n18287), .C2(n18286), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n16866), .ZN(n18288) );
  NAND4_X1 U21381 ( .A1(n18291), .A2(n18290), .A3(n18289), .A4(n18288), .ZN(
        P3_U2862) );
  INV_X1 U21382 ( .A(n18292), .ZN(n18293) );
  AOI211_X1 U21383 ( .C1(n18294), .C2(n18293), .A(n18926), .B(n18971), .ZN(
        n18811) );
  OAI21_X1 U21384 ( .B1(n18811), .B2(n18295), .A(n18304), .ZN(n18296) );
  OAI221_X1 U21385 ( .B1(n18607), .B2(n18956), .C1(n18607), .C2(n18304), .A(
        n18296), .ZN(P3_U2863) );
  NAND2_X1 U21386 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18541) );
  NOR2_X1 U21387 ( .A1(n18956), .A2(n18297), .ZN(n18299) );
  AOI221_X1 U21388 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18541), .C1(n18299), 
        .C2(n18541), .A(n18298), .ZN(n18303) );
  OAI221_X1 U21389 ( .B1(n18663), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18663), .C2(n18300), .A(n18304), .ZN(n18301) );
  AOI22_X1 U21390 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18303), .B1(
        n18301), .B2(n18798), .ZN(P3_U2865) );
  INV_X1 U21391 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20929) );
  NOR2_X1 U21392 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20929), .ZN(
        n18585) );
  NOR2_X1 U21393 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18798), .ZN(
        n18495) );
  NOR2_X1 U21394 ( .A1(n18585), .A2(n18495), .ZN(n18302) );
  OAI22_X1 U21395 ( .A1(n18303), .A2(n20929), .B1(n18302), .B2(n18301), .ZN(
        P3_U2866) );
  NOR2_X1 U21396 ( .A1(n18801), .A2(n18304), .ZN(P3_U2867) );
  NAND2_X1 U21397 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18792) );
  NAND2_X1 U21398 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18305) );
  NOR2_X2 U21399 ( .A1(n18792), .A2(n18305), .ZN(n18685) );
  NAND2_X1 U21400 ( .A1(n18793), .A2(n18607), .ZN(n18794) );
  NAND2_X1 U21401 ( .A1(n18798), .A2(n20929), .ZN(n18446) );
  NOR2_X1 U21402 ( .A1(n18794), .A2(n18446), .ZN(n18421) );
  CLKBUF_X1 U21403 ( .A(n18421), .Z(n18417) );
  NOR2_X1 U21404 ( .A1(n18685), .A2(n18417), .ZN(n18383) );
  OAI21_X1 U21405 ( .B1(n18607), .B2(n18935), .A(n18518), .ZN(n18470) );
  INV_X1 U21406 ( .A(n18305), .ZN(n18638) );
  NOR2_X1 U21407 ( .A1(n18793), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18562) );
  NOR2_X1 U21408 ( .A1(n18607), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18539) );
  OR2_X1 U21409 ( .A1(n18562), .A2(n18539), .ZN(n18614) );
  NAND2_X1 U21410 ( .A1(n18638), .A2(n18614), .ZN(n18660) );
  OAI22_X1 U21411 ( .A1(n18383), .A2(n18470), .B1(n18349), .B2(n18660), .ZN(
        n18352) );
  AND2_X1 U21412 ( .A1(n18692), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18693) );
  NAND2_X1 U21413 ( .A1(n18638), .A2(n18562), .ZN(n18684) );
  INV_X1 U21414 ( .A(n18684), .ZN(n18378) );
  AND2_X1 U21415 ( .A1(n18518), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18687) );
  NOR2_X1 U21416 ( .A1(n18819), .A2(n18383), .ZN(n18346) );
  AOI22_X1 U21417 ( .A1(n18693), .A2(n18378), .B1(n18687), .B2(n18346), .ZN(
        n18311) );
  NAND2_X1 U21418 ( .A1(n18307), .A2(n18306), .ZN(n18347) );
  NOR2_X1 U21419 ( .A1(n18308), .A2(n18347), .ZN(n18354) );
  NAND2_X1 U21420 ( .A1(n18638), .A2(n18793), .ZN(n18636) );
  NOR2_X2 U21421 ( .A1(n18607), .A2(n18636), .ZN(n18738) );
  NOR2_X2 U21422 ( .A1(n18309), .A2(n18349), .ZN(n18688) );
  AOI22_X1 U21423 ( .A1(n18417), .A2(n18354), .B1(n18738), .B2(n18688), .ZN(
        n18310) );
  OAI211_X1 U21424 ( .C1(n18312), .C2(n18352), .A(n18311), .B(n18310), .ZN(
        P3_U2868) );
  NOR2_X2 U21425 ( .A1(n18349), .A2(n19420), .ZN(n18699) );
  AND2_X1 U21426 ( .A1(n18518), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18697) );
  AOI22_X1 U21427 ( .A1(n18378), .A2(n18699), .B1(n18346), .B2(n18697), .ZN(
        n18315) );
  NOR2_X1 U21428 ( .A1(n18313), .A2(n18347), .ZN(n18358) );
  AND2_X1 U21429 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18692), .ZN(n18698) );
  AOI22_X1 U21430 ( .A1(n18417), .A2(n18358), .B1(n18738), .B2(n18698), .ZN(
        n18314) );
  OAI211_X1 U21431 ( .C1(n18316), .C2(n18352), .A(n18315), .B(n18314), .ZN(
        P3_U2869) );
  NOR2_X2 U21432 ( .A1(n18349), .A2(n20927), .ZN(n18704) );
  NOR2_X2 U21433 ( .A1(n18612), .A2(n18317), .ZN(n18703) );
  AOI22_X1 U21434 ( .A1(n18378), .A2(n18704), .B1(n18346), .B2(n18703), .ZN(
        n18320) );
  NOR2_X1 U21435 ( .A1(n18318), .A2(n18347), .ZN(n18361) );
  AND2_X1 U21436 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18692), .ZN(n18705) );
  AOI22_X1 U21437 ( .A1(n18417), .A2(n18361), .B1(n18738), .B2(n18705), .ZN(
        n18319) );
  OAI211_X1 U21438 ( .C1(n18321), .C2(n18352), .A(n18320), .B(n18319), .ZN(
        P3_U2870) );
  NOR2_X2 U21439 ( .A1(n19430), .A2(n18349), .ZN(n18711) );
  NOR2_X2 U21440 ( .A1(n18612), .A2(n18322), .ZN(n18709) );
  AOI22_X1 U21441 ( .A1(n18738), .A2(n18711), .B1(n18346), .B2(n18709), .ZN(
        n18325) );
  NOR2_X1 U21442 ( .A1(n18323), .A2(n18347), .ZN(n18364) );
  NOR2_X2 U21443 ( .A1(n18349), .A2(n21059), .ZN(n18710) );
  AOI22_X1 U21444 ( .A1(n18417), .A2(n18364), .B1(n18378), .B2(n18710), .ZN(
        n18324) );
  OAI211_X1 U21445 ( .C1(n18326), .C2(n18352), .A(n18325), .B(n18324), .ZN(
        P3_U2871) );
  NOR2_X2 U21446 ( .A1(n21060), .A2(n18349), .ZN(n18717) );
  NOR2_X2 U21447 ( .A1(n18612), .A2(n18327), .ZN(n18715) );
  AOI22_X1 U21448 ( .A1(n18738), .A2(n18717), .B1(n18346), .B2(n18715), .ZN(
        n18330) );
  NOR2_X1 U21449 ( .A1(n18328), .A2(n18347), .ZN(n18367) );
  NOR2_X2 U21450 ( .A1(n18349), .A2(n20915), .ZN(n18716) );
  AOI22_X1 U21451 ( .A1(n18417), .A2(n18367), .B1(n18378), .B2(n18716), .ZN(
        n18329) );
  OAI211_X1 U21452 ( .C1(n18331), .C2(n18352), .A(n18330), .B(n18329), .ZN(
        P3_U2872) );
  NOR2_X2 U21453 ( .A1(n18332), .A2(n18349), .ZN(n18723) );
  NOR2_X2 U21454 ( .A1(n18612), .A2(n18333), .ZN(n18721) );
  AOI22_X1 U21455 ( .A1(n18738), .A2(n18723), .B1(n18346), .B2(n18721), .ZN(
        n18336) );
  NOR2_X1 U21456 ( .A1(n18334), .A2(n18347), .ZN(n18370) );
  AND2_X1 U21457 ( .A1(n18692), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18722) );
  AOI22_X1 U21458 ( .A1(n18417), .A2(n18370), .B1(n18378), .B2(n18722), .ZN(
        n18335) );
  OAI211_X1 U21459 ( .C1(n18337), .C2(n18352), .A(n18336), .B(n18335), .ZN(
        P3_U2873) );
  AND2_X1 U21460 ( .A1(n18692), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18729) );
  NOR2_X2 U21461 ( .A1(n18612), .A2(n18338), .ZN(n18727) );
  AOI22_X1 U21462 ( .A1(n18378), .A2(n18729), .B1(n18346), .B2(n18727), .ZN(
        n18342) );
  NOR2_X1 U21463 ( .A1(n18339), .A2(n18347), .ZN(n18373) );
  NOR2_X2 U21464 ( .A1(n11079), .A2(n18340), .ZN(n18728) );
  AOI22_X1 U21465 ( .A1(n18417), .A2(n18373), .B1(n18738), .B2(n18728), .ZN(
        n18341) );
  OAI211_X1 U21466 ( .C1(n18343), .C2(n18352), .A(n18342), .B(n18341), .ZN(
        P3_U2874) );
  NOR2_X2 U21467 ( .A1(n18349), .A2(n18344), .ZN(n18734) );
  NOR2_X2 U21468 ( .A1(n18345), .A2(n18612), .ZN(n18736) );
  AOI22_X1 U21469 ( .A1(n18738), .A2(n18734), .B1(n18346), .B2(n18736), .ZN(
        n18351) );
  NOR2_X1 U21470 ( .A1(n18348), .A2(n18347), .ZN(n18376) );
  NOR2_X2 U21471 ( .A1(n19449), .A2(n18349), .ZN(n18737) );
  AOI22_X1 U21472 ( .A1(n18417), .A2(n18376), .B1(n18378), .B2(n18737), .ZN(
        n18350) );
  OAI211_X1 U21473 ( .C1(n18353), .C2(n18352), .A(n18351), .B(n18350), .ZN(
        P3_U2875) );
  INV_X1 U21474 ( .A(n18354), .ZN(n18696) );
  INV_X1 U21475 ( .A(n18446), .ZN(n18404) );
  NAND2_X1 U21476 ( .A1(n18404), .A2(n18539), .ZN(n18382) );
  NAND2_X1 U21477 ( .A1(n18793), .A2(n18686), .ZN(n18540) );
  NOR2_X1 U21478 ( .A1(n18446), .A2(n18540), .ZN(n18377) );
  AOI22_X1 U21479 ( .A1(n18688), .A2(n18378), .B1(n18687), .B2(n18377), .ZN(
        n18357) );
  NOR2_X1 U21480 ( .A1(n20929), .A2(n18541), .ZN(n18689) );
  NAND2_X1 U21481 ( .A1(n18518), .A2(n18355), .ZN(n18584) );
  NOR2_X1 U21482 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18584), .ZN(
        n18637) );
  AOI22_X1 U21483 ( .A1(n18692), .A2(n18689), .B1(n18404), .B2(n18637), .ZN(
        n18379) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18379), .B1(
        n18685), .B2(n18693), .ZN(n18356) );
  OAI211_X1 U21485 ( .C1(n18696), .C2(n18382), .A(n18357), .B(n18356), .ZN(
        P3_U2876) );
  INV_X1 U21486 ( .A(n18358), .ZN(n18702) );
  AOI22_X1 U21487 ( .A1(n18685), .A2(n18699), .B1(n18697), .B2(n18377), .ZN(
        n18360) );
  AOI22_X1 U21488 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18379), .B1(
        n18378), .B2(n18698), .ZN(n18359) );
  OAI211_X1 U21489 ( .C1(n18702), .C2(n18382), .A(n18360), .B(n18359), .ZN(
        P3_U2877) );
  INV_X1 U21490 ( .A(n18361), .ZN(n18708) );
  AOI22_X1 U21491 ( .A1(n18685), .A2(n18704), .B1(n18703), .B2(n18377), .ZN(
        n18363) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18379), .B1(
        n18378), .B2(n18705), .ZN(n18362) );
  OAI211_X1 U21493 ( .C1(n18708), .C2(n18382), .A(n18363), .B(n18362), .ZN(
        P3_U2878) );
  INV_X1 U21494 ( .A(n18364), .ZN(n18714) );
  AOI22_X1 U21495 ( .A1(n18378), .A2(n18711), .B1(n18709), .B2(n18377), .ZN(
        n18366) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18379), .B1(
        n18685), .B2(n18710), .ZN(n18365) );
  OAI211_X1 U21497 ( .C1(n18714), .C2(n18382), .A(n18366), .B(n18365), .ZN(
        P3_U2879) );
  INV_X1 U21498 ( .A(n18367), .ZN(n18720) );
  AOI22_X1 U21499 ( .A1(n18378), .A2(n18717), .B1(n18715), .B2(n18377), .ZN(
        n18369) );
  AOI22_X1 U21500 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18379), .B1(
        n18685), .B2(n18716), .ZN(n18368) );
  OAI211_X1 U21501 ( .C1(n18720), .C2(n18382), .A(n18369), .B(n18368), .ZN(
        P3_U2880) );
  INV_X1 U21502 ( .A(n18370), .ZN(n18726) );
  AOI22_X1 U21503 ( .A1(n18685), .A2(n18722), .B1(n18721), .B2(n18377), .ZN(
        n18372) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18379), .B1(
        n18378), .B2(n18723), .ZN(n18371) );
  OAI211_X1 U21505 ( .C1(n18726), .C2(n18382), .A(n18372), .B(n18371), .ZN(
        P3_U2881) );
  INV_X1 U21506 ( .A(n18373), .ZN(n18732) );
  AOI22_X1 U21507 ( .A1(n18378), .A2(n18728), .B1(n18727), .B2(n18377), .ZN(
        n18375) );
  AOI22_X1 U21508 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18379), .B1(
        n18685), .B2(n18729), .ZN(n18374) );
  OAI211_X1 U21509 ( .C1(n18732), .C2(n18382), .A(n18375), .B(n18374), .ZN(
        P3_U2882) );
  INV_X1 U21510 ( .A(n18376), .ZN(n18742) );
  AOI22_X1 U21511 ( .A1(n18685), .A2(n18737), .B1(n18736), .B2(n18377), .ZN(
        n18381) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18379), .B1(
        n18378), .B2(n18734), .ZN(n18380) );
  OAI211_X1 U21513 ( .C1(n18742), .C2(n18382), .A(n18381), .B(n18380), .ZN(
        P3_U2883) );
  NAND2_X1 U21514 ( .A1(n18404), .A2(n18562), .ZN(n18403) );
  INV_X1 U21515 ( .A(n18382), .ZN(n18441) );
  INV_X1 U21516 ( .A(n18403), .ZN(n18462) );
  NOR2_X1 U21517 ( .A1(n18441), .A2(n18462), .ZN(n18425) );
  NOR2_X1 U21518 ( .A1(n18819), .A2(n18425), .ZN(n18399) );
  AOI22_X1 U21519 ( .A1(n18685), .A2(n18688), .B1(n18687), .B2(n18399), .ZN(
        n18386) );
  AOI221_X1 U21520 ( .B1(n18425), .B2(n18611), .C1(n18425), .C2(n18383), .A(
        n18470), .ZN(n18384) );
  INV_X1 U21521 ( .A(n18384), .ZN(n18400) );
  AOI22_X1 U21522 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18400), .B1(
        n18417), .B2(n18693), .ZN(n18385) );
  OAI211_X1 U21523 ( .C1(n18696), .C2(n18403), .A(n18386), .B(n18385), .ZN(
        P3_U2884) );
  AOI22_X1 U21524 ( .A1(n18417), .A2(n18699), .B1(n18697), .B2(n18399), .ZN(
        n18388) );
  AOI22_X1 U21525 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18400), .B1(
        n18685), .B2(n18698), .ZN(n18387) );
  OAI211_X1 U21526 ( .C1(n18702), .C2(n18403), .A(n18388), .B(n18387), .ZN(
        P3_U2885) );
  AOI22_X1 U21527 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18400), .B1(
        n18703), .B2(n18399), .ZN(n18390) );
  AOI22_X1 U21528 ( .A1(n18685), .A2(n18705), .B1(n18417), .B2(n18704), .ZN(
        n18389) );
  OAI211_X1 U21529 ( .C1(n18708), .C2(n18403), .A(n18390), .B(n18389), .ZN(
        P3_U2886) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18400), .B1(
        n18709), .B2(n18399), .ZN(n18392) );
  AOI22_X1 U21531 ( .A1(n18685), .A2(n18711), .B1(n18417), .B2(n18710), .ZN(
        n18391) );
  OAI211_X1 U21532 ( .C1(n18714), .C2(n18403), .A(n18392), .B(n18391), .ZN(
        P3_U2887) );
  AOI22_X1 U21533 ( .A1(n18417), .A2(n18716), .B1(n18715), .B2(n18399), .ZN(
        n18394) );
  AOI22_X1 U21534 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18400), .B1(
        n18685), .B2(n18717), .ZN(n18393) );
  OAI211_X1 U21535 ( .C1(n18720), .C2(n18403), .A(n18394), .B(n18393), .ZN(
        P3_U2888) );
  AOI22_X1 U21536 ( .A1(n18421), .A2(n18722), .B1(n18721), .B2(n18399), .ZN(
        n18396) );
  AOI22_X1 U21537 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18400), .B1(
        n18685), .B2(n18723), .ZN(n18395) );
  OAI211_X1 U21538 ( .C1(n18726), .C2(n18403), .A(n18396), .B(n18395), .ZN(
        P3_U2889) );
  AOI22_X1 U21539 ( .A1(n18421), .A2(n18729), .B1(n18727), .B2(n18399), .ZN(
        n18398) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18400), .B1(
        n18685), .B2(n18728), .ZN(n18397) );
  OAI211_X1 U21541 ( .C1(n18732), .C2(n18403), .A(n18398), .B(n18397), .ZN(
        P3_U2890) );
  AOI22_X1 U21542 ( .A1(n18421), .A2(n18737), .B1(n18736), .B2(n18399), .ZN(
        n18402) );
  AOI22_X1 U21543 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18400), .B1(
        n18685), .B2(n18734), .ZN(n18401) );
  OAI211_X1 U21544 ( .C1(n18742), .C2(n18403), .A(n18402), .B(n18401), .ZN(
        P3_U2891) );
  NOR2_X2 U21545 ( .A1(n18792), .A2(n18446), .ZN(n18489) );
  INV_X1 U21546 ( .A(n18489), .ZN(n18469) );
  AOI22_X1 U21547 ( .A1(n18693), .A2(n18441), .B1(n18687), .B2(n18420), .ZN(
        n18406) );
  AOI21_X1 U21548 ( .B1(n18793), .B2(n18611), .A(n18584), .ZN(n18494) );
  NAND2_X1 U21549 ( .A1(n18404), .A2(n18494), .ZN(n18422) );
  AOI22_X1 U21550 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18422), .B1(
        n18417), .B2(n18688), .ZN(n18405) );
  OAI211_X1 U21551 ( .C1(n18696), .C2(n18469), .A(n18406), .B(n18405), .ZN(
        P3_U2892) );
  AOI22_X1 U21552 ( .A1(n18421), .A2(n18698), .B1(n18697), .B2(n18420), .ZN(
        n18408) );
  AOI22_X1 U21553 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18422), .B1(
        n18699), .B2(n18441), .ZN(n18407) );
  OAI211_X1 U21554 ( .C1(n18702), .C2(n18469), .A(n18408), .B(n18407), .ZN(
        P3_U2893) );
  AOI22_X1 U21555 ( .A1(n18421), .A2(n18705), .B1(n18703), .B2(n18420), .ZN(
        n18410) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18422), .B1(
        n18704), .B2(n18441), .ZN(n18409) );
  OAI211_X1 U21557 ( .C1(n18708), .C2(n18469), .A(n18410), .B(n18409), .ZN(
        P3_U2894) );
  AOI22_X1 U21558 ( .A1(n18710), .A2(n18441), .B1(n18709), .B2(n18420), .ZN(
        n18412) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18422), .B1(
        n18421), .B2(n18711), .ZN(n18411) );
  OAI211_X1 U21560 ( .C1(n18714), .C2(n18469), .A(n18412), .B(n18411), .ZN(
        P3_U2895) );
  AOI22_X1 U21561 ( .A1(n18716), .A2(n18441), .B1(n18715), .B2(n18420), .ZN(
        n18414) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18422), .B1(
        n18421), .B2(n18717), .ZN(n18413) );
  OAI211_X1 U21563 ( .C1(n18720), .C2(n18469), .A(n18414), .B(n18413), .ZN(
        P3_U2896) );
  AOI22_X1 U21564 ( .A1(n18722), .A2(n18441), .B1(n18721), .B2(n18420), .ZN(
        n18416) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18422), .B1(
        n18421), .B2(n18723), .ZN(n18415) );
  OAI211_X1 U21566 ( .C1(n18726), .C2(n18469), .A(n18416), .B(n18415), .ZN(
        P3_U2897) );
  AOI22_X1 U21567 ( .A1(n18417), .A2(n18728), .B1(n18727), .B2(n18420), .ZN(
        n18419) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18422), .B1(
        n18729), .B2(n18441), .ZN(n18418) );
  OAI211_X1 U21569 ( .C1(n18732), .C2(n18469), .A(n18419), .B(n18418), .ZN(
        P3_U2898) );
  AOI22_X1 U21570 ( .A1(n18737), .A2(n18441), .B1(n18736), .B2(n18420), .ZN(
        n18424) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18422), .B1(
        n18421), .B2(n18734), .ZN(n18423) );
  OAI211_X1 U21572 ( .C1(n18742), .C2(n18469), .A(n18424), .B(n18423), .ZN(
        P3_U2899) );
  INV_X1 U21573 ( .A(n18495), .ZN(n18493) );
  NOR2_X2 U21574 ( .A1(n18794), .A2(n18493), .ZN(n18510) );
  INV_X1 U21575 ( .A(n18510), .ZN(n18468) );
  AOI21_X1 U21576 ( .B1(n18469), .B2(n18468), .A(n18819), .ZN(n18442) );
  AOI22_X1 U21577 ( .A1(n18693), .A2(n18462), .B1(n18687), .B2(n18442), .ZN(
        n18428) );
  AOI221_X1 U21578 ( .B1(n18425), .B2(n18469), .C1(n18611), .C2(n18469), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18426) );
  OAI21_X1 U21579 ( .B1(n18510), .B2(n18426), .A(n18518), .ZN(n18443) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18443), .B1(
        n18688), .B2(n18441), .ZN(n18427) );
  OAI211_X1 U21581 ( .C1(n18696), .C2(n18468), .A(n18428), .B(n18427), .ZN(
        P3_U2900) );
  AOI22_X1 U21582 ( .A1(n18699), .A2(n18462), .B1(n18697), .B2(n18442), .ZN(
        n18430) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18443), .B1(
        n18698), .B2(n18441), .ZN(n18429) );
  OAI211_X1 U21584 ( .C1(n18702), .C2(n18468), .A(n18430), .B(n18429), .ZN(
        P3_U2901) );
  AOI22_X1 U21585 ( .A1(n18705), .A2(n18441), .B1(n18703), .B2(n18442), .ZN(
        n18432) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18443), .B1(
        n18704), .B2(n18462), .ZN(n18431) );
  OAI211_X1 U21587 ( .C1(n18708), .C2(n18468), .A(n18432), .B(n18431), .ZN(
        P3_U2902) );
  AOI22_X1 U21588 ( .A1(n18711), .A2(n18441), .B1(n18709), .B2(n18442), .ZN(
        n18434) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18443), .B1(
        n18710), .B2(n18462), .ZN(n18433) );
  OAI211_X1 U21590 ( .C1(n18714), .C2(n18468), .A(n18434), .B(n18433), .ZN(
        P3_U2903) );
  AOI22_X1 U21591 ( .A1(n18717), .A2(n18441), .B1(n18715), .B2(n18442), .ZN(
        n18436) );
  AOI22_X1 U21592 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18443), .B1(
        n18716), .B2(n18462), .ZN(n18435) );
  OAI211_X1 U21593 ( .C1(n18720), .C2(n18468), .A(n18436), .B(n18435), .ZN(
        P3_U2904) );
  AOI22_X1 U21594 ( .A1(n18723), .A2(n18441), .B1(n18721), .B2(n18442), .ZN(
        n18438) );
  AOI22_X1 U21595 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18443), .B1(
        n18722), .B2(n18462), .ZN(n18437) );
  OAI211_X1 U21596 ( .C1(n18726), .C2(n18468), .A(n18438), .B(n18437), .ZN(
        P3_U2905) );
  AOI22_X1 U21597 ( .A1(n18729), .A2(n18462), .B1(n18727), .B2(n18442), .ZN(
        n18440) );
  AOI22_X1 U21598 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18443), .B1(
        n18728), .B2(n18441), .ZN(n18439) );
  OAI211_X1 U21599 ( .C1(n18732), .C2(n18468), .A(n18440), .B(n18439), .ZN(
        P3_U2906) );
  AOI22_X1 U21600 ( .A1(n18736), .A2(n18442), .B1(n18734), .B2(n18441), .ZN(
        n18445) );
  AOI22_X1 U21601 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18443), .B1(
        n18737), .B2(n18462), .ZN(n18444) );
  OAI211_X1 U21602 ( .C1(n18742), .C2(n18468), .A(n18445), .B(n18444), .ZN(
        P3_U2907) );
  NAND2_X1 U21603 ( .A1(n18495), .A2(n18539), .ZN(n18467) );
  NOR2_X1 U21604 ( .A1(n18493), .A2(n18540), .ZN(n18463) );
  AOI22_X1 U21605 ( .A1(n18693), .A2(n18489), .B1(n18687), .B2(n18463), .ZN(
        n18449) );
  NOR2_X1 U21606 ( .A1(n18793), .A2(n18446), .ZN(n18447) );
  AOI22_X1 U21607 ( .A1(n18692), .A2(n18447), .B1(n18495), .B2(n18637), .ZN(
        n18464) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18464), .B1(
        n18688), .B2(n18462), .ZN(n18448) );
  OAI211_X1 U21609 ( .C1(n18696), .C2(n18467), .A(n18449), .B(n18448), .ZN(
        P3_U2908) );
  AOI22_X1 U21610 ( .A1(n18698), .A2(n18462), .B1(n18697), .B2(n18463), .ZN(
        n18451) );
  AOI22_X1 U21611 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18464), .B1(
        n18699), .B2(n18489), .ZN(n18450) );
  OAI211_X1 U21612 ( .C1(n18702), .C2(n18467), .A(n18451), .B(n18450), .ZN(
        P3_U2909) );
  AOI22_X1 U21613 ( .A1(n18704), .A2(n18489), .B1(n18703), .B2(n18463), .ZN(
        n18453) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18464), .B1(
        n18705), .B2(n18462), .ZN(n18452) );
  OAI211_X1 U21615 ( .C1(n18708), .C2(n18467), .A(n18453), .B(n18452), .ZN(
        P3_U2910) );
  AOI22_X1 U21616 ( .A1(n18711), .A2(n18462), .B1(n18709), .B2(n18463), .ZN(
        n18455) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18464), .B1(
        n18710), .B2(n18489), .ZN(n18454) );
  OAI211_X1 U21618 ( .C1(n18714), .C2(n18467), .A(n18455), .B(n18454), .ZN(
        P3_U2911) );
  AOI22_X1 U21619 ( .A1(n18716), .A2(n18489), .B1(n18715), .B2(n18463), .ZN(
        n18457) );
  AOI22_X1 U21620 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18464), .B1(
        n18717), .B2(n18462), .ZN(n18456) );
  OAI211_X1 U21621 ( .C1(n18720), .C2(n18467), .A(n18457), .B(n18456), .ZN(
        P3_U2912) );
  AOI22_X1 U21622 ( .A1(n18722), .A2(n18489), .B1(n18721), .B2(n18463), .ZN(
        n18459) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18464), .B1(
        n18723), .B2(n18462), .ZN(n18458) );
  OAI211_X1 U21624 ( .C1(n18726), .C2(n18467), .A(n18459), .B(n18458), .ZN(
        P3_U2913) );
  AOI22_X1 U21625 ( .A1(n18729), .A2(n18489), .B1(n18727), .B2(n18463), .ZN(
        n18461) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18464), .B1(
        n18728), .B2(n18462), .ZN(n18460) );
  OAI211_X1 U21627 ( .C1(n18732), .C2(n18467), .A(n18461), .B(n18460), .ZN(
        P3_U2914) );
  AOI22_X1 U21628 ( .A1(n18736), .A2(n18463), .B1(n18734), .B2(n18462), .ZN(
        n18466) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18464), .B1(
        n18737), .B2(n18489), .ZN(n18465) );
  OAI211_X1 U21630 ( .C1(n18742), .C2(n18467), .A(n18466), .B(n18465), .ZN(
        P3_U2915) );
  NAND2_X1 U21631 ( .A1(n18495), .A2(n18562), .ZN(n18492) );
  INV_X1 U21632 ( .A(n18467), .ZN(n18534) );
  INV_X1 U21633 ( .A(n18492), .ZN(n18557) );
  NOR2_X1 U21634 ( .A1(n18534), .A2(n18557), .ZN(n18516) );
  NOR2_X1 U21635 ( .A1(n18819), .A2(n18516), .ZN(n18487) );
  AOI22_X1 U21636 ( .A1(n18688), .A2(n18489), .B1(n18687), .B2(n18487), .ZN(
        n18474) );
  INV_X1 U21637 ( .A(n18516), .ZN(n18472) );
  NAND2_X1 U21638 ( .A1(n18469), .A2(n18468), .ZN(n18471) );
  INV_X1 U21639 ( .A(n18470), .ZN(n18661) );
  OAI221_X1 U21640 ( .B1(n18472), .B2(n18663), .C1(n18472), .C2(n18471), .A(
        n18661), .ZN(n18488) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18488), .B1(
        n18693), .B2(n18510), .ZN(n18473) );
  OAI211_X1 U21642 ( .C1(n18696), .C2(n18492), .A(n18474), .B(n18473), .ZN(
        P3_U2916) );
  AOI22_X1 U21643 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18488), .B1(
        n18697), .B2(n18487), .ZN(n18476) );
  AOI22_X1 U21644 ( .A1(n18698), .A2(n18489), .B1(n18699), .B2(n18510), .ZN(
        n18475) );
  OAI211_X1 U21645 ( .C1(n18702), .C2(n18492), .A(n18476), .B(n18475), .ZN(
        P3_U2917) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18488), .B1(
        n18703), .B2(n18487), .ZN(n18478) );
  AOI22_X1 U21647 ( .A1(n18705), .A2(n18489), .B1(n18704), .B2(n18510), .ZN(
        n18477) );
  OAI211_X1 U21648 ( .C1(n18708), .C2(n18492), .A(n18478), .B(n18477), .ZN(
        P3_U2918) );
  AOI22_X1 U21649 ( .A1(n18711), .A2(n18489), .B1(n18709), .B2(n18487), .ZN(
        n18480) );
  AOI22_X1 U21650 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18488), .B1(
        n18710), .B2(n18510), .ZN(n18479) );
  OAI211_X1 U21651 ( .C1(n18714), .C2(n18492), .A(n18480), .B(n18479), .ZN(
        P3_U2919) );
  AOI22_X1 U21652 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18488), .B1(
        n18715), .B2(n18487), .ZN(n18482) );
  AOI22_X1 U21653 ( .A1(n18716), .A2(n18510), .B1(n18717), .B2(n18489), .ZN(
        n18481) );
  OAI211_X1 U21654 ( .C1(n18720), .C2(n18492), .A(n18482), .B(n18481), .ZN(
        P3_U2920) );
  AOI22_X1 U21655 ( .A1(n18722), .A2(n18510), .B1(n18721), .B2(n18487), .ZN(
        n18484) );
  AOI22_X1 U21656 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18488), .B1(
        n18723), .B2(n18489), .ZN(n18483) );
  OAI211_X1 U21657 ( .C1(n18726), .C2(n18492), .A(n18484), .B(n18483), .ZN(
        P3_U2921) );
  AOI22_X1 U21658 ( .A1(n18728), .A2(n18489), .B1(n18727), .B2(n18487), .ZN(
        n18486) );
  AOI22_X1 U21659 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18488), .B1(
        n18729), .B2(n18510), .ZN(n18485) );
  OAI211_X1 U21660 ( .C1(n18732), .C2(n18492), .A(n18486), .B(n18485), .ZN(
        P3_U2922) );
  AOI22_X1 U21661 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18488), .B1(
        n18736), .B2(n18487), .ZN(n18491) );
  AOI22_X1 U21662 ( .A1(n18737), .A2(n18510), .B1(n18734), .B2(n18489), .ZN(
        n18490) );
  OAI211_X1 U21663 ( .C1(n18742), .C2(n18492), .A(n18491), .B(n18490), .ZN(
        P3_U2923) );
  NOR2_X2 U21664 ( .A1(n18792), .A2(n18493), .ZN(n18581) );
  INV_X1 U21665 ( .A(n18581), .ZN(n18515) );
  AOI22_X1 U21666 ( .A1(n18688), .A2(n18510), .B1(n18687), .B2(n18511), .ZN(
        n18497) );
  NAND2_X1 U21667 ( .A1(n18495), .A2(n18494), .ZN(n18512) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18512), .B1(
        n18693), .B2(n18534), .ZN(n18496) );
  OAI211_X1 U21669 ( .C1(n18696), .C2(n18515), .A(n18497), .B(n18496), .ZN(
        P3_U2924) );
  AOI22_X1 U21670 ( .A1(n18699), .A2(n18534), .B1(n18697), .B2(n18511), .ZN(
        n18499) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18512), .B1(
        n18698), .B2(n18510), .ZN(n18498) );
  OAI211_X1 U21672 ( .C1(n18702), .C2(n18515), .A(n18499), .B(n18498), .ZN(
        P3_U2925) );
  AOI22_X1 U21673 ( .A1(n18705), .A2(n18510), .B1(n18703), .B2(n18511), .ZN(
        n18501) );
  AOI22_X1 U21674 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18512), .B1(
        n18704), .B2(n18534), .ZN(n18500) );
  OAI211_X1 U21675 ( .C1(n18708), .C2(n18515), .A(n18501), .B(n18500), .ZN(
        P3_U2926) );
  AOI22_X1 U21676 ( .A1(n18710), .A2(n18534), .B1(n18709), .B2(n18511), .ZN(
        n18503) );
  AOI22_X1 U21677 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18512), .B1(
        n18711), .B2(n18510), .ZN(n18502) );
  OAI211_X1 U21678 ( .C1(n18714), .C2(n18515), .A(n18503), .B(n18502), .ZN(
        P3_U2927) );
  AOI22_X1 U21679 ( .A1(n18716), .A2(n18534), .B1(n18715), .B2(n18511), .ZN(
        n18505) );
  AOI22_X1 U21680 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18512), .B1(
        n18717), .B2(n18510), .ZN(n18504) );
  OAI211_X1 U21681 ( .C1(n18720), .C2(n18515), .A(n18505), .B(n18504), .ZN(
        P3_U2928) );
  AOI22_X1 U21682 ( .A1(n18723), .A2(n18510), .B1(n18721), .B2(n18511), .ZN(
        n18507) );
  AOI22_X1 U21683 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18512), .B1(
        n18722), .B2(n18534), .ZN(n18506) );
  OAI211_X1 U21684 ( .C1(n18726), .C2(n18515), .A(n18507), .B(n18506), .ZN(
        P3_U2929) );
  AOI22_X1 U21685 ( .A1(n18728), .A2(n18510), .B1(n18727), .B2(n18511), .ZN(
        n18509) );
  AOI22_X1 U21686 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18512), .B1(
        n18729), .B2(n18534), .ZN(n18508) );
  OAI211_X1 U21687 ( .C1(n18732), .C2(n18515), .A(n18509), .B(n18508), .ZN(
        P3_U2930) );
  AOI22_X1 U21688 ( .A1(n18736), .A2(n18511), .B1(n18734), .B2(n18510), .ZN(
        n18514) );
  AOI22_X1 U21689 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18512), .B1(
        n18737), .B2(n18534), .ZN(n18513) );
  OAI211_X1 U21690 ( .C1(n18742), .C2(n18515), .A(n18514), .B(n18513), .ZN(
        P3_U2931) );
  INV_X1 U21691 ( .A(n18585), .ZN(n18610) );
  NOR2_X2 U21692 ( .A1(n18794), .A2(n18610), .ZN(n18601) );
  INV_X1 U21693 ( .A(n18601), .ZN(n18538) );
  NOR2_X1 U21694 ( .A1(n18581), .A2(n18601), .ZN(n18563) );
  NOR2_X1 U21695 ( .A1(n18819), .A2(n18563), .ZN(n18533) );
  AOI22_X1 U21696 ( .A1(n18693), .A2(n18557), .B1(n18687), .B2(n18533), .ZN(
        n18520) );
  OAI21_X1 U21697 ( .B1(n18516), .B2(n18611), .A(n18563), .ZN(n18517) );
  OAI211_X1 U21698 ( .C1(n18601), .C2(n18935), .A(n18518), .B(n18517), .ZN(
        n18535) );
  AOI22_X1 U21699 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18535), .B1(
        n18688), .B2(n18534), .ZN(n18519) );
  OAI211_X1 U21700 ( .C1(n18696), .C2(n18538), .A(n18520), .B(n18519), .ZN(
        P3_U2932) );
  AOI22_X1 U21701 ( .A1(n18698), .A2(n18534), .B1(n18697), .B2(n18533), .ZN(
        n18522) );
  AOI22_X1 U21702 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18535), .B1(
        n18699), .B2(n18557), .ZN(n18521) );
  OAI211_X1 U21703 ( .C1(n18702), .C2(n18538), .A(n18522), .B(n18521), .ZN(
        P3_U2933) );
  AOI22_X1 U21704 ( .A1(n18705), .A2(n18534), .B1(n18703), .B2(n18533), .ZN(
        n18524) );
  AOI22_X1 U21705 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18535), .B1(
        n18704), .B2(n18557), .ZN(n18523) );
  OAI211_X1 U21706 ( .C1(n18708), .C2(n18538), .A(n18524), .B(n18523), .ZN(
        P3_U2934) );
  AOI22_X1 U21707 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18535), .B1(
        n18709), .B2(n18533), .ZN(n18526) );
  AOI22_X1 U21708 ( .A1(n18710), .A2(n18557), .B1(n18711), .B2(n18534), .ZN(
        n18525) );
  OAI211_X1 U21709 ( .C1(n18714), .C2(n18538), .A(n18526), .B(n18525), .ZN(
        P3_U2935) );
  AOI22_X1 U21710 ( .A1(n18717), .A2(n18534), .B1(n18715), .B2(n18533), .ZN(
        n18528) );
  AOI22_X1 U21711 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18535), .B1(
        n18716), .B2(n18557), .ZN(n18527) );
  OAI211_X1 U21712 ( .C1(n18720), .C2(n18538), .A(n18528), .B(n18527), .ZN(
        P3_U2936) );
  AOI22_X1 U21713 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18535), .B1(
        n18721), .B2(n18533), .ZN(n18530) );
  AOI22_X1 U21714 ( .A1(n18722), .A2(n18557), .B1(n18723), .B2(n18534), .ZN(
        n18529) );
  OAI211_X1 U21715 ( .C1(n18726), .C2(n18538), .A(n18530), .B(n18529), .ZN(
        P3_U2937) );
  AOI22_X1 U21716 ( .A1(n18728), .A2(n18534), .B1(n18727), .B2(n18533), .ZN(
        n18532) );
  AOI22_X1 U21717 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18535), .B1(
        n18729), .B2(n18557), .ZN(n18531) );
  OAI211_X1 U21718 ( .C1(n18732), .C2(n18538), .A(n18532), .B(n18531), .ZN(
        P3_U2938) );
  AOI22_X1 U21719 ( .A1(n18737), .A2(n18557), .B1(n18736), .B2(n18533), .ZN(
        n18537) );
  AOI22_X1 U21720 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18535), .B1(
        n18734), .B2(n18534), .ZN(n18536) );
  OAI211_X1 U21721 ( .C1(n18742), .C2(n18538), .A(n18537), .B(n18536), .ZN(
        P3_U2939) );
  NAND2_X1 U21722 ( .A1(n18585), .A2(n18539), .ZN(n18586) );
  NOR2_X1 U21723 ( .A1(n18610), .A2(n18540), .ZN(n18558) );
  AOI22_X1 U21724 ( .A1(n18693), .A2(n18581), .B1(n18687), .B2(n18558), .ZN(
        n18544) );
  NOR2_X1 U21725 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18541), .ZN(
        n18542) );
  AOI22_X1 U21726 ( .A1(n18692), .A2(n18542), .B1(n18585), .B2(n18637), .ZN(
        n18559) );
  AOI22_X1 U21727 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18559), .B1(
        n18688), .B2(n18557), .ZN(n18543) );
  OAI211_X1 U21728 ( .C1(n18696), .C2(n18586), .A(n18544), .B(n18543), .ZN(
        P3_U2940) );
  AOI22_X1 U21729 ( .A1(n18699), .A2(n18581), .B1(n18697), .B2(n18558), .ZN(
        n18546) );
  AOI22_X1 U21730 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18559), .B1(
        n18698), .B2(n18557), .ZN(n18545) );
  OAI211_X1 U21731 ( .C1(n18702), .C2(n18586), .A(n18546), .B(n18545), .ZN(
        P3_U2941) );
  AOI22_X1 U21732 ( .A1(n18704), .A2(n18581), .B1(n18703), .B2(n18558), .ZN(
        n18548) );
  AOI22_X1 U21733 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18559), .B1(
        n18705), .B2(n18557), .ZN(n18547) );
  OAI211_X1 U21734 ( .C1(n18708), .C2(n18586), .A(n18548), .B(n18547), .ZN(
        P3_U2942) );
  AOI22_X1 U21735 ( .A1(n18711), .A2(n18557), .B1(n18709), .B2(n18558), .ZN(
        n18550) );
  AOI22_X1 U21736 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18559), .B1(
        n18710), .B2(n18581), .ZN(n18549) );
  OAI211_X1 U21737 ( .C1(n18714), .C2(n18586), .A(n18550), .B(n18549), .ZN(
        P3_U2943) );
  AOI22_X1 U21738 ( .A1(n18716), .A2(n18581), .B1(n18715), .B2(n18558), .ZN(
        n18552) );
  AOI22_X1 U21739 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18559), .B1(
        n18717), .B2(n18557), .ZN(n18551) );
  OAI211_X1 U21740 ( .C1(n18720), .C2(n18586), .A(n18552), .B(n18551), .ZN(
        P3_U2944) );
  AOI22_X1 U21741 ( .A1(n18722), .A2(n18581), .B1(n18721), .B2(n18558), .ZN(
        n18554) );
  AOI22_X1 U21742 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18559), .B1(
        n18723), .B2(n18557), .ZN(n18553) );
  OAI211_X1 U21743 ( .C1(n18726), .C2(n18586), .A(n18554), .B(n18553), .ZN(
        P3_U2945) );
  AOI22_X1 U21744 ( .A1(n18729), .A2(n18581), .B1(n18727), .B2(n18558), .ZN(
        n18556) );
  AOI22_X1 U21745 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18559), .B1(
        n18728), .B2(n18557), .ZN(n18555) );
  OAI211_X1 U21746 ( .C1(n18732), .C2(n18586), .A(n18556), .B(n18555), .ZN(
        P3_U2946) );
  AOI22_X1 U21747 ( .A1(n18736), .A2(n18558), .B1(n18734), .B2(n18557), .ZN(
        n18561) );
  AOI22_X1 U21748 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18559), .B1(
        n18737), .B2(n18581), .ZN(n18560) );
  OAI211_X1 U21749 ( .C1(n18742), .C2(n18586), .A(n18561), .B(n18560), .ZN(
        P3_U2947) );
  NAND2_X1 U21750 ( .A1(n18585), .A2(n18562), .ZN(n18608) );
  AOI21_X1 U21751 ( .B1(n18586), .B2(n18608), .A(n18819), .ZN(n18579) );
  AOI22_X1 U21752 ( .A1(n18688), .A2(n18581), .B1(n18687), .B2(n18579), .ZN(
        n18566) );
  OAI211_X1 U21753 ( .C1(n18563), .C2(n18611), .A(n18586), .B(n18608), .ZN(
        n18564) );
  NAND2_X1 U21754 ( .A1(n18661), .A2(n18564), .ZN(n18580) );
  AOI22_X1 U21755 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18580), .B1(
        n18693), .B2(n18601), .ZN(n18565) );
  OAI211_X1 U21756 ( .C1(n18696), .C2(n18608), .A(n18566), .B(n18565), .ZN(
        P3_U2948) );
  AOI22_X1 U21757 ( .A1(n18699), .A2(n18601), .B1(n18697), .B2(n18579), .ZN(
        n18568) );
  AOI22_X1 U21758 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18580), .B1(
        n18698), .B2(n18581), .ZN(n18567) );
  OAI211_X1 U21759 ( .C1(n18702), .C2(n18608), .A(n18568), .B(n18567), .ZN(
        P3_U2949) );
  AOI22_X1 U21760 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18580), .B1(
        n18703), .B2(n18579), .ZN(n18570) );
  AOI22_X1 U21761 ( .A1(n18705), .A2(n18581), .B1(n18704), .B2(n18601), .ZN(
        n18569) );
  OAI211_X1 U21762 ( .C1(n18708), .C2(n18608), .A(n18570), .B(n18569), .ZN(
        P3_U2950) );
  AOI22_X1 U21763 ( .A1(n18711), .A2(n18581), .B1(n18709), .B2(n18579), .ZN(
        n18572) );
  AOI22_X1 U21764 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18580), .B1(
        n18710), .B2(n18601), .ZN(n18571) );
  OAI211_X1 U21765 ( .C1(n18714), .C2(n18608), .A(n18572), .B(n18571), .ZN(
        P3_U2951) );
  AOI22_X1 U21766 ( .A1(n18717), .A2(n18581), .B1(n18715), .B2(n18579), .ZN(
        n18574) );
  AOI22_X1 U21767 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18580), .B1(
        n18716), .B2(n18601), .ZN(n18573) );
  OAI211_X1 U21768 ( .C1(n18720), .C2(n18608), .A(n18574), .B(n18573), .ZN(
        P3_U2952) );
  AOI22_X1 U21769 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18580), .B1(
        n18721), .B2(n18579), .ZN(n18576) );
  AOI22_X1 U21770 ( .A1(n18722), .A2(n18601), .B1(n18723), .B2(n18581), .ZN(
        n18575) );
  OAI211_X1 U21771 ( .C1(n18726), .C2(n18608), .A(n18576), .B(n18575), .ZN(
        P3_U2953) );
  AOI22_X1 U21772 ( .A1(n18729), .A2(n18601), .B1(n18727), .B2(n18579), .ZN(
        n18578) );
  AOI22_X1 U21773 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18580), .B1(
        n18728), .B2(n18581), .ZN(n18577) );
  OAI211_X1 U21774 ( .C1(n18732), .C2(n18608), .A(n18578), .B(n18577), .ZN(
        P3_U2954) );
  AOI22_X1 U21775 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18580), .B1(
        n18736), .B2(n18579), .ZN(n18583) );
  AOI22_X1 U21776 ( .A1(n18737), .A2(n18601), .B1(n18734), .B2(n18581), .ZN(
        n18582) );
  OAI211_X1 U21777 ( .C1(n18742), .C2(n18608), .A(n18583), .B(n18582), .ZN(
        P3_U2955) );
  NOR2_X2 U21778 ( .A1(n18792), .A2(n18610), .ZN(n18679) );
  INV_X1 U21779 ( .A(n18679), .ZN(n18606) );
  NOR2_X1 U21780 ( .A1(n18793), .A2(n18610), .ZN(n18639) );
  AND2_X1 U21781 ( .A1(n18686), .A2(n18639), .ZN(n18602) );
  AOI22_X1 U21782 ( .A1(n18688), .A2(n18601), .B1(n18687), .B2(n18602), .ZN(
        n18588) );
  INV_X1 U21783 ( .A(n18584), .ZN(n18690) );
  OAI211_X1 U21784 ( .C1(n18692), .C2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n18690), .B(n18585), .ZN(n18603) );
  INV_X1 U21785 ( .A(n18586), .ZN(n18632) );
  AOI22_X1 U21786 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18603), .B1(
        n18693), .B2(n18632), .ZN(n18587) );
  OAI211_X1 U21787 ( .C1(n18696), .C2(n18606), .A(n18588), .B(n18587), .ZN(
        P3_U2956) );
  AOI22_X1 U21788 ( .A1(n18699), .A2(n18632), .B1(n18697), .B2(n18602), .ZN(
        n18590) );
  AOI22_X1 U21789 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18603), .B1(
        n18698), .B2(n18601), .ZN(n18589) );
  OAI211_X1 U21790 ( .C1(n18702), .C2(n18606), .A(n18590), .B(n18589), .ZN(
        P3_U2957) );
  AOI22_X1 U21791 ( .A1(n18704), .A2(n18632), .B1(n18703), .B2(n18602), .ZN(
        n18592) );
  AOI22_X1 U21792 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18603), .B1(
        n18705), .B2(n18601), .ZN(n18591) );
  OAI211_X1 U21793 ( .C1(n18708), .C2(n18606), .A(n18592), .B(n18591), .ZN(
        P3_U2958) );
  AOI22_X1 U21794 ( .A1(n18711), .A2(n18601), .B1(n18709), .B2(n18602), .ZN(
        n18594) );
  AOI22_X1 U21795 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18603), .B1(
        n18710), .B2(n18632), .ZN(n18593) );
  OAI211_X1 U21796 ( .C1(n18714), .C2(n18606), .A(n18594), .B(n18593), .ZN(
        P3_U2959) );
  AOI22_X1 U21797 ( .A1(n18716), .A2(n18632), .B1(n18715), .B2(n18602), .ZN(
        n18596) );
  AOI22_X1 U21798 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18603), .B1(
        n18717), .B2(n18601), .ZN(n18595) );
  OAI211_X1 U21799 ( .C1(n18720), .C2(n18606), .A(n18596), .B(n18595), .ZN(
        P3_U2960) );
  AOI22_X1 U21800 ( .A1(n18722), .A2(n18632), .B1(n18721), .B2(n18602), .ZN(
        n18598) );
  AOI22_X1 U21801 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18603), .B1(
        n18723), .B2(n18601), .ZN(n18597) );
  OAI211_X1 U21802 ( .C1(n18726), .C2(n18606), .A(n18598), .B(n18597), .ZN(
        P3_U2961) );
  AOI22_X1 U21803 ( .A1(n18729), .A2(n18632), .B1(n18727), .B2(n18602), .ZN(
        n18600) );
  AOI22_X1 U21804 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18603), .B1(
        n18728), .B2(n18601), .ZN(n18599) );
  OAI211_X1 U21805 ( .C1(n18732), .C2(n18606), .A(n18600), .B(n18599), .ZN(
        P3_U2962) );
  AOI22_X1 U21806 ( .A1(n18736), .A2(n18602), .B1(n18734), .B2(n18601), .ZN(
        n18605) );
  AOI22_X1 U21807 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18603), .B1(
        n18737), .B2(n18632), .ZN(n18604) );
  OAI211_X1 U21808 ( .C1(n18742), .C2(n18606), .A(n18605), .B(n18604), .ZN(
        P3_U2963) );
  INV_X1 U21809 ( .A(n18636), .ZN(n18691) );
  NAND2_X1 U21810 ( .A1(n18691), .A2(n18607), .ZN(n18635) );
  INV_X1 U21811 ( .A(n18608), .ZN(n18654) );
  INV_X1 U21812 ( .A(n18635), .ZN(n18733) );
  NOR2_X1 U21813 ( .A1(n18679), .A2(n18733), .ZN(n18609) );
  NOR2_X1 U21814 ( .A1(n18819), .A2(n18609), .ZN(n18630) );
  AOI22_X1 U21815 ( .A1(n18693), .A2(n18654), .B1(n18687), .B2(n18630), .ZN(
        n18617) );
  INV_X1 U21816 ( .A(n18609), .ZN(n18662) );
  NOR2_X1 U21817 ( .A1(n18611), .A2(n18610), .ZN(n18615) );
  AOI21_X1 U21818 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18635), .A(n18612), 
        .ZN(n18613) );
  OAI221_X1 U21819 ( .B1(n18662), .B2(n18615), .C1(n18662), .C2(n18614), .A(
        n18613), .ZN(n18631) );
  AOI22_X1 U21820 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18631), .B1(
        n18688), .B2(n18632), .ZN(n18616) );
  OAI211_X1 U21821 ( .C1(n18696), .C2(n18635), .A(n18617), .B(n18616), .ZN(
        P3_U2964) );
  AOI22_X1 U21822 ( .A1(n18699), .A2(n18654), .B1(n18697), .B2(n18630), .ZN(
        n18619) );
  AOI22_X1 U21823 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18631), .B1(
        n18698), .B2(n18632), .ZN(n18618) );
  OAI211_X1 U21824 ( .C1(n18702), .C2(n18635), .A(n18619), .B(n18618), .ZN(
        P3_U2965) );
  AOI22_X1 U21825 ( .A1(n18705), .A2(n18632), .B1(n18703), .B2(n18630), .ZN(
        n18621) );
  AOI22_X1 U21826 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18631), .B1(
        n18704), .B2(n18654), .ZN(n18620) );
  OAI211_X1 U21827 ( .C1(n18708), .C2(n18635), .A(n18621), .B(n18620), .ZN(
        P3_U2966) );
  AOI22_X1 U21828 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18631), .B1(
        n18709), .B2(n18630), .ZN(n18623) );
  AOI22_X1 U21829 ( .A1(n18710), .A2(n18654), .B1(n18711), .B2(n18632), .ZN(
        n18622) );
  OAI211_X1 U21830 ( .C1(n18714), .C2(n18635), .A(n18623), .B(n18622), .ZN(
        P3_U2967) );
  AOI22_X1 U21831 ( .A1(n18717), .A2(n18632), .B1(n18715), .B2(n18630), .ZN(
        n18625) );
  AOI22_X1 U21832 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18631), .B1(
        n18716), .B2(n18654), .ZN(n18624) );
  OAI211_X1 U21833 ( .C1(n18720), .C2(n18635), .A(n18625), .B(n18624), .ZN(
        P3_U2968) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18631), .B1(
        n18721), .B2(n18630), .ZN(n18627) );
  AOI22_X1 U21835 ( .A1(n18722), .A2(n18654), .B1(n18723), .B2(n18632), .ZN(
        n18626) );
  OAI211_X1 U21836 ( .C1(n18726), .C2(n18635), .A(n18627), .B(n18626), .ZN(
        P3_U2969) );
  AOI22_X1 U21837 ( .A1(n18729), .A2(n18654), .B1(n18727), .B2(n18630), .ZN(
        n18629) );
  AOI22_X1 U21838 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18631), .B1(
        n18728), .B2(n18632), .ZN(n18628) );
  OAI211_X1 U21839 ( .C1(n18732), .C2(n18635), .A(n18629), .B(n18628), .ZN(
        P3_U2970) );
  AOI22_X1 U21840 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18631), .B1(
        n18736), .B2(n18630), .ZN(n18634) );
  AOI22_X1 U21841 ( .A1(n18737), .A2(n18654), .B1(n18734), .B2(n18632), .ZN(
        n18633) );
  OAI211_X1 U21842 ( .C1(n18742), .C2(n18635), .A(n18634), .B(n18633), .ZN(
        P3_U2971) );
  INV_X1 U21843 ( .A(n18738), .ZN(n18659) );
  NOR2_X1 U21844 ( .A1(n18819), .A2(n18636), .ZN(n18655) );
  AOI22_X1 U21845 ( .A1(n18693), .A2(n18679), .B1(n18687), .B2(n18655), .ZN(
        n18641) );
  AOI22_X1 U21846 ( .A1(n18692), .A2(n18639), .B1(n18638), .B2(n18637), .ZN(
        n18656) );
  AOI22_X1 U21847 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18656), .B1(
        n18688), .B2(n18654), .ZN(n18640) );
  OAI211_X1 U21848 ( .C1(n18659), .C2(n18696), .A(n18641), .B(n18640), .ZN(
        P3_U2972) );
  AOI22_X1 U21849 ( .A1(n18698), .A2(n18654), .B1(n18697), .B2(n18655), .ZN(
        n18643) );
  AOI22_X1 U21850 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18656), .B1(
        n18699), .B2(n18679), .ZN(n18642) );
  OAI211_X1 U21851 ( .C1(n18659), .C2(n18702), .A(n18643), .B(n18642), .ZN(
        P3_U2973) );
  AOI22_X1 U21852 ( .A1(n18705), .A2(n18654), .B1(n18703), .B2(n18655), .ZN(
        n18645) );
  AOI22_X1 U21853 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18656), .B1(
        n18704), .B2(n18679), .ZN(n18644) );
  OAI211_X1 U21854 ( .C1(n18659), .C2(n18708), .A(n18645), .B(n18644), .ZN(
        P3_U2974) );
  AOI22_X1 U21855 ( .A1(n18710), .A2(n18679), .B1(n18709), .B2(n18655), .ZN(
        n18647) );
  AOI22_X1 U21856 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18656), .B1(
        n18711), .B2(n18654), .ZN(n18646) );
  OAI211_X1 U21857 ( .C1(n18659), .C2(n18714), .A(n18647), .B(n18646), .ZN(
        P3_U2975) );
  AOI22_X1 U21858 ( .A1(n18716), .A2(n18679), .B1(n18715), .B2(n18655), .ZN(
        n18649) );
  AOI22_X1 U21859 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18656), .B1(
        n18717), .B2(n18654), .ZN(n18648) );
  OAI211_X1 U21860 ( .C1(n18659), .C2(n18720), .A(n18649), .B(n18648), .ZN(
        P3_U2976) );
  AOI22_X1 U21861 ( .A1(n18722), .A2(n18679), .B1(n18721), .B2(n18655), .ZN(
        n18651) );
  AOI22_X1 U21862 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18656), .B1(
        n18723), .B2(n18654), .ZN(n18650) );
  OAI211_X1 U21863 ( .C1(n18659), .C2(n18726), .A(n18651), .B(n18650), .ZN(
        P3_U2977) );
  AOI22_X1 U21864 ( .A1(n18729), .A2(n18679), .B1(n18727), .B2(n18655), .ZN(
        n18653) );
  AOI22_X1 U21865 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18656), .B1(
        n18728), .B2(n18654), .ZN(n18652) );
  OAI211_X1 U21866 ( .C1(n18659), .C2(n18732), .A(n18653), .B(n18652), .ZN(
        P3_U2978) );
  AOI22_X1 U21867 ( .A1(n18736), .A2(n18655), .B1(n18734), .B2(n18654), .ZN(
        n18658) );
  AOI22_X1 U21868 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18656), .B1(
        n18737), .B2(n18679), .ZN(n18657) );
  OAI211_X1 U21869 ( .C1(n18659), .C2(n18742), .A(n18658), .B(n18657), .ZN(
        P3_U2979) );
  NOR2_X1 U21870 ( .A1(n18819), .A2(n18660), .ZN(n18680) );
  AOI22_X1 U21871 ( .A1(n18688), .A2(n18679), .B1(n18687), .B2(n18680), .ZN(
        n18666) );
  INV_X1 U21872 ( .A(n18660), .ZN(n18664) );
  OAI221_X1 U21873 ( .B1(n18664), .B2(n18663), .C1(n18664), .C2(n18662), .A(
        n18661), .ZN(n18681) );
  AOI22_X1 U21874 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18681), .B1(
        n18693), .B2(n18733), .ZN(n18665) );
  OAI211_X1 U21875 ( .C1(n18696), .C2(n18684), .A(n18666), .B(n18665), .ZN(
        P3_U2980) );
  AOI22_X1 U21876 ( .A1(n18699), .A2(n18733), .B1(n18697), .B2(n18680), .ZN(
        n18668) );
  AOI22_X1 U21877 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18681), .B1(
        n18698), .B2(n18679), .ZN(n18667) );
  OAI211_X1 U21878 ( .C1(n18684), .C2(n18702), .A(n18668), .B(n18667), .ZN(
        P3_U2981) );
  AOI22_X1 U21879 ( .A1(n18705), .A2(n18679), .B1(n18703), .B2(n18680), .ZN(
        n18670) );
  AOI22_X1 U21880 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18681), .B1(
        n18704), .B2(n18733), .ZN(n18669) );
  OAI211_X1 U21881 ( .C1(n18684), .C2(n18708), .A(n18670), .B(n18669), .ZN(
        P3_U2982) );
  AOI22_X1 U21882 ( .A1(n18710), .A2(n18733), .B1(n18709), .B2(n18680), .ZN(
        n18672) );
  AOI22_X1 U21883 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18681), .B1(
        n18711), .B2(n18679), .ZN(n18671) );
  OAI211_X1 U21884 ( .C1(n18684), .C2(n18714), .A(n18672), .B(n18671), .ZN(
        P3_U2983) );
  AOI22_X1 U21885 ( .A1(n18717), .A2(n18679), .B1(n18715), .B2(n18680), .ZN(
        n18674) );
  AOI22_X1 U21886 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18681), .B1(
        n18716), .B2(n18733), .ZN(n18673) );
  OAI211_X1 U21887 ( .C1(n18684), .C2(n18720), .A(n18674), .B(n18673), .ZN(
        P3_U2984) );
  AOI22_X1 U21888 ( .A1(n18722), .A2(n18733), .B1(n18721), .B2(n18680), .ZN(
        n18676) );
  AOI22_X1 U21889 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18681), .B1(
        n18723), .B2(n18679), .ZN(n18675) );
  OAI211_X1 U21890 ( .C1(n18684), .C2(n18726), .A(n18676), .B(n18675), .ZN(
        P3_U2985) );
  AOI22_X1 U21891 ( .A1(n18729), .A2(n18733), .B1(n18727), .B2(n18680), .ZN(
        n18678) );
  AOI22_X1 U21892 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18681), .B1(
        n18728), .B2(n18679), .ZN(n18677) );
  OAI211_X1 U21893 ( .C1(n18684), .C2(n18732), .A(n18678), .B(n18677), .ZN(
        P3_U2986) );
  AOI22_X1 U21894 ( .A1(n18736), .A2(n18680), .B1(n18734), .B2(n18679), .ZN(
        n18683) );
  AOI22_X1 U21895 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18681), .B1(
        n18737), .B2(n18733), .ZN(n18682) );
  OAI211_X1 U21896 ( .C1(n18684), .C2(n18742), .A(n18683), .B(n18682), .ZN(
        P3_U2987) );
  INV_X1 U21897 ( .A(n18685), .ZN(n18743) );
  AND2_X1 U21898 ( .A1(n18686), .A2(n18689), .ZN(n18735) );
  AOI22_X1 U21899 ( .A1(n18688), .A2(n18733), .B1(n18687), .B2(n18735), .ZN(
        n18695) );
  AOI22_X1 U21900 ( .A1(n18692), .A2(n18691), .B1(n18690), .B2(n18689), .ZN(
        n18739) );
  AOI22_X1 U21901 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18739), .B1(
        n18738), .B2(n18693), .ZN(n18694) );
  OAI211_X1 U21902 ( .C1(n18743), .C2(n18696), .A(n18695), .B(n18694), .ZN(
        P3_U2988) );
  AOI22_X1 U21903 ( .A1(n18698), .A2(n18733), .B1(n18697), .B2(n18735), .ZN(
        n18701) );
  AOI22_X1 U21904 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18739), .B1(
        n18738), .B2(n18699), .ZN(n18700) );
  OAI211_X1 U21905 ( .C1(n18743), .C2(n18702), .A(n18701), .B(n18700), .ZN(
        P3_U2989) );
  AOI22_X1 U21906 ( .A1(n18738), .A2(n18704), .B1(n18703), .B2(n18735), .ZN(
        n18707) );
  AOI22_X1 U21907 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18739), .B1(
        n18705), .B2(n18733), .ZN(n18706) );
  OAI211_X1 U21908 ( .C1(n18743), .C2(n18708), .A(n18707), .B(n18706), .ZN(
        P3_U2990) );
  AOI22_X1 U21909 ( .A1(n18738), .A2(n18710), .B1(n18709), .B2(n18735), .ZN(
        n18713) );
  AOI22_X1 U21910 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18739), .B1(
        n18711), .B2(n18733), .ZN(n18712) );
  OAI211_X1 U21911 ( .C1(n18743), .C2(n18714), .A(n18713), .B(n18712), .ZN(
        P3_U2991) );
  AOI22_X1 U21912 ( .A1(n18738), .A2(n18716), .B1(n18715), .B2(n18735), .ZN(
        n18719) );
  AOI22_X1 U21913 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18739), .B1(
        n18717), .B2(n18733), .ZN(n18718) );
  OAI211_X1 U21914 ( .C1(n18743), .C2(n18720), .A(n18719), .B(n18718), .ZN(
        P3_U2992) );
  AOI22_X1 U21915 ( .A1(n18738), .A2(n18722), .B1(n18721), .B2(n18735), .ZN(
        n18725) );
  AOI22_X1 U21916 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18739), .B1(
        n18723), .B2(n18733), .ZN(n18724) );
  OAI211_X1 U21917 ( .C1(n18743), .C2(n18726), .A(n18725), .B(n18724), .ZN(
        P3_U2993) );
  AOI22_X1 U21918 ( .A1(n18728), .A2(n18733), .B1(n18727), .B2(n18735), .ZN(
        n18731) );
  AOI22_X1 U21919 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18739), .B1(
        n18738), .B2(n18729), .ZN(n18730) );
  OAI211_X1 U21920 ( .C1(n18743), .C2(n18732), .A(n18731), .B(n18730), .ZN(
        P3_U2994) );
  AOI22_X1 U21921 ( .A1(n18736), .A2(n18735), .B1(n18734), .B2(n18733), .ZN(
        n18741) );
  AOI22_X1 U21922 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18739), .B1(
        n18738), .B2(n18737), .ZN(n18740) );
  OAI211_X1 U21923 ( .C1(n18743), .C2(n18742), .A(n18741), .B(n18740), .ZN(
        P3_U2995) );
  NOR2_X1 U21924 ( .A1(n18785), .A2(n18744), .ZN(n18746) );
  OAI222_X1 U21925 ( .A1(n18750), .A2(n18749), .B1(n18748), .B2(n18747), .C1(
        n18746), .C2(n18745), .ZN(n18952) );
  OAI21_X1 U21926 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(P3_MORE_REG_SCAN_IN), .A(
        n18751), .ZN(n18752) );
  OAI211_X1 U21927 ( .C1(n18754), .C2(n18786), .A(n18753), .B(n18752), .ZN(
        n18806) );
  OAI21_X1 U21928 ( .B1(n18940), .B2(n18755), .A(n18767), .ZN(n18777) );
  NOR2_X1 U21929 ( .A1(n18777), .A2(n18756), .ZN(n18790) );
  OAI22_X1 U21930 ( .A1(n18758), .A2(n18790), .B1(n18757), .B2(n18768), .ZN(
        n18759) );
  INV_X1 U21931 ( .A(n18759), .ZN(n18760) );
  NOR2_X1 U21932 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18760), .ZN(
        n18917) );
  INV_X1 U21933 ( .A(n18761), .ZN(n18763) );
  OAI21_X1 U21934 ( .B1(n18764), .B2(n18763), .A(n18762), .ZN(n18776) );
  AOI21_X1 U21935 ( .B1(n18767), .B2(n18766), .A(n18765), .ZN(n18769) );
  AOI211_X1 U21936 ( .C1(n18770), .C2(n18776), .A(n18769), .B(n18768), .ZN(
        n18918) );
  NAND2_X1 U21937 ( .A1(n18786), .A2(n18918), .ZN(n18771) );
  AOI22_X1 U21938 ( .A1(n18786), .A2(n18917), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18771), .ZN(n18804) );
  INV_X1 U21939 ( .A(n18931), .ZN(n18784) );
  AOI21_X1 U21940 ( .B1(n18778), .B2(n18773), .A(n18772), .ZN(n18783) );
  INV_X1 U21941 ( .A(n18773), .ZN(n18775) );
  AOI22_X1 U21942 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18776), .B1(
        n18775), .B2(n18774), .ZN(n18780) );
  INV_X1 U21943 ( .A(n18777), .ZN(n18779) );
  OAI22_X1 U21944 ( .A1(n18781), .A2(n18780), .B1(n18779), .B2(n18778), .ZN(
        n18782) );
  AOI211_X1 U21945 ( .C1(n18785), .C2(n18784), .A(n18783), .B(n18782), .ZN(
        n18929) );
  AOI22_X1 U21946 ( .A1(n18796), .A2(n18933), .B1(n18929), .B2(n18786), .ZN(
        n18800) );
  NOR2_X1 U21947 ( .A1(n18788), .A2(n18787), .ZN(n18791) );
  AOI22_X1 U21948 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18789), .B1(
        n18791), .B2(n18940), .ZN(n18934) );
  AOI222_X1 U21949 ( .A1(n18934), .A2(n21186), .B1(n18934), .B2(n18793), .C1(
        n21186), .C2(n18792), .ZN(n18795) );
  OAI21_X1 U21950 ( .B1(n18796), .B2(n18795), .A(n18794), .ZN(n18799) );
  AND2_X1 U21951 ( .A1(n18800), .A2(n18799), .ZN(n18797) );
  OAI221_X1 U21952 ( .B1(n18800), .B2(n18799), .C1(n18798), .C2(n18797), .A(
        n18801), .ZN(n18803) );
  AOI21_X1 U21953 ( .B1(n18801), .B2(n20929), .A(n18800), .ZN(n18802) );
  AOI222_X1 U21954 ( .A1(n18804), .A2(n18803), .B1(n18804), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18803), .C2(n18802), .ZN(
        n18805) );
  NOR4_X1 U21955 ( .A1(n18807), .A2(n18952), .A3(n18806), .A4(n18805), .ZN(
        n18818) );
  NOR2_X1 U21956 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18965) );
  AOI22_X1 U21957 ( .A1(n21184), .A2(n18965), .B1(n18960), .B2(n18954), .ZN(
        n18808) );
  INV_X1 U21958 ( .A(n18808), .ZN(n18813) );
  OAI211_X1 U21959 ( .C1(n18810), .C2(n18809), .A(n18957), .B(n18818), .ZN(
        n18914) );
  OAI21_X1 U21960 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18953), .A(n18914), 
        .ZN(n18820) );
  NOR2_X1 U21961 ( .A1(n18811), .A2(n18820), .ZN(n18812) );
  MUX2_X1 U21962 ( .A(n18813), .B(n18812), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18816) );
  INV_X1 U21963 ( .A(n18814), .ZN(n18815) );
  OAI211_X1 U21964 ( .C1(n18818), .C2(n18817), .A(n18816), .B(n18815), .ZN(
        P3_U2996) );
  NAND2_X1 U21965 ( .A1(n18960), .A2(n18954), .ZN(n18823) );
  NAND4_X1 U21966 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(n18960), .A4(n18971), .ZN(n18825) );
  OR3_X1 U21967 ( .A1(n18821), .A2(n18820), .A3(n18819), .ZN(n18822) );
  NAND4_X1 U21968 ( .A1(n18824), .A2(n18823), .A3(n18825), .A4(n18822), .ZN(
        P3_U2997) );
  INV_X1 U21969 ( .A(n18965), .ZN(n18827) );
  AND4_X1 U21970 ( .A1(n18827), .A2(n18826), .A3(n18825), .A4(n18913), .ZN(
        P3_U2998) );
  AND2_X1 U21971 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18908), .ZN(
        P3_U2999) );
  AND2_X1 U21972 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18908), .ZN(
        P3_U3000) );
  AND2_X1 U21973 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18908), .ZN(
        P3_U3001) );
  AND2_X1 U21974 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18908), .ZN(
        P3_U3002) );
  AND2_X1 U21975 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18908), .ZN(
        P3_U3003) );
  AND2_X1 U21976 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18908), .ZN(
        P3_U3004) );
  AND2_X1 U21977 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18908), .ZN(
        P3_U3005) );
  AND2_X1 U21978 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18908), .ZN(
        P3_U3006) );
  AND2_X1 U21979 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18908), .ZN(
        P3_U3007) );
  AND2_X1 U21980 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18908), .ZN(
        P3_U3008) );
  AND2_X1 U21981 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18908), .ZN(
        P3_U3009) );
  AND2_X1 U21982 ( .A1(n18908), .A2(P3_DATAWIDTH_REG_20__SCAN_IN), .ZN(
        P3_U3010) );
  AND2_X1 U21983 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18908), .ZN(
        P3_U3011) );
  AND2_X1 U21984 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18908), .ZN(
        P3_U3012) );
  AND2_X1 U21985 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18908), .ZN(
        P3_U3013) );
  AND2_X1 U21986 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18908), .ZN(
        P3_U3014) );
  AND2_X1 U21987 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18908), .ZN(
        P3_U3015) );
  AND2_X1 U21988 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18908), .ZN(
        P3_U3016) );
  AND2_X1 U21989 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18908), .ZN(
        P3_U3017) );
  AND2_X1 U21990 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18908), .ZN(
        P3_U3018) );
  AND2_X1 U21991 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18908), .ZN(
        P3_U3019) );
  AND2_X1 U21992 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18908), .ZN(
        P3_U3020) );
  AND2_X1 U21993 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18908), .ZN(P3_U3021) );
  AND2_X1 U21994 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18908), .ZN(P3_U3022) );
  AND2_X1 U21995 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18908), .ZN(P3_U3023) );
  AND2_X1 U21996 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18908), .ZN(P3_U3024) );
  AND2_X1 U21997 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18908), .ZN(P3_U3025) );
  AND2_X1 U21998 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18908), .ZN(P3_U3026) );
  AND2_X1 U21999 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18908), .ZN(P3_U3027) );
  AND2_X1 U22000 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18908), .ZN(P3_U3028) );
  NAND2_X1 U22001 ( .A1(n18960), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18836) );
  NAND2_X1 U22002 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18836), .ZN(n18839) );
  INV_X1 U22003 ( .A(n18839), .ZN(n18831) );
  INV_X1 U22004 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18967) );
  INV_X1 U22005 ( .A(NA), .ZN(n20737) );
  OAI22_X1 U22006 ( .A1(n18828), .A2(n20743), .B1(P3_STATE_REG_0__SCAN_IN), 
        .B2(n20737), .ZN(n18829) );
  OAI21_X1 U22007 ( .B1(n18967), .B2(n18829), .A(n18969), .ZN(n18830) );
  OAI21_X1 U22008 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n18831), .A(n18830), 
        .ZN(P3_U3029) );
  NOR2_X1 U22009 ( .A1(n21159), .A2(n20743), .ZN(n18838) );
  OAI22_X1 U22010 ( .A1(n18838), .A2(n18967), .B1(n20743), .B2(n18832), .ZN(
        n18833) );
  NAND2_X1 U22011 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18833), .ZN(n18835) );
  NAND3_X1 U22012 ( .A1(n18835), .A2(n18836), .A3(n18834), .ZN(P3_U3030) );
  OAI22_X1 U22013 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18836), .ZN(n18837) );
  OAI22_X1 U22014 ( .A1(n18838), .A2(n18837), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18841) );
  OAI211_X1 U22015 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(n20737), .A(
        P3_STATE_REG_2__SCAN_IN), .B(n18839), .ZN(n18840) );
  OAI21_X1 U22016 ( .B1(n20932), .B2(n18841), .A(n18840), .ZN(P3_U3031) );
  OAI222_X1 U22017 ( .A1(n18941), .A2(n18893), .B1(n18842), .B2(n18950), .C1(
        n18843), .C2(n18896), .ZN(P3_U3032) );
  OAI222_X1 U22018 ( .A1(n18896), .A2(n21047), .B1(n18844), .B2(n18950), .C1(
        n18843), .C2(n18893), .ZN(P3_U3033) );
  OAI222_X1 U22019 ( .A1(n21047), .A2(n18893), .B1(n18845), .B2(n18950), .C1(
        n18846), .C2(n18896), .ZN(P3_U3034) );
  INV_X1 U22020 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18849) );
  OAI222_X1 U22021 ( .A1(n18896), .A2(n18849), .B1(n18847), .B2(n18950), .C1(
        n18846), .C2(n18893), .ZN(P3_U3035) );
  OAI222_X1 U22022 ( .A1(n18849), .A2(n18893), .B1(n18848), .B2(n18950), .C1(
        n18850), .C2(n18896), .ZN(P3_U3036) );
  OAI222_X1 U22023 ( .A1(n18896), .A2(n18852), .B1(n18851), .B2(n18950), .C1(
        n18850), .C2(n18893), .ZN(P3_U3037) );
  OAI222_X1 U22024 ( .A1(n18896), .A2(n18855), .B1(n18853), .B2(n18950), .C1(
        n18852), .C2(n18893), .ZN(P3_U3038) );
  OAI222_X1 U22025 ( .A1(n18855), .A2(n18893), .B1(n18854), .B2(n18950), .C1(
        n18856), .C2(n18896), .ZN(P3_U3039) );
  OAI222_X1 U22026 ( .A1(n18896), .A2(n18858), .B1(n18857), .B2(n18950), .C1(
        n18856), .C2(n18893), .ZN(P3_U3040) );
  OAI222_X1 U22027 ( .A1(n18896), .A2(n18860), .B1(n18859), .B2(n18950), .C1(
        n18858), .C2(n18893), .ZN(P3_U3041) );
  OAI222_X1 U22028 ( .A1(n18896), .A2(n21045), .B1(n18861), .B2(n18950), .C1(
        n18860), .C2(n18893), .ZN(P3_U3042) );
  OAI222_X1 U22029 ( .A1(n18896), .A2(n18863), .B1(n18862), .B2(n18950), .C1(
        n21045), .C2(n18893), .ZN(P3_U3043) );
  OAI222_X1 U22030 ( .A1(n18896), .A2(n21089), .B1(n18864), .B2(n18950), .C1(
        n18863), .C2(n18893), .ZN(P3_U3044) );
  OAI222_X1 U22031 ( .A1(n21089), .A2(n18893), .B1(n18865), .B2(n18950), .C1(
        n18866), .C2(n18896), .ZN(P3_U3045) );
  OAI222_X1 U22032 ( .A1(n18896), .A2(n18868), .B1(n18867), .B2(n18950), .C1(
        n18866), .C2(n18900), .ZN(P3_U3046) );
  OAI222_X1 U22033 ( .A1(n18896), .A2(n21129), .B1(n18869), .B2(n18950), .C1(
        n18868), .C2(n18900), .ZN(P3_U3047) );
  OAI222_X1 U22034 ( .A1(n21129), .A2(n18893), .B1(n18870), .B2(n18950), .C1(
        n18871), .C2(n18896), .ZN(P3_U3048) );
  OAI222_X1 U22035 ( .A1(n18896), .A2(n18873), .B1(n18872), .B2(n18950), .C1(
        n18871), .C2(n18900), .ZN(P3_U3049) );
  INV_X1 U22036 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18875) );
  OAI222_X1 U22037 ( .A1(n18896), .A2(n18875), .B1(n18874), .B2(n18950), .C1(
        n18873), .C2(n18900), .ZN(P3_U3050) );
  OAI222_X1 U22038 ( .A1(n18896), .A2(n18877), .B1(n18876), .B2(n18950), .C1(
        n18875), .C2(n18900), .ZN(P3_U3051) );
  INV_X1 U22039 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18879) );
  OAI222_X1 U22040 ( .A1(n18896), .A2(n18879), .B1(n18878), .B2(n18950), .C1(
        n18877), .C2(n18900), .ZN(P3_U3052) );
  OAI222_X1 U22041 ( .A1(n18896), .A2(n18881), .B1(n18880), .B2(n18950), .C1(
        n18879), .C2(n18900), .ZN(P3_U3053) );
  OAI222_X1 U22042 ( .A1(n18896), .A2(n18883), .B1(n18882), .B2(n18950), .C1(
        n18881), .C2(n18900), .ZN(P3_U3054) );
  OAI222_X1 U22043 ( .A1(n18896), .A2(n18885), .B1(n18884), .B2(n18950), .C1(
        n18883), .C2(n18900), .ZN(P3_U3055) );
  INV_X1 U22044 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18887) );
  OAI222_X1 U22045 ( .A1(n18896), .A2(n18887), .B1(n18886), .B2(n18950), .C1(
        n18885), .C2(n18900), .ZN(P3_U3056) );
  OAI222_X1 U22046 ( .A1(n18896), .A2(n18889), .B1(n18888), .B2(n18950), .C1(
        n18887), .C2(n18893), .ZN(P3_U3057) );
  INV_X1 U22047 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18892) );
  OAI222_X1 U22048 ( .A1(n18896), .A2(n18892), .B1(n18890), .B2(n18950), .C1(
        n18889), .C2(n18893), .ZN(P3_U3058) );
  OAI222_X1 U22049 ( .A1(n18892), .A2(n18893), .B1(n18891), .B2(n18950), .C1(
        n18894), .C2(n18896), .ZN(P3_U3059) );
  OAI222_X1 U22050 ( .A1(n18896), .A2(n18899), .B1(n18895), .B2(n18950), .C1(
        n18894), .C2(n18893), .ZN(P3_U3060) );
  OAI222_X1 U22051 ( .A1(n18900), .A2(n18899), .B1(n18898), .B2(n18950), .C1(
        n18897), .C2(n18896), .ZN(P3_U3061) );
  INV_X1 U22052 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18901) );
  AOI22_X1 U22053 ( .A1(n18950), .A2(n18902), .B1(n18901), .B2(n18969), .ZN(
        P3_U3274) );
  INV_X1 U22054 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18944) );
  INV_X1 U22055 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18903) );
  AOI22_X1 U22056 ( .A1(n18950), .A2(n18944), .B1(n18903), .B2(n18969), .ZN(
        P3_U3275) );
  INV_X1 U22057 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18904) );
  AOI22_X1 U22058 ( .A1(n18950), .A2(n18905), .B1(n18904), .B2(n18969), .ZN(
        P3_U3276) );
  INV_X1 U22059 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18947) );
  INV_X1 U22060 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18906) );
  AOI22_X1 U22061 ( .A1(n18950), .A2(n18947), .B1(n18906), .B2(n18969), .ZN(
        P3_U3277) );
  INV_X1 U22062 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18909) );
  INV_X1 U22063 ( .A(n18910), .ZN(n18907) );
  AOI21_X1 U22064 ( .B1(n18909), .B2(n18908), .A(n18907), .ZN(P3_U3280) );
  OAI21_X1 U22065 ( .B1(n18912), .B2(n18911), .A(n18910), .ZN(P3_U3281) );
  OAI221_X1 U22066 ( .B1(n18935), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18935), 
        .C2(n18914), .A(n18913), .ZN(P3_U3282) );
  INV_X1 U22067 ( .A(n18915), .ZN(n18916) );
  AOI22_X1 U22068 ( .A1(n21185), .A2(n18917), .B1(n21184), .B2(n18916), .ZN(
        n18922) );
  INV_X1 U22069 ( .A(n18918), .ZN(n18919) );
  AOI21_X1 U22070 ( .B1(n21185), .B2(n18919), .A(n21190), .ZN(n18921) );
  OAI22_X1 U22071 ( .A1(n21190), .A2(n18922), .B1(n18921), .B2(n18920), .ZN(
        P3_U3285) );
  AOI22_X1 U22072 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18924), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18923), .ZN(n21182) );
  NOR2_X1 U22073 ( .A1(n18926), .A2(n18925), .ZN(n21181) );
  INV_X1 U22074 ( .A(n21181), .ZN(n18927) );
  OAI22_X1 U22075 ( .A1(n18929), .A2(n18928), .B1(n21182), .B2(n18927), .ZN(
        n18930) );
  AOI21_X1 U22076 ( .B1(n21184), .B2(n18931), .A(n18930), .ZN(n18932) );
  AOI22_X1 U22077 ( .A1(n21190), .A2(n18933), .B1(n18932), .B2(n21187), .ZN(
        P3_U3288) );
  AOI21_X1 U22078 ( .B1(n18935), .B2(n18934), .A(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n18936) );
  OAI22_X1 U22079 ( .A1(n18937), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n21181), .B2(n18936), .ZN(n18938) );
  INV_X1 U22080 ( .A(n18938), .ZN(n18939) );
  AOI22_X1 U22081 ( .A1(n21190), .A2(n18940), .B1(n18939), .B2(n21187), .ZN(
        P3_U3290) );
  AOI21_X1 U22082 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18942) );
  AOI22_X1 U22083 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18942), .B2(n18941), .ZN(n18945) );
  AOI22_X1 U22084 ( .A1(n18948), .A2(n18945), .B1(n18944), .B2(n18943), .ZN(
        P3_U3292) );
  OAI21_X1 U22085 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18948), .ZN(n18946) );
  OAI21_X1 U22086 ( .B1(n18948), .B2(n18947), .A(n18946), .ZN(P3_U3293) );
  INV_X1 U22087 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18949) );
  AOI22_X1 U22088 ( .A1(n18950), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18949), 
        .B2(n18969), .ZN(P3_U3294) );
  MUX2_X1 U22089 ( .A(P3_MORE_REG_SCAN_IN), .B(n18952), .S(n18951), .Z(
        P3_U3295) );
  AOI21_X1 U22090 ( .B1(n18954), .B2(n18953), .A(n18973), .ZN(n18955) );
  OAI21_X1 U22091 ( .B1(n18957), .B2(n18956), .A(n18955), .ZN(n18968) );
  OAI21_X1 U22092 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18959), .A(n18958), 
        .ZN(n18961) );
  AOI211_X1 U22093 ( .C1(n18972), .C2(n18961), .A(n18960), .B(n18971), .ZN(
        n18963) );
  NOR2_X1 U22094 ( .A1(n18963), .A2(n18962), .ZN(n18964) );
  OAI21_X1 U22095 ( .B1(n18965), .B2(n18964), .A(n18968), .ZN(n18966) );
  OAI21_X1 U22096 ( .B1(n18968), .B2(n18967), .A(n18966), .ZN(P3_U3296) );
  INV_X1 U22097 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18976) );
  INV_X1 U22098 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18970) );
  AOI22_X1 U22099 ( .A1(n18950), .A2(n18976), .B1(n18970), .B2(n18969), .ZN(
        P3_U3297) );
  AOI21_X1 U22100 ( .B1(n21185), .B2(n18971), .A(n18973), .ZN(n18977) );
  INV_X1 U22101 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18974) );
  AOI22_X1 U22102 ( .A1(n18977), .A2(n18974), .B1(n18973), .B2(n18972), .ZN(
        P3_U3298) );
  AOI21_X1 U22103 ( .B1(n18977), .B2(n18976), .A(n18975), .ZN(P3_U3299) );
  INV_X1 U22104 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n21094) );
  INV_X1 U22105 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18978) );
  NAND2_X1 U22106 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20958), .ZN(n19984) );
  NAND2_X1 U22107 ( .A1(n21094), .A2(n20966), .ZN(n19981) );
  OAI21_X1 U22108 ( .B1(n21094), .B2(n19984), .A(n19981), .ZN(n20059) );
  INV_X1 U22109 ( .A(n20059), .ZN(n19974) );
  OAI21_X1 U22110 ( .B1(n21094), .B2(n18978), .A(n19974), .ZN(P2_U2815) );
  INV_X1 U22111 ( .A(n20120), .ZN(n18980) );
  INV_X1 U22112 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18979) );
  OAI22_X1 U22113 ( .A1(n18980), .A2(n18979), .B1(n20061), .B2(n19968), .ZN(
        P2_U2816) );
  OR2_X1 U22114 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20966), .ZN(n20126) );
  INV_X2 U22115 ( .A(n20126), .ZN(n20129) );
  AOI21_X1 U22116 ( .B1(n21094), .B2(n20958), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18981) );
  AOI22_X1 U22117 ( .A1(n20129), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18981), 
        .B2(n20126), .ZN(P2_U2817) );
  OAI21_X1 U22118 ( .B1(n19975), .B2(BS16), .A(n20059), .ZN(n20057) );
  OAI21_X1 U22119 ( .B1(n20059), .B2(n20107), .A(n20057), .ZN(P2_U2818) );
  NOR4_X1 U22120 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18985) );
  NOR4_X1 U22121 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18984) );
  NOR4_X1 U22122 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18983) );
  NOR4_X1 U22123 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18982) );
  NAND4_X1 U22124 ( .A1(n18985), .A2(n18984), .A3(n18983), .A4(n18982), .ZN(
        n18991) );
  NOR4_X1 U22125 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18989) );
  AOI211_X1 U22126 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_4__SCAN_IN), .B(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18988) );
  NOR4_X1 U22127 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18987) );
  NOR4_X1 U22128 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18986) );
  NAND4_X1 U22129 ( .A1(n18989), .A2(n18988), .A3(n18987), .A4(n18986), .ZN(
        n18990) );
  NOR2_X1 U22130 ( .A1(n18991), .A2(n18990), .ZN(n18999) );
  INV_X1 U22131 ( .A(n18999), .ZN(n18998) );
  NOR2_X1 U22132 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18998), .ZN(n18992) );
  INV_X1 U22133 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20055) );
  AOI22_X1 U22134 ( .A1(n18992), .A2(n18993), .B1(n20055), .B2(n18998), .ZN(
        P2_U2820) );
  OR3_X1 U22135 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18997) );
  INV_X1 U22136 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20053) );
  AOI22_X1 U22137 ( .A1(n18992), .A2(n18997), .B1(n18998), .B2(n20053), .ZN(
        P2_U2821) );
  INV_X1 U22138 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20058) );
  NAND2_X1 U22139 ( .A1(n18992), .A2(n20058), .ZN(n18996) );
  INV_X1 U22140 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19993) );
  OAI21_X1 U22141 ( .B1(n18993), .B2(n19993), .A(n18999), .ZN(n18994) );
  OAI21_X1 U22142 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18999), .A(n18994), 
        .ZN(n18995) );
  OAI221_X1 U22143 ( .B1(n18996), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18996), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18995), .ZN(P2_U2822) );
  INV_X1 U22144 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20051) );
  OAI221_X1 U22145 ( .B1(n18999), .B2(n20051), .C1(n18998), .C2(n18997), .A(
        n18996), .ZN(P2_U2823) );
  AOI211_X1 U22146 ( .C1(n19001), .C2(n19000), .A(n9857), .B(n19972), .ZN(
        n19007) );
  AOI22_X1 U22147 ( .A1(n19002), .A2(n19202), .B1(P2_REIP_REG_20__SCAN_IN), 
        .B2(n19204), .ZN(n19004) );
  AOI22_X1 U22148 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n19167), .B1(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19166), .ZN(n19003) );
  OAI211_X1 U22149 ( .C1(n19005), .C2(n19182), .A(n19004), .B(n19003), .ZN(
        n19006) );
  AOI211_X1 U22150 ( .C1(n19187), .C2(n19008), .A(n19007), .B(n19006), .ZN(
        n19009) );
  INV_X1 U22151 ( .A(n19009), .ZN(P2_U2835) );
  AOI211_X1 U22152 ( .C1(n19012), .C2(n19011), .A(n19010), .B(n19972), .ZN(
        n19019) );
  INV_X1 U22153 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19014) );
  AOI22_X1 U22154 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(n19167), .B1(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19166), .ZN(n19013) );
  OAI211_X1 U22155 ( .C1(n19154), .C2(n19014), .A(n19013), .B(n13196), .ZN(
        n19015) );
  INV_X1 U22156 ( .A(n19015), .ZN(n19016) );
  OAI21_X1 U22157 ( .B1(n19017), .B2(n19169), .A(n19016), .ZN(n19018) );
  AOI211_X1 U22158 ( .C1(n19203), .C2(n19020), .A(n19019), .B(n19018), .ZN(
        n19021) );
  OAI21_X1 U22159 ( .B1(n19022), .B2(n19199), .A(n19021), .ZN(P2_U2836) );
  AOI211_X1 U22160 ( .C1(n19025), .C2(n19023), .A(n19024), .B(n19972), .ZN(
        n19030) );
  AOI21_X1 U22161 ( .B1(P2_REIP_REG_18__SCAN_IN), .B2(n19204), .A(n19185), 
        .ZN(n19028) );
  AOI22_X1 U22162 ( .A1(n19026), .A2(n19202), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19166), .ZN(n19027) );
  OAI211_X1 U22163 ( .C1(n19207), .C2(n11598), .A(n19028), .B(n19027), .ZN(
        n19029) );
  AOI211_X1 U22164 ( .C1(n19187), .C2(n19031), .A(n19030), .B(n19029), .ZN(
        n19032) );
  OAI21_X1 U22165 ( .B1(n19033), .B2(n19182), .A(n19032), .ZN(P2_U2837) );
  AOI211_X1 U22166 ( .C1(n19036), .C2(n19035), .A(n19034), .B(n19972), .ZN(
        n19043) );
  INV_X1 U22167 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19038) );
  AOI22_X1 U22168 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19166), .B1(
        P2_EBX_REG_17__SCAN_IN), .B2(n19167), .ZN(n19037) );
  OAI211_X1 U22169 ( .C1(n19154), .C2(n19038), .A(n19037), .B(n13196), .ZN(
        n19039) );
  INV_X1 U22170 ( .A(n19039), .ZN(n19040) );
  OAI21_X1 U22171 ( .B1(n19041), .B2(n19169), .A(n19040), .ZN(n19042) );
  AOI211_X1 U22172 ( .C1(n19203), .C2(n19044), .A(n19043), .B(n19042), .ZN(
        n19045) );
  OAI21_X1 U22173 ( .B1(n19046), .B2(n19199), .A(n19045), .ZN(P2_U2838) );
  INV_X1 U22174 ( .A(n19047), .ZN(n19048) );
  OAI22_X1 U22175 ( .A1(n19048), .A2(n19169), .B1(n19207), .B2(n11588), .ZN(
        n19049) );
  AOI211_X1 U22176 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n19204), .A(n19185), 
        .B(n19049), .ZN(n19058) );
  OAI21_X1 U22177 ( .B1(n19051), .B2(n19050), .A(n19198), .ZN(n19053) );
  OAI22_X1 U22178 ( .A1(n19054), .A2(n19053), .B1(n19052), .B2(n19182), .ZN(
        n19055) );
  AOI21_X1 U22179 ( .B1(n19056), .B2(n19187), .A(n19055), .ZN(n19057) );
  OAI211_X1 U22180 ( .C1(n19059), .C2(n19144), .A(n19058), .B(n19057), .ZN(
        P2_U2839) );
  OAI21_X1 U22181 ( .B1(n11032), .B2(n19154), .A(n13196), .ZN(n19062) );
  OAI22_X1 U22182 ( .A1(n19060), .A2(n19169), .B1(n11585), .B2(n19207), .ZN(
        n19061) );
  AOI211_X1 U22183 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n19166), .A(
        n19062), .B(n19061), .ZN(n19069) );
  NAND2_X1 U22184 ( .A1(n19173), .A2(n19063), .ZN(n19064) );
  XNOR2_X1 U22185 ( .A(n19065), .B(n19064), .ZN(n19066) );
  AOI22_X1 U22186 ( .A1(n19067), .A2(n19187), .B1(n19198), .B2(n19066), .ZN(
        n19068) );
  OAI211_X1 U22187 ( .C1(n19221), .C2(n19182), .A(n19069), .B(n19068), .ZN(
        P2_U2840) );
  INV_X1 U22188 ( .A(n19070), .ZN(n19072) );
  AOI22_X1 U22189 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19211), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n19167), .ZN(n19071) );
  OAI21_X1 U22190 ( .B1(n19072), .B2(n19169), .A(n19071), .ZN(n19073) );
  AOI211_X1 U22191 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19204), .A(n19185), 
        .B(n19073), .ZN(n19080) );
  NOR2_X1 U22192 ( .A1(n10058), .A2(n19074), .ZN(n19076) );
  XNOR2_X1 U22193 ( .A(n19076), .B(n19075), .ZN(n19077) );
  AOI22_X1 U22194 ( .A1(n19187), .A2(n19078), .B1(n19198), .B2(n19077), .ZN(
        n19079) );
  OAI211_X1 U22195 ( .C1(n19182), .C2(n19223), .A(n19080), .B(n19079), .ZN(
        P2_U2841) );
  AOI22_X1 U22196 ( .A1(n19081), .A2(n19202), .B1(P2_EBX_REG_13__SCAN_IN), 
        .B2(n19167), .ZN(n19082) );
  OAI211_X1 U22197 ( .C1(n11025), .C2(n19154), .A(n19082), .B(n13196), .ZN(
        n19083) );
  AOI21_X1 U22198 ( .B1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19166), .A(
        n19083), .ZN(n19089) );
  NAND2_X1 U22199 ( .A1(n19173), .A2(n19084), .ZN(n19085) );
  XNOR2_X1 U22200 ( .A(n19086), .B(n19085), .ZN(n19087) );
  AOI22_X1 U22201 ( .A1(n19198), .A2(n19087), .B1(n19203), .B2(n19224), .ZN(
        n19088) );
  OAI211_X1 U22202 ( .C1(n19199), .C2(n19090), .A(n19089), .B(n19088), .ZN(
        P2_U2842) );
  NOR2_X1 U22203 ( .A1(n10058), .A2(n19091), .ZN(n19106) );
  XOR2_X1 U22204 ( .A(n19106), .B(n19092), .Z(n19099) );
  AOI22_X1 U22205 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19211), .B1(
        P2_EBX_REG_12__SCAN_IN), .B2(n19167), .ZN(n19093) );
  OAI21_X1 U22206 ( .B1(n19094), .B2(n19169), .A(n19093), .ZN(n19095) );
  AOI211_X1 U22207 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19204), .A(n19185), 
        .B(n19095), .ZN(n19098) );
  AOI22_X1 U22208 ( .A1(n19187), .A2(n19096), .B1(n19203), .B2(n19226), .ZN(
        n19097) );
  OAI211_X1 U22209 ( .C1(n19972), .C2(n19099), .A(n19098), .B(n19097), .ZN(
        P2_U2843) );
  AOI22_X1 U22210 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19211), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n19204), .ZN(n19102) );
  AOI22_X1 U22211 ( .A1(n19100), .A2(n19202), .B1(n19203), .B2(n19230), .ZN(
        n19101) );
  NAND3_X1 U22212 ( .A1(n19102), .A2(n19101), .A3(n13196), .ZN(n19103) );
  AOI21_X1 U22213 ( .B1(P2_EBX_REG_11__SCAN_IN), .B2(n19167), .A(n19103), .ZN(
        n19110) );
  AOI21_X1 U22214 ( .B1(n19108), .B2(n19104), .A(n19972), .ZN(n19105) );
  AOI22_X1 U22215 ( .A1(n19108), .A2(n19107), .B1(n19106), .B2(n19105), .ZN(
        n19109) );
  OAI211_X1 U22216 ( .C1(n19199), .C2(n19111), .A(n19110), .B(n19109), .ZN(
        P2_U2844) );
  OAI21_X1 U22217 ( .B1(n20011), .B2(n19154), .A(n13196), .ZN(n19114) );
  OAI22_X1 U22218 ( .A1(n19112), .A2(n19169), .B1(n11570), .B2(n19207), .ZN(
        n19113) );
  AOI211_X1 U22219 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n19166), .A(
        n19114), .B(n19113), .ZN(n19120) );
  NOR2_X1 U22220 ( .A1(n10058), .A2(n19115), .ZN(n19117) );
  XNOR2_X1 U22221 ( .A(n19117), .B(n19116), .ZN(n19118) );
  AOI22_X1 U22222 ( .A1(n19187), .A2(n9846), .B1(n19198), .B2(n19118), .ZN(
        n19119) );
  OAI211_X1 U22223 ( .C1(n19182), .C2(n19233), .A(n19120), .B(n19119), .ZN(
        P2_U2845) );
  AOI22_X1 U22224 ( .A1(n19121), .A2(n19202), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n19167), .ZN(n19122) );
  OAI21_X1 U22225 ( .B1(n19123), .B2(n19144), .A(n19122), .ZN(n19124) );
  AOI211_X1 U22226 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n19204), .A(n19185), .B(
        n19124), .ZN(n19130) );
  NAND2_X1 U22227 ( .A1(n19173), .A2(n19125), .ZN(n19126) );
  XNOR2_X1 U22228 ( .A(n19127), .B(n19126), .ZN(n19128) );
  AOI22_X1 U22229 ( .A1(n19198), .A2(n19128), .B1(n19203), .B2(n19234), .ZN(
        n19129) );
  OAI211_X1 U22230 ( .C1(n19199), .C2(n19131), .A(n19130), .B(n19129), .ZN(
        P2_U2846) );
  AOI22_X1 U22231 ( .A1(n19132), .A2(n19202), .B1(P2_EBX_REG_8__SCAN_IN), .B2(
        n19167), .ZN(n19133) );
  OAI21_X1 U22232 ( .B1(n21066), .B2(n19144), .A(n19133), .ZN(n19134) );
  AOI211_X1 U22233 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n19204), .A(n19185), .B(
        n19134), .ZN(n19141) );
  NOR2_X1 U22234 ( .A1(n10058), .A2(n19135), .ZN(n19137) );
  XNOR2_X1 U22235 ( .A(n19137), .B(n19136), .ZN(n19138) );
  AOI22_X1 U22236 ( .A1(n19187), .A2(n19139), .B1(n19198), .B2(n19138), .ZN(
        n19140) );
  OAI211_X1 U22237 ( .C1(n19182), .C2(n19239), .A(n19141), .B(n19140), .ZN(
        P2_U2847) );
  AOI22_X1 U22238 ( .A1(n19142), .A2(n19202), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19167), .ZN(n19143) );
  OAI21_X1 U22239 ( .B1(n19145), .B2(n19144), .A(n19143), .ZN(n19146) );
  AOI211_X1 U22240 ( .C1(P2_REIP_REG_7__SCAN_IN), .C2(n19204), .A(n19185), .B(
        n19146), .ZN(n19152) );
  NAND2_X1 U22241 ( .A1(n19173), .A2(n19147), .ZN(n19148) );
  XNOR2_X1 U22242 ( .A(n19149), .B(n19148), .ZN(n19150) );
  AOI22_X1 U22243 ( .A1(n19198), .A2(n19150), .B1(n19203), .B2(n19241), .ZN(
        n19151) );
  OAI211_X1 U22244 ( .C1(n19199), .C2(n19153), .A(n19152), .B(n19151), .ZN(
        P2_U2848) );
  OAI21_X1 U22245 ( .B1(n20003), .B2(n19154), .A(n13196), .ZN(n19158) );
  OAI22_X1 U22246 ( .A1(n19156), .A2(n19169), .B1(n19207), .B2(n19155), .ZN(
        n19157) );
  AOI211_X1 U22247 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19211), .A(
        n19158), .B(n19157), .ZN(n19164) );
  NOR2_X1 U22248 ( .A1(n10058), .A2(n19159), .ZN(n19161) );
  XNOR2_X1 U22249 ( .A(n19161), .B(n19160), .ZN(n19162) );
  AOI22_X1 U22250 ( .A1(n19198), .A2(n19162), .B1(n19203), .B2(n9848), .ZN(
        n19163) );
  OAI211_X1 U22251 ( .C1(n19199), .C2(n19165), .A(n19164), .B(n19163), .ZN(
        P2_U2849) );
  AOI22_X1 U22252 ( .A1(P2_EBX_REG_5__SCAN_IN), .A2(n19167), .B1(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19166), .ZN(n19168) );
  OAI21_X1 U22253 ( .B1(n19170), .B2(n19169), .A(n19168), .ZN(n19171) );
  AOI211_X1 U22254 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19204), .A(n19185), .B(
        n19171), .ZN(n19178) );
  NAND2_X1 U22255 ( .A1(n19173), .A2(n19172), .ZN(n19174) );
  XNOR2_X1 U22256 ( .A(n19175), .B(n19174), .ZN(n19176) );
  AOI22_X1 U22257 ( .A1(n19198), .A2(n19176), .B1(n19203), .B2(n19245), .ZN(
        n19177) );
  OAI211_X1 U22258 ( .C1(n19199), .C2(n19179), .A(n19178), .B(n19177), .ZN(
        P2_U2850) );
  AOI22_X1 U22259 ( .A1(n19180), .A2(n19202), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19211), .ZN(n19196) );
  OAI22_X1 U22260 ( .A1(n19207), .A2(n19183), .B1(n19182), .B2(n19181), .ZN(
        n19184) );
  AOI211_X1 U22261 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19204), .A(n19185), .B(
        n19184), .ZN(n19195) );
  INV_X1 U22262 ( .A(n19186), .ZN(n19246) );
  AOI22_X1 U22263 ( .A1(n19246), .A2(n19210), .B1(n19370), .B2(n19187), .ZN(
        n19194) );
  INV_X1 U22264 ( .A(n19373), .ZN(n19192) );
  NOR2_X1 U22265 ( .A1(n10058), .A2(n19188), .ZN(n19191) );
  AOI21_X1 U22266 ( .B1(n19192), .B2(n19191), .A(n19972), .ZN(n19190) );
  OAI21_X1 U22267 ( .B1(n19192), .B2(n19191), .A(n19190), .ZN(n19193) );
  NAND4_X1 U22268 ( .A1(n19196), .A2(n19195), .A3(n19194), .A4(n19193), .ZN(
        P2_U2851) );
  INV_X1 U22269 ( .A(n19197), .ZN(n19214) );
  NOR2_X1 U22270 ( .A1(n19200), .A2(n19199), .ZN(n19209) );
  AOI22_X1 U22271 ( .A1(n19203), .A2(n19273), .B1(n19202), .B2(n19201), .ZN(
        n19206) );
  NAND2_X1 U22272 ( .A1(n19204), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n19205) );
  OAI211_X1 U22273 ( .C1(n19207), .C2(n11203), .A(n19206), .B(n19205), .ZN(
        n19208) );
  AOI211_X1 U22274 ( .C1(n19274), .C2(n19210), .A(n19209), .B(n19208), .ZN(
        n19213) );
  NAND2_X1 U22275 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19211), .ZN(
        n19212) );
  OAI211_X1 U22276 ( .C1(n19214), .C2(n19972), .A(n19213), .B(n19212), .ZN(
        P2_U2855) );
  AOI22_X1 U22277 ( .A1(n19216), .A2(n19263), .B1(n19215), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19219) );
  AOI22_X1 U22278 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19217), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19262), .ZN(n19218) );
  NAND2_X1 U22279 ( .A1(n19219), .A2(n19218), .ZN(P2_U2888) );
  INV_X1 U22280 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19322) );
  OAI222_X1 U22281 ( .A1(n19322), .A2(n19270), .B1(n19221), .B2(n19238), .C1(
        n19220), .C2(n19269), .ZN(P2_U2904) );
  AOI22_X1 U22282 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19262), .B1(n19356), 
        .B2(n19280), .ZN(n19222) );
  OAI21_X1 U22283 ( .B1(n19238), .B2(n19223), .A(n19222), .ZN(P2_U2905) );
  INV_X1 U22284 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19326) );
  INV_X1 U22285 ( .A(n19238), .ZN(n19244) );
  AOI22_X1 U22286 ( .A1(n19224), .A2(n19244), .B1(n19354), .B2(n19280), .ZN(
        n19225) );
  OAI21_X1 U22287 ( .B1(n19270), .B2(n19326), .A(n19225), .ZN(P2_U2906) );
  AOI22_X1 U22288 ( .A1(n19226), .A2(n19244), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n19262), .ZN(n19227) );
  OAI21_X1 U22289 ( .B1(n19228), .B2(n19269), .A(n19227), .ZN(P2_U2907) );
  AOI22_X1 U22290 ( .A1(n19230), .A2(n19244), .B1(n19229), .B2(n19280), .ZN(
        n19231) );
  OAI21_X1 U22291 ( .B1(n19270), .B2(n20917), .A(n19231), .ZN(P2_U2908) );
  INV_X1 U22292 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19330) );
  OAI222_X1 U22293 ( .A1(n19330), .A2(n19270), .B1(n19233), .B2(n19238), .C1(
        n19269), .C2(n19232), .ZN(P2_U2909) );
  AOI22_X1 U22294 ( .A1(n19234), .A2(n19244), .B1(P2_EAX_REG_9__SCAN_IN), .B2(
        n19262), .ZN(n19235) );
  OAI21_X1 U22295 ( .B1(n19236), .B2(n19269), .A(n19235), .ZN(P2_U2910) );
  INV_X1 U22296 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19334) );
  OAI222_X1 U22297 ( .A1(n19334), .A2(n19270), .B1(n19239), .B2(n19238), .C1(
        n19269), .C2(n19237), .ZN(P2_U2911) );
  INV_X1 U22298 ( .A(n19240), .ZN(n19455) );
  AOI22_X1 U22299 ( .A1(n19241), .A2(n19244), .B1(P2_EAX_REG_7__SCAN_IN), .B2(
        n19262), .ZN(n19242) );
  OAI21_X1 U22300 ( .B1(n19455), .B2(n19269), .A(n19242), .ZN(P2_U2912) );
  AOI22_X1 U22301 ( .A1(n9848), .A2(n19244), .B1(P2_EAX_REG_6__SCAN_IN), .B2(
        n19262), .ZN(n19243) );
  OAI21_X1 U22302 ( .B1(n19443), .B2(n19269), .A(n19243), .ZN(P2_U2913) );
  AOI22_X1 U22303 ( .A1(n19245), .A2(n19244), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19262), .ZN(n19249) );
  NAND3_X1 U22304 ( .A1(n19247), .A2(n19246), .A3(n10867), .ZN(n19248) );
  OAI211_X1 U22305 ( .C1(n19439), .C2(n19269), .A(n19249), .B(n19248), .ZN(
        P2_U2914) );
  AOI22_X1 U22306 ( .A1(n19263), .A2(n20065), .B1(n19262), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n19255) );
  AOI21_X1 U22307 ( .B1(n19252), .B2(n19251), .A(n19250), .ZN(n19253) );
  OR2_X1 U22308 ( .A1(n19253), .A2(n19275), .ZN(n19254) );
  OAI211_X1 U22309 ( .C1(n19432), .C2(n19269), .A(n19255), .B(n19254), .ZN(
        P2_U2916) );
  AOI22_X1 U22310 ( .A1(n20074), .A2(n19263), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19262), .ZN(n19261) );
  AOI21_X1 U22311 ( .B1(n19258), .B2(n19257), .A(n19256), .ZN(n19259) );
  OR2_X1 U22312 ( .A1(n19259), .A2(n19275), .ZN(n19260) );
  OAI211_X1 U22313 ( .C1(n19427), .C2(n19269), .A(n19261), .B(n19260), .ZN(
        P2_U2917) );
  AOI22_X1 U22314 ( .A1(n19263), .A2(n20083), .B1(n19262), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19268) );
  AOI21_X1 U22315 ( .B1(n19277), .B2(n19265), .A(n19264), .ZN(n19266) );
  OR2_X1 U22316 ( .A1(n19266), .A2(n19275), .ZN(n19267) );
  OAI211_X1 U22317 ( .C1(n19423), .C2(n19269), .A(n19268), .B(n19267), .ZN(
        P2_U2918) );
  INV_X1 U22318 ( .A(n19273), .ZN(n19271) );
  INV_X1 U22319 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19353) );
  OAI22_X1 U22320 ( .A1(n19272), .A2(n19271), .B1(n19270), .B2(n19353), .ZN(
        n19279) );
  NOR2_X1 U22321 ( .A1(n19274), .A2(n19273), .ZN(n19276) );
  NOR3_X1 U22322 ( .A1(n19277), .A2(n19276), .A3(n19275), .ZN(n19278) );
  AOI211_X1 U22323 ( .C1(n19281), .C2(n19280), .A(n19279), .B(n19278), .ZN(
        n19282) );
  INV_X1 U22324 ( .A(n19282), .ZN(P2_U2919) );
  OR2_X1 U22325 ( .A1(n10850), .A2(n9755), .ZN(n19284) );
  OAI21_X1 U22326 ( .B1(n19285), .B2(n19284), .A(n19283), .ZN(n19286) );
  NAND2_X1 U22327 ( .A1(n19287), .A2(n19352), .ZN(n19294) );
  NOR2_X1 U22328 ( .A1(n19294), .A2(n19288), .ZN(P2_U2920) );
  NOR2_X1 U22329 ( .A1(n19352), .A2(n19289), .ZN(n19293) );
  AOI22_X1 U22330 ( .A1(P2_EAX_REG_30__SCAN_IN), .A2(n19293), .B1(n19350), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19290) );
  OAI21_X1 U22331 ( .B1(n20891), .B2(n19294), .A(n19290), .ZN(P2_U2921) );
  AOI22_X1 U22332 ( .A1(P2_EAX_REG_29__SCAN_IN), .A2(n19293), .B1(n19350), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n19291) );
  OAI21_X1 U22333 ( .B1(n19294), .B2(n19292), .A(n19291), .ZN(P2_U2922) );
  INV_X1 U22334 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n19296) );
  INV_X2 U22335 ( .A(n19294), .ZN(n19339) );
  AOI22_X1 U22336 ( .A1(n19350), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19295) );
  OAI21_X1 U22337 ( .B1(n19296), .B2(n19319), .A(n19295), .ZN(P2_U2923) );
  AOI22_X1 U22338 ( .A1(n19350), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n19297) );
  OAI21_X1 U22339 ( .B1(n21123), .B2(n19319), .A(n19297), .ZN(P2_U2924) );
  INV_X1 U22340 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n19299) );
  AOI22_X1 U22341 ( .A1(n19350), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19298) );
  OAI21_X1 U22342 ( .B1(n19299), .B2(n19319), .A(n19298), .ZN(P2_U2925) );
  INV_X1 U22343 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n19301) );
  AOI22_X1 U22344 ( .A1(n19350), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n19300) );
  OAI21_X1 U22345 ( .B1(n19301), .B2(n19319), .A(n19300), .ZN(P2_U2926) );
  INV_X1 U22346 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n19303) );
  AOI22_X1 U22347 ( .A1(n19350), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19302) );
  OAI21_X1 U22348 ( .B1(n19303), .B2(n19319), .A(n19302), .ZN(P2_U2927) );
  INV_X1 U22349 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19305) );
  AOI22_X1 U22350 ( .A1(n19350), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19304) );
  OAI21_X1 U22351 ( .B1(n19305), .B2(n19319), .A(n19304), .ZN(P2_U2928) );
  AOI22_X1 U22352 ( .A1(n19350), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n19306) );
  OAI21_X1 U22353 ( .B1(n19307), .B2(n19319), .A(n19306), .ZN(P2_U2929) );
  INV_X1 U22354 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n19309) );
  AOI22_X1 U22355 ( .A1(n19350), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n19308) );
  OAI21_X1 U22356 ( .B1(n19309), .B2(n19319), .A(n19308), .ZN(P2_U2930) );
  INV_X1 U22357 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19311) );
  AOI22_X1 U22358 ( .A1(n19350), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19310) );
  OAI21_X1 U22359 ( .B1(n19311), .B2(n19319), .A(n19310), .ZN(P2_U2931) );
  INV_X1 U22360 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n19313) );
  AOI22_X1 U22361 ( .A1(n19350), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19312) );
  OAI21_X1 U22362 ( .B1(n19313), .B2(n19319), .A(n19312), .ZN(P2_U2932) );
  INV_X1 U22363 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19315) );
  AOI22_X1 U22364 ( .A1(n19350), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19314) );
  OAI21_X1 U22365 ( .B1(n19315), .B2(n19319), .A(n19314), .ZN(P2_U2933) );
  INV_X1 U22366 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n19317) );
  AOI22_X1 U22367 ( .A1(n19350), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n19316) );
  OAI21_X1 U22368 ( .B1(n19317), .B2(n19319), .A(n19316), .ZN(P2_U2934) );
  INV_X1 U22369 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19320) );
  AOI22_X1 U22370 ( .A1(n19350), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n19318) );
  OAI21_X1 U22371 ( .B1(n19320), .B2(n19319), .A(n19318), .ZN(P2_U2935) );
  AOI22_X1 U22372 ( .A1(n19350), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19321) );
  OAI21_X1 U22373 ( .B1(n19322), .B2(n19352), .A(n19321), .ZN(P2_U2936) );
  INV_X1 U22374 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19324) );
  AOI22_X1 U22375 ( .A1(n19350), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19323) );
  OAI21_X1 U22376 ( .B1(n19324), .B2(n19352), .A(n19323), .ZN(P2_U2937) );
  AOI22_X1 U22377 ( .A1(n19350), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19325) );
  OAI21_X1 U22378 ( .B1(n19326), .B2(n19352), .A(n19325), .ZN(P2_U2938) );
  INV_X1 U22379 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n21138) );
  AOI22_X1 U22380 ( .A1(n19350), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19327) );
  OAI21_X1 U22381 ( .B1(n21138), .B2(n19352), .A(n19327), .ZN(P2_U2939) );
  AOI22_X1 U22382 ( .A1(n19350), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19328) );
  OAI21_X1 U22383 ( .B1(n20917), .B2(n19352), .A(n19328), .ZN(P2_U2940) );
  AOI22_X1 U22384 ( .A1(n19350), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19329) );
  OAI21_X1 U22385 ( .B1(n19330), .B2(n19352), .A(n19329), .ZN(P2_U2941) );
  INV_X1 U22386 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19332) );
  AOI22_X1 U22387 ( .A1(n19350), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19331) );
  OAI21_X1 U22388 ( .B1(n19332), .B2(n19352), .A(n19331), .ZN(P2_U2942) );
  AOI22_X1 U22389 ( .A1(n19350), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19333) );
  OAI21_X1 U22390 ( .B1(n19334), .B2(n19352), .A(n19333), .ZN(P2_U2943) );
  INV_X1 U22391 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19336) );
  AOI22_X1 U22392 ( .A1(n19350), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19335) );
  OAI21_X1 U22393 ( .B1(n19336), .B2(n19352), .A(n19335), .ZN(P2_U2944) );
  INV_X1 U22394 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19338) );
  AOI22_X1 U22395 ( .A1(n19350), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19337) );
  OAI21_X1 U22396 ( .B1(n19338), .B2(n19352), .A(n19337), .ZN(P2_U2945) );
  INV_X1 U22397 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19341) );
  AOI22_X1 U22398 ( .A1(n19350), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19340) );
  OAI21_X1 U22399 ( .B1(n19341), .B2(n19352), .A(n19340), .ZN(P2_U2946) );
  INV_X1 U22400 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19343) );
  AOI22_X1 U22401 ( .A1(n19350), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19342) );
  OAI21_X1 U22402 ( .B1(n19343), .B2(n19352), .A(n19342), .ZN(P2_U2947) );
  INV_X1 U22403 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19345) );
  AOI22_X1 U22404 ( .A1(n19350), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19344) );
  OAI21_X1 U22405 ( .B1(n19345), .B2(n19352), .A(n19344), .ZN(P2_U2948) );
  INV_X1 U22406 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19347) );
  AOI22_X1 U22407 ( .A1(n19350), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19346) );
  OAI21_X1 U22408 ( .B1(n19347), .B2(n19352), .A(n19346), .ZN(P2_U2949) );
  INV_X1 U22409 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19349) );
  AOI22_X1 U22410 ( .A1(n19350), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19348) );
  OAI21_X1 U22411 ( .B1(n19349), .B2(n19352), .A(n19348), .ZN(P2_U2950) );
  AOI22_X1 U22412 ( .A1(n19350), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19351) );
  OAI21_X1 U22413 ( .B1(n19353), .B2(n19352), .A(n19351), .ZN(P2_U2951) );
  AOI22_X1 U22414 ( .A1(P2_EAX_REG_29__SCAN_IN), .A2(n19362), .B1(n19361), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n19355) );
  NAND2_X1 U22415 ( .A1(n19357), .A2(n19354), .ZN(n19359) );
  NAND2_X1 U22416 ( .A1(n19355), .A2(n19359), .ZN(P2_U2965) );
  AOI22_X1 U22417 ( .A1(P2_EAX_REG_30__SCAN_IN), .A2(n19362), .B1(n19361), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19358) );
  NAND2_X1 U22418 ( .A1(n19357), .A2(n19356), .ZN(n19363) );
  NAND2_X1 U22419 ( .A1(n19358), .A2(n19363), .ZN(P2_U2966) );
  AOI22_X1 U22420 ( .A1(n19362), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n19361), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n19360) );
  NAND2_X1 U22421 ( .A1(n19360), .A2(n19359), .ZN(P2_U2980) );
  AOI22_X1 U22422 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19362), .B1(n19361), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19364) );
  NAND2_X1 U22423 ( .A1(n19364), .A2(n19363), .ZN(P2_U2981) );
  AOI22_X1 U22424 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19376), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19365), .ZN(n19372) );
  INV_X1 U22425 ( .A(n19366), .ZN(n19368) );
  OAI22_X1 U22426 ( .A1(n19368), .A2(n19385), .B1(n19367), .B2(n9780), .ZN(
        n19369) );
  AOI21_X1 U22427 ( .B1(n19382), .B2(n19370), .A(n19369), .ZN(n19371) );
  OAI211_X1 U22428 ( .C1(n19374), .C2(n19373), .A(n19372), .B(n19371), .ZN(
        P2_U3010) );
  NOR2_X1 U22429 ( .A1(n19376), .A2(n19375), .ZN(n19390) );
  OAI21_X1 U22430 ( .B1(n19379), .B2(n19378), .A(n19377), .ZN(n19380) );
  INV_X1 U22431 ( .A(n19380), .ZN(n19384) );
  NAND2_X1 U22432 ( .A1(n19382), .A2(n19381), .ZN(n19383) );
  OAI211_X1 U22433 ( .C1(n19386), .C2(n19385), .A(n19384), .B(n19383), .ZN(
        n19387) );
  INV_X1 U22434 ( .A(n19387), .ZN(n19388) );
  OAI21_X1 U22435 ( .B1(n19390), .B2(n19389), .A(n19388), .ZN(P2_U3014) );
  AOI22_X1 U22436 ( .A1(n19392), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19391), .B2(n20083), .ZN(n19393) );
  OAI21_X1 U22437 ( .B1(n19395), .B2(n19394), .A(n19393), .ZN(n19401) );
  AOI211_X1 U22438 ( .C1(n19399), .C2(n19398), .A(n19397), .B(n19396), .ZN(
        n19400) );
  AOI211_X1 U22439 ( .C1(n19402), .C2(n11087), .A(n19401), .B(n19400), .ZN(
        n19404) );
  OAI211_X1 U22440 ( .C1(n19406), .C2(n19405), .A(n19404), .B(n19403), .ZN(
        P2_U3045) );
  NAND2_X1 U22441 ( .A1(n20069), .A2(n20076), .ZN(n19518) );
  OR2_X1 U22442 ( .A1(n19518), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19462) );
  NOR2_X1 U22443 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19462), .ZN(
        n19454) );
  AOI22_X1 U22444 ( .A1(n19886), .A2(n19960), .B1(n19876), .B2(n19454), .ZN(
        n19419) );
  NAND3_X1 U22445 ( .A1(n19409), .A2(n20064), .A3(n19485), .ZN(n19410) );
  NAND2_X1 U22446 ( .A1(n20064), .A2(n20107), .ZN(n19871) );
  NAND2_X1 U22447 ( .A1(n19410), .A2(n19871), .ZN(n19414) );
  OAI21_X1 U22448 ( .B1(n19415), .B2(n20113), .A(n19879), .ZN(n19411) );
  AOI21_X1 U22449 ( .B1(n19414), .B2(n19412), .A(n19411), .ZN(n19413) );
  OAI21_X1 U22450 ( .B1(n19413), .B2(n19454), .A(n19883), .ZN(n19457) );
  OAI21_X1 U22451 ( .B1(n19954), .B2(n19454), .A(n19414), .ZN(n19417) );
  OAI21_X1 U22452 ( .B1(n19415), .B2(n19454), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19416) );
  NAND2_X1 U22453 ( .A1(n19417), .A2(n19416), .ZN(n19456) );
  AOI22_X1 U22454 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19457), .B1(
        n19833), .B2(n19456), .ZN(n19418) );
  OAI211_X1 U22455 ( .C1(n19803), .C2(n19485), .A(n19419), .B(n19418), .ZN(
        P2_U3048) );
  OAI22_X1 U22456 ( .A1(n19421), .A2(n19446), .B1(n19420), .B2(n19448), .ZN(
        n19918) );
  AOI22_X1 U22457 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19451), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19450), .ZN(n19847) );
  NOR2_X2 U22458 ( .A1(n19453), .A2(n19422), .ZN(n19915) );
  AOI22_X1 U22459 ( .A1(n19917), .A2(n19960), .B1(n19915), .B2(n19454), .ZN(
        n19425) );
  NOR2_X2 U22460 ( .A1(n19423), .A2(n19796), .ZN(n19916) );
  AOI22_X1 U22461 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19457), .B1(
        n19916), .B2(n19456), .ZN(n19424) );
  OAI211_X1 U22462 ( .C1(n19806), .C2(n19485), .A(n19425), .B(n19424), .ZN(
        P2_U3049) );
  AOI22_X1 U22463 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19451), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19450), .ZN(n19850) );
  NOR2_X2 U22464 ( .A1(n19453), .A2(n10317), .ZN(n19921) );
  AOI22_X1 U22465 ( .A1(n19923), .A2(n19960), .B1(n19921), .B2(n19454), .ZN(
        n19429) );
  NOR2_X2 U22466 ( .A1(n19427), .A2(n19796), .ZN(n19922) );
  AOI22_X1 U22467 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19457), .B1(
        n19922), .B2(n19456), .ZN(n19428) );
  OAI211_X1 U22468 ( .C1(n19809), .C2(n19485), .A(n19429), .B(n19428), .ZN(
        P2_U3050) );
  AOI22_X1 U22469 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19451), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19450), .ZN(n19812) );
  OAI22_X2 U22470 ( .A1(n19431), .A2(n19446), .B1(n19430), .B2(n19448), .ZN(
        n19931) );
  NOR2_X2 U22471 ( .A1(n19453), .A2(n10345), .ZN(n19928) );
  AOI22_X1 U22472 ( .A1(n19931), .A2(n19960), .B1(n19928), .B2(n19454), .ZN(
        n19434) );
  NOR2_X2 U22473 ( .A1(n19432), .A2(n19796), .ZN(n19929) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19457), .B1(
        n19929), .B2(n19456), .ZN(n19433) );
  OAI211_X1 U22475 ( .C1(n19812), .C2(n19485), .A(n19434), .B(n19433), .ZN(
        P2_U3051) );
  AOI22_X1 U22476 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19451), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19450), .ZN(n19856) );
  AOI22_X1 U22477 ( .A1(n19936), .A2(n19960), .B1(n19934), .B2(n19454), .ZN(
        n19438) );
  NAND2_X1 U22478 ( .A1(n19436), .A2(n19883), .ZN(n19901) );
  AOI22_X1 U22479 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19457), .B1(
        n19935), .B2(n19456), .ZN(n19437) );
  OAI211_X1 U22480 ( .C1(n19815), .C2(n19485), .A(n19438), .B(n19437), .ZN(
        P2_U3052) );
  AOI22_X1 U22481 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19451), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19450), .ZN(n19818) );
  AOI22_X1 U22482 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19450), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19451), .ZN(n19859) );
  NOR2_X2 U22483 ( .A1(n19453), .A2(n11394), .ZN(n19941) );
  AOI22_X1 U22484 ( .A1(n19944), .A2(n19960), .B1(n19941), .B2(n19454), .ZN(
        n19441) );
  NOR2_X2 U22485 ( .A1(n19439), .A2(n19796), .ZN(n19942) );
  AOI22_X1 U22486 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19457), .B1(
        n19942), .B2(n19456), .ZN(n19440) );
  OAI211_X1 U22487 ( .C1(n19818), .C2(n19485), .A(n19441), .B(n19440), .ZN(
        P2_U3053) );
  AOI22_X1 U22488 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19451), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19450), .ZN(n19821) );
  AOI22_X1 U22489 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19450), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19451), .ZN(n19862) );
  NOR2_X2 U22490 ( .A1(n19453), .A2(n19442), .ZN(n19947) );
  AOI22_X1 U22491 ( .A1(n19950), .A2(n19960), .B1(n19947), .B2(n19454), .ZN(
        n19445) );
  NOR2_X2 U22492 ( .A1(n19443), .A2(n19796), .ZN(n19948) );
  AOI22_X1 U22493 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19457), .B1(
        n19948), .B2(n19456), .ZN(n19444) );
  OAI211_X1 U22494 ( .C1(n19821), .C2(n19485), .A(n19445), .B(n19444), .ZN(
        P2_U3054) );
  OAI22_X1 U22495 ( .A1(n19449), .A2(n19448), .B1(n19447), .B2(n19446), .ZN(
        n19959) );
  AOI22_X1 U22496 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19451), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19450), .ZN(n19868) );
  NOR2_X2 U22497 ( .A1(n19453), .A2(n19452), .ZN(n19953) );
  AOI22_X1 U22498 ( .A1(n19957), .A2(n19960), .B1(n19953), .B2(n19454), .ZN(
        n19459) );
  NOR2_X2 U22499 ( .A1(n19455), .A2(n19796), .ZN(n19955) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19457), .B1(
        n19955), .B2(n19456), .ZN(n19458) );
  OAI211_X1 U22501 ( .C1(n19828), .C2(n19485), .A(n19459), .B(n19458), .ZN(
        P2_U3055) );
  NAND2_X1 U22502 ( .A1(n19695), .A2(n19580), .ZN(n19490) );
  INV_X1 U22503 ( .A(n20064), .ZN(n19694) );
  NOR2_X1 U22504 ( .A1(n19693), .A2(n19518), .ZN(n19480) );
  OAI21_X1 U22505 ( .B1(n19460), .B2(n19480), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19461) );
  OAI21_X1 U22506 ( .B1(n19462), .B2(n19694), .A(n19461), .ZN(n19481) );
  AOI22_X1 U22507 ( .A1(n19481), .A2(n19833), .B1(n19876), .B2(n19480), .ZN(
        n19466) );
  AOI21_X1 U22508 ( .B1(n11257), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19464) );
  OAI21_X1 U22509 ( .B1(n19581), .B2(n19692), .A(n19462), .ZN(n19463) );
  OAI211_X1 U22510 ( .C1(n19480), .C2(n19464), .A(n19463), .B(n19883), .ZN(
        n19482) );
  INV_X1 U22511 ( .A(n19485), .ZN(n19477) );
  AOI22_X1 U22512 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19482), .B1(
        n19477), .B2(n19886), .ZN(n19465) );
  OAI211_X1 U22513 ( .C1(n19803), .C2(n19490), .A(n19466), .B(n19465), .ZN(
        P2_U3056) );
  AOI22_X1 U22514 ( .A1(n19481), .A2(n19916), .B1(n19915), .B2(n19480), .ZN(
        n19468) );
  AOI22_X1 U22515 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19482), .B1(
        n19513), .B2(n19918), .ZN(n19467) );
  OAI211_X1 U22516 ( .C1(n19847), .C2(n19485), .A(n19468), .B(n19467), .ZN(
        P2_U3057) );
  AOI22_X1 U22517 ( .A1(n19481), .A2(n19922), .B1(n19921), .B2(n19480), .ZN(
        n19470) );
  AOI22_X1 U22518 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19482), .B1(
        n19477), .B2(n19923), .ZN(n19469) );
  OAI211_X1 U22519 ( .C1(n19809), .C2(n19490), .A(n19470), .B(n19469), .ZN(
        P2_U3058) );
  AOI22_X1 U22520 ( .A1(n19481), .A2(n19929), .B1(n19928), .B2(n19480), .ZN(
        n19472) );
  AOI22_X1 U22521 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19482), .B1(
        n19477), .B2(n19931), .ZN(n19471) );
  OAI211_X1 U22522 ( .C1(n19812), .C2(n19490), .A(n19472), .B(n19471), .ZN(
        P2_U3059) );
  AOI22_X1 U22523 ( .A1(n19481), .A2(n19935), .B1(n19934), .B2(n19480), .ZN(
        n19474) );
  AOI22_X1 U22524 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19482), .B1(
        n19477), .B2(n19936), .ZN(n19473) );
  OAI211_X1 U22525 ( .C1(n19815), .C2(n19490), .A(n19474), .B(n19473), .ZN(
        P2_U3060) );
  AOI22_X1 U22526 ( .A1(n19481), .A2(n19942), .B1(n19941), .B2(n19480), .ZN(
        n19476) );
  INV_X1 U22527 ( .A(n19818), .ZN(n19943) );
  AOI22_X1 U22528 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19482), .B1(
        n19513), .B2(n19943), .ZN(n19475) );
  OAI211_X1 U22529 ( .C1(n19859), .C2(n19485), .A(n19476), .B(n19475), .ZN(
        P2_U3061) );
  AOI22_X1 U22530 ( .A1(n19481), .A2(n19948), .B1(n19947), .B2(n19480), .ZN(
        n19479) );
  AOI22_X1 U22531 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19482), .B1(
        n19477), .B2(n19950), .ZN(n19478) );
  OAI211_X1 U22532 ( .C1(n19821), .C2(n19490), .A(n19479), .B(n19478), .ZN(
        P2_U3062) );
  AOI22_X1 U22533 ( .A1(n19481), .A2(n19955), .B1(n19953), .B2(n19480), .ZN(
        n19484) );
  AOI22_X1 U22534 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19482), .B1(
        n19513), .B2(n19959), .ZN(n19483) );
  OAI211_X1 U22535 ( .C1(n19868), .C2(n19485), .A(n19484), .B(n19483), .ZN(
        P2_U3063) );
  INV_X1 U22536 ( .A(n19486), .ZN(n19489) );
  NOR2_X1 U22537 ( .A1(n19726), .A2(n19518), .ZN(n19511) );
  OAI21_X1 U22538 ( .B1(n19489), .B2(n19511), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19488) );
  NOR2_X1 U22539 ( .A1(n19729), .A2(n19518), .ZN(n19491) );
  INV_X1 U22540 ( .A(n19491), .ZN(n19487) );
  NAND2_X1 U22541 ( .A1(n19488), .A2(n19487), .ZN(n19512) );
  AOI22_X1 U22542 ( .A1(n19833), .A2(n19512), .B1(n19876), .B2(n19511), .ZN(
        n19498) );
  INV_X1 U22543 ( .A(n19511), .ZN(n19495) );
  OAI21_X1 U22544 ( .B1(n19489), .B2(n20113), .A(n19879), .ZN(n19494) );
  AOI21_X1 U22545 ( .B1(n19540), .B2(n19490), .A(n20107), .ZN(n19492) );
  NOR3_X1 U22546 ( .A1(n19492), .A2(n19491), .A3(n19694), .ZN(n19493) );
  AOI211_X1 U22547 ( .C1(n19495), .C2(n19494), .A(n19796), .B(n19493), .ZN(
        n19496) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19886), .ZN(n19497) );
  OAI211_X1 U22549 ( .C1(n19803), .C2(n19540), .A(n19498), .B(n19497), .ZN(
        P2_U3064) );
  AOI22_X1 U22550 ( .A1(n19512), .A2(n19916), .B1(n19915), .B2(n19511), .ZN(
        n19500) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19917), .ZN(n19499) );
  OAI211_X1 U22552 ( .C1(n19806), .C2(n19540), .A(n19500), .B(n19499), .ZN(
        P2_U3065) );
  AOI22_X1 U22553 ( .A1(n19512), .A2(n19922), .B1(n19921), .B2(n19511), .ZN(
        n19502) );
  AOI22_X1 U22554 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19923), .ZN(n19501) );
  OAI211_X1 U22555 ( .C1(n19809), .C2(n19540), .A(n19502), .B(n19501), .ZN(
        P2_U3066) );
  AOI22_X1 U22556 ( .A1(n19512), .A2(n19929), .B1(n19928), .B2(n19511), .ZN(
        n19504) );
  AOI22_X1 U22557 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19931), .ZN(n19503) );
  OAI211_X1 U22558 ( .C1(n19812), .C2(n19540), .A(n19504), .B(n19503), .ZN(
        P2_U3067) );
  AOI22_X1 U22559 ( .A1(n19935), .A2(n19512), .B1(n19934), .B2(n19511), .ZN(
        n19506) );
  AOI22_X1 U22560 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19936), .ZN(n19505) );
  OAI211_X1 U22561 ( .C1(n19815), .C2(n19540), .A(n19506), .B(n19505), .ZN(
        P2_U3068) );
  AOI22_X1 U22562 ( .A1(n19512), .A2(n19942), .B1(n19941), .B2(n19511), .ZN(
        n19508) );
  AOI22_X1 U22563 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19944), .ZN(n19507) );
  OAI211_X1 U22564 ( .C1(n19818), .C2(n19540), .A(n19508), .B(n19507), .ZN(
        P2_U3069) );
  AOI22_X1 U22565 ( .A1(n19512), .A2(n19948), .B1(n19947), .B2(n19511), .ZN(
        n19510) );
  AOI22_X1 U22566 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19950), .ZN(n19509) );
  OAI211_X1 U22567 ( .C1(n19821), .C2(n19540), .A(n19510), .B(n19509), .ZN(
        P2_U3070) );
  AOI22_X1 U22568 ( .A1(n19512), .A2(n19955), .B1(n19953), .B2(n19511), .ZN(
        n19516) );
  AOI22_X1 U22569 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19957), .ZN(n19515) );
  OAI211_X1 U22570 ( .C1(n19828), .C2(n19540), .A(n19516), .B(n19515), .ZN(
        P2_U3071) );
  INV_X1 U22571 ( .A(n19886), .ZN(n19844) );
  NOR2_X1 U22572 ( .A1(n19517), .A2(n19518), .ZN(n19543) );
  AOI22_X1 U22573 ( .A1(n19877), .A2(n19576), .B1(n19876), .B2(n19543), .ZN(
        n19529) );
  INV_X1 U22574 ( .A(n20060), .ZN(n19761) );
  OAI21_X1 U22575 ( .B1(n19581), .B2(n19761), .A(n20064), .ZN(n19527) );
  NOR2_X1 U22576 ( .A1(n20085), .A2(n19518), .ZN(n19523) );
  INV_X1 U22577 ( .A(n19519), .ZN(n19524) );
  OAI21_X1 U22578 ( .B1(n19524), .B2(n20113), .A(n19879), .ZN(n19521) );
  INV_X1 U22579 ( .A(n19543), .ZN(n19520) );
  AOI21_X1 U22580 ( .B1(n19521), .B2(n19520), .A(n19796), .ZN(n19522) );
  OAI21_X1 U22581 ( .B1(n19527), .B2(n19523), .A(n19522), .ZN(n19546) );
  INV_X1 U22582 ( .A(n19523), .ZN(n19526) );
  OAI21_X1 U22583 ( .B1(n19524), .B2(n19543), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19525) );
  OAI21_X1 U22584 ( .B1(n19527), .B2(n19526), .A(n19525), .ZN(n19545) );
  AOI22_X1 U22585 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19546), .B1(
        n19833), .B2(n19545), .ZN(n19528) );
  OAI211_X1 U22586 ( .C1(n19844), .C2(n19540), .A(n19529), .B(n19528), .ZN(
        P2_U3072) );
  INV_X1 U22587 ( .A(n19540), .ZN(n19544) );
  AOI22_X1 U22588 ( .A1(n19917), .A2(n19544), .B1(n19543), .B2(n19915), .ZN(
        n19531) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19546), .B1(
        n19916), .B2(n19545), .ZN(n19530) );
  OAI211_X1 U22590 ( .C1(n19806), .C2(n19554), .A(n19531), .B(n19530), .ZN(
        P2_U3073) );
  AOI22_X1 U22591 ( .A1(n19923), .A2(n19544), .B1(n19543), .B2(n19921), .ZN(
        n19533) );
  AOI22_X1 U22592 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19546), .B1(
        n19922), .B2(n19545), .ZN(n19532) );
  OAI211_X1 U22593 ( .C1(n19809), .C2(n19554), .A(n19533), .B(n19532), .ZN(
        P2_U3074) );
  INV_X1 U22594 ( .A(n19931), .ZN(n19853) );
  INV_X1 U22595 ( .A(n19812), .ZN(n19930) );
  AOI22_X1 U22596 ( .A1(n19930), .A2(n19576), .B1(n19543), .B2(n19928), .ZN(
        n19535) );
  AOI22_X1 U22597 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19546), .B1(
        n19929), .B2(n19545), .ZN(n19534) );
  OAI211_X1 U22598 ( .C1(n19853), .C2(n19540), .A(n19535), .B(n19534), .ZN(
        P2_U3075) );
  AOI22_X1 U22599 ( .A1(n19936), .A2(n19544), .B1(n19543), .B2(n19934), .ZN(
        n19537) );
  AOI22_X1 U22600 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19546), .B1(
        n19935), .B2(n19545), .ZN(n19536) );
  OAI211_X1 U22601 ( .C1(n19815), .C2(n19554), .A(n19537), .B(n19536), .ZN(
        P2_U3076) );
  AOI22_X1 U22602 ( .A1(n19943), .A2(n19576), .B1(n19543), .B2(n19941), .ZN(
        n19539) );
  AOI22_X1 U22603 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19546), .B1(
        n19942), .B2(n19545), .ZN(n19538) );
  OAI211_X1 U22604 ( .C1(n19859), .C2(n19540), .A(n19539), .B(n19538), .ZN(
        P2_U3077) );
  AOI22_X1 U22605 ( .A1(n19950), .A2(n19544), .B1(n19543), .B2(n19947), .ZN(
        n19542) );
  AOI22_X1 U22606 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19546), .B1(
        n19948), .B2(n19545), .ZN(n19541) );
  OAI211_X1 U22607 ( .C1(n19821), .C2(n19554), .A(n19542), .B(n19541), .ZN(
        P2_U3078) );
  AOI22_X1 U22608 ( .A1(n19957), .A2(n19544), .B1(n19543), .B2(n19953), .ZN(
        n19548) );
  AOI22_X1 U22609 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19546), .B1(
        n19955), .B2(n19545), .ZN(n19547) );
  OAI211_X1 U22610 ( .C1(n19828), .C2(n19554), .A(n19548), .B(n19547), .ZN(
        P2_U3079) );
  NAND3_X1 U22611 ( .A1(n19611), .A2(n20085), .A3(n20092), .ZN(n19555) );
  AND3_X1 U22612 ( .A1(n19556), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19555), 
        .ZN(n19553) );
  NAND2_X1 U22613 ( .A1(n19551), .A2(n19550), .ZN(n19792) );
  NOR2_X1 U22614 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19792), .ZN(
        n19559) );
  AOI21_X1 U22615 ( .B1(n19559), .B2(n19879), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19552) );
  NOR2_X1 U22616 ( .A1(n19553), .A2(n19552), .ZN(n19575) );
  INV_X1 U22617 ( .A(n19555), .ZN(n19574) );
  AOI22_X1 U22618 ( .A1(n19575), .A2(n19833), .B1(n19876), .B2(n19574), .ZN(
        n19561) );
  AOI21_X1 U22619 ( .B1(n19554), .B2(n19610), .A(n20107), .ZN(n19558) );
  OAI211_X1 U22620 ( .C1(n19556), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19555), 
        .B(n19694), .ZN(n19557) );
  OAI211_X1 U22621 ( .C1(n19559), .C2(n19558), .A(n19883), .B(n19557), .ZN(
        n19577) );
  AOI22_X1 U22622 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19577), .B1(
        n19576), .B2(n19886), .ZN(n19560) );
  OAI211_X1 U22623 ( .C1(n19803), .C2(n19610), .A(n19561), .B(n19560), .ZN(
        P2_U3080) );
  AOI22_X1 U22624 ( .A1(n19575), .A2(n19916), .B1(n19915), .B2(n19574), .ZN(
        n19563) );
  AOI22_X1 U22625 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19577), .B1(
        n19576), .B2(n19917), .ZN(n19562) );
  OAI211_X1 U22626 ( .C1(n19806), .C2(n19610), .A(n19563), .B(n19562), .ZN(
        P2_U3081) );
  AOI22_X1 U22627 ( .A1(n19575), .A2(n19922), .B1(n19921), .B2(n19574), .ZN(
        n19565) );
  AOI22_X1 U22628 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19577), .B1(
        n19576), .B2(n19923), .ZN(n19564) );
  OAI211_X1 U22629 ( .C1(n19809), .C2(n19610), .A(n19565), .B(n19564), .ZN(
        P2_U3082) );
  AOI22_X1 U22630 ( .A1(n19575), .A2(n19929), .B1(n19928), .B2(n19574), .ZN(
        n19567) );
  AOI22_X1 U22631 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19577), .B1(
        n19576), .B2(n19931), .ZN(n19566) );
  OAI211_X1 U22632 ( .C1(n19812), .C2(n19610), .A(n19567), .B(n19566), .ZN(
        P2_U3083) );
  AOI22_X1 U22633 ( .A1(n19575), .A2(n19935), .B1(n19934), .B2(n19574), .ZN(
        n19569) );
  AOI22_X1 U22634 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19577), .B1(
        n19576), .B2(n19936), .ZN(n19568) );
  OAI211_X1 U22635 ( .C1(n19815), .C2(n19610), .A(n19569), .B(n19568), .ZN(
        P2_U3084) );
  AOI22_X1 U22636 ( .A1(n19575), .A2(n19942), .B1(n19941), .B2(n19574), .ZN(
        n19571) );
  AOI22_X1 U22637 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19577), .B1(
        n19576), .B2(n19944), .ZN(n19570) );
  OAI211_X1 U22638 ( .C1(n19818), .C2(n19610), .A(n19571), .B(n19570), .ZN(
        P2_U3085) );
  AOI22_X1 U22639 ( .A1(n19575), .A2(n19948), .B1(n19947), .B2(n19574), .ZN(
        n19573) );
  AOI22_X1 U22640 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19577), .B1(
        n19576), .B2(n19950), .ZN(n19572) );
  OAI211_X1 U22641 ( .C1(n19821), .C2(n19610), .A(n19573), .B(n19572), .ZN(
        P2_U3086) );
  AOI22_X1 U22642 ( .A1(n19575), .A2(n19955), .B1(n19953), .B2(n19574), .ZN(
        n19579) );
  AOI22_X1 U22643 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19577), .B1(
        n19576), .B2(n19957), .ZN(n19578) );
  OAI211_X1 U22644 ( .C1(n19828), .C2(n19610), .A(n19579), .B(n19578), .ZN(
        P2_U3087) );
  INV_X1 U22645 ( .A(n19611), .ZN(n19613) );
  NOR2_X1 U22646 ( .A1(n19693), .A2(n19613), .ZN(n19605) );
  AOI22_X1 U22647 ( .A1(n19877), .A2(n19637), .B1(n19876), .B2(n19605), .ZN(
        n19591) );
  OAI21_X1 U22648 ( .B1(n19581), .B2(n19840), .A(n20064), .ZN(n19589) );
  NAND2_X1 U22649 ( .A1(n20085), .A2(n19611), .ZN(n19588) );
  INV_X1 U22650 ( .A(n19588), .ZN(n19584) );
  INV_X1 U22651 ( .A(n19605), .ZN(n19582) );
  OAI211_X1 U22652 ( .C1(n19585), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19694), 
        .B(n19582), .ZN(n19583) );
  OAI211_X1 U22653 ( .C1(n19589), .C2(n19584), .A(n19883), .B(n19583), .ZN(
        n19607) );
  INV_X1 U22654 ( .A(n19585), .ZN(n19586) );
  OAI21_X1 U22655 ( .B1(n19586), .B2(n19605), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19587) );
  OAI21_X1 U22656 ( .B1(n19589), .B2(n19588), .A(n19587), .ZN(n19606) );
  AOI22_X1 U22657 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19607), .B1(
        n19833), .B2(n19606), .ZN(n19590) );
  OAI211_X1 U22658 ( .C1(n19844), .C2(n19610), .A(n19591), .B(n19590), .ZN(
        P2_U3088) );
  INV_X1 U22659 ( .A(n19610), .ZN(n19598) );
  AOI22_X1 U22660 ( .A1(n19917), .A2(n19598), .B1(n19915), .B2(n19605), .ZN(
        n19593) );
  AOI22_X1 U22661 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19607), .B1(
        n19916), .B2(n19606), .ZN(n19592) );
  OAI211_X1 U22662 ( .C1(n19806), .C2(n19634), .A(n19593), .B(n19592), .ZN(
        P2_U3089) );
  AOI22_X1 U22663 ( .A1(n19924), .A2(n19637), .B1(n19921), .B2(n19605), .ZN(
        n19595) );
  AOI22_X1 U22664 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19607), .B1(
        n19922), .B2(n19606), .ZN(n19594) );
  OAI211_X1 U22665 ( .C1(n19850), .C2(n19610), .A(n19595), .B(n19594), .ZN(
        P2_U3090) );
  AOI22_X1 U22666 ( .A1(n19930), .A2(n19637), .B1(n19928), .B2(n19605), .ZN(
        n19597) );
  AOI22_X1 U22667 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19607), .B1(
        n19929), .B2(n19606), .ZN(n19596) );
  OAI211_X1 U22668 ( .C1(n19853), .C2(n19610), .A(n19597), .B(n19596), .ZN(
        P2_U3091) );
  AOI22_X1 U22669 ( .A1(n19936), .A2(n19598), .B1(n19934), .B2(n19605), .ZN(
        n19600) );
  AOI22_X1 U22670 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19607), .B1(
        n19935), .B2(n19606), .ZN(n19599) );
  OAI211_X1 U22671 ( .C1(n19815), .C2(n19634), .A(n19600), .B(n19599), .ZN(
        P2_U3092) );
  AOI22_X1 U22672 ( .A1(n19943), .A2(n19637), .B1(n19941), .B2(n19605), .ZN(
        n19602) );
  AOI22_X1 U22673 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19607), .B1(
        n19942), .B2(n19606), .ZN(n19601) );
  OAI211_X1 U22674 ( .C1(n19859), .C2(n19610), .A(n19602), .B(n19601), .ZN(
        P2_U3093) );
  INV_X1 U22675 ( .A(n19821), .ZN(n19949) );
  AOI22_X1 U22676 ( .A1(n19949), .A2(n19637), .B1(n19947), .B2(n19605), .ZN(
        n19604) );
  AOI22_X1 U22677 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19607), .B1(
        n19948), .B2(n19606), .ZN(n19603) );
  OAI211_X1 U22678 ( .C1(n19862), .C2(n19610), .A(n19604), .B(n19603), .ZN(
        P2_U3094) );
  AOI22_X1 U22679 ( .A1(n19959), .A2(n19637), .B1(n19953), .B2(n19605), .ZN(
        n19609) );
  AOI22_X1 U22680 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19607), .B1(
        n19955), .B2(n19606), .ZN(n19608) );
  OAI211_X1 U22681 ( .C1(n19868), .C2(n19610), .A(n19609), .B(n19608), .ZN(
        P2_U3095) );
  NAND2_X1 U22682 ( .A1(n19612), .A2(n19611), .ZN(n19617) );
  INV_X1 U22683 ( .A(n11184), .ZN(n19614) );
  NOR2_X1 U22684 ( .A1(n19726), .A2(n19613), .ZN(n19635) );
  NOR3_X1 U22685 ( .A1(n19614), .A2(n19635), .A3(n20113), .ZN(n19616) );
  AOI211_X2 U22686 ( .C1(n20113), .C2(n19617), .A(n19615), .B(n19616), .ZN(
        n19636) );
  AOI22_X1 U22687 ( .A1(n19636), .A2(n19833), .B1(n19876), .B2(n19635), .ZN(
        n19621) );
  OAI21_X1 U22688 ( .B1(n19637), .B2(n19658), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19618) );
  AOI211_X1 U22689 ( .C1(n19618), .C2(n19617), .A(n19796), .B(n19616), .ZN(
        n19619) );
  AOI22_X1 U22690 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19638), .B1(
        n19637), .B2(n19886), .ZN(n19620) );
  OAI211_X1 U22691 ( .C1(n19803), .C2(n19645), .A(n19621), .B(n19620), .ZN(
        P2_U3096) );
  AOI22_X1 U22692 ( .A1(n19636), .A2(n19916), .B1(n19915), .B2(n19635), .ZN(
        n19623) );
  AOI22_X1 U22693 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19638), .B1(
        n19637), .B2(n19917), .ZN(n19622) );
  OAI211_X1 U22694 ( .C1(n19806), .C2(n19645), .A(n19623), .B(n19622), .ZN(
        P2_U3097) );
  AOI22_X1 U22695 ( .A1(n19636), .A2(n19922), .B1(n19921), .B2(n19635), .ZN(
        n19625) );
  AOI22_X1 U22696 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19638), .B1(
        n19658), .B2(n19924), .ZN(n19624) );
  OAI211_X1 U22697 ( .C1(n19850), .C2(n19634), .A(n19625), .B(n19624), .ZN(
        P2_U3098) );
  AOI22_X1 U22698 ( .A1(n19636), .A2(n19929), .B1(n19928), .B2(n19635), .ZN(
        n19627) );
  AOI22_X1 U22699 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19638), .B1(
        n19637), .B2(n19931), .ZN(n19626) );
  OAI211_X1 U22700 ( .C1(n19812), .C2(n19645), .A(n19627), .B(n19626), .ZN(
        P2_U3099) );
  AOI22_X1 U22701 ( .A1(n19636), .A2(n19935), .B1(n19934), .B2(n19635), .ZN(
        n19629) );
  AOI22_X1 U22702 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19638), .B1(
        n19658), .B2(n19937), .ZN(n19628) );
  OAI211_X1 U22703 ( .C1(n19856), .C2(n19634), .A(n19629), .B(n19628), .ZN(
        P2_U3100) );
  AOI22_X1 U22704 ( .A1(n19636), .A2(n19942), .B1(n19941), .B2(n19635), .ZN(
        n19631) );
  AOI22_X1 U22705 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19638), .B1(
        n19658), .B2(n19943), .ZN(n19630) );
  OAI211_X1 U22706 ( .C1(n19859), .C2(n19634), .A(n19631), .B(n19630), .ZN(
        P2_U3101) );
  AOI22_X1 U22707 ( .A1(n19636), .A2(n19948), .B1(n19947), .B2(n19635), .ZN(
        n19633) );
  AOI22_X1 U22708 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19638), .B1(
        n19658), .B2(n19949), .ZN(n19632) );
  OAI211_X1 U22709 ( .C1(n19862), .C2(n19634), .A(n19633), .B(n19632), .ZN(
        P2_U3102) );
  AOI22_X1 U22710 ( .A1(n19636), .A2(n19955), .B1(n19953), .B2(n19635), .ZN(
        n19640) );
  AOI22_X1 U22711 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19638), .B1(
        n19637), .B2(n19957), .ZN(n19639) );
  OAI211_X1 U22712 ( .C1(n19828), .C2(n19645), .A(n19640), .B(n19639), .ZN(
        P2_U3103) );
  INV_X1 U22713 ( .A(n19664), .ZN(n19667) );
  AOI22_X1 U22714 ( .A1(n19657), .A2(n19916), .B1(n19667), .B2(n19915), .ZN(
        n19642) );
  AOI22_X1 U22715 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19659), .B1(
        n19683), .B2(n19918), .ZN(n19641) );
  OAI211_X1 U22716 ( .C1(n19847), .C2(n19645), .A(n19642), .B(n19641), .ZN(
        P2_U3105) );
  AOI22_X1 U22717 ( .A1(n19657), .A2(n19922), .B1(n19667), .B2(n19921), .ZN(
        n19644) );
  AOI22_X1 U22718 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19659), .B1(
        n19683), .B2(n19924), .ZN(n19643) );
  OAI211_X1 U22719 ( .C1(n19850), .C2(n19645), .A(n19644), .B(n19643), .ZN(
        P2_U3106) );
  AOI22_X1 U22720 ( .A1(n19657), .A2(n19929), .B1(n19667), .B2(n19928), .ZN(
        n19647) );
  AOI22_X1 U22721 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19659), .B1(
        n19658), .B2(n19931), .ZN(n19646) );
  OAI211_X1 U22722 ( .C1(n19812), .C2(n19691), .A(n19647), .B(n19646), .ZN(
        P2_U3107) );
  INV_X1 U22723 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n19650) );
  AOI22_X1 U22724 ( .A1(n19657), .A2(n19935), .B1(n19667), .B2(n19934), .ZN(
        n19649) );
  AOI22_X1 U22725 ( .A1(n19683), .A2(n19937), .B1(n19658), .B2(n19936), .ZN(
        n19648) );
  OAI211_X1 U22726 ( .C1(n19656), .C2(n19650), .A(n19649), .B(n19648), .ZN(
        P2_U3108) );
  AOI22_X1 U22727 ( .A1(n19657), .A2(n19942), .B1(n19667), .B2(n19941), .ZN(
        n19652) );
  AOI22_X1 U22728 ( .A1(n19683), .A2(n19943), .B1(n19658), .B2(n19944), .ZN(
        n19651) );
  OAI211_X1 U22729 ( .C1(n19656), .C2(n11176), .A(n19652), .B(n19651), .ZN(
        P2_U3109) );
  INV_X1 U22730 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n19655) );
  AOI22_X1 U22731 ( .A1(n19657), .A2(n19948), .B1(n19667), .B2(n19947), .ZN(
        n19654) );
  AOI22_X1 U22732 ( .A1(n19683), .A2(n19949), .B1(n19658), .B2(n19950), .ZN(
        n19653) );
  OAI211_X1 U22733 ( .C1(n19656), .C2(n19655), .A(n19654), .B(n19653), .ZN(
        P2_U3110) );
  AOI22_X1 U22734 ( .A1(n19657), .A2(n19955), .B1(n19667), .B2(n19953), .ZN(
        n19661) );
  AOI22_X1 U22735 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19659), .B1(
        n19658), .B2(n19957), .ZN(n19660) );
  OAI211_X1 U22736 ( .C1(n19828), .C2(n19691), .A(n19661), .B(n19660), .ZN(
        P2_U3111) );
  NAND2_X1 U22737 ( .A1(n20076), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19763) );
  OR2_X1 U22738 ( .A1(n19763), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19702) );
  NOR2_X1 U22739 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19702), .ZN(
        n19686) );
  AOI22_X1 U22740 ( .A1(n19886), .A2(n19683), .B1(n19876), .B2(n19686), .ZN(
        n19672) );
  NAND3_X1 U22741 ( .A1(n19691), .A2(n20064), .A3(n19718), .ZN(n19662) );
  NAND2_X1 U22742 ( .A1(n19662), .A2(n19871), .ZN(n19666) );
  INV_X1 U22743 ( .A(n11177), .ZN(n19668) );
  OAI21_X1 U22744 ( .B1(n19668), .B2(n20113), .A(n19879), .ZN(n19663) );
  AOI21_X1 U22745 ( .B1(n19666), .B2(n19664), .A(n19663), .ZN(n19665) );
  OAI21_X1 U22746 ( .B1(n19667), .B2(n19686), .A(n19666), .ZN(n19670) );
  OAI21_X1 U22747 ( .B1(n19668), .B2(n19686), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19669) );
  NAND2_X1 U22748 ( .A1(n19670), .A2(n19669), .ZN(n19687) );
  AOI22_X1 U22749 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19688), .B1(
        n19833), .B2(n19687), .ZN(n19671) );
  OAI211_X1 U22750 ( .C1(n19803), .C2(n19718), .A(n19672), .B(n19671), .ZN(
        P2_U3112) );
  AOI22_X1 U22751 ( .A1(n19918), .A2(n19719), .B1(n19686), .B2(n19915), .ZN(
        n19674) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19688), .B1(
        n19916), .B2(n19687), .ZN(n19673) );
  OAI211_X1 U22753 ( .C1(n19847), .C2(n19691), .A(n19674), .B(n19673), .ZN(
        P2_U3113) );
  AOI22_X1 U22754 ( .A1(n19924), .A2(n19719), .B1(n19686), .B2(n19921), .ZN(
        n19676) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19688), .B1(
        n19922), .B2(n19687), .ZN(n19675) );
  OAI211_X1 U22756 ( .C1(n19850), .C2(n19691), .A(n19676), .B(n19675), .ZN(
        P2_U3114) );
  AOI22_X1 U22757 ( .A1(n19931), .A2(n19683), .B1(n19686), .B2(n19928), .ZN(
        n19678) );
  AOI22_X1 U22758 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19688), .B1(
        n19929), .B2(n19687), .ZN(n19677) );
  OAI211_X1 U22759 ( .C1(n19812), .C2(n19718), .A(n19678), .B(n19677), .ZN(
        P2_U3115) );
  AOI22_X1 U22760 ( .A1(n19937), .A2(n19719), .B1(n19686), .B2(n19934), .ZN(
        n19680) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19688), .B1(
        n19935), .B2(n19687), .ZN(n19679) );
  OAI211_X1 U22762 ( .C1(n19856), .C2(n19691), .A(n19680), .B(n19679), .ZN(
        P2_U3116) );
  AOI22_X1 U22763 ( .A1(n19944), .A2(n19683), .B1(n19686), .B2(n19941), .ZN(
        n19682) );
  AOI22_X1 U22764 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19688), .B1(
        n19942), .B2(n19687), .ZN(n19681) );
  OAI211_X1 U22765 ( .C1(n19818), .C2(n19718), .A(n19682), .B(n19681), .ZN(
        P2_U3117) );
  AOI22_X1 U22766 ( .A1(n19950), .A2(n19683), .B1(n19686), .B2(n19947), .ZN(
        n19685) );
  AOI22_X1 U22767 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19688), .B1(
        n19948), .B2(n19687), .ZN(n19684) );
  OAI211_X1 U22768 ( .C1(n19821), .C2(n19718), .A(n19685), .B(n19684), .ZN(
        P2_U3118) );
  AOI22_X1 U22769 ( .A1(n19959), .A2(n19719), .B1(n19686), .B2(n19953), .ZN(
        n19690) );
  AOI22_X1 U22770 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19688), .B1(
        n19955), .B2(n19687), .ZN(n19689) );
  OAI211_X1 U22771 ( .C1(n19868), .C2(n19691), .A(n19690), .B(n19689), .ZN(
        P2_U3119) );
  NOR2_X1 U22772 ( .A1(n19693), .A2(n19763), .ZN(n19730) );
  AOI22_X1 U22773 ( .A1(n19886), .A2(n19719), .B1(n19876), .B2(n19730), .ZN(
        n19705) );
  AOI21_X1 U22774 ( .B1(n19699), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19697) );
  AOI21_X1 U22775 ( .B1(n19835), .B2(n19695), .A(n19694), .ZN(n19698) );
  NAND2_X1 U22776 ( .A1(n19698), .A2(n19702), .ZN(n19696) );
  OAI211_X1 U22777 ( .C1(n19730), .C2(n19697), .A(n19696), .B(n19883), .ZN(
        n19721) );
  INV_X1 U22778 ( .A(n19698), .ZN(n19703) );
  INV_X1 U22779 ( .A(n19699), .ZN(n19700) );
  OAI21_X1 U22780 ( .B1(n19700), .B2(n19730), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19701) );
  OAI21_X1 U22781 ( .B1(n19703), .B2(n19702), .A(n19701), .ZN(n19720) );
  AOI22_X1 U22782 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19721), .B1(
        n19833), .B2(n19720), .ZN(n19704) );
  OAI211_X1 U22783 ( .C1(n19803), .C2(n19724), .A(n19705), .B(n19704), .ZN(
        P2_U3120) );
  AOI22_X1 U22784 ( .A1(n19917), .A2(n19719), .B1(n19915), .B2(n19730), .ZN(
        n19707) );
  AOI22_X1 U22785 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19721), .B1(
        n19916), .B2(n19720), .ZN(n19706) );
  OAI211_X1 U22786 ( .C1(n19806), .C2(n19724), .A(n19707), .B(n19706), .ZN(
        P2_U3121) );
  AOI22_X1 U22787 ( .A1(n19924), .A2(n19751), .B1(n19921), .B2(n19730), .ZN(
        n19709) );
  AOI22_X1 U22788 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19721), .B1(
        n19922), .B2(n19720), .ZN(n19708) );
  OAI211_X1 U22789 ( .C1(n19850), .C2(n19718), .A(n19709), .B(n19708), .ZN(
        P2_U3122) );
  AOI22_X1 U22790 ( .A1(n19930), .A2(n19751), .B1(n19730), .B2(n19928), .ZN(
        n19711) );
  AOI22_X1 U22791 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19721), .B1(
        n19929), .B2(n19720), .ZN(n19710) );
  OAI211_X1 U22792 ( .C1(n19853), .C2(n19718), .A(n19711), .B(n19710), .ZN(
        P2_U3123) );
  AOI22_X1 U22793 ( .A1(n19937), .A2(n19751), .B1(n19934), .B2(n19730), .ZN(
        n19713) );
  AOI22_X1 U22794 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19721), .B1(
        n19935), .B2(n19720), .ZN(n19712) );
  OAI211_X1 U22795 ( .C1(n19856), .C2(n19718), .A(n19713), .B(n19712), .ZN(
        P2_U3124) );
  AOI22_X1 U22796 ( .A1(n19943), .A2(n19751), .B1(n19730), .B2(n19941), .ZN(
        n19715) );
  AOI22_X1 U22797 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19721), .B1(
        n19942), .B2(n19720), .ZN(n19714) );
  OAI211_X1 U22798 ( .C1(n19859), .C2(n19718), .A(n19715), .B(n19714), .ZN(
        P2_U3125) );
  AOI22_X1 U22799 ( .A1(n19949), .A2(n19751), .B1(n19730), .B2(n19947), .ZN(
        n19717) );
  AOI22_X1 U22800 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19721), .B1(
        n19948), .B2(n19720), .ZN(n19716) );
  OAI211_X1 U22801 ( .C1(n19862), .C2(n19718), .A(n19717), .B(n19716), .ZN(
        P2_U3126) );
  AOI22_X1 U22802 ( .A1(n19957), .A2(n19719), .B1(n19953), .B2(n19730), .ZN(
        n19723) );
  AOI22_X1 U22803 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19721), .B1(
        n19955), .B2(n19720), .ZN(n19722) );
  OAI211_X1 U22804 ( .C1(n19828), .C2(n19724), .A(n19723), .B(n19722), .ZN(
        P2_U3127) );
  INV_X1 U22805 ( .A(n19731), .ZN(n19727) );
  NOR2_X1 U22806 ( .A1(n19726), .A2(n19763), .ZN(n19749) );
  OAI21_X1 U22807 ( .B1(n19727), .B2(n19749), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19728) );
  OAI21_X1 U22808 ( .B1(n19763), .B2(n19729), .A(n19728), .ZN(n19750) );
  AOI22_X1 U22809 ( .A1(n19833), .A2(n19750), .B1(n19876), .B2(n19749), .ZN(
        n19736) );
  AOI221_X1 U22810 ( .B1(n19751), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19780), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19730), .ZN(n19732) );
  MUX2_X1 U22811 ( .A(n19732), .B(n19731), .S(P2_STATE2_REG_2__SCAN_IN), .Z(
        n19733) );
  NOR2_X1 U22812 ( .A1(n19733), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19734) );
  AOI22_X1 U22813 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19752), .B1(
        n19751), .B2(n19886), .ZN(n19735) );
  OAI211_X1 U22814 ( .C1(n19803), .C2(n19788), .A(n19736), .B(n19735), .ZN(
        P2_U3128) );
  AOI22_X1 U22815 ( .A1(n19750), .A2(n19916), .B1(n19915), .B2(n19749), .ZN(
        n19738) );
  AOI22_X1 U22816 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19752), .B1(
        n19751), .B2(n19917), .ZN(n19737) );
  OAI211_X1 U22817 ( .C1(n19806), .C2(n19788), .A(n19738), .B(n19737), .ZN(
        P2_U3129) );
  AOI22_X1 U22818 ( .A1(n19750), .A2(n19922), .B1(n19921), .B2(n19749), .ZN(
        n19740) );
  AOI22_X1 U22819 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19752), .B1(
        n19751), .B2(n19923), .ZN(n19739) );
  OAI211_X1 U22820 ( .C1(n19809), .C2(n19788), .A(n19740), .B(n19739), .ZN(
        P2_U3130) );
  AOI22_X1 U22821 ( .A1(n19750), .A2(n19929), .B1(n19928), .B2(n19749), .ZN(
        n19742) );
  AOI22_X1 U22822 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19752), .B1(
        n19751), .B2(n19931), .ZN(n19741) );
  OAI211_X1 U22823 ( .C1(n19812), .C2(n19788), .A(n19742), .B(n19741), .ZN(
        P2_U3131) );
  AOI22_X1 U22824 ( .A1(n19935), .A2(n19750), .B1(n19934), .B2(n19749), .ZN(
        n19744) );
  AOI22_X1 U22825 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19752), .B1(
        n19751), .B2(n19936), .ZN(n19743) );
  OAI211_X1 U22826 ( .C1(n19815), .C2(n19788), .A(n19744), .B(n19743), .ZN(
        P2_U3132) );
  AOI22_X1 U22827 ( .A1(n19750), .A2(n19942), .B1(n19941), .B2(n19749), .ZN(
        n19746) );
  AOI22_X1 U22828 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19752), .B1(
        n19751), .B2(n19944), .ZN(n19745) );
  OAI211_X1 U22829 ( .C1(n19818), .C2(n19788), .A(n19746), .B(n19745), .ZN(
        P2_U3133) );
  AOI22_X1 U22830 ( .A1(n19750), .A2(n19948), .B1(n19947), .B2(n19749), .ZN(
        n19748) );
  AOI22_X1 U22831 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19752), .B1(
        n19751), .B2(n19950), .ZN(n19747) );
  OAI211_X1 U22832 ( .C1(n19821), .C2(n19788), .A(n19748), .B(n19747), .ZN(
        P2_U3134) );
  AOI22_X1 U22833 ( .A1(n19750), .A2(n19955), .B1(n19953), .B2(n19749), .ZN(
        n19754) );
  AOI22_X1 U22834 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19752), .B1(
        n19751), .B2(n19957), .ZN(n19753) );
  OAI211_X1 U22835 ( .C1(n19828), .C2(n19788), .A(n19754), .B(n19753), .ZN(
        P2_U3135) );
  OR3_X1 U22836 ( .A1(n20085), .A2(n19763), .A3(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n19759) );
  INV_X1 U22837 ( .A(n19763), .ZN(n19755) );
  NAND2_X1 U22838 ( .A1(n19756), .A2(n19755), .ZN(n19760) );
  NAND3_X1 U22839 ( .A1(n19757), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19760), 
        .ZN(n19764) );
  INV_X1 U22840 ( .A(n19764), .ZN(n19758) );
  AOI21_X1 U22841 ( .B1(n19759), .B2(n20113), .A(n19758), .ZN(n19784) );
  INV_X1 U22842 ( .A(n19760), .ZN(n19783) );
  AOI22_X1 U22843 ( .A1(n19784), .A2(n19833), .B1(n19876), .B2(n19783), .ZN(
        n19769) );
  INV_X1 U22844 ( .A(n19835), .ZN(n19762) );
  NOR3_X1 U22845 ( .A1(n19762), .A2(P2_STATE2_REG_3__SCAN_IN), .A3(n19761), 
        .ZN(n19766) );
  AOI211_X1 U22846 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20092), .A(n20085), 
        .B(n19763), .ZN(n19765) );
  OAI211_X1 U22847 ( .C1(n19766), .C2(n19765), .A(n19883), .B(n19764), .ZN(
        n19785) );
  INV_X1 U22848 ( .A(n19841), .ZN(n19767) );
  NAND2_X1 U22849 ( .A1(n19767), .A2(n20060), .ZN(n19794) );
  AOI22_X1 U22850 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19785), .B1(
        n19824), .B2(n19877), .ZN(n19768) );
  OAI211_X1 U22851 ( .C1(n19844), .C2(n19788), .A(n19769), .B(n19768), .ZN(
        P2_U3136) );
  AOI22_X1 U22852 ( .A1(n19784), .A2(n19916), .B1(n19915), .B2(n19783), .ZN(
        n19771) );
  AOI22_X1 U22853 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19785), .B1(
        n19780), .B2(n19917), .ZN(n19770) );
  OAI211_X1 U22854 ( .C1(n19806), .C2(n19794), .A(n19771), .B(n19770), .ZN(
        P2_U3137) );
  AOI22_X1 U22855 ( .A1(n19784), .A2(n19922), .B1(n19921), .B2(n19783), .ZN(
        n19773) );
  AOI22_X1 U22856 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19785), .B1(
        n19824), .B2(n19924), .ZN(n19772) );
  OAI211_X1 U22857 ( .C1(n19850), .C2(n19788), .A(n19773), .B(n19772), .ZN(
        P2_U3138) );
  AOI22_X1 U22858 ( .A1(n19784), .A2(n19929), .B1(n19928), .B2(n19783), .ZN(
        n19775) );
  AOI22_X1 U22859 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19785), .B1(
        n19824), .B2(n19930), .ZN(n19774) );
  OAI211_X1 U22860 ( .C1(n19853), .C2(n19788), .A(n19775), .B(n19774), .ZN(
        P2_U3139) );
  AOI22_X1 U22861 ( .A1(n19784), .A2(n19935), .B1(n19934), .B2(n19783), .ZN(
        n19777) );
  AOI22_X1 U22862 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19785), .B1(
        n19824), .B2(n19937), .ZN(n19776) );
  OAI211_X1 U22863 ( .C1(n19856), .C2(n19788), .A(n19777), .B(n19776), .ZN(
        P2_U3140) );
  AOI22_X1 U22864 ( .A1(n19784), .A2(n19942), .B1(n19941), .B2(n19783), .ZN(
        n19779) );
  AOI22_X1 U22865 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19785), .B1(
        n19780), .B2(n19944), .ZN(n19778) );
  OAI211_X1 U22866 ( .C1(n19818), .C2(n19794), .A(n19779), .B(n19778), .ZN(
        P2_U3141) );
  AOI22_X1 U22867 ( .A1(n19784), .A2(n19948), .B1(n19947), .B2(n19783), .ZN(
        n19782) );
  AOI22_X1 U22868 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19785), .B1(
        n19780), .B2(n19950), .ZN(n19781) );
  OAI211_X1 U22869 ( .C1(n19821), .C2(n19794), .A(n19782), .B(n19781), .ZN(
        P2_U3142) );
  AOI22_X1 U22870 ( .A1(n19784), .A2(n19955), .B1(n19953), .B2(n19783), .ZN(
        n19787) );
  AOI22_X1 U22871 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19785), .B1(
        n19824), .B2(n19959), .ZN(n19786) );
  OAI211_X1 U22872 ( .C1(n19868), .C2(n19788), .A(n19787), .B(n19786), .ZN(
        P2_U3143) );
  INV_X1 U22873 ( .A(n19790), .ZN(n19791) );
  NAND3_X1 U22874 ( .A1(n20085), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19837) );
  NOR2_X1 U22875 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19837), .ZN(
        n19822) );
  NOR3_X1 U22876 ( .A1(n19791), .A2(n19822), .A3(n20113), .ZN(n19795) );
  NOR2_X1 U22877 ( .A1(n20069), .A2(n19792), .ZN(n19800) );
  AOI21_X1 U22878 ( .B1(n19800), .B2(n19879), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19793) );
  NOR2_X1 U22879 ( .A1(n19795), .A2(n19793), .ZN(n19823) );
  AOI22_X1 U22880 ( .A1(n19823), .A2(n19833), .B1(n19876), .B2(n19822), .ZN(
        n19802) );
  AOI21_X1 U22881 ( .B1(n19867), .B2(n19794), .A(n20107), .ZN(n19799) );
  INV_X1 U22882 ( .A(n19822), .ZN(n19797) );
  AOI211_X1 U22883 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19797), .A(n19796), 
        .B(n19795), .ZN(n19798) );
  OAI21_X1 U22884 ( .B1(n19800), .B2(n19799), .A(n19798), .ZN(n19825) );
  AOI22_X1 U22885 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19825), .B1(
        n19824), .B2(n19886), .ZN(n19801) );
  OAI211_X1 U22886 ( .C1(n19803), .C2(n19867), .A(n19802), .B(n19801), .ZN(
        P2_U3144) );
  AOI22_X1 U22887 ( .A1(n19823), .A2(n19916), .B1(n19915), .B2(n19822), .ZN(
        n19805) );
  AOI22_X1 U22888 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19825), .B1(
        n19824), .B2(n19917), .ZN(n19804) );
  OAI211_X1 U22889 ( .C1(n19806), .C2(n19867), .A(n19805), .B(n19804), .ZN(
        P2_U3145) );
  AOI22_X1 U22890 ( .A1(n19823), .A2(n19922), .B1(n19921), .B2(n19822), .ZN(
        n19808) );
  AOI22_X1 U22891 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19825), .B1(
        n19824), .B2(n19923), .ZN(n19807) );
  OAI211_X1 U22892 ( .C1(n19809), .C2(n19867), .A(n19808), .B(n19807), .ZN(
        P2_U3146) );
  AOI22_X1 U22893 ( .A1(n19823), .A2(n19929), .B1(n19928), .B2(n19822), .ZN(
        n19811) );
  AOI22_X1 U22894 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19825), .B1(
        n19824), .B2(n19931), .ZN(n19810) );
  OAI211_X1 U22895 ( .C1(n19812), .C2(n19867), .A(n19811), .B(n19810), .ZN(
        P2_U3147) );
  AOI22_X1 U22896 ( .A1(n19823), .A2(n19935), .B1(n19934), .B2(n19822), .ZN(
        n19814) );
  AOI22_X1 U22897 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19825), .B1(
        n19824), .B2(n19936), .ZN(n19813) );
  OAI211_X1 U22898 ( .C1(n19815), .C2(n19867), .A(n19814), .B(n19813), .ZN(
        P2_U3148) );
  AOI22_X1 U22899 ( .A1(n19823), .A2(n19942), .B1(n19941), .B2(n19822), .ZN(
        n19817) );
  AOI22_X1 U22900 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19825), .B1(
        n19824), .B2(n19944), .ZN(n19816) );
  OAI211_X1 U22901 ( .C1(n19818), .C2(n19867), .A(n19817), .B(n19816), .ZN(
        P2_U3149) );
  AOI22_X1 U22902 ( .A1(n19823), .A2(n19948), .B1(n19947), .B2(n19822), .ZN(
        n19820) );
  AOI22_X1 U22903 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19825), .B1(
        n19824), .B2(n19950), .ZN(n19819) );
  OAI211_X1 U22904 ( .C1(n19821), .C2(n19867), .A(n19820), .B(n19819), .ZN(
        P2_U3150) );
  AOI22_X1 U22905 ( .A1(n19823), .A2(n19955), .B1(n19953), .B2(n19822), .ZN(
        n19827) );
  AOI22_X1 U22906 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19825), .B1(
        n19824), .B2(n19957), .ZN(n19826) );
  OAI211_X1 U22907 ( .C1(n19828), .C2(n19867), .A(n19827), .B(n19826), .ZN(
        P2_U3151) );
  INV_X1 U22908 ( .A(n19829), .ZN(n19830) );
  NOR2_X1 U22909 ( .A1(n20092), .A2(n19837), .ZN(n19874) );
  NOR3_X1 U22910 ( .A1(n19830), .A2(n19874), .A3(n20113), .ZN(n19836) );
  INV_X1 U22911 ( .A(n19837), .ZN(n19831) );
  AOI21_X1 U22912 ( .B1(n19879), .B2(n19831), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19832) );
  NOR2_X1 U22913 ( .A1(n19836), .A2(n19832), .ZN(n19863) );
  AOI22_X1 U22914 ( .A1(n19863), .A2(n19833), .B1(n19876), .B2(n19874), .ZN(
        n19843) );
  NAND2_X1 U22915 ( .A1(n19835), .A2(n19834), .ZN(n19838) );
  AOI21_X1 U22916 ( .B1(n19838), .B2(n19837), .A(n19836), .ZN(n19839) );
  OAI211_X1 U22917 ( .C1(n19874), .C2(n19879), .A(n19883), .B(n19839), .ZN(
        n19864) );
  AOI22_X1 U22918 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19864), .B1(
        n19909), .B2(n19877), .ZN(n19842) );
  OAI211_X1 U22919 ( .C1(n19844), .C2(n19867), .A(n19843), .B(n19842), .ZN(
        P2_U3152) );
  AOI22_X1 U22920 ( .A1(n19863), .A2(n19916), .B1(n19915), .B2(n19874), .ZN(
        n19846) );
  AOI22_X1 U22921 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19864), .B1(
        n19909), .B2(n19918), .ZN(n19845) );
  OAI211_X1 U22922 ( .C1(n19847), .C2(n19867), .A(n19846), .B(n19845), .ZN(
        P2_U3153) );
  AOI22_X1 U22923 ( .A1(n19863), .A2(n19922), .B1(n19921), .B2(n19874), .ZN(
        n19849) );
  AOI22_X1 U22924 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19864), .B1(
        n19909), .B2(n19924), .ZN(n19848) );
  OAI211_X1 U22925 ( .C1(n19850), .C2(n19867), .A(n19849), .B(n19848), .ZN(
        P2_U3154) );
  AOI22_X1 U22926 ( .A1(n19863), .A2(n19929), .B1(n19928), .B2(n19874), .ZN(
        n19852) );
  AOI22_X1 U22927 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19864), .B1(
        n19909), .B2(n19930), .ZN(n19851) );
  OAI211_X1 U22928 ( .C1(n19853), .C2(n19867), .A(n19852), .B(n19851), .ZN(
        P2_U3155) );
  AOI22_X1 U22929 ( .A1(n19863), .A2(n19935), .B1(n19934), .B2(n19874), .ZN(
        n19855) );
  AOI22_X1 U22930 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19864), .B1(
        n19909), .B2(n19937), .ZN(n19854) );
  OAI211_X1 U22931 ( .C1(n19856), .C2(n19867), .A(n19855), .B(n19854), .ZN(
        P2_U3156) );
  AOI22_X1 U22932 ( .A1(n19863), .A2(n19942), .B1(n19941), .B2(n19874), .ZN(
        n19858) );
  AOI22_X1 U22933 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19864), .B1(
        n19909), .B2(n19943), .ZN(n19857) );
  OAI211_X1 U22934 ( .C1(n19859), .C2(n19867), .A(n19858), .B(n19857), .ZN(
        P2_U3157) );
  AOI22_X1 U22935 ( .A1(n19863), .A2(n19948), .B1(n19947), .B2(n19874), .ZN(
        n19861) );
  AOI22_X1 U22936 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19864), .B1(
        n19909), .B2(n19949), .ZN(n19860) );
  OAI211_X1 U22937 ( .C1(n19862), .C2(n19867), .A(n19861), .B(n19860), .ZN(
        P2_U3158) );
  AOI22_X1 U22938 ( .A1(n19863), .A2(n19955), .B1(n19953), .B2(n19874), .ZN(
        n19866) );
  AOI22_X1 U22939 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19864), .B1(
        n19909), .B2(n19959), .ZN(n19865) );
  OAI211_X1 U22940 ( .C1(n19868), .C2(n19867), .A(n19866), .B(n19865), .ZN(
        P2_U3159) );
  NAND3_X1 U22941 ( .A1(n19870), .A2(n19869), .A3(n20064), .ZN(n19872) );
  NAND2_X1 U22942 ( .A1(n19872), .A2(n19871), .ZN(n19878) );
  NOR2_X1 U22943 ( .A1(n19873), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19908) );
  OR2_X1 U22944 ( .A1(n19908), .A2(n19874), .ZN(n19884) );
  INV_X1 U22945 ( .A(n19908), .ZN(n19880) );
  AOI21_X1 U22946 ( .B1(n11171), .B2(n19880), .A(n20113), .ZN(n19875) );
  AOI22_X1 U22947 ( .A1(n19877), .A2(n19958), .B1(n19876), .B2(n19908), .ZN(
        n19888) );
  INV_X1 U22948 ( .A(n19878), .ZN(n19885) );
  OAI21_X1 U22949 ( .B1(n11120), .B2(n20113), .A(n19879), .ZN(n19881) );
  NAND2_X1 U22950 ( .A1(n19881), .A2(n19880), .ZN(n19882) );
  OAI211_X1 U22951 ( .C1(n19885), .C2(n19884), .A(n19883), .B(n19882), .ZN(
        n19910) );
  AOI22_X1 U22952 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19910), .B1(
        n19909), .B2(n19886), .ZN(n19887) );
  OAI211_X1 U22953 ( .C1(n19914), .C2(n19889), .A(n19888), .B(n19887), .ZN(
        P2_U3160) );
  INV_X1 U22954 ( .A(n19916), .ZN(n19892) );
  AOI22_X1 U22955 ( .A1(n19917), .A2(n19909), .B1(n19915), .B2(n19908), .ZN(
        n19891) );
  AOI22_X1 U22956 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19910), .B1(
        n19958), .B2(n19918), .ZN(n19890) );
  OAI211_X1 U22957 ( .C1(n19914), .C2(n19892), .A(n19891), .B(n19890), .ZN(
        P2_U3161) );
  INV_X1 U22958 ( .A(n19922), .ZN(n19895) );
  AOI22_X1 U22959 ( .A1(n19924), .A2(n19958), .B1(n19921), .B2(n19908), .ZN(
        n19894) );
  AOI22_X1 U22960 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19910), .B1(
        n19909), .B2(n19923), .ZN(n19893) );
  OAI211_X1 U22961 ( .C1(n19914), .C2(n19895), .A(n19894), .B(n19893), .ZN(
        P2_U3162) );
  INV_X1 U22962 ( .A(n19929), .ZN(n19898) );
  AOI22_X1 U22963 ( .A1(n19930), .A2(n19958), .B1(n19908), .B2(n19928), .ZN(
        n19897) );
  AOI22_X1 U22964 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19910), .B1(
        n19909), .B2(n19931), .ZN(n19896) );
  OAI211_X1 U22965 ( .C1(n19914), .C2(n19898), .A(n19897), .B(n19896), .ZN(
        P2_U3163) );
  AOI22_X1 U22966 ( .A1(n19936), .A2(n19909), .B1(n19934), .B2(n19908), .ZN(
        n19900) );
  AOI22_X1 U22967 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19910), .B1(
        n19958), .B2(n19937), .ZN(n19899) );
  OAI211_X1 U22968 ( .C1(n19914), .C2(n19901), .A(n19900), .B(n19899), .ZN(
        P2_U3164) );
  INV_X1 U22969 ( .A(n19942), .ZN(n19904) );
  AOI22_X1 U22970 ( .A1(n19944), .A2(n19909), .B1(n19908), .B2(n19941), .ZN(
        n19903) );
  AOI22_X1 U22971 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19910), .B1(
        n19958), .B2(n19943), .ZN(n19902) );
  OAI211_X1 U22972 ( .C1(n19914), .C2(n19904), .A(n19903), .B(n19902), .ZN(
        P2_U3165) );
  INV_X1 U22973 ( .A(n19948), .ZN(n19907) );
  AOI22_X1 U22974 ( .A1(n19949), .A2(n19958), .B1(n19908), .B2(n19947), .ZN(
        n19906) );
  AOI22_X1 U22975 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19910), .B1(
        n19909), .B2(n19950), .ZN(n19905) );
  OAI211_X1 U22976 ( .C1(n19914), .C2(n19907), .A(n19906), .B(n19905), .ZN(
        P2_U3166) );
  INV_X1 U22977 ( .A(n19955), .ZN(n19913) );
  AOI22_X1 U22978 ( .A1(n19959), .A2(n19958), .B1(n19953), .B2(n19908), .ZN(
        n19912) );
  AOI22_X1 U22979 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19910), .B1(
        n19909), .B2(n19957), .ZN(n19911) );
  OAI211_X1 U22980 ( .C1(n19914), .C2(n19913), .A(n19912), .B(n19911), .ZN(
        P2_U3167) );
  AOI22_X1 U22981 ( .A1(n19956), .A2(n19916), .B1(n19954), .B2(n19915), .ZN(
        n19920) );
  AOI22_X1 U22982 ( .A1(n19960), .A2(n19918), .B1(n19958), .B2(n19917), .ZN(
        n19919) );
  OAI211_X1 U22983 ( .C1(n19964), .C2(n11095), .A(n19920), .B(n19919), .ZN(
        P2_U3169) );
  INV_X1 U22984 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n19927) );
  AOI22_X1 U22985 ( .A1(n19956), .A2(n19922), .B1(n19954), .B2(n19921), .ZN(
        n19926) );
  AOI22_X1 U22986 ( .A1(n19960), .A2(n19924), .B1(n19958), .B2(n19923), .ZN(
        n19925) );
  OAI211_X1 U22987 ( .C1(n19964), .C2(n19927), .A(n19926), .B(n19925), .ZN(
        P2_U3170) );
  AOI22_X1 U22988 ( .A1(n19956), .A2(n19929), .B1(n19954), .B2(n19928), .ZN(
        n19933) );
  AOI22_X1 U22989 ( .A1(n19958), .A2(n19931), .B1(n19960), .B2(n19930), .ZN(
        n19932) );
  OAI211_X1 U22990 ( .C1(n19964), .C2(n11144), .A(n19933), .B(n19932), .ZN(
        P2_U3171) );
  INV_X1 U22991 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n19940) );
  AOI22_X1 U22992 ( .A1(n19935), .A2(n19956), .B1(n19954), .B2(n19934), .ZN(
        n19939) );
  AOI22_X1 U22993 ( .A1(n19960), .A2(n19937), .B1(n19958), .B2(n19936), .ZN(
        n19938) );
  OAI211_X1 U22994 ( .C1(n19964), .C2(n19940), .A(n19939), .B(n19938), .ZN(
        P2_U3172) );
  AOI22_X1 U22995 ( .A1(n19956), .A2(n19942), .B1(n19954), .B2(n19941), .ZN(
        n19946) );
  AOI22_X1 U22996 ( .A1(n19958), .A2(n19944), .B1(n19960), .B2(n19943), .ZN(
        n19945) );
  OAI211_X1 U22997 ( .C1(n19964), .C2(n11166), .A(n19946), .B(n19945), .ZN(
        P2_U3173) );
  AOI22_X1 U22998 ( .A1(n19956), .A2(n19948), .B1(n19954), .B2(n19947), .ZN(
        n19952) );
  AOI22_X1 U22999 ( .A1(n19958), .A2(n19950), .B1(n19960), .B2(n19949), .ZN(
        n19951) );
  OAI211_X1 U23000 ( .C1(n19964), .C2(n11245), .A(n19952), .B(n19951), .ZN(
        P2_U3174) );
  INV_X1 U23001 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n19963) );
  AOI22_X1 U23002 ( .A1(n19956), .A2(n19955), .B1(n19954), .B2(n19953), .ZN(
        n19962) );
  AOI22_X1 U23003 ( .A1(n19960), .A2(n19959), .B1(n19958), .B2(n19957), .ZN(
        n19961) );
  OAI211_X1 U23004 ( .C1(n19964), .C2(n19963), .A(n19962), .B(n19961), .ZN(
        P2_U3175) );
  NOR2_X1 U23005 ( .A1(n19350), .A2(n19965), .ZN(n19971) );
  OAI21_X1 U23006 ( .B1(n20061), .B2(n19966), .A(n9755), .ZN(n19970) );
  NAND2_X1 U23007 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n20114), .ZN(n19967) );
  AOI21_X1 U23008 ( .B1(n19968), .B2(n19971), .A(n19967), .ZN(n19969) );
  AOI21_X1 U23009 ( .B1(n19971), .B2(n19970), .A(n19969), .ZN(n19973) );
  NAND2_X1 U23010 ( .A1(n19973), .A2(n19972), .ZN(P2_U3177) );
  AND2_X1 U23011 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19974), .ZN(
        P2_U3179) );
  AND2_X1 U23012 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19974), .ZN(
        P2_U3180) );
  AND2_X1 U23013 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19974), .ZN(
        P2_U3181) );
  AND2_X1 U23014 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19974), .ZN(
        P2_U3182) );
  AND2_X1 U23015 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19974), .ZN(
        P2_U3183) );
  AND2_X1 U23016 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19974), .ZN(
        P2_U3184) );
  AND2_X1 U23017 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19974), .ZN(
        P2_U3185) );
  AND2_X1 U23018 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19974), .ZN(
        P2_U3186) );
  AND2_X1 U23019 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19974), .ZN(
        P2_U3187) );
  AND2_X1 U23020 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19974), .ZN(
        P2_U3188) );
  AND2_X1 U23021 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19974), .ZN(
        P2_U3189) );
  AND2_X1 U23022 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19974), .ZN(
        P2_U3190) );
  AND2_X1 U23023 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19974), .ZN(
        P2_U3191) );
  AND2_X1 U23024 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19974), .ZN(
        P2_U3192) );
  AND2_X1 U23025 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19974), .ZN(
        P2_U3193) );
  AND2_X1 U23026 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19974), .ZN(
        P2_U3194) );
  AND2_X1 U23027 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19974), .ZN(
        P2_U3195) );
  AND2_X1 U23028 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19974), .ZN(
        P2_U3196) );
  AND2_X1 U23029 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19974), .ZN(
        P2_U3197) );
  AND2_X1 U23030 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19974), .ZN(
        P2_U3198) );
  AND2_X1 U23031 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19974), .ZN(
        P2_U3199) );
  AND2_X1 U23032 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19974), .ZN(
        P2_U3200) );
  AND2_X1 U23033 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19974), .ZN(P2_U3201) );
  AND2_X1 U23034 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19974), .ZN(P2_U3202) );
  AND2_X1 U23035 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19974), .ZN(P2_U3203) );
  AND2_X1 U23036 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19974), .ZN(P2_U3204) );
  AND2_X1 U23037 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19974), .ZN(P2_U3205) );
  AND2_X1 U23038 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19974), .ZN(P2_U3206) );
  AND2_X1 U23039 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19974), .ZN(P2_U3207) );
  AND2_X1 U23040 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19974), .ZN(P2_U3208) );
  NAND2_X1 U23041 ( .A1(n20114), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19987) );
  NAND3_X1 U23042 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19987), .ZN(n19977) );
  AOI211_X1 U23043 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20743), .A(
        n19975), .B(n20129), .ZN(n19976) );
  NOR2_X1 U23044 ( .A1(n20737), .A2(n19981), .ZN(n19992) );
  AOI211_X1 U23045 ( .C1(n20958), .C2(n19977), .A(n19976), .B(n19992), .ZN(
        n19978) );
  INV_X1 U23046 ( .A(n19978), .ZN(P2_U3209) );
  INV_X1 U23047 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19979) );
  AOI21_X1 U23048 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20743), .A(n20958), 
        .ZN(n19985) );
  NOR2_X1 U23049 ( .A1(n19979), .A2(n19985), .ZN(n19982) );
  AOI21_X1 U23050 ( .B1(n19982), .B2(n19981), .A(n19980), .ZN(n19983) );
  OAI211_X1 U23051 ( .C1(n20743), .C2(n19984), .A(n19983), .B(n19987), .ZN(
        P2_U3210) );
  AOI21_X1 U23052 ( .B1(n19986), .B2(n20114), .A(n19985), .ZN(n19991) );
  OAI22_X1 U23053 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19988), .B1(NA), 
        .B2(n19987), .ZN(n19989) );
  OAI211_X1 U23054 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19989), .ZN(n19990) );
  OAI21_X1 U23055 ( .B1(n19992), .B2(n19991), .A(n19990), .ZN(P2_U3211) );
  NAND2_X1 U23056 ( .A1(n20129), .A2(n20958), .ZN(n20049) );
  CLKBUF_X1 U23057 ( .A(n20049), .Z(n20045) );
  OAI222_X1 U23058 ( .A1(n20045), .A2(n19996), .B1(n19994), .B2(n20129), .C1(
        n19993), .C2(n20046), .ZN(P2_U3212) );
  OAI222_X1 U23059 ( .A1(n20046), .A2(n19996), .B1(n19995), .B2(n20129), .C1(
        n19998), .C2(n20045), .ZN(P2_U3213) );
  OAI222_X1 U23060 ( .A1(n20046), .A2(n19998), .B1(n19997), .B2(n20129), .C1(
        n19999), .C2(n20045), .ZN(P2_U3214) );
  INV_X1 U23061 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n20001) );
  OAI222_X1 U23062 ( .A1(n20049), .A2(n20001), .B1(n20000), .B2(n20129), .C1(
        n19999), .C2(n20046), .ZN(P2_U3215) );
  OAI222_X1 U23063 ( .A1(n20049), .A2(n20003), .B1(n20002), .B2(n20129), .C1(
        n20001), .C2(n20046), .ZN(P2_U3216) );
  INV_X1 U23064 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20005) );
  OAI222_X1 U23065 ( .A1(n20049), .A2(n20005), .B1(n20004), .B2(n20129), .C1(
        n20003), .C2(n20046), .ZN(P2_U3217) );
  INV_X1 U23066 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20007) );
  OAI222_X1 U23067 ( .A1(n20049), .A2(n20007), .B1(n20006), .B2(n20129), .C1(
        n20005), .C2(n20046), .ZN(P2_U3218) );
  INV_X1 U23068 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20009) );
  OAI222_X1 U23069 ( .A1(n20049), .A2(n20009), .B1(n20008), .B2(n20129), .C1(
        n20007), .C2(n20046), .ZN(P2_U3219) );
  OAI222_X1 U23070 ( .A1(n20045), .A2(n20011), .B1(n20010), .B2(n20129), .C1(
        n20009), .C2(n20046), .ZN(P2_U3220) );
  OAI222_X1 U23071 ( .A1(n20045), .A2(n11018), .B1(n20012), .B2(n20129), .C1(
        n20011), .C2(n20046), .ZN(P2_U3221) );
  OAI222_X1 U23072 ( .A1(n20045), .A2(n20014), .B1(n20013), .B2(n20129), .C1(
        n11018), .C2(n20046), .ZN(P2_U3222) );
  OAI222_X1 U23073 ( .A1(n20045), .A2(n11025), .B1(n20015), .B2(n20129), .C1(
        n20014), .C2(n20046), .ZN(P2_U3223) );
  OAI222_X1 U23074 ( .A1(n20045), .A2(n20017), .B1(n20016), .B2(n20129), .C1(
        n11025), .C2(n20046), .ZN(P2_U3224) );
  OAI222_X1 U23075 ( .A1(n20045), .A2(n11032), .B1(n20018), .B2(n20129), .C1(
        n20017), .C2(n20046), .ZN(P2_U3225) );
  INV_X1 U23076 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20020) );
  OAI222_X1 U23077 ( .A1(n20049), .A2(n20020), .B1(n20019), .B2(n20129), .C1(
        n11032), .C2(n20046), .ZN(P2_U3226) );
  OAI222_X1 U23078 ( .A1(n20049), .A2(n19038), .B1(n20888), .B2(n20129), .C1(
        n20020), .C2(n20046), .ZN(P2_U3227) );
  INV_X1 U23079 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20022) );
  OAI222_X1 U23080 ( .A1(n20049), .A2(n20022), .B1(n20021), .B2(n20129), .C1(
        n19038), .C2(n20046), .ZN(P2_U3228) );
  OAI222_X1 U23081 ( .A1(n20049), .A2(n19014), .B1(n20023), .B2(n20129), .C1(
        n20022), .C2(n20046), .ZN(P2_U3229) );
  OAI222_X1 U23082 ( .A1(n20049), .A2(n20025), .B1(n20024), .B2(n20129), .C1(
        n19014), .C2(n20046), .ZN(P2_U3230) );
  OAI222_X1 U23083 ( .A1(n20049), .A2(n20027), .B1(n20026), .B2(n20129), .C1(
        n20025), .C2(n20046), .ZN(P2_U3231) );
  OAI222_X1 U23084 ( .A1(n20045), .A2(n20029), .B1(n20028), .B2(n20129), .C1(
        n20027), .C2(n20046), .ZN(P2_U3232) );
  INV_X1 U23085 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20031) );
  OAI222_X1 U23086 ( .A1(n20045), .A2(n20031), .B1(n20030), .B2(n20129), .C1(
        n20029), .C2(n20046), .ZN(P2_U3233) );
  OAI222_X1 U23087 ( .A1(n20045), .A2(n20033), .B1(n20032), .B2(n20129), .C1(
        n20031), .C2(n20046), .ZN(P2_U3234) );
  INV_X1 U23088 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20035) );
  OAI222_X1 U23089 ( .A1(n20045), .A2(n20035), .B1(n20034), .B2(n20129), .C1(
        n20033), .C2(n20046), .ZN(P2_U3235) );
  INV_X1 U23090 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20037) );
  OAI222_X1 U23091 ( .A1(n20045), .A2(n20037), .B1(n20036), .B2(n20129), .C1(
        n20035), .C2(n20046), .ZN(P2_U3236) );
  INV_X1 U23092 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20040) );
  OAI222_X1 U23093 ( .A1(n20045), .A2(n20040), .B1(n20038), .B2(n20129), .C1(
        n20037), .C2(n20046), .ZN(P2_U3237) );
  OAI222_X1 U23094 ( .A1(n20046), .A2(n20040), .B1(n20039), .B2(n20129), .C1(
        n20041), .C2(n20045), .ZN(P2_U3238) );
  OAI222_X1 U23095 ( .A1(n20045), .A2(n20043), .B1(n20042), .B2(n20129), .C1(
        n20041), .C2(n20046), .ZN(P2_U3239) );
  OAI222_X1 U23096 ( .A1(n20045), .A2(n15458), .B1(n20044), .B2(n20129), .C1(
        n20043), .C2(n20046), .ZN(P2_U3240) );
  OAI222_X1 U23097 ( .A1(n20049), .A2(n20048), .B1(n20047), .B2(n20129), .C1(
        n15458), .C2(n20046), .ZN(P2_U3241) );
  INV_X1 U23098 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20050) );
  AOI22_X1 U23099 ( .A1(n20129), .A2(n20051), .B1(n20050), .B2(n20126), .ZN(
        P2_U3585) );
  MUX2_X1 U23100 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20129), .Z(P2_U3586) );
  INV_X1 U23101 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20052) );
  AOI22_X1 U23102 ( .A1(n20129), .A2(n20053), .B1(n20052), .B2(n20126), .ZN(
        P2_U3587) );
  INV_X1 U23103 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20054) );
  AOI22_X1 U23104 ( .A1(n20129), .A2(n20055), .B1(n20054), .B2(n20126), .ZN(
        P2_U3588) );
  OAI21_X1 U23105 ( .B1(n20059), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20057), 
        .ZN(n20056) );
  INV_X1 U23106 ( .A(n20056), .ZN(P2_U3591) );
  OAI21_X1 U23107 ( .B1(n20059), .B2(n20058), .A(n20057), .ZN(P2_U3592) );
  AND2_X1 U23108 ( .A1(n20064), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20081) );
  NAND2_X1 U23109 ( .A1(n20060), .A2(n20081), .ZN(n20070) );
  NAND3_X1 U23110 ( .A1(n20079), .A2(n20061), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20062) );
  NAND2_X1 U23111 ( .A1(n20062), .A2(n20077), .ZN(n20071) );
  NAND2_X1 U23112 ( .A1(n20070), .A2(n20071), .ZN(n20067) );
  AOI222_X1 U23113 ( .A1(n20067), .A2(n20066), .B1(n20065), .B2(
        P2_STATE2_REG_3__SCAN_IN), .C1(n20064), .C2(n20063), .ZN(n20068) );
  AOI22_X1 U23114 ( .A1(n20093), .A2(n20069), .B1(n20068), .B2(n20090), .ZN(
        P2_U3602) );
  OAI21_X1 U23115 ( .B1(n20072), .B2(n20071), .A(n20070), .ZN(n20073) );
  AOI21_X1 U23116 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20074), .A(n20073), 
        .ZN(n20075) );
  AOI22_X1 U23117 ( .A1(n20093), .A2(n20076), .B1(n20075), .B2(n20090), .ZN(
        P2_U3603) );
  INV_X1 U23118 ( .A(n20077), .ZN(n20122) );
  NOR2_X1 U23119 ( .A1(n20122), .A2(n20078), .ZN(n20080) );
  MUX2_X1 U23120 ( .A(n20081), .B(n20080), .S(n20079), .Z(n20082) );
  AOI21_X1 U23121 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20083), .A(n20082), 
        .ZN(n20084) );
  AOI22_X1 U23122 ( .A1(n20093), .A2(n20085), .B1(n20084), .B2(n20090), .ZN(
        P2_U3604) );
  OAI22_X1 U23123 ( .A1(n20086), .A2(n20122), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19879), .ZN(n20087) );
  AOI21_X1 U23124 ( .B1(n20089), .B2(n20088), .A(n20087), .ZN(n20091) );
  AOI22_X1 U23125 ( .A1(n20093), .A2(n20092), .B1(n20091), .B2(n20090), .ZN(
        P2_U3605) );
  INV_X1 U23126 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20094) );
  AOI22_X1 U23127 ( .A1(n20129), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20094), 
        .B2(n20126), .ZN(P2_U3608) );
  INV_X1 U23128 ( .A(n20095), .ZN(n20096) );
  AOI21_X1 U23129 ( .B1(n20098), .B2(n20097), .A(n20096), .ZN(n20100) );
  AOI211_X1 U23130 ( .C1(n20102), .C2(n20101), .A(n20100), .B(n20099), .ZN(
        n20103) );
  INV_X1 U23131 ( .A(n20103), .ZN(n20105) );
  MUX2_X1 U23132 ( .A(P2_MORE_REG_SCAN_IN), .B(n20105), .S(n20104), .Z(
        P2_U3609) );
  OAI21_X1 U23133 ( .B1(n20107), .B2(n20108), .A(n20106), .ZN(n20112) );
  NAND3_X1 U23134 ( .A1(n9748), .A2(n20109), .A3(n20108), .ZN(n20111) );
  AND2_X1 U23135 ( .A1(n20112), .A2(n20111), .ZN(n20117) );
  NOR2_X1 U23136 ( .A1(n20114), .A2(n20113), .ZN(n20116) );
  OAI22_X1 U23137 ( .A1(n20117), .A2(n20119), .B1(n20116), .B2(n20115), .ZN(
        n20125) );
  NAND4_X1 U23138 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .A3(n20119), .A4(n20118), .ZN(n20121) );
  OAI211_X1 U23139 ( .C1(n20123), .C2(n20122), .A(n20121), .B(n20120), .ZN(
        n20124) );
  MUX2_X1 U23140 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n20125), .S(n20124), 
        .Z(P2_U3610) );
  INV_X1 U23141 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n20127) );
  AOI22_X1 U23142 ( .A1(n20129), .A2(n20128), .B1(n20127), .B2(n20126), .ZN(
        P2_U3611) );
  AOI21_X1 U23143 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n11789), .A(n20738), 
        .ZN(n20741) );
  INV_X1 U23144 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20131) );
  OR2_X1 U23145 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20130), .ZN(n20836) );
  INV_X2 U23146 ( .A(n20836), .ZN(n20850) );
  AOI21_X1 U23147 ( .B1(n20741), .B2(n20131), .A(n20850), .ZN(P1_U2802) );
  INV_X1 U23148 ( .A(n20132), .ZN(n20134) );
  OAI21_X1 U23149 ( .B1(n20134), .B2(n20133), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20135) );
  OAI21_X1 U23150 ( .B1(n20136), .B2(n9918), .A(n20135), .ZN(P1_U2803) );
  NOR2_X1 U23151 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20138) );
  OAI21_X1 U23152 ( .B1(n20138), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20836), .ZN(
        n20137) );
  OAI21_X1 U23153 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20836), .A(n20137), 
        .ZN(P1_U2804) );
  NOR2_X1 U23154 ( .A1(n20850), .A2(n20741), .ZN(n20731) );
  OAI21_X1 U23155 ( .B1(BS16), .B2(n20138), .A(n20731), .ZN(n20798) );
  OAI21_X1 U23156 ( .B1(n20731), .B2(n20840), .A(n20798), .ZN(P1_U2805) );
  INV_X1 U23157 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20140) );
  OAI21_X1 U23158 ( .B1(n20141), .B2(n20140), .A(n20139), .ZN(P1_U2806) );
  NOR4_X1 U23159 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20145) );
  NOR4_X1 U23160 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20144) );
  NOR4_X1 U23161 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20143) );
  NOR4_X1 U23162 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20142) );
  NAND4_X1 U23163 ( .A1(n20145), .A2(n20144), .A3(n20143), .A4(n20142), .ZN(
        n20151) );
  NOR4_X1 U23164 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_2__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n20149) );
  AOI211_X1 U23165 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_5__SCAN_IN), .B(
        P1_DATAWIDTH_REG_21__SCAN_IN), .ZN(n20148) );
  NOR4_X1 U23166 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20147) );
  NOR4_X1 U23167 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20146) );
  NAND4_X1 U23168 ( .A1(n20149), .A2(n20148), .A3(n20147), .A4(n20146), .ZN(
        n20150) );
  NOR2_X1 U23169 ( .A1(n20151), .A2(n20150), .ZN(n20835) );
  INV_X1 U23170 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20796) );
  NOR3_X1 U23171 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20153) );
  OAI21_X1 U23172 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20153), .A(n20835), .ZN(
        n20152) );
  OAI21_X1 U23173 ( .B1(n20835), .B2(n20796), .A(n20152), .ZN(P1_U2807) );
  INV_X1 U23174 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20793) );
  NOR2_X1 U23175 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20829) );
  OAI21_X1 U23176 ( .B1(n20153), .B2(n20829), .A(n20835), .ZN(n20154) );
  OAI21_X1 U23177 ( .B1(n20835), .B2(n20793), .A(n20154), .ZN(P1_U2808) );
  AOI22_X1 U23178 ( .A1(n20206), .A2(P1_EBX_REG_9__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n20193), .ZN(n20155) );
  OAI211_X1 U23179 ( .C1(n20156), .C2(n20191), .A(n20155), .B(n20207), .ZN(
        n20157) );
  AOI221_X1 U23180 ( .B1(n20159), .B2(P1_REIP_REG_9__SCAN_IN), .C1(n20158), 
        .C2(n14294), .A(n20157), .ZN(n20165) );
  INV_X1 U23181 ( .A(n20160), .ZN(n20163) );
  AOI22_X1 U23182 ( .A1(n20163), .A2(n20185), .B1(n20162), .B2(n20161), .ZN(
        n20164) );
  NAND2_X1 U23183 ( .A1(n20165), .A2(n20164), .ZN(P1_U2831) );
  NAND2_X1 U23184 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20166) );
  OAI21_X1 U23185 ( .B1(n20166), .B2(n20188), .A(n20189), .ZN(n20182) );
  OAI22_X1 U23186 ( .A1(n20191), .A2(n20167), .B1(n20756), .B2(n20182), .ZN(
        n20173) );
  NAND4_X1 U23187 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n20179), .A4(n20756), .ZN(n20168) );
  NAND2_X1 U23188 ( .A1(n20207), .A2(n20168), .ZN(n20169) );
  AOI21_X1 U23189 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n20193), .A(
        n20169), .ZN(n20170) );
  OAI21_X1 U23190 ( .B1(n20194), .B2(n20171), .A(n20170), .ZN(n20172) );
  NOR2_X1 U23191 ( .A1(n20173), .A2(n20172), .ZN(n20176) );
  NAND2_X1 U23192 ( .A1(n20174), .A2(n20185), .ZN(n20175) );
  AND2_X1 U23193 ( .A1(n20176), .A2(n20175), .ZN(n20177) );
  OAI21_X1 U23194 ( .B1(n20178), .B2(n20216), .A(n20177), .ZN(P1_U2833) );
  INV_X1 U23195 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20226) );
  NAND2_X1 U23196 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n20179), .ZN(n20180) );
  OAI22_X1 U23197 ( .A1(n20194), .A2(n20226), .B1(P1_REIP_REG_6__SCAN_IN), 
        .B2(n20180), .ZN(n20184) );
  INV_X1 U23198 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20754) );
  AOI22_X1 U23199 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20193), .B1(
        n20205), .B2(n20221), .ZN(n20181) );
  OAI211_X1 U23200 ( .C1(n20754), .C2(n20182), .A(n20181), .B(n20207), .ZN(
        n20183) );
  AOI211_X1 U23201 ( .C1(n20224), .C2(n20185), .A(n20184), .B(n20183), .ZN(
        n20186) );
  OAI21_X1 U23202 ( .B1(n20187), .B2(n20216), .A(n20186), .ZN(P1_U2834) );
  INV_X1 U23203 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20752) );
  NAND2_X1 U23204 ( .A1(n20189), .A2(n20188), .ZN(n20220) );
  OAI22_X1 U23205 ( .A1(n20191), .A2(n20190), .B1(n20752), .B2(n20220), .ZN(
        n20192) );
  AOI211_X1 U23206 ( .C1(n20193), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n20299), .B(n20192), .ZN(n20200) );
  OAI22_X1 U23207 ( .A1(n20196), .A2(P1_REIP_REG_5__SCAN_IN), .B1(n20195), 
        .B2(n20194), .ZN(n20197) );
  AOI21_X1 U23208 ( .B1(n20218), .B2(n20198), .A(n20197), .ZN(n20199) );
  OAI211_X1 U23209 ( .C1(n20201), .C2(n20216), .A(n20200), .B(n20199), .ZN(
        P1_U2835) );
  NOR3_X1 U23210 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20203), .A3(n20202), .ZN(
        n20204) );
  AOI21_X1 U23211 ( .B1(n20300), .B2(n20205), .A(n20204), .ZN(n20215) );
  INV_X1 U23212 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20209) );
  NAND2_X1 U23213 ( .A1(n20206), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n20208) );
  OAI211_X1 U23214 ( .C1(n20210), .C2(n20209), .A(n20208), .B(n20207), .ZN(
        n20211) );
  AOI21_X1 U23215 ( .B1(n20213), .B2(n20212), .A(n20211), .ZN(n20214) );
  OAI211_X1 U23216 ( .C1(n20216), .C2(n20297), .A(n20215), .B(n20214), .ZN(
        n20217) );
  AOI21_X1 U23217 ( .B1(n20292), .B2(n20218), .A(n20217), .ZN(n20219) );
  OAI21_X1 U23218 ( .B1(n20750), .B2(n20220), .A(n20219), .ZN(P1_U2836) );
  AOI22_X1 U23219 ( .A1(n20224), .A2(n20223), .B1(n20222), .B2(n20221), .ZN(
        n20225) );
  OAI21_X1 U23220 ( .B1(n20227), .B2(n20226), .A(n20225), .ZN(P1_U2866) );
  AOI22_X1 U23221 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20228), .B1(n20248), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20229) );
  OAI21_X1 U23222 ( .B1(n20231), .B2(n20230), .A(n20229), .ZN(P1_U2921) );
  AOI22_X1 U23223 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20232) );
  OAI21_X1 U23224 ( .B1(n14291), .B2(n20250), .A(n20232), .ZN(P1_U2922) );
  AOI22_X1 U23225 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20233) );
  OAI21_X1 U23226 ( .B1(n14317), .B2(n20250), .A(n20233), .ZN(P1_U2923) );
  AOI22_X1 U23227 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20234) );
  OAI21_X1 U23228 ( .B1(n14330), .B2(n20250), .A(n20234), .ZN(P1_U2924) );
  AOI22_X1 U23229 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20847), .B1(n20239), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20235) );
  OAI21_X1 U23230 ( .B1(n14301), .B2(n20250), .A(n20235), .ZN(P1_U2925) );
  AOI22_X1 U23231 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20847), .B1(n20239), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20236) );
  OAI21_X1 U23232 ( .B1(n14227), .B2(n20250), .A(n20236), .ZN(P1_U2926) );
  AOI22_X1 U23233 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20237) );
  OAI21_X1 U23234 ( .B1(n14237), .B2(n20250), .A(n20237), .ZN(P1_U2927) );
  AOI22_X1 U23235 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20847), .B1(n20239), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20238) );
  OAI21_X1 U23236 ( .B1(n14192), .B2(n20250), .A(n20238), .ZN(P1_U2928) );
  AOI22_X1 U23237 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20847), .B1(n20239), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20240) );
  OAI21_X1 U23238 ( .B1(n12238), .B2(n20250), .A(n20240), .ZN(P1_U2929) );
  AOI22_X1 U23239 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20241) );
  OAI21_X1 U23240 ( .B1(n12198), .B2(n20250), .A(n20241), .ZN(P1_U2930) );
  AOI22_X1 U23241 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20242) );
  OAI21_X1 U23242 ( .B1(n12188), .B2(n20250), .A(n20242), .ZN(P1_U2931) );
  AOI22_X1 U23243 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20243) );
  OAI21_X1 U23244 ( .B1(n20244), .B2(n20250), .A(n20243), .ZN(P1_U2932) );
  AOI22_X1 U23245 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20245) );
  OAI21_X1 U23246 ( .B1(n12172), .B2(n20250), .A(n20245), .ZN(P1_U2933) );
  AOI22_X1 U23247 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20246) );
  OAI21_X1 U23248 ( .B1(n12143), .B2(n20250), .A(n20246), .ZN(P1_U2934) );
  AOI22_X1 U23249 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20247) );
  OAI21_X1 U23250 ( .B1(n12153), .B2(n20250), .A(n20247), .ZN(P1_U2935) );
  AOI22_X1 U23251 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20847), .B1(n20248), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20249) );
  OAI21_X1 U23252 ( .B1(n21053), .B2(n20250), .A(n20249), .ZN(P1_U2936) );
  AOI22_X1 U23253 ( .A1(n20281), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20257), .ZN(n20253) );
  INV_X1 U23254 ( .A(n20251), .ZN(n20252) );
  NAND2_X1 U23255 ( .A1(n20269), .A2(n20252), .ZN(n20271) );
  NAND2_X1 U23256 ( .A1(n20253), .A2(n20271), .ZN(P1_U2945) );
  AOI22_X1 U23257 ( .A1(n20281), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20257), .ZN(n20256) );
  INV_X1 U23258 ( .A(n20254), .ZN(n20255) );
  NAND2_X1 U23259 ( .A1(n20269), .A2(n20255), .ZN(n20275) );
  NAND2_X1 U23260 ( .A1(n20256), .A2(n20275), .ZN(P1_U2947) );
  AOI22_X1 U23261 ( .A1(n20281), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20257), .ZN(n20260) );
  INV_X1 U23262 ( .A(n20258), .ZN(n20259) );
  NAND2_X1 U23263 ( .A1(n20269), .A2(n20259), .ZN(n20277) );
  NAND2_X1 U23264 ( .A1(n20260), .A2(n20277), .ZN(P1_U2948) );
  AOI22_X1 U23265 ( .A1(n20281), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20284), .ZN(n20263) );
  INV_X1 U23266 ( .A(n20261), .ZN(n20262) );
  NAND2_X1 U23267 ( .A1(n20269), .A2(n20262), .ZN(n20279) );
  NAND2_X1 U23268 ( .A1(n20263), .A2(n20279), .ZN(P1_U2949) );
  AOI22_X1 U23269 ( .A1(n20281), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20284), .ZN(n20266) );
  INV_X1 U23270 ( .A(n20264), .ZN(n20265) );
  NAND2_X1 U23271 ( .A1(n20269), .A2(n20265), .ZN(n20282) );
  NAND2_X1 U23272 ( .A1(n20266), .A2(n20282), .ZN(P1_U2950) );
  AOI22_X1 U23273 ( .A1(n20281), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20284), .ZN(n20270) );
  INV_X1 U23274 ( .A(n20267), .ZN(n20268) );
  NAND2_X1 U23275 ( .A1(n20269), .A2(n20268), .ZN(n20285) );
  NAND2_X1 U23276 ( .A1(n20270), .A2(n20285), .ZN(P1_U2951) );
  AOI22_X1 U23277 ( .A1(n20281), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20257), .ZN(n20272) );
  NAND2_X1 U23278 ( .A1(n20272), .A2(n20271), .ZN(P1_U2960) );
  AOI22_X1 U23279 ( .A1(n20281), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20284), .ZN(n20274) );
  NAND2_X1 U23280 ( .A1(n20274), .A2(n20273), .ZN(P1_U2961) );
  AOI22_X1 U23281 ( .A1(n20281), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20257), .ZN(n20276) );
  NAND2_X1 U23282 ( .A1(n20276), .A2(n20275), .ZN(P1_U2962) );
  AOI22_X1 U23283 ( .A1(n20281), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20284), .ZN(n20278) );
  NAND2_X1 U23284 ( .A1(n20278), .A2(n20277), .ZN(P1_U2963) );
  AOI22_X1 U23285 ( .A1(n20281), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20257), .ZN(n20280) );
  NAND2_X1 U23286 ( .A1(n20280), .A2(n20279), .ZN(P1_U2964) );
  AOI22_X1 U23287 ( .A1(n20281), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20284), .ZN(n20283) );
  NAND2_X1 U23288 ( .A1(n20283), .A2(n20282), .ZN(P1_U2965) );
  AOI22_X1 U23289 ( .A1(n20281), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20284), .ZN(n20286) );
  NAND2_X1 U23290 ( .A1(n20286), .A2(n20285), .ZN(P1_U2966) );
  AOI22_X1 U23291 ( .A1(n20287), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20299), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20296) );
  OAI21_X1 U23292 ( .B1(n20288), .B2(n20290), .A(n20289), .ZN(n20291) );
  INV_X1 U23293 ( .A(n20291), .ZN(n20302) );
  AOI22_X1 U23294 ( .A1(n20302), .A2(n20294), .B1(n20293), .B2(n20292), .ZN(
        n20295) );
  OAI211_X1 U23295 ( .C1(n20298), .C2(n20297), .A(n20296), .B(n20295), .ZN(
        P1_U2995) );
  AOI22_X1 U23296 ( .A1(n20312), .A2(n20300), .B1(n20299), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n20307) );
  AOI22_X1 U23297 ( .A1(n20302), .A2(n20318), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n20301), .ZN(n20306) );
  OAI211_X1 U23298 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20304), .B(n20303), .ZN(n20305) );
  NAND3_X1 U23299 ( .A1(n20307), .A2(n20306), .A3(n20305), .ZN(P1_U3027) );
  INV_X1 U23300 ( .A(n20308), .ZN(n20311) );
  INV_X1 U23301 ( .A(n20309), .ZN(n20310) );
  AOI21_X1 U23302 ( .B1(n20312), .B2(n20311), .A(n20310), .ZN(n20325) );
  NAND2_X1 U23303 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20315) );
  OAI21_X1 U23304 ( .B1(n20315), .B2(n20314), .A(n20313), .ZN(n20319) );
  INV_X1 U23305 ( .A(n20316), .ZN(n20317) );
  AOI22_X1 U23306 ( .A1(n20319), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20318), .B2(n20317), .ZN(n20324) );
  NAND3_X1 U23307 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20321), .A3(
        n20320), .ZN(n20322) );
  NAND4_X1 U23308 ( .A1(n20325), .A2(n20324), .A3(n20323), .A4(n20322), .ZN(
        P1_U3029) );
  NOR2_X1 U23309 ( .A1(n20326), .A2(n20823), .ZN(P1_U3032) );
  INV_X1 U23310 ( .A(n20493), .ZN(n20327) );
  INV_X1 U23311 ( .A(n20679), .ZN(n20643) );
  NOR2_X1 U23312 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20328), .ZN(
        n20351) );
  AOI22_X1 U23313 ( .A1(n20721), .A2(n20643), .B1(n20351), .B2(n20669), .ZN(
        n20338) );
  INV_X1 U23314 ( .A(n20721), .ZN(n20329) );
  NAND2_X1 U23315 ( .A1(n20329), .A2(n20372), .ZN(n20330) );
  AOI21_X1 U23316 ( .B1(n20330), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20667), 
        .ZN(n20334) );
  NAND2_X1 U23317 ( .A1(n9847), .A2(n20518), .ZN(n20335) );
  NAND2_X1 U23318 ( .A1(n20332), .A2(n20331), .ZN(n20433) );
  AOI22_X1 U23319 ( .A1(n20334), .A2(n20335), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20433), .ZN(n20333) );
  OAI211_X1 U23320 ( .C1(n20351), .C2(n20526), .A(n20525), .B(n20333), .ZN(
        n20353) );
  INV_X1 U23321 ( .A(n20334), .ZN(n20336) );
  AOI22_X1 U23322 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20353), .B1(
        n20670), .B2(n20352), .ZN(n20337) );
  OAI211_X1 U23323 ( .C1(n20646), .C2(n20372), .A(n20338), .B(n20337), .ZN(
        P1_U3033) );
  AOI22_X1 U23324 ( .A1(n20721), .A2(n20647), .B1(n20351), .B2(n20680), .ZN(
        n20340) );
  AOI22_X1 U23325 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20353), .B1(
        n20681), .B2(n20352), .ZN(n20339) );
  OAI211_X1 U23326 ( .C1(n20650), .C2(n20372), .A(n20340), .B(n20339), .ZN(
        P1_U3034) );
  AOI22_X1 U23327 ( .A1(n20721), .A2(n20651), .B1(n20351), .B2(n20686), .ZN(
        n20342) );
  AOI22_X1 U23328 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20353), .B1(
        n20687), .B2(n20352), .ZN(n20341) );
  OAI211_X1 U23329 ( .C1(n20654), .C2(n20372), .A(n20342), .B(n20341), .ZN(
        P1_U3035) );
  AOI22_X1 U23330 ( .A1(n20721), .A2(n20608), .B1(n20692), .B2(n20351), .ZN(
        n20344) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20353), .B1(
        n20693), .B2(n20352), .ZN(n20343) );
  OAI211_X1 U23332 ( .C1(n20611), .C2(n20372), .A(n20344), .B(n20343), .ZN(
        P1_U3036) );
  AOI22_X1 U23333 ( .A1(n20721), .A2(n20578), .B1(n20351), .B2(n20698), .ZN(
        n20346) );
  AOI22_X1 U23334 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20353), .B1(
        n20699), .B2(n20352), .ZN(n20345) );
  OAI211_X1 U23335 ( .C1(n20581), .C2(n20372), .A(n20346), .B(n20345), .ZN(
        P1_U3037) );
  AOI22_X1 U23336 ( .A1(n20721), .A2(n20614), .B1(n20351), .B2(n20704), .ZN(
        n20348) );
  AOI22_X1 U23337 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20353), .B1(
        n20705), .B2(n20352), .ZN(n20347) );
  OAI211_X1 U23338 ( .C1(n20617), .C2(n20372), .A(n20348), .B(n20347), .ZN(
        P1_U3038) );
  AOI22_X1 U23339 ( .A1(n20721), .A2(n20657), .B1(n20351), .B2(n20710), .ZN(
        n20350) );
  AOI22_X1 U23340 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20353), .B1(
        n20711), .B2(n20352), .ZN(n20349) );
  OAI211_X1 U23341 ( .C1(n20662), .C2(n20372), .A(n20350), .B(n20349), .ZN(
        P1_U3039) );
  AOI22_X1 U23342 ( .A1(n20721), .A2(n20587), .B1(n20351), .B2(n20716), .ZN(
        n20355) );
  AOI22_X1 U23343 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20353), .B1(
        n20719), .B2(n20352), .ZN(n20354) );
  OAI211_X1 U23344 ( .C1(n20593), .C2(n20372), .A(n20355), .B(n20354), .ZN(
        P1_U3040) );
  AOI22_X1 U23345 ( .A1(n20670), .A2(n20367), .B1(n20669), .B2(n20366), .ZN(
        n20357) );
  AOI22_X1 U23346 ( .A1(n20369), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n20368), .B2(n20676), .ZN(n20356) );
  OAI211_X1 U23347 ( .C1(n20679), .C2(n20372), .A(n20357), .B(n20356), .ZN(
        P1_U3041) );
  AOI22_X1 U23348 ( .A1(n20681), .A2(n20367), .B1(n20680), .B2(n20366), .ZN(
        n20359) );
  AOI22_X1 U23349 ( .A1(n20369), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n20368), .B2(n20682), .ZN(n20358) );
  OAI211_X1 U23350 ( .C1(n20685), .C2(n20372), .A(n20359), .B(n20358), .ZN(
        P1_U3042) );
  AOI22_X1 U23351 ( .A1(n20693), .A2(n20367), .B1(n20692), .B2(n20366), .ZN(
        n20361) );
  AOI22_X1 U23352 ( .A1(n20369), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n20368), .B2(n20694), .ZN(n20360) );
  OAI211_X1 U23353 ( .C1(n20697), .C2(n20372), .A(n20361), .B(n20360), .ZN(
        P1_U3044) );
  AOI22_X1 U23354 ( .A1(n20699), .A2(n20367), .B1(n20698), .B2(n20366), .ZN(
        n20363) );
  AOI22_X1 U23355 ( .A1(n20369), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n20368), .B2(n20700), .ZN(n20362) );
  OAI211_X1 U23356 ( .C1(n20703), .C2(n20372), .A(n20363), .B(n20362), .ZN(
        P1_U3045) );
  AOI22_X1 U23357 ( .A1(n20705), .A2(n20367), .B1(n20704), .B2(n20366), .ZN(
        n20365) );
  AOI22_X1 U23358 ( .A1(n20369), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n20368), .B2(n20706), .ZN(n20364) );
  OAI211_X1 U23359 ( .C1(n20709), .C2(n20372), .A(n20365), .B(n20364), .ZN(
        P1_U3046) );
  AOI22_X1 U23360 ( .A1(n20711), .A2(n20367), .B1(n20710), .B2(n20366), .ZN(
        n20371) );
  AOI22_X1 U23361 ( .A1(n20369), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n20368), .B2(n20712), .ZN(n20370) );
  OAI211_X1 U23362 ( .C1(n20715), .C2(n20372), .A(n20371), .B(n20370), .ZN(
        P1_U3047) );
  INV_X1 U23363 ( .A(n20669), .ZN(n20373) );
  OAI22_X1 U23364 ( .A1(n20385), .A2(n20679), .B1(n20373), .B2(n20384), .ZN(
        n20374) );
  INV_X1 U23365 ( .A(n20374), .ZN(n20376) );
  AOI22_X1 U23366 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20388), .B1(
        n20670), .B2(n20387), .ZN(n20375) );
  OAI211_X1 U23367 ( .C1(n20646), .C2(n20425), .A(n20376), .B(n20375), .ZN(
        P1_U3049) );
  INV_X1 U23368 ( .A(n20686), .ZN(n20406) );
  OAI22_X1 U23369 ( .A1(n20385), .A2(n20691), .B1(n20406), .B2(n20384), .ZN(
        n20377) );
  INV_X1 U23370 ( .A(n20377), .ZN(n20379) );
  AOI22_X1 U23371 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20388), .B1(
        n20687), .B2(n20387), .ZN(n20378) );
  OAI211_X1 U23372 ( .C1(n20654), .C2(n20425), .A(n20379), .B(n20378), .ZN(
        P1_U3051) );
  INV_X1 U23373 ( .A(n20698), .ZN(n20380) );
  OAI22_X1 U23374 ( .A1(n20385), .A2(n20703), .B1(n20380), .B2(n20384), .ZN(
        n20381) );
  INV_X1 U23375 ( .A(n20381), .ZN(n20383) );
  AOI22_X1 U23376 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20388), .B1(
        n20699), .B2(n20387), .ZN(n20382) );
  OAI211_X1 U23377 ( .C1(n20581), .C2(n20425), .A(n20383), .B(n20382), .ZN(
        P1_U3053) );
  OAI22_X1 U23378 ( .A1(n20385), .A2(n20715), .B1(n20419), .B2(n20384), .ZN(
        n20386) );
  INV_X1 U23379 ( .A(n20386), .ZN(n20390) );
  AOI22_X1 U23380 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20388), .B1(
        n20711), .B2(n20387), .ZN(n20389) );
  OAI211_X1 U23381 ( .C1(n20662), .C2(n20425), .A(n20390), .B(n20389), .ZN(
        P1_U3055) );
  OR2_X1 U23382 ( .A1(n20594), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20423) );
  INV_X1 U23383 ( .A(n20423), .ZN(n20416) );
  AOI22_X1 U23384 ( .A1(n20452), .A2(n20676), .B1(n20416), .B2(n20669), .ZN(
        n20401) );
  NOR2_X1 U23385 ( .A1(n20393), .A2(n20392), .ZN(n20664) );
  AOI21_X1 U23386 ( .B1(n9847), .B2(n20664), .A(n20416), .ZN(n20398) );
  AOI21_X1 U23387 ( .B1(n20394), .B2(n20809), .A(n20598), .ZN(n20399) );
  INV_X1 U23388 ( .A(n20399), .ZN(n20395) );
  AOI22_X1 U23389 ( .A1(n20398), .A2(n20395), .B1(n20667), .B2(n20397), .ZN(
        n20396) );
  NAND2_X1 U23390 ( .A1(n20673), .A2(n20396), .ZN(n20428) );
  OAI22_X1 U23391 ( .A1(n20399), .A2(n20398), .B1(n20839), .B2(n20397), .ZN(
        n20427) );
  AOI22_X1 U23392 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20428), .B1(
        n20670), .B2(n20427), .ZN(n20400) );
  OAI211_X1 U23393 ( .C1(n20679), .C2(n20425), .A(n20401), .B(n20400), .ZN(
        P1_U3057) );
  OAI22_X1 U23394 ( .A1(n20425), .A2(n20685), .B1(n20402), .B2(n20423), .ZN(
        n20403) );
  INV_X1 U23395 ( .A(n20403), .ZN(n20405) );
  AOI22_X1 U23396 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20428), .B1(
        n20681), .B2(n20427), .ZN(n20404) );
  OAI211_X1 U23397 ( .C1(n20650), .C2(n20461), .A(n20405), .B(n20404), .ZN(
        P1_U3058) );
  OAI22_X1 U23398 ( .A1(n20425), .A2(n20691), .B1(n20406), .B2(n20423), .ZN(
        n20407) );
  INV_X1 U23399 ( .A(n20407), .ZN(n20409) );
  AOI22_X1 U23400 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20428), .B1(
        n20687), .B2(n20427), .ZN(n20408) );
  OAI211_X1 U23401 ( .C1(n20654), .C2(n20461), .A(n20409), .B(n20408), .ZN(
        P1_U3059) );
  OAI22_X1 U23402 ( .A1(n20425), .A2(n20697), .B1(n20410), .B2(n20423), .ZN(
        n20411) );
  INV_X1 U23403 ( .A(n20411), .ZN(n20413) );
  AOI22_X1 U23404 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20428), .B1(
        n20693), .B2(n20427), .ZN(n20412) );
  OAI211_X1 U23405 ( .C1(n20611), .C2(n20461), .A(n20413), .B(n20412), .ZN(
        P1_U3060) );
  AOI22_X1 U23406 ( .A1(n20452), .A2(n20700), .B1(n20416), .B2(n20698), .ZN(
        n20415) );
  AOI22_X1 U23407 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20428), .B1(
        n20699), .B2(n20427), .ZN(n20414) );
  OAI211_X1 U23408 ( .C1(n20703), .C2(n20425), .A(n20415), .B(n20414), .ZN(
        P1_U3061) );
  AOI22_X1 U23409 ( .A1(n20452), .A2(n20706), .B1(n20416), .B2(n20704), .ZN(
        n20418) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20428), .B1(
        n20705), .B2(n20427), .ZN(n20417) );
  OAI211_X1 U23411 ( .C1(n20709), .C2(n20425), .A(n20418), .B(n20417), .ZN(
        P1_U3062) );
  OAI22_X1 U23412 ( .A1(n20425), .A2(n20715), .B1(n20419), .B2(n20423), .ZN(
        n20420) );
  INV_X1 U23413 ( .A(n20420), .ZN(n20422) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20428), .B1(
        n20711), .B2(n20427), .ZN(n20421) );
  OAI211_X1 U23415 ( .C1(n20662), .C2(n20461), .A(n20422), .B(n20421), .ZN(
        P1_U3063) );
  OAI22_X1 U23416 ( .A1(n20425), .A2(n20726), .B1(n20424), .B2(n20423), .ZN(
        n20426) );
  INV_X1 U23417 ( .A(n20426), .ZN(n20430) );
  AOI22_X1 U23418 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20428), .B1(
        n20719), .B2(n20427), .ZN(n20429) );
  OAI211_X1 U23419 ( .C1(n20593), .C2(n20461), .A(n20430), .B(n20429), .ZN(
        P1_U3064) );
  NAND3_X1 U23420 ( .A1(n20487), .A2(n20518), .A3(n20809), .ZN(n20431) );
  OAI21_X1 U23421 ( .B1(n20433), .B2(n20432), .A(n20431), .ZN(n20456) );
  NOR2_X1 U23422 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20434), .ZN(
        n20455) );
  AOI22_X1 U23423 ( .A1(n20670), .A2(n20456), .B1(n20669), .B2(n20455), .ZN(
        n20441) );
  INV_X1 U23424 ( .A(n20487), .ZN(n20436) );
  OAI21_X1 U23425 ( .B1(n20452), .B2(n20457), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20435) );
  OAI21_X1 U23426 ( .B1(n20437), .B2(n20436), .A(n20435), .ZN(n20439) );
  OAI221_X1 U23427 ( .B1(n20455), .B2(n20526), .C1(n20455), .C2(n20439), .A(
        n20438), .ZN(n20458) );
  AOI22_X1 U23428 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20458), .B1(
        n20452), .B2(n20643), .ZN(n20440) );
  OAI211_X1 U23429 ( .C1(n20646), .C2(n20473), .A(n20441), .B(n20440), .ZN(
        P1_U3065) );
  AOI22_X1 U23430 ( .A1(n20681), .A2(n20456), .B1(n20680), .B2(n20455), .ZN(
        n20443) );
  AOI22_X1 U23431 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20682), .ZN(n20442) );
  OAI211_X1 U23432 ( .C1(n20685), .C2(n20461), .A(n20443), .B(n20442), .ZN(
        P1_U3066) );
  AOI22_X1 U23433 ( .A1(n20687), .A2(n20456), .B1(n20686), .B2(n20455), .ZN(
        n20445) );
  AOI22_X1 U23434 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20458), .B1(
        n20452), .B2(n20651), .ZN(n20444) );
  OAI211_X1 U23435 ( .C1(n20654), .C2(n20473), .A(n20445), .B(n20444), .ZN(
        P1_U3067) );
  AOI22_X1 U23436 ( .A1(n20693), .A2(n20456), .B1(n20692), .B2(n20455), .ZN(
        n20447) );
  AOI22_X1 U23437 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20694), .ZN(n20446) );
  OAI211_X1 U23438 ( .C1(n20697), .C2(n20461), .A(n20447), .B(n20446), .ZN(
        P1_U3068) );
  AOI22_X1 U23439 ( .A1(n20699), .A2(n20456), .B1(n20698), .B2(n20455), .ZN(
        n20449) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20458), .B1(
        n20452), .B2(n20578), .ZN(n20448) );
  OAI211_X1 U23441 ( .C1(n20581), .C2(n20473), .A(n20449), .B(n20448), .ZN(
        P1_U3069) );
  AOI22_X1 U23442 ( .A1(n20705), .A2(n20456), .B1(n20704), .B2(n20455), .ZN(
        n20451) );
  AOI22_X1 U23443 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20706), .ZN(n20450) );
  OAI211_X1 U23444 ( .C1(n20709), .C2(n20461), .A(n20451), .B(n20450), .ZN(
        P1_U3070) );
  AOI22_X1 U23445 ( .A1(n20711), .A2(n20456), .B1(n20710), .B2(n20455), .ZN(
        n20454) );
  AOI22_X1 U23446 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20458), .B1(
        n20452), .B2(n20657), .ZN(n20453) );
  OAI211_X1 U23447 ( .C1(n20662), .C2(n20473), .A(n20454), .B(n20453), .ZN(
        P1_U3071) );
  AOI22_X1 U23448 ( .A1(n20719), .A2(n20456), .B1(n20716), .B2(n20455), .ZN(
        n20460) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20720), .ZN(n20459) );
  OAI211_X1 U23450 ( .C1(n20726), .C2(n20461), .A(n20460), .B(n20459), .ZN(
        P1_U3072) );
  AOI22_X1 U23451 ( .A1(n20670), .A2(n20469), .B1(n20669), .B2(n20468), .ZN(
        n20463) );
  AOI22_X1 U23452 ( .A1(n20470), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n20481), .B2(n20676), .ZN(n20462) );
  OAI211_X1 U23453 ( .C1(n20679), .C2(n20473), .A(n20463), .B(n20462), .ZN(
        P1_U3073) );
  AOI22_X1 U23454 ( .A1(n20681), .A2(n20469), .B1(n20680), .B2(n20468), .ZN(
        n20465) );
  AOI22_X1 U23455 ( .A1(n20470), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n20481), .B2(n20682), .ZN(n20464) );
  OAI211_X1 U23456 ( .C1(n20685), .C2(n20473), .A(n20465), .B(n20464), .ZN(
        P1_U3074) );
  AOI22_X1 U23457 ( .A1(n20699), .A2(n20469), .B1(n20698), .B2(n20468), .ZN(
        n20467) );
  AOI22_X1 U23458 ( .A1(n20470), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n20481), .B2(n20700), .ZN(n20466) );
  OAI211_X1 U23459 ( .C1(n20703), .C2(n20473), .A(n20467), .B(n20466), .ZN(
        P1_U3077) );
  AOI22_X1 U23460 ( .A1(n20719), .A2(n20469), .B1(n20716), .B2(n20468), .ZN(
        n20472) );
  AOI22_X1 U23461 ( .A1(n20470), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n20481), .B2(n20720), .ZN(n20471) );
  OAI211_X1 U23462 ( .C1(n20726), .C2(n20473), .A(n20472), .B(n20471), .ZN(
        P1_U3080) );
  AOI22_X1 U23463 ( .A1(n20481), .A2(n20643), .B1(n20480), .B2(n20669), .ZN(
        n20475) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20483), .B1(
        n20670), .B2(n20482), .ZN(n20474) );
  OAI211_X1 U23465 ( .C1(n20646), .C2(n20508), .A(n20475), .B(n20474), .ZN(
        P1_U3081) );
  AOI22_X1 U23466 ( .A1(n20481), .A2(n20651), .B1(n20480), .B2(n20686), .ZN(
        n20477) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20483), .B1(
        n20687), .B2(n20482), .ZN(n20476) );
  OAI211_X1 U23468 ( .C1(n20654), .C2(n20508), .A(n20477), .B(n20476), .ZN(
        P1_U3083) );
  AOI22_X1 U23469 ( .A1(n20481), .A2(n20578), .B1(n20480), .B2(n20698), .ZN(
        n20479) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20483), .B1(
        n20699), .B2(n20482), .ZN(n20478) );
  OAI211_X1 U23471 ( .C1(n20581), .C2(n20508), .A(n20479), .B(n20478), .ZN(
        P1_U3085) );
  AOI22_X1 U23472 ( .A1(n20481), .A2(n20587), .B1(n20480), .B2(n20716), .ZN(
        n20485) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20483), .B1(
        n20719), .B2(n20482), .ZN(n20484) );
  OAI211_X1 U23474 ( .C1(n20593), .C2(n20508), .A(n20485), .B(n20484), .ZN(
        P1_U3088) );
  INV_X1 U23475 ( .A(n20486), .ZN(n20509) );
  AOI21_X1 U23476 ( .B1(n20487), .B2(n20664), .A(n20509), .ZN(n20489) );
  OAI22_X1 U23477 ( .A1(n20489), .A2(n20667), .B1(n20488), .B2(n20839), .ZN(
        n20510) );
  AOI22_X1 U23478 ( .A1(n20670), .A2(n20510), .B1(n20509), .B2(n20669), .ZN(
        n20495) );
  NOR2_X1 U23479 ( .A1(n20817), .A2(n20667), .ZN(n20490) );
  OAI21_X1 U23480 ( .B1(n20490), .B2(n20598), .A(n20489), .ZN(n20491) );
  OAI211_X1 U23481 ( .C1(n20492), .C2(n20809), .A(n20673), .B(n20491), .ZN(
        n20512) );
  NAND2_X1 U23482 ( .A1(n20817), .A2(n20493), .ZN(n20515) );
  AOI22_X1 U23483 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20512), .B1(
        n20543), .B2(n20676), .ZN(n20494) );
  OAI211_X1 U23484 ( .C1(n20679), .C2(n20508), .A(n20495), .B(n20494), .ZN(
        P1_U3089) );
  AOI22_X1 U23485 ( .A1(n20681), .A2(n20510), .B1(n20509), .B2(n20680), .ZN(
        n20497) );
  AOI22_X1 U23486 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20512), .B1(
        n20511), .B2(n20647), .ZN(n20496) );
  OAI211_X1 U23487 ( .C1(n20650), .C2(n20515), .A(n20497), .B(n20496), .ZN(
        P1_U3090) );
  AOI22_X1 U23488 ( .A1(n20687), .A2(n20510), .B1(n20509), .B2(n20686), .ZN(
        n20499) );
  AOI22_X1 U23489 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20512), .B1(
        n20511), .B2(n20651), .ZN(n20498) );
  OAI211_X1 U23490 ( .C1(n20654), .C2(n20515), .A(n20499), .B(n20498), .ZN(
        P1_U3091) );
  AOI22_X1 U23491 ( .A1(n20693), .A2(n20510), .B1(n20509), .B2(n20692), .ZN(
        n20501) );
  AOI22_X1 U23492 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20512), .B1(
        n20511), .B2(n20608), .ZN(n20500) );
  OAI211_X1 U23493 ( .C1(n20611), .C2(n20515), .A(n20501), .B(n20500), .ZN(
        P1_U3092) );
  AOI22_X1 U23494 ( .A1(n20699), .A2(n20510), .B1(n20509), .B2(n20698), .ZN(
        n20503) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20512), .B1(
        n20543), .B2(n20700), .ZN(n20502) );
  OAI211_X1 U23496 ( .C1(n20703), .C2(n20508), .A(n20503), .B(n20502), .ZN(
        P1_U3093) );
  AOI22_X1 U23497 ( .A1(n20705), .A2(n20510), .B1(n20509), .B2(n20704), .ZN(
        n20505) );
  AOI22_X1 U23498 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20512), .B1(
        n20511), .B2(n20614), .ZN(n20504) );
  OAI211_X1 U23499 ( .C1(n20617), .C2(n20515), .A(n20505), .B(n20504), .ZN(
        P1_U3094) );
  AOI22_X1 U23500 ( .A1(n20711), .A2(n20510), .B1(n20509), .B2(n20710), .ZN(
        n20507) );
  AOI22_X1 U23501 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20512), .B1(
        n20543), .B2(n20712), .ZN(n20506) );
  OAI211_X1 U23502 ( .C1(n20715), .C2(n20508), .A(n20507), .B(n20506), .ZN(
        P1_U3095) );
  AOI22_X1 U23503 ( .A1(n20719), .A2(n20510), .B1(n20509), .B2(n20716), .ZN(
        n20514) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20512), .B1(
        n20511), .B2(n20587), .ZN(n20513) );
  OAI211_X1 U23505 ( .C1(n20593), .C2(n20515), .A(n20514), .B(n20513), .ZN(
        P1_U3096) );
  NAND3_X1 U23506 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12111), .A3(
        n20517), .ZN(n20549) );
  NOR2_X1 U23507 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20549), .ZN(
        n20541) );
  AOI21_X1 U23508 ( .B1(n20595), .B2(n20518), .A(n20541), .ZN(n20522) );
  OAI22_X1 U23509 ( .A1(n20522), .A2(n20667), .B1(n20520), .B2(n20519), .ZN(
        n20542) );
  AOI22_X1 U23510 ( .A1(n20670), .A2(n20542), .B1(n20669), .B2(n20541), .ZN(
        n20528) );
  INV_X1 U23511 ( .A(n20573), .ZN(n20521) );
  OAI21_X1 U23512 ( .B1(n20521), .B2(n20543), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20523) );
  NAND2_X1 U23513 ( .A1(n20523), .A2(n20522), .ZN(n20524) );
  AOI22_X1 U23514 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20643), .ZN(n20527) );
  OAI211_X1 U23515 ( .C1(n20646), .C2(n20573), .A(n20528), .B(n20527), .ZN(
        P1_U3097) );
  AOI22_X1 U23516 ( .A1(n20681), .A2(n20542), .B1(n20680), .B2(n20541), .ZN(
        n20530) );
  AOI22_X1 U23517 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20647), .ZN(n20529) );
  OAI211_X1 U23518 ( .C1(n20650), .C2(n20573), .A(n20530), .B(n20529), .ZN(
        P1_U3098) );
  AOI22_X1 U23519 ( .A1(n20687), .A2(n20542), .B1(n20686), .B2(n20541), .ZN(
        n20532) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20651), .ZN(n20531) );
  OAI211_X1 U23521 ( .C1(n20654), .C2(n20573), .A(n20532), .B(n20531), .ZN(
        P1_U3099) );
  AOI22_X1 U23522 ( .A1(n20693), .A2(n20542), .B1(n20692), .B2(n20541), .ZN(
        n20534) );
  AOI22_X1 U23523 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20608), .ZN(n20533) );
  OAI211_X1 U23524 ( .C1(n20611), .C2(n20573), .A(n20534), .B(n20533), .ZN(
        P1_U3100) );
  AOI22_X1 U23525 ( .A1(n20699), .A2(n20542), .B1(n20698), .B2(n20541), .ZN(
        n20536) );
  AOI22_X1 U23526 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20578), .ZN(n20535) );
  OAI211_X1 U23527 ( .C1(n20581), .C2(n20573), .A(n20536), .B(n20535), .ZN(
        P1_U3101) );
  AOI22_X1 U23528 ( .A1(n20705), .A2(n20542), .B1(n20704), .B2(n20541), .ZN(
        n20538) );
  AOI22_X1 U23529 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20614), .ZN(n20537) );
  OAI211_X1 U23530 ( .C1(n20617), .C2(n20573), .A(n20538), .B(n20537), .ZN(
        P1_U3102) );
  AOI22_X1 U23531 ( .A1(n20711), .A2(n20542), .B1(n20710), .B2(n20541), .ZN(
        n20540) );
  AOI22_X1 U23532 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20657), .ZN(n20539) );
  OAI211_X1 U23533 ( .C1(n20662), .C2(n20573), .A(n20540), .B(n20539), .ZN(
        P1_U3103) );
  AOI22_X1 U23534 ( .A1(n20719), .A2(n20542), .B1(n20716), .B2(n20541), .ZN(
        n20546) );
  AOI22_X1 U23535 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20587), .ZN(n20545) );
  OAI211_X1 U23536 ( .C1(n20593), .C2(n20573), .A(n20546), .B(n20545), .ZN(
        P1_U3104) );
  NOR2_X1 U23537 ( .A1(n20547), .A2(n20549), .ZN(n20568) );
  AOI21_X1 U23538 ( .B1(n20595), .B2(n20548), .A(n20568), .ZN(n20550) );
  OAI22_X1 U23539 ( .A1(n20550), .A2(n20667), .B1(n20549), .B2(n20839), .ZN(
        n20569) );
  AOI22_X1 U23540 ( .A1(n20670), .A2(n20569), .B1(n20669), .B2(n20568), .ZN(
        n20555) );
  INV_X1 U23541 ( .A(n20549), .ZN(n20553) );
  INV_X1 U23542 ( .A(n20812), .ZN(n20551) );
  OAI211_X1 U23543 ( .C1(n20551), .C2(n20840), .A(n20550), .B(n20809), .ZN(
        n20552) );
  OAI211_X1 U23544 ( .C1(n20553), .C2(n20809), .A(n20552), .B(n20673), .ZN(
        n20570) );
  AOI22_X1 U23545 ( .A1(n20570), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n20588), .B2(n20676), .ZN(n20554) );
  OAI211_X1 U23546 ( .C1(n20679), .C2(n20573), .A(n20555), .B(n20554), .ZN(
        P1_U3105) );
  AOI22_X1 U23547 ( .A1(n20681), .A2(n20569), .B1(n20680), .B2(n20568), .ZN(
        n20557) );
  AOI22_X1 U23548 ( .A1(n20570), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n20588), .B2(n20682), .ZN(n20556) );
  OAI211_X1 U23549 ( .C1(n20685), .C2(n20573), .A(n20557), .B(n20556), .ZN(
        P1_U3106) );
  AOI22_X1 U23550 ( .A1(n20687), .A2(n20569), .B1(n20686), .B2(n20568), .ZN(
        n20559) );
  AOI22_X1 U23551 ( .A1(n20570), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n20588), .B2(n20688), .ZN(n20558) );
  OAI211_X1 U23552 ( .C1(n20691), .C2(n20573), .A(n20559), .B(n20558), .ZN(
        P1_U3107) );
  AOI22_X1 U23553 ( .A1(n20693), .A2(n20569), .B1(n20692), .B2(n20568), .ZN(
        n20561) );
  AOI22_X1 U23554 ( .A1(n20570), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n20588), .B2(n20694), .ZN(n20560) );
  OAI211_X1 U23555 ( .C1(n20697), .C2(n20573), .A(n20561), .B(n20560), .ZN(
        P1_U3108) );
  AOI22_X1 U23556 ( .A1(n20699), .A2(n20569), .B1(n20698), .B2(n20568), .ZN(
        n20563) );
  AOI22_X1 U23557 ( .A1(n20570), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n20588), .B2(n20700), .ZN(n20562) );
  OAI211_X1 U23558 ( .C1(n20703), .C2(n20573), .A(n20563), .B(n20562), .ZN(
        P1_U3109) );
  AOI22_X1 U23559 ( .A1(n20705), .A2(n20569), .B1(n20704), .B2(n20568), .ZN(
        n20565) );
  AOI22_X1 U23560 ( .A1(n20570), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n20588), .B2(n20706), .ZN(n20564) );
  OAI211_X1 U23561 ( .C1(n20709), .C2(n20573), .A(n20565), .B(n20564), .ZN(
        P1_U3110) );
  AOI22_X1 U23562 ( .A1(n20711), .A2(n20569), .B1(n20710), .B2(n20568), .ZN(
        n20567) );
  AOI22_X1 U23563 ( .A1(n20570), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n20588), .B2(n20712), .ZN(n20566) );
  OAI211_X1 U23564 ( .C1(n20715), .C2(n20573), .A(n20567), .B(n20566), .ZN(
        P1_U3111) );
  AOI22_X1 U23565 ( .A1(n20719), .A2(n20569), .B1(n20716), .B2(n20568), .ZN(
        n20572) );
  AOI22_X1 U23566 ( .A1(n20570), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n20588), .B2(n20720), .ZN(n20571) );
  OAI211_X1 U23567 ( .C1(n20726), .C2(n20573), .A(n20572), .B(n20571), .ZN(
        P1_U3112) );
  AOI22_X1 U23568 ( .A1(n20588), .A2(n20643), .B1(n20586), .B2(n20669), .ZN(
        n20575) );
  AOI22_X1 U23569 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20590), .B1(
        n20670), .B2(n20589), .ZN(n20574) );
  OAI211_X1 U23570 ( .C1(n20646), .C2(n20627), .A(n20575), .B(n20574), .ZN(
        P1_U3113) );
  AOI22_X1 U23571 ( .A1(n20588), .A2(n20647), .B1(n20586), .B2(n20680), .ZN(
        n20577) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20590), .B1(
        n20681), .B2(n20589), .ZN(n20576) );
  OAI211_X1 U23573 ( .C1(n20650), .C2(n20627), .A(n20577), .B(n20576), .ZN(
        P1_U3114) );
  AOI22_X1 U23574 ( .A1(n20588), .A2(n20578), .B1(n20586), .B2(n20698), .ZN(
        n20580) );
  AOI22_X1 U23575 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20590), .B1(
        n20699), .B2(n20589), .ZN(n20579) );
  OAI211_X1 U23576 ( .C1(n20581), .C2(n20627), .A(n20580), .B(n20579), .ZN(
        P1_U3117) );
  AOI22_X1 U23577 ( .A1(n20588), .A2(n20614), .B1(n20586), .B2(n20704), .ZN(
        n20583) );
  AOI22_X1 U23578 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20590), .B1(
        n20705), .B2(n20589), .ZN(n20582) );
  OAI211_X1 U23579 ( .C1(n20617), .C2(n20627), .A(n20583), .B(n20582), .ZN(
        P1_U3118) );
  AOI22_X1 U23580 ( .A1(n20588), .A2(n20657), .B1(n20586), .B2(n20710), .ZN(
        n20585) );
  AOI22_X1 U23581 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20590), .B1(
        n20711), .B2(n20589), .ZN(n20584) );
  OAI211_X1 U23582 ( .C1(n20662), .C2(n20627), .A(n20585), .B(n20584), .ZN(
        P1_U3119) );
  AOI22_X1 U23583 ( .A1(n20588), .A2(n20587), .B1(n20586), .B2(n20716), .ZN(
        n20592) );
  AOI22_X1 U23584 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20590), .B1(
        n20719), .B2(n20589), .ZN(n20591) );
  OAI211_X1 U23585 ( .C1(n20593), .C2(n20627), .A(n20592), .B(n20591), .ZN(
        P1_U3120) );
  NOR2_X1 U23586 ( .A1(n20594), .A2(n20825), .ZN(n20621) );
  AOI21_X1 U23587 ( .B1(n20595), .B2(n20664), .A(n20621), .ZN(n20597) );
  OAI22_X1 U23588 ( .A1(n20597), .A2(n20667), .B1(n20596), .B2(n20839), .ZN(
        n20622) );
  AOI22_X1 U23589 ( .A1(n20670), .A2(n20622), .B1(n20669), .B2(n20621), .ZN(
        n20603) );
  INV_X1 U23590 ( .A(n20596), .ZN(n20601) );
  NOR2_X1 U23591 ( .A1(n20812), .A2(n20667), .ZN(n20599) );
  OAI21_X1 U23592 ( .B1(n20599), .B2(n20598), .A(n20597), .ZN(n20600) );
  OAI211_X1 U23593 ( .C1(n20809), .C2(n20601), .A(n20673), .B(n20600), .ZN(
        n20624) );
  AOI22_X1 U23594 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20624), .B1(
        n20623), .B2(n20676), .ZN(n20602) );
  OAI211_X1 U23595 ( .C1(n20679), .C2(n20627), .A(n20603), .B(n20602), .ZN(
        P1_U3121) );
  AOI22_X1 U23596 ( .A1(n20681), .A2(n20622), .B1(n20680), .B2(n20621), .ZN(
        n20605) );
  AOI22_X1 U23597 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20624), .B1(
        n20623), .B2(n20682), .ZN(n20604) );
  OAI211_X1 U23598 ( .C1(n20685), .C2(n20627), .A(n20605), .B(n20604), .ZN(
        P1_U3122) );
  AOI22_X1 U23599 ( .A1(n20687), .A2(n20622), .B1(n20686), .B2(n20621), .ZN(
        n20607) );
  AOI22_X1 U23600 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20624), .B1(
        n20623), .B2(n20688), .ZN(n20606) );
  OAI211_X1 U23601 ( .C1(n20691), .C2(n20627), .A(n20607), .B(n20606), .ZN(
        P1_U3123) );
  AOI22_X1 U23602 ( .A1(n20693), .A2(n20622), .B1(n20692), .B2(n20621), .ZN(
        n20610) );
  AOI22_X1 U23603 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20624), .B1(
        n20618), .B2(n20608), .ZN(n20609) );
  OAI211_X1 U23604 ( .C1(n20611), .C2(n20636), .A(n20610), .B(n20609), .ZN(
        P1_U3124) );
  AOI22_X1 U23605 ( .A1(n20699), .A2(n20622), .B1(n20698), .B2(n20621), .ZN(
        n20613) );
  AOI22_X1 U23606 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20624), .B1(
        n20623), .B2(n20700), .ZN(n20612) );
  OAI211_X1 U23607 ( .C1(n20703), .C2(n20627), .A(n20613), .B(n20612), .ZN(
        P1_U3125) );
  AOI22_X1 U23608 ( .A1(n20705), .A2(n20622), .B1(n20704), .B2(n20621), .ZN(
        n20616) );
  AOI22_X1 U23609 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20624), .B1(
        n20618), .B2(n20614), .ZN(n20615) );
  OAI211_X1 U23610 ( .C1(n20617), .C2(n20636), .A(n20616), .B(n20615), .ZN(
        P1_U3126) );
  AOI22_X1 U23611 ( .A1(n20711), .A2(n20622), .B1(n20710), .B2(n20621), .ZN(
        n20620) );
  AOI22_X1 U23612 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20624), .B1(
        n20618), .B2(n20657), .ZN(n20619) );
  OAI211_X1 U23613 ( .C1(n20662), .C2(n20636), .A(n20620), .B(n20619), .ZN(
        P1_U3127) );
  AOI22_X1 U23614 ( .A1(n20719), .A2(n20622), .B1(n20716), .B2(n20621), .ZN(
        n20626) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20624), .B1(
        n20623), .B2(n20720), .ZN(n20625) );
  OAI211_X1 U23616 ( .C1(n20726), .C2(n20627), .A(n20626), .B(n20625), .ZN(
        P1_U3128) );
  AOI22_X1 U23617 ( .A1(n20639), .A2(n20694), .B1(n20631), .B2(n20692), .ZN(
        n20630) );
  INV_X1 U23618 ( .A(n20628), .ZN(n20633) );
  AOI22_X1 U23619 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20633), .B1(
        n20693), .B2(n20632), .ZN(n20629) );
  OAI211_X1 U23620 ( .C1(n20697), .C2(n20636), .A(n20630), .B(n20629), .ZN(
        P1_U3132) );
  AOI22_X1 U23621 ( .A1(n20639), .A2(n20700), .B1(n20631), .B2(n20698), .ZN(
        n20635) );
  AOI22_X1 U23622 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20633), .B1(
        n20699), .B2(n20632), .ZN(n20634) );
  OAI211_X1 U23623 ( .C1(n20703), .C2(n20636), .A(n20635), .B(n20634), .ZN(
        P1_U3133) );
  INV_X1 U23624 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n20885) );
  AOI22_X1 U23625 ( .A1(n20670), .A2(n20638), .B1(n20669), .B2(n20637), .ZN(
        n20641) );
  AOI22_X1 U23626 ( .A1(n20639), .A2(n20643), .B1(n20658), .B2(n20676), .ZN(
        n20640) );
  OAI211_X1 U23627 ( .C1(n20642), .C2(n20885), .A(n20641), .B(n20640), .ZN(
        P1_U3137) );
  AOI22_X1 U23628 ( .A1(n20670), .A2(n20656), .B1(n20669), .B2(n20655), .ZN(
        n20645) );
  AOI22_X1 U23629 ( .A1(n20659), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n20658), .B2(n20643), .ZN(n20644) );
  OAI211_X1 U23630 ( .C1(n20646), .C2(n20725), .A(n20645), .B(n20644), .ZN(
        P1_U3145) );
  AOI22_X1 U23631 ( .A1(n20681), .A2(n20656), .B1(n20680), .B2(n20655), .ZN(
        n20649) );
  AOI22_X1 U23632 ( .A1(n20659), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n20658), .B2(n20647), .ZN(n20648) );
  OAI211_X1 U23633 ( .C1(n20650), .C2(n20725), .A(n20649), .B(n20648), .ZN(
        P1_U3146) );
  AOI22_X1 U23634 ( .A1(n20687), .A2(n20656), .B1(n20686), .B2(n20655), .ZN(
        n20653) );
  AOI22_X1 U23635 ( .A1(n20659), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n20658), .B2(n20651), .ZN(n20652) );
  OAI211_X1 U23636 ( .C1(n20654), .C2(n20725), .A(n20653), .B(n20652), .ZN(
        P1_U3147) );
  AOI22_X1 U23637 ( .A1(n20711), .A2(n20656), .B1(n20710), .B2(n20655), .ZN(
        n20661) );
  AOI22_X1 U23638 ( .A1(n20659), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n20658), .B2(n20657), .ZN(n20660) );
  OAI211_X1 U23639 ( .C1(n20662), .C2(n20725), .A(n20661), .B(n20660), .ZN(
        P1_U3151) );
  INV_X1 U23640 ( .A(n20663), .ZN(n20717) );
  AOI21_X1 U23641 ( .B1(n20665), .B2(n20664), .A(n20717), .ZN(n20668) );
  OAI22_X1 U23642 ( .A1(n20668), .A2(n20667), .B1(n20666), .B2(n20839), .ZN(
        n20718) );
  AOI22_X1 U23643 ( .A1(n20670), .A2(n20718), .B1(n20717), .B2(n20669), .ZN(
        n20678) );
  INV_X1 U23644 ( .A(n20816), .ZN(n20671) );
  NOR2_X1 U23645 ( .A1(n20672), .A2(n20671), .ZN(n20674) );
  OAI21_X1 U23646 ( .B1(n20675), .B2(n20674), .A(n20673), .ZN(n20722) );
  AOI22_X1 U23647 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20722), .B1(
        n20721), .B2(n20676), .ZN(n20677) );
  OAI211_X1 U23648 ( .C1(n20679), .C2(n20725), .A(n20678), .B(n20677), .ZN(
        P1_U3153) );
  AOI22_X1 U23649 ( .A1(n20681), .A2(n20718), .B1(n20717), .B2(n20680), .ZN(
        n20684) );
  AOI22_X1 U23650 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20722), .B1(
        n20721), .B2(n20682), .ZN(n20683) );
  OAI211_X1 U23651 ( .C1(n20685), .C2(n20725), .A(n20684), .B(n20683), .ZN(
        P1_U3154) );
  AOI22_X1 U23652 ( .A1(n20687), .A2(n20718), .B1(n20717), .B2(n20686), .ZN(
        n20690) );
  AOI22_X1 U23653 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20722), .B1(
        n20721), .B2(n20688), .ZN(n20689) );
  OAI211_X1 U23654 ( .C1(n20691), .C2(n20725), .A(n20690), .B(n20689), .ZN(
        P1_U3155) );
  AOI22_X1 U23655 ( .A1(n20693), .A2(n20718), .B1(n20717), .B2(n20692), .ZN(
        n20696) );
  AOI22_X1 U23656 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20722), .B1(
        n20721), .B2(n20694), .ZN(n20695) );
  OAI211_X1 U23657 ( .C1(n20697), .C2(n20725), .A(n20696), .B(n20695), .ZN(
        P1_U3156) );
  AOI22_X1 U23658 ( .A1(n20699), .A2(n20718), .B1(n20717), .B2(n20698), .ZN(
        n20702) );
  AOI22_X1 U23659 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20722), .B1(
        n20721), .B2(n20700), .ZN(n20701) );
  OAI211_X1 U23660 ( .C1(n20703), .C2(n20725), .A(n20702), .B(n20701), .ZN(
        P1_U3157) );
  AOI22_X1 U23661 ( .A1(n20705), .A2(n20718), .B1(n20717), .B2(n20704), .ZN(
        n20708) );
  AOI22_X1 U23662 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20722), .B1(
        n20721), .B2(n20706), .ZN(n20707) );
  OAI211_X1 U23663 ( .C1(n20709), .C2(n20725), .A(n20708), .B(n20707), .ZN(
        P1_U3158) );
  AOI22_X1 U23664 ( .A1(n20711), .A2(n20718), .B1(n20717), .B2(n20710), .ZN(
        n20714) );
  AOI22_X1 U23665 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20722), .B1(
        n20721), .B2(n20712), .ZN(n20713) );
  OAI211_X1 U23666 ( .C1(n20715), .C2(n20725), .A(n20714), .B(n20713), .ZN(
        P1_U3159) );
  AOI22_X1 U23667 ( .A1(n20719), .A2(n20718), .B1(n20717), .B2(n20716), .ZN(
        n20724) );
  AOI22_X1 U23668 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20722), .B1(
        n20721), .B2(n20720), .ZN(n20723) );
  OAI211_X1 U23669 ( .C1(n20726), .C2(n20725), .A(n20724), .B(n20723), .ZN(
        P1_U3160) );
  NOR2_X1 U23670 ( .A1(n9918), .A2(n20727), .ZN(n20730) );
  INV_X1 U23671 ( .A(n20728), .ZN(n20729) );
  OAI21_X1 U23672 ( .B1(n20730), .B2(n20839), .A(n20729), .ZN(P1_U3163) );
  INV_X1 U23673 ( .A(n20731), .ZN(n20800) );
  AND2_X1 U23674 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20800), .ZN(
        P1_U3164) );
  AND2_X1 U23675 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20800), .ZN(
        P1_U3165) );
  AND2_X1 U23676 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20800), .ZN(
        P1_U3166) );
  AND2_X1 U23677 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20800), .ZN(
        P1_U3167) );
  AND2_X1 U23678 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20800), .ZN(
        P1_U3168) );
  AND2_X1 U23679 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20800), .ZN(
        P1_U3169) );
  AND2_X1 U23680 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20800), .ZN(
        P1_U3170) );
  AND2_X1 U23681 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20800), .ZN(
        P1_U3171) );
  AND2_X1 U23682 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20800), .ZN(
        P1_U3172) );
  AND2_X1 U23683 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20800), .ZN(
        P1_U3173) );
  AND2_X1 U23684 ( .A1(n20800), .A2(P1_DATAWIDTH_REG_21__SCAN_IN), .ZN(
        P1_U3174) );
  AND2_X1 U23685 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20800), .ZN(
        P1_U3175) );
  AND2_X1 U23686 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20800), .ZN(
        P1_U3176) );
  AND2_X1 U23687 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20800), .ZN(
        P1_U3177) );
  AND2_X1 U23688 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20800), .ZN(
        P1_U3178) );
  AND2_X1 U23689 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20800), .ZN(
        P1_U3179) );
  AND2_X1 U23690 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20800), .ZN(
        P1_U3180) );
  AND2_X1 U23691 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20800), .ZN(
        P1_U3181) );
  AND2_X1 U23692 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20800), .ZN(
        P1_U3182) );
  AND2_X1 U23693 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20800), .ZN(
        P1_U3183) );
  AND2_X1 U23694 ( .A1(n20800), .A2(P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(
        P1_U3184) );
  AND2_X1 U23695 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20800), .ZN(
        P1_U3185) );
  AND2_X1 U23696 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20800), .ZN(P1_U3186) );
  AND2_X1 U23697 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20800), .ZN(P1_U3187) );
  AND2_X1 U23698 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20800), .ZN(P1_U3188) );
  AND2_X1 U23699 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20800), .ZN(P1_U3189) );
  AND2_X1 U23700 ( .A1(n20800), .A2(P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(P1_U3190) );
  AND2_X1 U23701 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20800), .ZN(P1_U3191) );
  AND2_X1 U23702 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20800), .ZN(P1_U3192) );
  AND2_X1 U23703 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20800), .ZN(P1_U3193) );
  AOI21_X1 U23704 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20732), .A(n20738), 
        .ZN(n20745) );
  NOR2_X1 U23705 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20733) );
  OAI22_X1 U23706 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20737), .B1(n20733), 
        .B2(n20743), .ZN(n20734) );
  NOR2_X1 U23707 ( .A1(n20739), .A2(n20734), .ZN(n20735) );
  OAI22_X1 U23708 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20745), .B1(n20850), 
        .B2(n20735), .ZN(P1_U3194) );
  AOI222_X1 U23709 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20737), .B1(
        P1_STATE_REG_2__SCAN_IN), .B2(P1_STATE_REG_1__SCAN_IN), .C1(n20737), 
        .C2(n20736), .ZN(n20744) );
  NOR3_X1 U23710 ( .A1(NA), .A2(n20738), .A3(n20846), .ZN(n20740) );
  OAI22_X1 U23711 ( .A1(n20741), .A2(n20740), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20739), .ZN(n20742) );
  OAI22_X1 U23712 ( .A1(n20745), .A2(n20744), .B1(n20743), .B2(n20742), .ZN(
        P1_U3196) );
  NAND2_X1 U23713 ( .A1(n20850), .A2(n11789), .ZN(n20784) );
  INV_X1 U23714 ( .A(n20784), .ZN(n20789) );
  NAND2_X1 U23715 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20850), .ZN(n20787) );
  INV_X1 U23716 ( .A(n20787), .ZN(n20790) );
  AOI222_X1 U23717 ( .A1(n20789), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20836), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20790), .ZN(n20746) );
  INV_X1 U23718 ( .A(n20746), .ZN(P1_U3197) );
  AOI222_X1 U23719 ( .A1(n20790), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20836), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20789), .ZN(n20747) );
  INV_X1 U23720 ( .A(n20747), .ZN(P1_U3198) );
  OAI222_X1 U23721 ( .A1(n20787), .A2(n20749), .B1(n20748), .B2(n20850), .C1(
        n20750), .C2(n20784), .ZN(P1_U3199) );
  INV_X1 U23722 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20877) );
  OAI222_X1 U23723 ( .A1(n20784), .A2(n20752), .B1(n20877), .B2(n20850), .C1(
        n20750), .C2(n20787), .ZN(P1_U3200) );
  INV_X1 U23724 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20751) );
  OAI222_X1 U23725 ( .A1(n20787), .A2(n20752), .B1(n20751), .B2(n20850), .C1(
        n20754), .C2(n20784), .ZN(P1_U3201) );
  INV_X1 U23726 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20753) );
  OAI222_X1 U23727 ( .A1(n20787), .A2(n20754), .B1(n20753), .B2(n20850), .C1(
        n20756), .C2(n20784), .ZN(P1_U3202) );
  AOI22_X1 U23728 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20836), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n20789), .ZN(n20755) );
  OAI21_X1 U23729 ( .B1(n20756), .B2(n20787), .A(n20755), .ZN(P1_U3203) );
  AOI22_X1 U23730 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n20836), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n20790), .ZN(n20757) );
  OAI21_X1 U23731 ( .B1(n14294), .B2(n20784), .A(n20757), .ZN(P1_U3204) );
  INV_X1 U23732 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20758) );
  OAI222_X1 U23733 ( .A1(n20784), .A2(n14949), .B1(n20758), .B2(n20850), .C1(
        n14294), .C2(n20787), .ZN(P1_U3205) );
  INV_X1 U23734 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20759) );
  OAI222_X1 U23735 ( .A1(n20787), .A2(n14949), .B1(n20759), .B2(n20850), .C1(
        n15146), .C2(n20784), .ZN(P1_U3206) );
  AOI22_X1 U23736 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20836), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20789), .ZN(n20760) );
  OAI21_X1 U23737 ( .B1(n15146), .B2(n20787), .A(n20760), .ZN(P1_U3207) );
  AOI22_X1 U23738 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20836), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20790), .ZN(n20761) );
  OAI21_X1 U23739 ( .B1(n14939), .B2(n20784), .A(n20761), .ZN(P1_U3208) );
  AOI22_X1 U23740 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20836), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20789), .ZN(n20762) );
  OAI21_X1 U23741 ( .B1(n14939), .B2(n20787), .A(n20762), .ZN(P1_U3209) );
  AOI22_X1 U23742 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20836), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20790), .ZN(n20763) );
  OAI21_X1 U23743 ( .B1(n20764), .B2(n20784), .A(n20763), .ZN(P1_U3210) );
  AOI222_X1 U23744 ( .A1(n20790), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20836), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20789), .ZN(n20765) );
  INV_X1 U23745 ( .A(n20765), .ZN(P1_U3211) );
  AOI222_X1 U23746 ( .A1(n20790), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20836), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20789), .ZN(n20766) );
  INV_X1 U23747 ( .A(n20766), .ZN(P1_U3212) );
  INV_X1 U23748 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21096) );
  INV_X1 U23749 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20768) );
  OAI222_X1 U23750 ( .A1(n20784), .A2(n21096), .B1(n20768), .B2(n20850), .C1(
        n20767), .C2(n20787), .ZN(P1_U3213) );
  INV_X1 U23751 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20769) );
  OAI222_X1 U23752 ( .A1(n20784), .A2(n20771), .B1(n20769), .B2(n20850), .C1(
        n21096), .C2(n20787), .ZN(P1_U3214) );
  AOI22_X1 U23753 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20836), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20789), .ZN(n20770) );
  OAI21_X1 U23754 ( .B1(n20771), .B2(n20787), .A(n20770), .ZN(P1_U3215) );
  INV_X1 U23755 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20773) );
  AOI22_X1 U23756 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20836), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20790), .ZN(n20772) );
  OAI21_X1 U23757 ( .B1(n20773), .B2(n20784), .A(n20772), .ZN(P1_U3216) );
  INV_X1 U23758 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20774) );
  OAI222_X1 U23759 ( .A1(n20784), .A2(n20776), .B1(n20774), .B2(n20850), .C1(
        n20773), .C2(n20787), .ZN(P1_U3217) );
  INV_X1 U23760 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20775) );
  OAI222_X1 U23761 ( .A1(n20787), .A2(n20776), .B1(n20775), .B2(n20850), .C1(
        n20778), .C2(n20784), .ZN(P1_U3218) );
  INV_X1 U23762 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20777) );
  OAI222_X1 U23763 ( .A1(n20787), .A2(n20778), .B1(n20777), .B2(n20850), .C1(
        n20780), .C2(n20784), .ZN(P1_U3219) );
  AOI22_X1 U23764 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n20789), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20836), .ZN(n20779) );
  OAI21_X1 U23765 ( .B1(n20780), .B2(n20787), .A(n20779), .ZN(P1_U3220) );
  INV_X1 U23766 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20855) );
  OAI222_X1 U23767 ( .A1(n20787), .A2(n14636), .B1(n20855), .B2(n20850), .C1(
        n20782), .C2(n20784), .ZN(P1_U3221) );
  INV_X1 U23768 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20781) );
  OAI222_X1 U23769 ( .A1(n20787), .A2(n20782), .B1(n20781), .B2(n20850), .C1(
        n21163), .C2(n20784), .ZN(P1_U3222) );
  INV_X1 U23770 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20783) );
  INV_X1 U23771 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20786) );
  OAI222_X1 U23772 ( .A1(n20787), .A2(n21163), .B1(n20783), .B2(n20850), .C1(
        n20786), .C2(n20784), .ZN(P1_U3223) );
  INV_X1 U23773 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20785) );
  OAI222_X1 U23774 ( .A1(n20787), .A2(n20786), .B1(n20785), .B2(n20850), .C1(
        n21141), .C2(n20784), .ZN(P1_U3224) );
  AOI222_X1 U23775 ( .A1(n20789), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20836), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20790), .ZN(n20788) );
  INV_X1 U23776 ( .A(n20788), .ZN(P1_U3225) );
  AOI222_X1 U23777 ( .A1(n20790), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20836), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20789), .ZN(n20791) );
  INV_X1 U23778 ( .A(n20791), .ZN(P1_U3226) );
  INV_X1 U23779 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20792) );
  AOI22_X1 U23780 ( .A1(n20850), .A2(n20793), .B1(n20792), .B2(n20836), .ZN(
        P1_U3458) );
  INV_X1 U23781 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20830) );
  INV_X1 U23782 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20794) );
  AOI22_X1 U23783 ( .A1(n20850), .A2(n20830), .B1(n20794), .B2(n20836), .ZN(
        P1_U3459) );
  INV_X1 U23784 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20795) );
  AOI22_X1 U23785 ( .A1(n20850), .A2(n20796), .B1(n20795), .B2(n20836), .ZN(
        P1_U3460) );
  INV_X1 U23786 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20833) );
  INV_X1 U23787 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20797) );
  AOI22_X1 U23788 ( .A1(n20850), .A2(n20833), .B1(n20797), .B2(n20836), .ZN(
        P1_U3461) );
  INV_X1 U23789 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20828) );
  INV_X1 U23790 ( .A(n20798), .ZN(n20799) );
  AOI21_X1 U23791 ( .B1(n20828), .B2(n20800), .A(n20799), .ZN(P1_U3464) );
  AOI21_X1 U23792 ( .B1(n20800), .B2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n20799), 
        .ZN(n20801) );
  INV_X1 U23793 ( .A(n20801), .ZN(P1_U3465) );
  AOI22_X1 U23794 ( .A1(n20805), .A2(n20804), .B1(n20803), .B2(n20802), .ZN(
        n20806) );
  INV_X1 U23795 ( .A(n20806), .ZN(n20808) );
  MUX2_X1 U23796 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20808), .S(
        n20807), .Z(P1_U3469) );
  INV_X1 U23797 ( .A(n20823), .ZN(n20826) );
  NAND2_X1 U23798 ( .A1(n20809), .A2(n20840), .ZN(n20821) );
  OAI21_X1 U23799 ( .B1(n20812), .B2(n20811), .A(n20810), .ZN(n20819) );
  INV_X1 U23800 ( .A(n20813), .ZN(n20814) );
  AOI22_X1 U23801 ( .A1(n20817), .A2(n20816), .B1(n20815), .B2(n20814), .ZN(
        n20818) );
  OAI211_X1 U23802 ( .C1(n20821), .C2(n20820), .A(n20819), .B(n20818), .ZN(
        n20822) );
  INV_X1 U23803 ( .A(n20822), .ZN(n20824) );
  AOI22_X1 U23804 ( .A1(n20826), .A2(n20825), .B1(n20824), .B2(n20823), .ZN(
        P1_U3475) );
  NOR3_X1 U23805 ( .A1(n20828), .A2(P1_REIP_REG_0__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .ZN(n20827) );
  AOI221_X1 U23806 ( .B1(n20829), .B2(n20828), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n20827), .ZN(n20831) );
  INV_X1 U23807 ( .A(n20835), .ZN(n20832) );
  AOI22_X1 U23808 ( .A1(n20835), .A2(n20831), .B1(n20830), .B2(n20832), .ZN(
        P1_U3481) );
  NOR2_X1 U23809 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20834) );
  AOI22_X1 U23810 ( .A1(n20835), .A2(n20834), .B1(n20833), .B2(n20832), .ZN(
        P1_U3482) );
  AOI22_X1 U23811 ( .A1(n20850), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20837), 
        .B2(n20836), .ZN(P1_U3483) );
  AOI211_X1 U23812 ( .C1(n20841), .C2(n20840), .A(n20839), .B(n20838), .ZN(
        n20842) );
  AOI21_X1 U23813 ( .B1(n20843), .B2(n9918), .A(n20842), .ZN(n20849) );
  AOI211_X1 U23814 ( .C1(n20847), .C2(n20846), .A(n20845), .B(n20844), .ZN(
        n20848) );
  MUX2_X1 U23815 ( .A(n20849), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20848), 
        .Z(P1_U3485) );
  MUX2_X1 U23816 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20850), .Z(P1_U3486) );
  INV_X1 U23817 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n20852) );
  AOI22_X1 U23818 ( .A1(n20852), .A2(keyinput108), .B1(keyinput6), .B2(n11176), 
        .ZN(n20851) );
  OAI221_X1 U23819 ( .B1(n20852), .B2(keyinput108), .C1(n11176), .C2(keyinput6), .A(n20851), .ZN(n20865) );
  INV_X1 U23820 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n20854) );
  AOI22_X1 U23821 ( .A1(n20855), .A2(keyinput1), .B1(keyinput15), .B2(n20854), 
        .ZN(n20853) );
  OAI221_X1 U23822 ( .B1(n20855), .B2(keyinput1), .C1(n20854), .C2(keyinput15), 
        .A(n20853), .ZN(n20864) );
  AOI22_X1 U23823 ( .A1(n20858), .A2(keyinput47), .B1(n20857), .B2(keyinput68), 
        .ZN(n20856) );
  OAI221_X1 U23824 ( .B1(n20858), .B2(keyinput47), .C1(n20857), .C2(keyinput68), .A(n20856), .ZN(n20863) );
  INV_X1 U23825 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n20861) );
  AOI22_X1 U23826 ( .A1(n20861), .A2(keyinput121), .B1(keyinput76), .B2(n20860), .ZN(n20859) );
  OAI221_X1 U23827 ( .B1(n20861), .B2(keyinput121), .C1(n20860), .C2(
        keyinput76), .A(n20859), .ZN(n20862) );
  NOR4_X1 U23828 ( .A1(n20865), .A2(n20864), .A3(n20863), .A4(n20862), .ZN(
        n21179) );
  AOI22_X1 U23829 ( .A1(n13853), .A2(keyinput62), .B1(n20867), .B2(keyinput2), 
        .ZN(n20866) );
  OAI221_X1 U23830 ( .B1(n13853), .B2(keyinput62), .C1(n20867), .C2(keyinput2), 
        .A(n20866), .ZN(n20871) );
  XNOR2_X1 U23831 ( .A(n20868), .B(keyinput8), .ZN(n20870) );
  XNOR2_X1 U23832 ( .A(n9930), .B(keyinput49), .ZN(n20869) );
  OR3_X1 U23833 ( .A1(n20871), .A2(n20870), .A3(n20869), .ZN(n20880) );
  INV_X1 U23834 ( .A(keyinput69), .ZN(n20874) );
  INV_X1 U23835 ( .A(keyinput58), .ZN(n20873) );
  AOI22_X1 U23836 ( .A1(n20874), .A2(P3_ADDRESS_REG_23__SCAN_IN), .B1(
        P2_CODEFETCH_REG_SCAN_IN), .B2(n20873), .ZN(n20872) );
  OAI221_X1 U23837 ( .B1(n20874), .B2(P3_ADDRESS_REG_23__SCAN_IN), .C1(n20873), 
        .C2(P2_CODEFETCH_REG_SCAN_IN), .A(n20872), .ZN(n20879) );
  INV_X1 U23838 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n20876) );
  AOI22_X1 U23839 ( .A1(n20877), .A2(keyinput48), .B1(n20876), .B2(keyinput106), .ZN(n20875) );
  OAI221_X1 U23840 ( .B1(n20877), .B2(keyinput48), .C1(n20876), .C2(
        keyinput106), .A(n20875), .ZN(n20878) );
  NOR3_X1 U23841 ( .A1(n20880), .A2(n20879), .A3(n20878), .ZN(n21178) );
  AOI22_X1 U23842 ( .A1(n20882), .A2(keyinput35), .B1(n11186), .B2(keyinput96), 
        .ZN(n20881) );
  OAI221_X1 U23843 ( .B1(n20882), .B2(keyinput35), .C1(n11186), .C2(keyinput96), .A(n20881), .ZN(n20978) );
  INV_X1 U23844 ( .A(DATAI_20_), .ZN(n20884) );
  AOI22_X1 U23845 ( .A1(n20885), .A2(keyinput41), .B1(keyinput16), .B2(n20884), 
        .ZN(n20883) );
  OAI221_X1 U23846 ( .B1(n20885), .B2(keyinput41), .C1(n20884), .C2(keyinput16), .A(n20883), .ZN(n20977) );
  INV_X1 U23847 ( .A(keyinput64), .ZN(n20887) );
  OAI22_X1 U23848 ( .A1(n20888), .A2(keyinput60), .B1(n20887), .B2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .ZN(n20886) );
  AOI221_X1 U23849 ( .B1(n20888), .B2(keyinput60), .C1(
        P1_DATAWIDTH_REG_21__SCAN_IN), .C2(n20887), .A(n20886), .ZN(n20909) );
  INV_X1 U23850 ( .A(keyinput11), .ZN(n20890) );
  OAI22_X1 U23851 ( .A1(keyinput52), .A2(n20891), .B1(n20890), .B2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20889) );
  AOI221_X1 U23852 ( .B1(n20891), .B2(keyinput52), .C1(n20890), .C2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A(n20889), .ZN(n20908) );
  INV_X1 U23853 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n20894) );
  INV_X1 U23854 ( .A(keyinput112), .ZN(n20893) );
  AOI22_X1 U23855 ( .A1(n20894), .A2(keyinput73), .B1(
        P2_DATAWIDTH_REG_11__SCAN_IN), .B2(n20893), .ZN(n20892) );
  OAI221_X1 U23856 ( .B1(n20894), .B2(keyinput73), .C1(n20893), .C2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A(n20892), .ZN(n20906) );
  INV_X1 U23857 ( .A(keyinput13), .ZN(n20896) );
  AOI22_X1 U23858 ( .A1(n12467), .A2(keyinput3), .B1(P3_LWORD_REG_4__SCAN_IN), 
        .B2(n20896), .ZN(n20895) );
  OAI221_X1 U23859 ( .B1(n12467), .B2(keyinput3), .C1(n20896), .C2(
        P3_LWORD_REG_4__SCAN_IN), .A(n20895), .ZN(n20905) );
  INV_X1 U23860 ( .A(DATAI_7_), .ZN(n20899) );
  AOI22_X1 U23861 ( .A1(n20899), .A2(keyinput28), .B1(keyinput111), .B2(n20898), .ZN(n20897) );
  OAI221_X1 U23862 ( .B1(n20899), .B2(keyinput28), .C1(n20898), .C2(
        keyinput111), .A(n20897), .ZN(n20904) );
  INV_X1 U23863 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n20902) );
  INV_X1 U23864 ( .A(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n20901) );
  AOI22_X1 U23865 ( .A1(n20902), .A2(keyinput61), .B1(keyinput127), .B2(n20901), .ZN(n20900) );
  OAI221_X1 U23866 ( .B1(n20902), .B2(keyinput61), .C1(n20901), .C2(
        keyinput127), .A(n20900), .ZN(n20903) );
  NOR4_X1 U23867 ( .A1(n20906), .A2(n20905), .A3(n20904), .A4(n20903), .ZN(
        n20907) );
  NAND3_X1 U23868 ( .A1(n20909), .A2(n20908), .A3(n20907), .ZN(n20976) );
  INV_X1 U23869 ( .A(keyinput84), .ZN(n20911) );
  AOI22_X1 U23870 ( .A1(n20912), .A2(keyinput55), .B1(P2_UWORD_REG_5__SCAN_IN), 
        .B2(n20911), .ZN(n20910) );
  OAI221_X1 U23871 ( .B1(n20912), .B2(keyinput55), .C1(n20911), .C2(
        P2_UWORD_REG_5__SCAN_IN), .A(n20910), .ZN(n20924) );
  INV_X1 U23872 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n20914) );
  AOI22_X1 U23873 ( .A1(n20915), .A2(keyinput43), .B1(n20914), .B2(keyinput21), 
        .ZN(n20913) );
  OAI221_X1 U23874 ( .B1(n20915), .B2(keyinput43), .C1(n20914), .C2(keyinput21), .A(n20913), .ZN(n20923) );
  INV_X1 U23875 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n20916) );
  XOR2_X1 U23876 ( .A(keyinput87), .B(n20916), .Z(n20921) );
  XOR2_X1 U23877 ( .A(n20917), .B(keyinput56), .Z(n20920) );
  XNOR2_X1 U23878 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B(keyinput90), .ZN(
        n20919) );
  XNOR2_X1 U23879 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput20), 
        .ZN(n20918) );
  NAND4_X1 U23880 ( .A1(n20921), .A2(n20920), .A3(n20919), .A4(n20918), .ZN(
        n20922) );
  NOR3_X1 U23881 ( .A1(n20924), .A2(n20923), .A3(n20922), .ZN(n20974) );
  AOI22_X1 U23882 ( .A1(n20927), .A2(keyinput125), .B1(n20926), .B2(keyinput46), .ZN(n20925) );
  OAI221_X1 U23883 ( .B1(n20927), .B2(keyinput125), .C1(n20926), .C2(
        keyinput46), .A(n20925), .ZN(n20940) );
  AOI22_X1 U23884 ( .A1(n20930), .A2(keyinput67), .B1(keyinput65), .B2(n20929), 
        .ZN(n20928) );
  OAI221_X1 U23885 ( .B1(n20930), .B2(keyinput67), .C1(n20929), .C2(keyinput65), .A(n20928), .ZN(n20939) );
  INV_X1 U23886 ( .A(READY21_REG_SCAN_IN), .ZN(n20933) );
  AOI22_X1 U23887 ( .A1(n20933), .A2(keyinput59), .B1(keyinput63), .B2(n20932), 
        .ZN(n20931) );
  OAI221_X1 U23888 ( .B1(n20933), .B2(keyinput59), .C1(n20932), .C2(keyinput63), .A(n20931), .ZN(n20938) );
  AOI22_X1 U23889 ( .A1(n20936), .A2(keyinput116), .B1(keyinput118), .B2(
        n20935), .ZN(n20934) );
  OAI221_X1 U23890 ( .B1(n20936), .B2(keyinput116), .C1(n20935), .C2(
        keyinput118), .A(n20934), .ZN(n20937) );
  NOR4_X1 U23891 ( .A1(n20940), .A2(n20939), .A3(n20938), .A4(n20937), .ZN(
        n20973) );
  INV_X1 U23892 ( .A(keyinput83), .ZN(n20942) );
  AOI22_X1 U23893 ( .A1(n14294), .A2(keyinput103), .B1(
        P2_LWORD_REG_13__SCAN_IN), .B2(n20942), .ZN(n20941) );
  OAI221_X1 U23894 ( .B1(n14294), .B2(keyinput103), .C1(n20942), .C2(
        P2_LWORD_REG_13__SCAN_IN), .A(n20941), .ZN(n20955) );
  INV_X1 U23895 ( .A(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n20944) );
  AOI22_X1 U23896 ( .A1(n20945), .A2(keyinput33), .B1(n20944), .B2(keyinput19), 
        .ZN(n20943) );
  OAI221_X1 U23897 ( .B1(n20945), .B2(keyinput33), .C1(n20944), .C2(keyinput19), .A(n20943), .ZN(n20954) );
  INV_X1 U23898 ( .A(keyinput95), .ZN(n20947) );
  AOI22_X1 U23899 ( .A1(n20948), .A2(keyinput30), .B1(P2_UWORD_REG_14__SCAN_IN), .B2(n20947), .ZN(n20946) );
  OAI221_X1 U23900 ( .B1(n20948), .B2(keyinput30), .C1(n20947), .C2(
        P2_UWORD_REG_14__SCAN_IN), .A(n20946), .ZN(n20953) );
  AOI22_X1 U23901 ( .A1(n20951), .A2(keyinput82), .B1(n20950), .B2(keyinput104), .ZN(n20949) );
  OAI221_X1 U23902 ( .B1(n20951), .B2(keyinput82), .C1(n20950), .C2(
        keyinput104), .A(n20949), .ZN(n20952) );
  NOR4_X1 U23903 ( .A1(n20955), .A2(n20954), .A3(n20953), .A4(n20952), .ZN(
        n20972) );
  AOI22_X1 U23904 ( .A1(n20958), .A2(keyinput75), .B1(keyinput7), .B2(n20957), 
        .ZN(n20956) );
  OAI221_X1 U23905 ( .B1(n20958), .B2(keyinput75), .C1(n20957), .C2(keyinput7), 
        .A(n20956), .ZN(n20970) );
  AOI22_X1 U23906 ( .A1(n20960), .A2(keyinput14), .B1(n13642), .B2(keyinput45), 
        .ZN(n20959) );
  OAI221_X1 U23907 ( .B1(n20960), .B2(keyinput14), .C1(n13642), .C2(keyinput45), .A(n20959), .ZN(n20969) );
  AOI22_X1 U23908 ( .A1(n20963), .A2(keyinput70), .B1(n20962), .B2(keyinput74), 
        .ZN(n20961) );
  OAI221_X1 U23909 ( .B1(n20963), .B2(keyinput70), .C1(n20962), .C2(keyinput74), .A(n20961), .ZN(n20968) );
  INV_X1 U23910 ( .A(keyinput5), .ZN(n20965) );
  AOI22_X1 U23911 ( .A1(n20966), .A2(keyinput107), .B1(P1_UWORD_REG_2__SCAN_IN), .B2(n20965), .ZN(n20964) );
  OAI221_X1 U23912 ( .B1(n20966), .B2(keyinput107), .C1(n20965), .C2(
        P1_UWORD_REG_2__SCAN_IN), .A(n20964), .ZN(n20967) );
  NOR4_X1 U23913 ( .A1(n20970), .A2(n20969), .A3(n20968), .A4(n20967), .ZN(
        n20971) );
  NAND4_X1 U23914 ( .A1(n20974), .A2(n20973), .A3(n20972), .A4(n20971), .ZN(
        n20975) );
  NOR4_X1 U23915 ( .A1(n20978), .A2(n20977), .A3(n20976), .A4(n20975), .ZN(
        n21177) );
  NOR4_X1 U23916 ( .A1(keyinput35), .A2(keyinput96), .A3(keyinput3), .A4(
        keyinput13), .ZN(n20979) );
  NAND3_X1 U23917 ( .A1(keyinput73), .A2(keyinput112), .A3(n20979), .ZN(n20991) );
  NAND2_X1 U23918 ( .A1(keyinput58), .A2(keyinput106), .ZN(n20980) );
  NOR3_X1 U23919 ( .A1(keyinput48), .A2(keyinput69), .A3(n20980), .ZN(n20989)
         );
  NAND2_X1 U23920 ( .A1(keyinput2), .A2(keyinput49), .ZN(n20981) );
  NOR3_X1 U23921 ( .A1(keyinput8), .A2(keyinput62), .A3(n20981), .ZN(n20988)
         );
  NOR2_X1 U23922 ( .A1(keyinput64), .A2(keyinput127), .ZN(n20982) );
  NAND3_X1 U23923 ( .A1(keyinput60), .A2(keyinput61), .A3(n20982), .ZN(n20986)
         );
  NAND4_X1 U23924 ( .A1(keyinput52), .A2(keyinput11), .A3(keyinput28), .A4(
        keyinput111), .ZN(n20985) );
  NAND4_X1 U23925 ( .A1(keyinput121), .A2(keyinput76), .A3(keyinput47), .A4(
        keyinput68), .ZN(n20984) );
  NAND4_X1 U23926 ( .A1(keyinput1), .A2(keyinput15), .A3(keyinput108), .A4(
        keyinput6), .ZN(n20983) );
  NOR4_X1 U23927 ( .A1(n20986), .A2(n20985), .A3(n20984), .A4(n20983), .ZN(
        n20987) );
  NAND3_X1 U23928 ( .A1(n20989), .A2(n20988), .A3(n20987), .ZN(n20990) );
  NOR4_X1 U23929 ( .A1(keyinput41), .A2(keyinput16), .A3(n20991), .A4(n20990), 
        .ZN(n21175) );
  INV_X1 U23930 ( .A(keyinput116), .ZN(n20992) );
  NAND4_X1 U23931 ( .A1(keyinput118), .A2(keyinput59), .A3(keyinput63), .A4(
        n20992), .ZN(n21042) );
  NOR2_X1 U23932 ( .A1(keyinput125), .A2(keyinput65), .ZN(n20993) );
  NAND3_X1 U23933 ( .A1(keyinput67), .A2(keyinput46), .A3(n20993), .ZN(n21041)
         );
  NOR2_X1 U23934 ( .A1(keyinput84), .A2(keyinput21), .ZN(n20994) );
  NAND3_X1 U23935 ( .A1(keyinput43), .A2(keyinput55), .A3(n20994), .ZN(n20995)
         );
  NOR3_X1 U23936 ( .A1(keyinput56), .A2(keyinput20), .A3(n20995), .ZN(n21004)
         );
  NOR2_X1 U23937 ( .A1(keyinput5), .A2(keyinput74), .ZN(n20996) );
  NAND3_X1 U23938 ( .A1(keyinput107), .A2(keyinput70), .A3(n20996), .ZN(n21002) );
  INV_X1 U23939 ( .A(keyinput7), .ZN(n20997) );
  NAND4_X1 U23940 ( .A1(keyinput45), .A2(keyinput14), .A3(keyinput75), .A4(
        n20997), .ZN(n21001) );
  NAND4_X1 U23941 ( .A1(keyinput103), .A2(keyinput83), .A3(keyinput95), .A4(
        keyinput30), .ZN(n21000) );
  NOR2_X1 U23942 ( .A1(keyinput33), .A2(keyinput82), .ZN(n20998) );
  NAND3_X1 U23943 ( .A1(keyinput19), .A2(keyinput104), .A3(n20998), .ZN(n20999) );
  NOR4_X1 U23944 ( .A1(n21002), .A2(n21001), .A3(n21000), .A4(n20999), .ZN(
        n21003) );
  NAND4_X1 U23945 ( .A1(keyinput87), .A2(keyinput90), .A3(n21004), .A4(n21003), 
        .ZN(n21040) );
  NAND4_X1 U23946 ( .A1(keyinput81), .A2(keyinput92), .A3(keyinput18), .A4(
        keyinput78), .ZN(n21020) );
  INV_X1 U23947 ( .A(keyinput88), .ZN(n21005) );
  NAND4_X1 U23948 ( .A1(keyinput57), .A2(keyinput98), .A3(keyinput44), .A4(
        n21005), .ZN(n21019) );
  NOR2_X1 U23949 ( .A1(keyinput40), .A2(keyinput53), .ZN(n21006) );
  NAND3_X1 U23950 ( .A1(keyinput102), .A2(keyinput36), .A3(n21006), .ZN(n21007) );
  NOR3_X1 U23951 ( .A1(keyinput17), .A2(keyinput110), .A3(n21007), .ZN(n21008)
         );
  NAND3_X1 U23952 ( .A1(keyinput27), .A2(keyinput85), .A3(n21008), .ZN(n21018)
         );
  INV_X1 U23953 ( .A(keyinput105), .ZN(n21009) );
  NOR4_X1 U23954 ( .A1(keyinput99), .A2(keyinput119), .A3(keyinput31), .A4(
        n21009), .ZN(n21016) );
  NAND2_X1 U23955 ( .A1(keyinput124), .A2(keyinput101), .ZN(n21010) );
  NOR3_X1 U23956 ( .A1(keyinput79), .A2(keyinput66), .A3(n21010), .ZN(n21015)
         );
  NAND2_X1 U23957 ( .A1(keyinput0), .A2(keyinput123), .ZN(n21011) );
  NOR3_X1 U23958 ( .A1(keyinput10), .A2(keyinput91), .A3(n21011), .ZN(n21014)
         );
  NAND2_X1 U23959 ( .A1(keyinput100), .A2(keyinput89), .ZN(n21012) );
  NOR3_X1 U23960 ( .A1(keyinput115), .A2(keyinput42), .A3(n21012), .ZN(n21013)
         );
  NAND4_X1 U23961 ( .A1(n21016), .A2(n21015), .A3(n21014), .A4(n21013), .ZN(
        n21017) );
  NOR4_X1 U23962 ( .A1(n21020), .A2(n21019), .A3(n21018), .A4(n21017), .ZN(
        n21038) );
  INV_X1 U23963 ( .A(keyinput72), .ZN(n21021) );
  NOR4_X1 U23964 ( .A1(keyinput50), .A2(keyinput113), .A3(keyinput32), .A4(
        n21021), .ZN(n21037) );
  NAND2_X1 U23965 ( .A1(keyinput23), .A2(keyinput122), .ZN(n21022) );
  NOR3_X1 U23966 ( .A1(keyinput22), .A2(keyinput80), .A3(n21022), .ZN(n21036)
         );
  INV_X1 U23967 ( .A(keyinput39), .ZN(n21023) );
  NAND4_X1 U23968 ( .A1(keyinput54), .A2(keyinput34), .A3(keyinput77), .A4(
        n21023), .ZN(n21030) );
  NOR2_X1 U23969 ( .A1(keyinput120), .A2(keyinput86), .ZN(n21024) );
  NAND3_X1 U23970 ( .A1(keyinput9), .A2(keyinput126), .A3(n21024), .ZN(n21029)
         );
  INV_X1 U23971 ( .A(keyinput71), .ZN(n21025) );
  NAND4_X1 U23972 ( .A1(keyinput29), .A2(keyinput51), .A3(keyinput97), .A4(
        n21025), .ZN(n21028) );
  NOR2_X1 U23973 ( .A1(keyinput94), .A2(keyinput12), .ZN(n21026) );
  NAND3_X1 U23974 ( .A1(keyinput24), .A2(keyinput117), .A3(n21026), .ZN(n21027) );
  NOR4_X1 U23975 ( .A1(n21030), .A2(n21029), .A3(n21028), .A4(n21027), .ZN(
        n21033) );
  NAND4_X1 U23976 ( .A1(keyinput4), .A2(keyinput26), .A3(keyinput25), .A4(
        keyinput109), .ZN(n21031) );
  NOR3_X1 U23977 ( .A1(keyinput38), .A2(keyinput114), .A3(n21031), .ZN(n21032)
         );
  NAND3_X1 U23978 ( .A1(n21033), .A2(n21032), .A3(keyinput37), .ZN(n21034) );
  NOR2_X1 U23979 ( .A1(keyinput93), .A2(n21034), .ZN(n21035) );
  NAND4_X1 U23980 ( .A1(n21038), .A2(n21037), .A3(n21036), .A4(n21035), .ZN(
        n21039) );
  NOR4_X1 U23981 ( .A1(n21042), .A2(n21041), .A3(n21040), .A4(n21039), .ZN(
        n21174) );
  AOI22_X1 U23982 ( .A1(n21045), .A2(keyinput98), .B1(n21044), .B2(keyinput57), 
        .ZN(n21043) );
  OAI221_X1 U23983 ( .B1(n21045), .B2(keyinput98), .C1(n21044), .C2(keyinput57), .A(n21043), .ZN(n21057) );
  AOI22_X1 U23984 ( .A1(n21048), .A2(keyinput88), .B1(keyinput44), .B2(n21047), 
        .ZN(n21046) );
  OAI221_X1 U23985 ( .B1(n21048), .B2(keyinput88), .C1(n21047), .C2(keyinput44), .A(n21046), .ZN(n21056) );
  AOI22_X1 U23986 ( .A1(n21050), .A2(keyinput81), .B1(n11242), .B2(keyinput92), 
        .ZN(n21049) );
  OAI221_X1 U23987 ( .B1(n21050), .B2(keyinput81), .C1(n11242), .C2(keyinput92), .A(n21049), .ZN(n21055) );
  INV_X1 U23988 ( .A(keyinput18), .ZN(n21052) );
  AOI22_X1 U23989 ( .A1(n21053), .A2(keyinput78), .B1(
        P1_DATAWIDTH_REG_11__SCAN_IN), .B2(n21052), .ZN(n21051) );
  OAI221_X1 U23990 ( .B1(n21053), .B2(keyinput78), .C1(n21052), .C2(
        P1_DATAWIDTH_REG_11__SCAN_IN), .A(n21051), .ZN(n21054) );
  NOR4_X1 U23991 ( .A1(n21057), .A2(n21056), .A3(n21055), .A4(n21054), .ZN(
        n21104) );
  AOI22_X1 U23992 ( .A1(n21060), .A2(keyinput101), .B1(keyinput79), .B2(n21059), .ZN(n21058) );
  OAI221_X1 U23993 ( .B1(n21060), .B2(keyinput101), .C1(n21059), .C2(
        keyinput79), .A(n21058), .ZN(n21071) );
  AOI22_X1 U23994 ( .A1(n21062), .A2(keyinput124), .B1(n11018), .B2(keyinput66), .ZN(n21061) );
  OAI221_X1 U23995 ( .B1(n21062), .B2(keyinput124), .C1(n11018), .C2(
        keyinput66), .A(n21061), .ZN(n21070) );
  AOI22_X1 U23996 ( .A1(n21064), .A2(keyinput99), .B1(keyinput119), .B2(n12238), .ZN(n21063) );
  OAI221_X1 U23997 ( .B1(n21064), .B2(keyinput99), .C1(n12238), .C2(
        keyinput119), .A(n21063), .ZN(n21069) );
  AOI22_X1 U23998 ( .A1(n21067), .A2(keyinput31), .B1(n21066), .B2(keyinput105), .ZN(n21065) );
  OAI221_X1 U23999 ( .B1(n21067), .B2(keyinput31), .C1(n21066), .C2(
        keyinput105), .A(n21065), .ZN(n21068) );
  NOR4_X1 U24000 ( .A1(n21071), .A2(n21070), .A3(n21069), .A4(n21068), .ZN(
        n21103) );
  INV_X1 U24001 ( .A(keyinput89), .ZN(n21073) );
  AOI22_X1 U24002 ( .A1(n21074), .A2(keyinput115), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n21073), .ZN(n21072) );
  OAI221_X1 U24003 ( .B1(n21074), .B2(keyinput115), .C1(n21073), .C2(
        P1_DATAO_REG_18__SCAN_IN), .A(n21072), .ZN(n21086) );
  AOI22_X1 U24004 ( .A1(n21077), .A2(keyinput100), .B1(n21076), .B2(keyinput42), .ZN(n21075) );
  OAI221_X1 U24005 ( .B1(n21077), .B2(keyinput100), .C1(n21076), .C2(
        keyinput42), .A(n21075), .ZN(n21085) );
  INV_X1 U24006 ( .A(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n21080) );
  INV_X1 U24007 ( .A(keyinput10), .ZN(n21079) );
  AOI22_X1 U24008 ( .A1(n21080), .A2(keyinput123), .B1(
        P2_BYTEENABLE_REG_0__SCAN_IN), .B2(n21079), .ZN(n21078) );
  OAI221_X1 U24009 ( .B1(n21080), .B2(keyinput123), .C1(n21079), .C2(
        P2_BYTEENABLE_REG_0__SCAN_IN), .A(n21078), .ZN(n21084) );
  AOI22_X1 U24010 ( .A1(n21082), .A2(keyinput91), .B1(n13158), .B2(keyinput0), 
        .ZN(n21081) );
  OAI221_X1 U24011 ( .B1(n21082), .B2(keyinput91), .C1(n13158), .C2(keyinput0), 
        .A(n21081), .ZN(n21083) );
  NOR4_X1 U24012 ( .A1(n21086), .A2(n21085), .A3(n21084), .A4(n21083), .ZN(
        n21102) );
  INV_X1 U24013 ( .A(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n21088) );
  AOI22_X1 U24014 ( .A1(n21089), .A2(keyinput27), .B1(n21088), .B2(keyinput85), 
        .ZN(n21087) );
  OAI221_X1 U24015 ( .B1(n21089), .B2(keyinput27), .C1(n21088), .C2(keyinput85), .A(n21087), .ZN(n21100) );
  INV_X1 U24016 ( .A(keyinput40), .ZN(n21091) );
  AOI22_X1 U24017 ( .A1(n21092), .A2(keyinput102), .B1(
        P3_DATAO_REG_23__SCAN_IN), .B2(n21091), .ZN(n21090) );
  OAI221_X1 U24018 ( .B1(n21092), .B2(keyinput102), .C1(n21091), .C2(
        P3_DATAO_REG_23__SCAN_IN), .A(n21090), .ZN(n21099) );
  AOI22_X1 U24019 ( .A1(n10736), .A2(keyinput17), .B1(keyinput110), .B2(n21094), .ZN(n21093) );
  OAI221_X1 U24020 ( .B1(n10736), .B2(keyinput17), .C1(n21094), .C2(
        keyinput110), .A(n21093), .ZN(n21098) );
  AOI22_X1 U24021 ( .A1(n21096), .A2(keyinput53), .B1(n11610), .B2(keyinput36), 
        .ZN(n21095) );
  OAI221_X1 U24022 ( .B1(n21096), .B2(keyinput53), .C1(n11610), .C2(keyinput36), .A(n21095), .ZN(n21097) );
  NOR4_X1 U24023 ( .A1(n21100), .A2(n21099), .A3(n21098), .A4(n21097), .ZN(
        n21101) );
  NAND4_X1 U24024 ( .A1(n21104), .A2(n21103), .A3(n21102), .A4(n21101), .ZN(
        n21173) );
  INV_X1 U24025 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n21106) );
  AOI22_X1 U24026 ( .A1(n21107), .A2(keyinput22), .B1(keyinput122), .B2(n21106), .ZN(n21105) );
  OAI221_X1 U24027 ( .B1(n21107), .B2(keyinput22), .C1(n21106), .C2(
        keyinput122), .A(n21105), .ZN(n21120) );
  INV_X1 U24028 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n21110) );
  AOI22_X1 U24029 ( .A1(n21110), .A2(keyinput80), .B1(keyinput23), .B2(n21109), 
        .ZN(n21108) );
  OAI221_X1 U24030 ( .B1(n21110), .B2(keyinput80), .C1(n21109), .C2(keyinput23), .A(n21108), .ZN(n21119) );
  INV_X1 U24031 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n21113) );
  INV_X1 U24032 ( .A(keyinput50), .ZN(n21112) );
  AOI22_X1 U24033 ( .A1(n21113), .A2(keyinput72), .B1(P1_UWORD_REG_8__SCAN_IN), 
        .B2(n21112), .ZN(n21111) );
  OAI221_X1 U24034 ( .B1(n21113), .B2(keyinput72), .C1(n21112), .C2(
        P1_UWORD_REG_8__SCAN_IN), .A(n21111), .ZN(n21118) );
  INV_X1 U24035 ( .A(keyinput32), .ZN(n21115) );
  AOI22_X1 U24036 ( .A1(n21116), .A2(keyinput113), .B1(
        P3_DATAWIDTH_REG_20__SCAN_IN), .B2(n21115), .ZN(n21114) );
  OAI221_X1 U24037 ( .B1(n21116), .B2(keyinput113), .C1(n21115), .C2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A(n21114), .ZN(n21117) );
  NOR4_X1 U24038 ( .A1(n21120), .A2(n21119), .A3(n21118), .A4(n21117), .ZN(
        n21171) );
  AOI22_X1 U24039 ( .A1(n21123), .A2(keyinput120), .B1(keyinput9), .B2(n21122), 
        .ZN(n21121) );
  OAI221_X1 U24040 ( .B1(n21123), .B2(keyinput120), .C1(n21122), .C2(keyinput9), .A(n21121), .ZN(n21136) );
  AOI22_X1 U24041 ( .A1(n21126), .A2(keyinput126), .B1(keyinput86), .B2(n21125), .ZN(n21124) );
  OAI221_X1 U24042 ( .B1(n21126), .B2(keyinput126), .C1(n21125), .C2(
        keyinput86), .A(n21124), .ZN(n21135) );
  INV_X1 U24043 ( .A(keyinput54), .ZN(n21128) );
  AOI22_X1 U24044 ( .A1(n21129), .A2(keyinput39), .B1(
        P2_READREQUEST_REG_SCAN_IN), .B2(n21128), .ZN(n21127) );
  OAI221_X1 U24045 ( .B1(n21129), .B2(keyinput39), .C1(n21128), .C2(
        P2_READREQUEST_REG_SCAN_IN), .A(n21127), .ZN(n21134) );
  AOI22_X1 U24046 ( .A1(n21132), .A2(keyinput34), .B1(keyinput77), .B2(n21131), 
        .ZN(n21130) );
  OAI221_X1 U24047 ( .B1(n21132), .B2(keyinput34), .C1(n21131), .C2(keyinput77), .A(n21130), .ZN(n21133) );
  NOR4_X1 U24048 ( .A1(n21136), .A2(n21135), .A3(n21134), .A4(n21133), .ZN(
        n21170) );
  AOI22_X1 U24049 ( .A1(n21139), .A2(keyinput94), .B1(n21138), .B2(keyinput24), 
        .ZN(n21137) );
  OAI221_X1 U24050 ( .B1(n21139), .B2(keyinput94), .C1(n21138), .C2(keyinput24), .A(n21137), .ZN(n21152) );
  INV_X1 U24051 ( .A(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n21142) );
  AOI22_X1 U24052 ( .A1(n21142), .A2(keyinput12), .B1(keyinput117), .B2(n21141), .ZN(n21140) );
  OAI221_X1 U24053 ( .B1(n21142), .B2(keyinput12), .C1(n21141), .C2(
        keyinput117), .A(n21140), .ZN(n21151) );
  INV_X1 U24054 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n21145) );
  INV_X1 U24055 ( .A(keyinput29), .ZN(n21144) );
  AOI22_X1 U24056 ( .A1(n21145), .A2(keyinput51), .B1(P3_DATAO_REG_7__SCAN_IN), 
        .B2(n21144), .ZN(n21143) );
  OAI221_X1 U24057 ( .B1(n21145), .B2(keyinput51), .C1(n21144), .C2(
        P3_DATAO_REG_7__SCAN_IN), .A(n21143), .ZN(n21150) );
  INV_X1 U24058 ( .A(DATAI_24_), .ZN(n21147) );
  AOI22_X1 U24059 ( .A1(n21148), .A2(keyinput71), .B1(n21147), .B2(keyinput97), 
        .ZN(n21146) );
  OAI221_X1 U24060 ( .B1(n21148), .B2(keyinput71), .C1(n21147), .C2(keyinput97), .A(n21146), .ZN(n21149) );
  NOR4_X1 U24061 ( .A1(n21152), .A2(n21151), .A3(n21150), .A4(n21149), .ZN(
        n21169) );
  INV_X1 U24062 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n21155) );
  AOI22_X1 U24063 ( .A1(n21155), .A2(keyinput4), .B1(keyinput26), .B2(n21154), 
        .ZN(n21153) );
  OAI221_X1 U24064 ( .B1(n21155), .B2(keyinput4), .C1(n21154), .C2(keyinput26), 
        .A(n21153), .ZN(n21167) );
  INV_X1 U24065 ( .A(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n21157) );
  AOI22_X1 U24066 ( .A1(n11638), .A2(keyinput38), .B1(keyinput114), .B2(n21157), .ZN(n21156) );
  OAI221_X1 U24067 ( .B1(n11638), .B2(keyinput38), .C1(n21157), .C2(
        keyinput114), .A(n21156), .ZN(n21166) );
  INV_X1 U24068 ( .A(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n21160) );
  AOI22_X1 U24069 ( .A1(n21160), .A2(keyinput25), .B1(keyinput109), .B2(n21159), .ZN(n21158) );
  OAI221_X1 U24070 ( .B1(n21160), .B2(keyinput25), .C1(n21159), .C2(
        keyinput109), .A(n21158), .ZN(n21165) );
  INV_X1 U24071 ( .A(keyinput93), .ZN(n21162) );
  AOI22_X1 U24072 ( .A1(n21163), .A2(keyinput37), .B1(
        P2_DATAWIDTH_REG_4__SCAN_IN), .B2(n21162), .ZN(n21161) );
  OAI221_X1 U24073 ( .B1(n21163), .B2(keyinput37), .C1(n21162), .C2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A(n21161), .ZN(n21164) );
  NOR4_X1 U24074 ( .A1(n21167), .A2(n21166), .A3(n21165), .A4(n21164), .ZN(
        n21168) );
  NAND4_X1 U24075 ( .A1(n21171), .A2(n21170), .A3(n21169), .A4(n21168), .ZN(
        n21172) );
  AOI211_X1 U24076 ( .C1(n21175), .C2(n21174), .A(n21173), .B(n21172), .ZN(
        n21176) );
  NAND4_X1 U24077 ( .A1(n21179), .A2(n21178), .A3(n21177), .A4(n21176), .ZN(
        n21192) );
  INV_X1 U24078 ( .A(n21180), .ZN(n21183) );
  AOI222_X1 U24079 ( .A1(n21186), .A2(n21185), .B1(n21184), .B2(n21183), .C1(
        n21182), .C2(n21181), .ZN(n21188) );
  AOI22_X1 U24080 ( .A1(n21190), .A2(n21189), .B1(n21188), .B2(n21187), .ZN(
        n21191) );
  XNOR2_X1 U24081 ( .A(n21192), .B(n21191), .ZN(P3_U3289) );
  OR2_X2 U11193 ( .A1(n16259), .A2(n16260), .ZN(n16257) );
  AND2_X2 U12413 ( .A1(n13175), .A2(n13135), .ZN(n13176) );
  INV_X2 U11299 ( .A(n19173), .ZN(n10058) );
  NOR2_X2 U12460 ( .A1(n13161), .A2(n14411), .ZN(n13156) );
  NOR2_X2 U12462 ( .A1(n13167), .A2(n16347), .ZN(n13168) );
  NOR2_X2 U12463 ( .A1(n13165), .A2(n16340), .ZN(n13166) );
  NOR2_X2 U16331 ( .A1(n16272), .A2(n16273), .ZN(n16271) );
  NOR2_X2 U12026 ( .A1(n13283), .A2(n13285), .ZN(n13284) );
  INV_X1 U11203 ( .A(n18313), .ZN(n18959) );
  OR2_X1 U13966 ( .A1(n11102), .A2(n15847), .ZN(n19699) );
  AND2_X1 U12667 ( .A1(n10060), .A2(n10059), .ZN(n16299) );
  AND2_X2 U13244 ( .A1(n10794), .A2(n10456), .ZN(n10469) );
  OR2_X1 U13764 ( .A1(n11493), .A2(n11394), .ZN(n11205) );
  NAND2_X1 U11534 ( .A1(n11205), .A2(n11204), .ZN(n11225) );
  NOR2_X1 U12595 ( .A1(n9893), .A2(n9850), .ZN(n11294) );
  CLKBUF_X2 U11197 ( .A(n11695), .Z(n12559) );
  XNOR2_X1 U11213 ( .A(n11921), .B(n11920), .ZN(n12157) );
  OR2_X1 U11236 ( .A1(n15952), .A2(n10058), .ZN(n10060) );
  OR2_X1 U11238 ( .A1(n19035), .A2(n9836), .ZN(n10071) );
  CLKBUF_X2 U11246 ( .A(n11635), .Z(n11644) );
  NOR2_X1 U11247 ( .A1(n13162), .A2(n13164), .ZN(n13163) );
  CLKBUF_X1 U11262 ( .A(n13006), .Z(n9773) );
  INV_X1 U11302 ( .A(n15138), .ZN(n15089) );
  CLKBUF_X1 U11320 ( .A(n12157), .Z(n15167) );
  NOR2_X1 U11345 ( .A1(n10058), .A2(n16252), .ZN(n13184) );
  NOR2_X1 U11430 ( .A1(n16271), .A2(n10058), .ZN(n16259) );
  CLKBUF_X1 U11437 ( .A(n16696), .Z(n17029) );
  CLKBUF_X1 U11586 ( .A(n20239), .Z(n20248) );
  AND2_X1 U11755 ( .A1(n10056), .A2(n10054), .ZN(n13240) );
  CLKBUF_X1 U11757 ( .A(n13356), .Z(n19361) );
  CLKBUF_X1 U11815 ( .A(n10331), .Z(n9748) );
  NOR2_X1 U12173 ( .A1(n16254), .A2(n16253), .ZN(n16252) );
  CLKBUF_X1 U12341 ( .A(n16655), .Z(n16654) );
endmodule

