

module b21_C_SARLock_k_128_6 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4393, n4396, n4397, n4398, n4399, n4400, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265;

  NAND2_X1 U4899 ( .A1(n9575), .A2(n9348), .ZN(n9576) );
  AND2_X1 U4901 ( .A1(n9362), .A2(n9361), .ZN(n9423) );
  AND2_X2 U4903 ( .A1(n6100), .A2(n6093), .ZN(n8307) );
  INV_X1 U4904 ( .A(n5996), .ZN(n8421) );
  AND2_X1 U4905 ( .A1(n8435), .A2(n5103), .ZN(n5241) );
  INV_X2 U4906 ( .A(n5412), .ZN(n5604) );
  NOR2_X1 U4907 ( .A1(n5933), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5935) );
  NOR2_X2 U4908 ( .A1(n6022), .A2(n5772), .ZN(n6123) );
  INV_X1 U4909 ( .A(n7777), .ZN(n4393) );
  INV_X1 U4911 ( .A(n4393), .ZN(P2_U3152) );
  NAND2_X1 U4912 ( .A1(n9594), .A2(n9340), .ZN(n9575) );
  NAND2_X1 U4913 ( .A1(n5872), .A2(n10150), .ZN(n5656) );
  INV_X1 U4914 ( .A(n8307), .ZN(n8298) );
  OAI21_X1 U4915 ( .B1(n9632), .B2(n4710), .A(n4492), .ZN(n9594) );
  INV_X1 U4916 ( .A(n9154), .ZN(n8150) );
  AND2_X1 U4917 ( .A1(n9403), .A2(n9402), .ZN(n9163) );
  NOR2_X1 U4918 ( .A1(n4590), .A2(n6022), .ZN(n4730) );
  NAND2_X1 U4919 ( .A1(n5105), .A2(n5103), .ZN(n5412) );
  INV_X1 U4920 ( .A(n7480), .ZN(n8297) );
  OAI21_X1 U4921 ( .B1(n8236), .B2(n4551), .A(n4548), .ZN(n9077) );
  INV_X1 U4922 ( .A(n8425), .ZN(n6030) );
  NOR2_X1 U4923 ( .A1(n9520), .A2(n9682), .ZN(n9511) );
  INV_X1 U4924 ( .A(n9590), .ZN(n9709) );
  INV_X1 U4925 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6320) );
  INV_X1 U4926 ( .A(n8367), .ZN(n5743) );
  NAND2_X1 U4927 ( .A1(n5729), .A2(n5572), .ZN(n8683) );
  AOI21_X1 U4928 ( .B1(n8811), .B2(n8634), .A(n8633), .ZN(n8798) );
  AOI21_X1 U4929 ( .B1(n4732), .B2(n9870), .A(n4731), .ZN(n9684) );
  INV_X1 U4930 ( .A(n5458), .ZN(n6980) );
  AND4_X1 U4931 ( .A1(n5774), .A2(n5773), .A3(n6232), .A4(n6680), .ZN(n4396)
         );
  INV_X1 U4932 ( .A(n5637), .ZN(n5294) );
  BUF_X4 U4933 ( .A(n5625), .Z(n4397) );
  NAND2_X1 U4934 ( .A1(n5210), .A2(n4402), .ZN(n5625) );
  AOI22_X2 U4935 ( .A1(n8748), .A2(n8761), .B1(n8641), .B2(n8755), .ZN(n8737)
         );
  NOR2_X2 U4936 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5949) );
  INV_X2 U4937 ( .A(n8365), .ZN(n5886) );
  INV_X1 U4938 ( .A(n4402), .ZN(n4398) );
  NAND2_X2 U4939 ( .A1(n4501), .A2(n4500), .ZN(n4960) );
  BUF_X8 U4940 ( .A(n4960), .Z(n4402) );
  INV_X1 U4941 ( .A(n8324), .ZN(n8300) );
  OR2_X1 U4942 ( .A1(n8899), .A2(n8697), .ZN(n5729) );
  OR2_X1 U4943 ( .A1(n7685), .A2(n4828), .ZN(n4835) );
  AND2_X1 U4944 ( .A1(n5491), .A2(n5490), .ZN(n8773) );
  NAND2_X1 U4945 ( .A1(n6787), .A2(n6786), .ZN(n6788) );
  NAND2_X1 U4946 ( .A1(n8473), .A2(n8474), .ZN(n8472) );
  INV_X2 U4947 ( .A(n9610), .ZN(n4399) );
  NAND2_X2 U4948 ( .A1(n5657), .A2(n5656), .ZN(n5806) );
  OR2_X1 U4949 ( .A1(n8568), .A2(n10156), .ZN(n5679) );
  INV_X1 U4950 ( .A(n4639), .ZN(n10156) );
  INV_X2 U4951 ( .A(n4637), .ZN(n10150) );
  OAI211_X1 U4952 ( .C1(n5219), .C2(n6180), .A(n5211), .B(n4638), .ZN(n4637)
         );
  AOI21_X1 U4953 ( .B1(n5163), .B2(n4975), .A(n4949), .ZN(n5149) );
  INV_X1 U4954 ( .A(n5965), .ZN(n8149) );
  INV_X2 U4955 ( .A(n4402), .ZN(n6179) );
  AND4_X1 U4956 ( .A1(n4634), .A2(n4448), .A3(n5077), .A4(n5076), .ZN(n4591)
         );
  CLKBUF_X2 U4957 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n10129) );
  AOI211_X1 U4958 ( .C1(n5749), .C2(n5748), .A(n5747), .B(n5746), .ZN(n5767)
         );
  NOR3_X1 U4959 ( .A1(n5749), .A2(n10145), .A3(n5677), .ZN(n5747) );
  OAI21_X1 U4960 ( .B1(n9436), .B2(n9435), .A(n9434), .ZN(n9446) );
  NAND2_X1 U4961 ( .A1(n4612), .A2(n4611), .ZN(n5749) );
  AOI21_X1 U4962 ( .B1(n9773), .B2(n10107), .A(n4701), .ZN(n4700) );
  AOI21_X1 U4963 ( .B1(n4613), .B2(n4615), .A(n5855), .ZN(n4611) );
  INV_X1 U4964 ( .A(n4614), .ZN(n4613) );
  AOI211_X1 U4965 ( .C1(n9687), .C2(n9884), .A(n9531), .B(n9530), .ZN(n9532)
         );
  OAI21_X1 U4966 ( .B1(n5635), .B2(n5634), .A(n4416), .ZN(n4615) );
  XNOR2_X1 U4967 ( .A(n8507), .B(n4517), .ZN(n8511) );
  OAI211_X1 U4968 ( .C1(n4471), .C2(n9187), .A(n4903), .B(n4902), .ZN(n9686)
         );
  AOI21_X1 U4969 ( .B1(n5591), .B2(n8684), .A(n5590), .ZN(n5594) );
  AOI21_X1 U4970 ( .B1(n4498), .B2(n9870), .A(n4495), .ZN(n9690) );
  OR2_X1 U4971 ( .A1(n9517), .A2(n4904), .ZN(n4903) );
  NOR2_X1 U4972 ( .A1(n9518), .A2(n9527), .ZN(n9517) );
  NAND2_X1 U4973 ( .A1(n4519), .A2(n4518), .ZN(n8450) );
  NAND2_X1 U4974 ( .A1(n4486), .A2(n5732), .ZN(n5733) );
  OAI21_X1 U4975 ( .B1(n8737), .B2(n4842), .A(n4841), .ZN(n4843) );
  NAND2_X1 U4976 ( .A1(n8357), .A2(n8356), .ZN(n8449) );
  OR2_X1 U4977 ( .A1(n8879), .A2(n6611), .ZN(n5638) );
  OR2_X1 U4978 ( .A1(n9158), .A2(n9192), .ZN(n9394) );
  NAND2_X1 U4979 ( .A1(n9150), .A2(n9149), .ZN(n9192) );
  OAI21_X1 U4980 ( .B1(n9559), .B2(n4924), .A(n4922), .ZN(n9533) );
  NAND2_X1 U4981 ( .A1(n5627), .A2(n5626), .ZN(n8879) );
  NAND2_X1 U4982 ( .A1(n8402), .A2(n8401), .ZN(n9559) );
  NAND2_X1 U4983 ( .A1(n8713), .A2(n8714), .ZN(n5725) );
  NAND2_X1 U4984 ( .A1(n5602), .A2(n5601), .ZN(n8623) );
  NAND2_X1 U4985 ( .A1(n4531), .A2(n4530), .ZN(n9132) );
  NAND2_X1 U4986 ( .A1(n8637), .A2(n4948), .ZN(n8785) );
  OR2_X1 U4987 ( .A1(n9583), .A2(n4762), .ZN(n9520) );
  AND2_X1 U4988 ( .A1(n4891), .A2(n5724), .ZN(n4890) );
  NAND2_X1 U4989 ( .A1(n8366), .A2(n8698), .ZN(n8699) );
  XNOR2_X1 U4990 ( .A(n5614), .B(SI_30_), .ZN(n9152) );
  AOI21_X1 U4991 ( .B1(n4925), .B2(n4923), .A(n4433), .ZN(n4922) );
  INV_X1 U4992 ( .A(n9423), .ZN(n9540) );
  OR2_X1 U4993 ( .A1(n9688), .A2(n8429), .ZN(n9365) );
  INV_X1 U4994 ( .A(n4844), .ZN(n4842) );
  AOI21_X1 U4995 ( .B1(n4844), .B2(n5516), .A(n4418), .ZN(n4841) );
  INV_X1 U4996 ( .A(n5729), .ZN(n4887) );
  NAND2_X1 U4997 ( .A1(n8306), .A2(n8305), .ZN(n9688) );
  AND2_X1 U4998 ( .A1(n5724), .A2(n5534), .ZN(n8714) );
  NAND2_X1 U4999 ( .A1(n4428), .A2(n4544), .ZN(n4543) );
  OR2_X1 U5000 ( .A1(n8910), .A2(n8696), .ZN(n5724) );
  NAND2_X1 U5001 ( .A1(n5087), .A2(n5086), .ZN(n8906) );
  AND2_X1 U5002 ( .A1(n5722), .A2(n5535), .ZN(n8725) );
  OR2_X1 U5003 ( .A1(n9703), .A2(n9582), .ZN(n9254) );
  XNOR2_X1 U5004 ( .A(n5576), .B(n5575), .ZN(n8303) );
  NAND2_X1 U5005 ( .A1(n5114), .A2(n5113), .ZN(n8910) );
  NAND2_X1 U5006 ( .A1(n8257), .A2(n8256), .ZN(n9703) );
  NAND2_X1 U5007 ( .A1(n4663), .A2(n5558), .ZN(n5576) );
  OR2_X1 U5008 ( .A1(n8914), .A2(n8642), .ZN(n5722) );
  XNOR2_X1 U5009 ( .A(n5542), .B(n5541), .ZN(n8270) );
  NAND2_X1 U5010 ( .A1(n4835), .A2(n4832), .ZN(n7871) );
  NAND2_X1 U5011 ( .A1(n7885), .A2(n5703), .ZN(n7863) );
  XNOR2_X1 U5012 ( .A(n5556), .B(n5557), .ZN(n8287) );
  NAND2_X1 U5013 ( .A1(n5556), .A2(n5557), .ZN(n4663) );
  NAND2_X1 U5014 ( .A1(n5544), .A2(n5543), .ZN(n5556) );
  NAND2_X1 U5015 ( .A1(n8921), .A2(n8763), .ZN(n5721) );
  XNOR2_X1 U5016 ( .A(n5112), .B(n5111), .ZN(n8254) );
  NAND2_X1 U5017 ( .A1(n7682), .A2(n4893), .ZN(n7885) );
  NAND2_X1 U5018 ( .A1(n4912), .A2(n4911), .ZN(n7747) );
  INV_X1 U5019 ( .A(n9608), .ZN(n9714) );
  NAND2_X1 U5020 ( .A1(n4688), .A2(n4692), .ZN(n5544) );
  OAI21_X1 U5021 ( .B1(n5522), .B2(n5062), .A(n5061), .ZN(n5112) );
  AND2_X1 U5022 ( .A1(n5652), .A2(n8790), .ZN(n8804) );
  INV_X1 U5023 ( .A(n9617), .ZN(n9717) );
  OR2_X1 U5024 ( .A1(n8926), .A2(n8641), .ZN(n5649) );
  AND2_X1 U5025 ( .A1(n8225), .A2(n8224), .ZN(n9608) );
  NAND2_X1 U5026 ( .A1(n5138), .A2(n5137), .ZN(n8921) );
  NAND2_X1 U5027 ( .A1(n8171), .A2(n8170), .ZN(n9728) );
  INV_X1 U5028 ( .A(n8773), .ZN(n8931) );
  AND2_X1 U5029 ( .A1(n8211), .A2(n8210), .ZN(n9617) );
  NAND2_X1 U5030 ( .A1(n5501), .A2(n5500), .ZN(n8926) );
  NAND2_X1 U5031 ( .A1(n8192), .A2(n8191), .ZN(n9723) );
  NOR2_X1 U5032 ( .A1(n4957), .A2(n8962), .ZN(n8864) );
  OR2_X1 U5033 ( .A1(n7791), .A2(n7790), .ZN(n7793) );
  XNOR2_X1 U5034 ( .A(n5475), .B(n5474), .ZN(n8168) );
  NAND2_X1 U5035 ( .A1(n7326), .A2(n4633), .ZN(n7329) );
  OAI21_X1 U5036 ( .B1(n5499), .B2(n5498), .A(n5052), .ZN(n5136) );
  NAND2_X1 U5037 ( .A1(n8008), .A2(n8007), .ZN(n9105) );
  NAND2_X1 U5038 ( .A1(n5443), .A2(n5442), .ZN(n8946) );
  INV_X4 U5039 ( .A(n9568), .ZN(n8404) );
  INV_X1 U5040 ( .A(n4829), .ZN(n4836) );
  AND2_X1 U5041 ( .A1(n5043), .A2(n5472), .ZN(n5489) );
  AOI21_X1 U5042 ( .B1(n4740), .B2(n4743), .A(n4738), .ZN(n4737) );
  OAI21_X1 U5043 ( .B1(n7686), .B2(n4830), .A(n4452), .ZN(n4829) );
  AND2_X1 U5044 ( .A1(n4821), .A2(n7599), .ZN(n7985) );
  NAND2_X1 U5045 ( .A1(n7906), .A2(n7905), .ZN(n9745) );
  AOI21_X1 U5046 ( .B1(n4866), .B2(n4865), .A(n4864), .ZN(n4863) );
  AND2_X1 U5047 ( .A1(n5386), .A2(n5702), .ZN(n7686) );
  AOI21_X1 U5048 ( .B1(n4721), .B2(n4720), .A(n4719), .ZN(n4718) );
  AND2_X1 U5049 ( .A1(n4741), .A2(n7628), .ZN(n4740) );
  NAND2_X1 U5050 ( .A1(n5814), .A2(n5813), .ZN(n7526) );
  OR2_X1 U5051 ( .A1(n7979), .A2(n9136), .ZN(n9310) );
  OR2_X1 U5052 ( .A1(n8967), .A2(n7898), .ZN(n5703) );
  NAND2_X1 U5053 ( .A1(n7831), .A2(n7830), .ZN(n9750) );
  NAND2_X1 U5054 ( .A1(n7750), .A2(n7749), .ZN(n9754) );
  NAND2_X1 U5055 ( .A1(n5378), .A2(n5377), .ZN(n8967) );
  NAND2_X1 U5056 ( .A1(n5365), .A2(n5364), .ZN(n8972) );
  NAND2_X1 U5057 ( .A1(n7569), .A2(n7568), .ZN(n7979) );
  NOR2_X1 U5058 ( .A1(n7394), .A2(n7393), .ZN(n4742) );
  NAND2_X1 U5059 ( .A1(n7557), .A2(n7556), .ZN(n9759) );
  NAND2_X1 U5060 ( .A1(n5344), .A2(n5343), .ZN(n10193) );
  OAI21_X2 U5061 ( .B1(n7378), .B2(n7368), .A(n8846), .ZN(n8849) );
  NAND2_X1 U5062 ( .A1(n7279), .A2(n7278), .ZN(n9765) );
  NAND2_X1 U5063 ( .A1(n5327), .A2(n5326), .ZN(n7730) );
  NAND2_X1 U5064 ( .A1(n7188), .A2(n7187), .ZN(n7492) );
  NOR2_X1 U5065 ( .A1(n4795), .A2(n6013), .ZN(n4794) );
  NAND2_X1 U5066 ( .A1(n8472), .A2(n4734), .ZN(n7143) );
  NAND2_X1 U5067 ( .A1(n5285), .A2(n5284), .ZN(n7598) );
  NAND2_X1 U5068 ( .A1(n7183), .A2(n7182), .ZN(n7451) );
  AND3_X1 U5069 ( .A1(n5257), .A2(n5256), .A3(n5255), .ZN(n7468) );
  NAND2_X2 U5070 ( .A1(n6902), .A2(n10042), .ZN(n9610) );
  NAND2_X1 U5071 ( .A1(n6059), .A2(n4493), .ZN(n7051) );
  NAND2_X1 U5072 ( .A1(n4670), .A2(n4981), .ZN(n5251) );
  OR2_X1 U5073 ( .A1(n6191), .A2(n5219), .ZN(n5196) );
  AND2_X2 U5074 ( .A1(n8307), .A2(n6626), .ZN(n8324) );
  AND3_X2 U5075 ( .A1(n4642), .A2(n5180), .A3(n5181), .ZN(n7004) );
  NAND2_X1 U5076 ( .A1(n5855), .A2(n5762), .ZN(n5864) );
  AND2_X1 U5077 ( .A1(n4623), .A2(n4622), .ZN(n6807) );
  NAND2_X1 U5078 ( .A1(n10145), .A2(n5861), .ZN(n8367) );
  NAND4_X1 U5079 ( .A1(n5216), .A2(n5215), .A3(n5214), .A4(n5213), .ZN(n8568)
         );
  INV_X2 U5080 ( .A(n5219), .ZN(n5623) );
  NAND4_X1 U5081 ( .A1(n5175), .A2(n5174), .A3(n5173), .A4(n5172), .ZN(n8566)
         );
  AND4_X1 U5082 ( .A1(n6001), .A2(n6000), .A3(n5999), .A4(n5998), .ZN(n6966)
         );
  AND4_X1 U5083 ( .A1(n6021), .A2(n6020), .A3(n6019), .A4(n6018), .ZN(n7027)
         );
  CLKBUF_X2 U5084 ( .A(n5973), .Z(n4400) );
  OR2_X1 U5085 ( .A1(n6831), .A2(n4475), .ZN(n4623) );
  AND4_X1 U5086 ( .A1(n6057), .A2(n6056), .A3(n6055), .A4(n6054), .ZN(n7064)
         );
  OR2_X1 U5087 ( .A1(n5625), .A2(n6190), .ZN(n4640) );
  AND4_X1 U5088 ( .A1(n6036), .A2(n6035), .A3(n6034), .A4(n6033), .ZN(n7021)
         );
  NAND2_X1 U5089 ( .A1(n6998), .A2(n6980), .ZN(n5863) );
  NAND2_X2 U5090 ( .A1(n5105), .A2(n5104), .ZN(n5628) );
  INV_X2 U5091 ( .A(n6003), .ZN(n9151) );
  INV_X1 U5092 ( .A(n8333), .ZN(n5995) );
  AND2_X1 U5093 ( .A1(n5948), .A2(n7142), .ZN(n6625) );
  AND2_X1 U5094 ( .A1(n4855), .A2(n4668), .ZN(n4667) );
  AOI21_X1 U5095 ( .B1(n4696), .B2(n4694), .A(n4693), .ZN(n4692) );
  NAND2_X1 U5096 ( .A1(n5128), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5640) );
  AND2_X1 U5097 ( .A1(n4619), .A2(n4616), .ZN(n5100) );
  INV_X1 U5098 ( .A(n4426), .ZN(n4619) );
  OR2_X1 U5099 ( .A1(n5935), .A2(n6320), .ZN(n5932) );
  MUX2_X1 U5100 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5934), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5936) );
  XNOR2_X1 U5101 ( .A(n4973), .B(SI_4_), .ZN(n5164) );
  XNOR2_X1 U5102 ( .A(n4979), .B(SI_6_), .ZN(n5193) );
  XNOR2_X1 U5103 ( .A(n4976), .B(SI_5_), .ZN(n5148) );
  INV_X2 U5104 ( .A(n9000), .ZN(n8438) );
  AND3_X1 U5105 ( .A1(n4804), .A2(n4440), .A3(n4730), .ZN(n5803) );
  AND3_X1 U5106 ( .A1(n4396), .A2(n4950), .A3(n4447), .ZN(n4804) );
  NAND2_X1 U5107 ( .A1(n4457), .A2(n4802), .ZN(n4945) );
  NOR2_X1 U5108 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(n5129), .ZN(n5130) );
  NOR2_X1 U5109 ( .A1(n4896), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n4760) );
  NAND4_X1 U5110 ( .A1(n5190), .A2(n5254), .A3(n4746), .A4(n4745), .ZN(n5072)
         );
  OR2_X1 U5111 ( .A1(n4403), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4410) );
  INV_X1 U5112 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5769) );
  INV_X1 U5113 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5791) );
  INV_X1 U5114 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5768) );
  INV_X1 U5115 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5770) );
  INV_X1 U5116 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6038) );
  INV_X1 U5117 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6236) );
  INV_X1 U5118 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6680) );
  INV_X1 U5119 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6232) );
  INV_X1 U5120 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6908) );
  NOR2_X1 U5121 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5773) );
  INV_X1 U5122 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5771) );
  NOR2_X1 U5123 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5071) );
  INV_X2 U5124 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U5125 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5254) );
  INV_X1 U5126 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4745) );
  INV_X1 U5127 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4746) );
  AOI211_X1 U5128 ( .C1(n9681), .C2(n9884), .A(n8433), .B(n8432), .ZN(n8434)
         );
  OAI21_X2 U5129 ( .B1(n8817), .B2(n5711), .A(n5710), .ZN(n8774) );
  OAI21_X2 U5130 ( .B1(n7526), .B2(n5816), .A(n5815), .ZN(n7597) );
  NOR2_X2 U5131 ( .A1(n7535), .A2(n7412), .ZN(n7411) );
  XNOR2_X2 U5132 ( .A(n4627), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9803) );
  NAND2_X1 U5133 ( .A1(n5210), .A2(n6179), .ZN(n5219) );
  XNOR2_X2 U5134 ( .A(n5932), .B(n9790), .ZN(n5938) );
  NAND2_X1 U5135 ( .A1(n5580), .A2(n5579), .ZN(n5600) );
  NAND2_X1 U5136 ( .A1(n5576), .A2(n5575), .ZN(n5580) );
  INV_X1 U5137 ( .A(n8356), .ZN(n4518) );
  INV_X1 U5138 ( .A(n8357), .ZN(n4519) );
  OR2_X1 U5139 ( .A1(n4882), .A2(n5708), .ZN(n4881) );
  NAND2_X1 U5140 ( .A1(n9353), .A2(n9369), .ZN(n4579) );
  NAND2_X1 U5141 ( .A1(n7531), .A2(n5686), .ZN(n4892) );
  INV_X1 U5142 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5124) );
  NOR2_X1 U5143 ( .A1(n4813), .A2(n4541), .ZN(n4540) );
  INV_X1 U5144 ( .A(n4543), .ZN(n4541) );
  NAND2_X1 U5145 ( .A1(n4540), .A2(n4546), .ZN(n4538) );
  NAND2_X1 U5146 ( .A1(n4992), .A2(n4991), .ZN(n4995) );
  INV_X1 U5147 ( .A(n5633), .ZN(n5609) );
  NAND2_X1 U5148 ( .A1(n5075), .A2(n4897), .ZN(n4896) );
  INV_X1 U5149 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n4897) );
  OR2_X1 U5150 ( .A1(n8041), .A2(n8555), .ZN(n5645) );
  OR2_X1 U5151 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4403) );
  INV_X1 U5152 ( .A(n8235), .ZN(n4552) );
  AND2_X1 U5153 ( .A1(n9608), .A2(n8399), .ZN(n9264) );
  AOI21_X1 U5154 ( .B1(n4932), .B2(n8394), .A(n4459), .ZN(n4930) );
  INV_X1 U5155 ( .A(n4932), .ZN(n4931) );
  OR2_X1 U5156 ( .A1(n9750), .A2(n8131), .ZN(n9323) );
  INV_X1 U5157 ( .A(n9292), .ZN(n4723) );
  NAND2_X1 U5158 ( .A1(n4682), .A2(n4681), .ZN(n5391) );
  AOI21_X1 U5159 ( .B1(n4683), .B2(n4686), .A(n4451), .ZN(n4681) );
  INV_X1 U5160 ( .A(n4661), .ZN(n4660) );
  OAI21_X1 U5161 ( .B1(n4951), .B2(n4662), .A(n4946), .ZN(n4661) );
  NAND2_X1 U5162 ( .A1(n5194), .A2(n5193), .ZN(n4670) );
  NAND2_X1 U5163 ( .A1(n7857), .A2(n7856), .ZN(n7894) );
  NOR2_X1 U5164 ( .A1(n8542), .A2(n4754), .ZN(n4753) );
  INV_X1 U5165 ( .A(n4751), .ZN(n4750) );
  OAI21_X1 U5166 ( .B1(n8542), .B2(n4752), .A(n8372), .ZN(n4751) );
  NAND2_X1 U5167 ( .A1(n8492), .A2(n8496), .ZN(n4752) );
  AND2_X1 U5168 ( .A1(n4735), .A2(n4734), .ZN(n8473) );
  NAND2_X1 U5169 ( .A1(n4529), .A2(n4736), .ZN(n4735) );
  INV_X1 U5170 ( .A(n5873), .ZN(n4736) );
  INV_X1 U5171 ( .A(n5874), .ZN(n4529) );
  INV_X1 U5172 ( .A(n7395), .ZN(n4744) );
  NAND2_X1 U5173 ( .A1(n7623), .A2(n4742), .ZN(n4741) );
  OR2_X1 U5174 ( .A1(n8508), .A2(n8510), .ZN(n8359) );
  NAND2_X1 U5175 ( .A1(n8449), .A2(n8358), .ZN(n8360) );
  INV_X1 U5176 ( .A(n5241), .ZN(n5629) );
  INV_X1 U5177 ( .A(n5628), .ZN(n5603) );
  NAND2_X1 U5178 ( .A1(n7221), .A2(n7222), .ZN(n7326) );
  NOR2_X1 U5179 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4878) );
  AND2_X1 U5180 ( .A1(n7869), .A2(n5702), .ZN(n4893) );
  INV_X1 U5181 ( .A(n4397), .ZN(n5459) );
  INV_X1 U5182 ( .A(n5210), .ZN(n6592) );
  NAND2_X1 U5183 ( .A1(n7432), .A2(n5679), .ZN(n7005) );
  OR2_X1 U5184 ( .A1(n10139), .A2(n5835), .ZN(n7150) );
  OR2_X1 U5185 ( .A1(n10045), .A2(n8298), .ZN(n5953) );
  NAND2_X1 U5186 ( .A1(n4818), .A2(n4558), .ZN(n4557) );
  INV_X1 U5187 ( .A(n7457), .ZN(n4558) );
  OAI21_X1 U5188 ( .B1(n9528), .B2(n8420), .A(n9365), .ZN(n4733) );
  NOR2_X1 U5189 ( .A1(n8400), .A2(n4938), .ZN(n4937) );
  INV_X1 U5190 ( .A(n8397), .ZN(n4938) );
  OR2_X1 U5191 ( .A1(n9181), .A2(n8020), .ZN(n8017) );
  NAND2_X1 U5192 ( .A1(n4499), .A2(n4703), .ZN(n7751) );
  AOI21_X1 U5193 ( .B1(n4706), .B2(n4705), .A(n4704), .ZN(n4703) );
  INV_X1 U5194 ( .A(n4708), .ZN(n4705) );
  NAND2_X1 U5195 ( .A1(n9863), .A2(n9214), .ZN(n7578) );
  NAND2_X1 U5196 ( .A1(n8410), .A2(n8409), .ZN(n9682) );
  NAND2_X1 U5197 ( .A1(n6068), .A2(n4820), .ZN(n6093) );
  NOR2_X1 U5198 ( .A1(n7646), .A2(n7403), .ZN(n4820) );
  NOR2_X1 U5199 ( .A1(n6833), .A2(n6832), .ZN(n6831) );
  OAI21_X1 U5200 ( .B1(n8073), .B2(n10122), .A(n4632), .ZN(n4631) );
  AOI21_X1 U5201 ( .B1(n8074), .B2(n10119), .A(n9815), .ZN(n4632) );
  INV_X1 U5202 ( .A(n9686), .ZN(n4901) );
  OR2_X1 U5203 ( .A1(n4609), .A2(n5352), .ZN(n4605) );
  INV_X1 U5204 ( .A(n5700), .ZN(n4608) );
  AND2_X1 U5205 ( .A1(n5663), .A2(n5637), .ZN(n4610) );
  NAND2_X1 U5206 ( .A1(n4585), .A2(n9349), .ZN(n9359) );
  OAI21_X1 U5207 ( .B1(n5540), .B2(n5294), .A(n5539), .ZN(n4600) );
  AND2_X1 U5208 ( .A1(n6182), .A2(n6190), .ZN(n4641) );
  NAND2_X1 U5209 ( .A1(n4816), .A2(n9086), .ZN(n4814) );
  INV_X1 U5210 ( .A(n9369), .ZN(n4578) );
  OAI21_X1 U5211 ( .B1(n4579), .B2(n8404), .A(n4577), .ZN(n4576) );
  INV_X1 U5212 ( .A(n9368), .ZN(n4577) );
  INV_X1 U5213 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4592) );
  AND2_X1 U5214 ( .A1(n4800), .A2(n8147), .ZN(n4799) );
  NAND2_X1 U5215 ( .A1(n9068), .A2(n4801), .ZN(n4800) );
  OAI21_X1 U5216 ( .B1(n5600), .B2(n5599), .A(n5598), .ZN(n5617) );
  NAND2_X1 U5217 ( .A1(n4986), .A2(n4985), .ZN(n4989) );
  NAND2_X1 U5218 ( .A1(n4597), .A2(n4595), .ZN(n5591) );
  NOR2_X1 U5219 ( .A1(n4596), .A2(n5731), .ZN(n4595) );
  INV_X1 U5220 ( .A(n5574), .ZN(n4596) );
  NAND2_X1 U5221 ( .A1(n4414), .A2(n4827), .ZN(n4649) );
  NAND2_X1 U5222 ( .A1(n4891), .A2(n8645), .ZN(n4825) );
  NAND2_X1 U5223 ( .A1(n5093), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5463) );
  OR2_X1 U5224 ( .A1(n8953), .A2(n8820), .ZN(n8631) );
  INV_X1 U5225 ( .A(n4852), .ZN(n4851) );
  AND2_X1 U5226 ( .A1(n8816), .A2(n8805), .ZN(n5711) );
  INV_X1 U5227 ( .A(n7982), .ZN(n4858) );
  OR2_X1 U5228 ( .A1(n5305), .A2(n5304), .ZN(n5329) );
  NAND2_X1 U5229 ( .A1(n4491), .A2(n4892), .ZN(n5825) );
  AND2_X1 U5230 ( .A1(n4760), .A2(n5124), .ZN(n4759) );
  INV_X1 U5231 ( .A(n5146), .ZN(n4879) );
  OAI21_X1 U5232 ( .B1(n4535), .B2(n6047), .A(n6117), .ZN(n4534) );
  NAND2_X1 U5233 ( .A1(n6050), .A2(n4536), .ZN(n4535) );
  INV_X1 U5234 ( .A(n6118), .ZN(n4536) );
  INV_X1 U5235 ( .A(n8167), .ZN(n4544) );
  NAND2_X1 U5236 ( .A1(n4922), .A2(n4924), .ZN(n4919) );
  NOR2_X1 U5237 ( .A1(n9423), .A2(n4921), .ZN(n4920) );
  INV_X1 U5238 ( .A(n4922), .ZN(n4921) );
  NAND2_X1 U5239 ( .A1(n8405), .A2(n9568), .ZN(n9422) );
  INV_X1 U5240 ( .A(n9216), .ZN(n4709) );
  INV_X1 U5241 ( .A(n4914), .ZN(n4913) );
  OAI21_X1 U5242 ( .B1(n7552), .B2(n4915), .A(n7566), .ZN(n4914) );
  INV_X1 U5243 ( .A(n7554), .ZN(n4915) );
  OR2_X1 U5244 ( .A1(n9880), .A2(n9759), .ZN(n7589) );
  NAND2_X1 U5245 ( .A1(n7291), .A2(n4776), .ZN(n4775) );
  NOR2_X1 U5246 ( .A1(n7492), .A2(n7451), .ZN(n4776) );
  NAND2_X1 U5247 ( .A1(n7184), .A2(n4942), .ZN(n4941) );
  INV_X1 U5248 ( .A(n7178), .ZN(n4942) );
  INV_X1 U5249 ( .A(n9171), .ZN(n4943) );
  XNOR2_X1 U5250 ( .A(n4728), .B(n4400), .ZN(n4571) );
  XNOR2_X1 U5251 ( .A(n5617), .B(n5616), .ZN(n5614) );
  INV_X1 U5252 ( .A(n4945), .ZN(n4944) );
  NOR2_X1 U5253 ( .A1(n5111), .A2(n4699), .ZN(n4698) );
  INV_X1 U5254 ( .A(n5061), .ZN(n4699) );
  AOI21_X1 U5255 ( .B1(n4698), .B2(n5062), .A(n4697), .ZN(n4696) );
  INV_X1 U5256 ( .A(n5066), .ZN(n4697) );
  INV_X1 U5257 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5785) );
  NOR2_X1 U5258 ( .A1(n5456), .A2(n4678), .ZN(n4677) );
  INV_X1 U5259 ( .A(n5036), .ZN(n4678) );
  NAND2_X1 U5260 ( .A1(n5439), .A2(n5034), .ZN(n4679) );
  NAND2_X1 U5261 ( .A1(n5021), .A2(n5020), .ZN(n5390) );
  OR2_X1 U5262 ( .A1(n4685), .A2(n5012), .ZN(n4684) );
  INV_X1 U5263 ( .A(n5356), .ZN(n4685) );
  NAND2_X1 U5264 ( .A1(n4687), .A2(n5356), .ZN(n4686) );
  INV_X1 U5265 ( .A(n5340), .ZN(n4687) );
  NAND2_X1 U5266 ( .A1(n4997), .A2(n4996), .ZN(n5320) );
  XNOR2_X1 U5267 ( .A(n5001), .B(SI_11_), .ZN(n5322) );
  INV_X1 U5268 ( .A(n4995), .ZN(n4662) );
  AND2_X1 U5269 ( .A1(n4995), .A2(n4994), .ZN(n4951) );
  AND2_X1 U5270 ( .A1(n7950), .A2(n7942), .ZN(n4758) );
  NAND2_X1 U5271 ( .A1(n7938), .A2(n7937), .ZN(n7943) );
  AND2_X1 U5272 ( .A1(n5741), .A2(n6980), .ZN(n5861) );
  AND2_X1 U5273 ( .A1(n8092), .A2(n8087), .ZN(n4757) );
  INV_X1 U5274 ( .A(n7671), .ZN(n4738) );
  INV_X1 U5275 ( .A(n4740), .ZN(n4522) );
  OR2_X1 U5276 ( .A1(n5504), .A2(n5095), .ZN(n5505) );
  INV_X1 U5277 ( .A(n4758), .ZN(n4516) );
  AOI21_X1 U5278 ( .B1(n4758), .B2(n4515), .A(n4514), .ZN(n4513) );
  INV_X1 U5279 ( .A(n7937), .ZN(n4515) );
  INV_X1 U5280 ( .A(n8077), .ZN(n4514) );
  AND2_X1 U5281 ( .A1(n8082), .A2(n8081), .ZN(n8528) );
  OR2_X1 U5282 ( .A1(n7130), .A2(n7127), .ZN(n4528) );
  NAND2_X1 U5283 ( .A1(n7894), .A2(n7893), .ZN(n7930) );
  INV_X1 U5284 ( .A(n5733), .ZN(n5735) );
  AND4_X1 U5285 ( .A1(n5486), .A2(n5485), .A3(n5484), .A4(n5483), .ZN(n8487)
         );
  NAND2_X1 U5286 ( .A1(n7327), .A2(n7328), .ZN(n4633) );
  NOR3_X1 U5287 ( .A1(n8699), .A2(n4649), .A3(n8623), .ZN(n8622) );
  NAND2_X1 U5288 ( .A1(n5583), .A2(n5582), .ZN(n8041) );
  AND2_X1 U5289 ( .A1(n5645), .A2(n5732), .ZN(n8647) );
  AND2_X1 U5290 ( .A1(n5122), .A2(n5121), .ZN(n8696) );
  OAI21_X1 U5291 ( .B1(n8724), .B2(n5723), .A(n5722), .ZN(n8713) );
  OR2_X1 U5292 ( .A1(n8744), .A2(n8763), .ZN(n4947) );
  NOR2_X1 U5293 ( .A1(n8725), .A2(n4845), .ZN(n4844) );
  INV_X1 U5294 ( .A(n4947), .ZN(n4845) );
  INV_X1 U5295 ( .A(n8728), .ZN(n8763) );
  OR2_X1 U5296 ( .A1(n4646), .A2(n8636), .ZN(n4948) );
  OR2_X1 U5297 ( .A1(n8942), .A2(n8822), .ZN(n8635) );
  NAND2_X1 U5298 ( .A1(n8828), .A2(n4853), .ZN(n4852) );
  INV_X1 U5299 ( .A(n4854), .ZN(n4853) );
  NOR2_X1 U5300 ( .A1(n8856), .A2(n8855), .ZN(n8858) );
  NOR2_X1 U5301 ( .A1(n8967), .A2(n8556), .ZN(n4833) );
  AND4_X1 U5302 ( .A1(n5403), .A2(n5402), .A3(n5401), .A4(n5400), .ZN(n8854)
         );
  OR2_X1 U5303 ( .A1(n7685), .A2(n7684), .ZN(n4839) );
  NAND2_X1 U5304 ( .A1(n7681), .A2(n7686), .ZN(n7682) );
  AND2_X1 U5305 ( .A1(n5663), .A2(n5700), .ZN(n7684) );
  INV_X1 U5306 ( .A(n5696), .ZN(n4864) );
  OR2_X1 U5307 ( .A1(n6591), .A2(n5827), .ZN(n8851) );
  INV_X1 U5308 ( .A(n8819), .ZN(n8853) );
  AND3_X1 U5309 ( .A1(n5679), .A2(n5654), .A3(n5656), .ZN(n4870) );
  NAND2_X1 U5310 ( .A1(n5679), .A2(n5654), .ZN(n7425) );
  AND2_X1 U5311 ( .A1(n6708), .A2(n5827), .ZN(n8819) );
  NAND2_X1 U5312 ( .A1(n8303), .A2(n5623), .ZN(n5560) );
  AND2_X1 U5313 ( .A1(n10145), .A2(n5741), .ZN(n10195) );
  INV_X1 U5314 ( .A(n10186), .ZN(n10194) );
  OR2_X1 U5315 ( .A1(n4397), .A2(n6195), .ZN(n4642) );
  AND2_X1 U5316 ( .A1(n8108), .A2(n7160), .ZN(n10145) );
  AND2_X1 U5317 ( .A1(n5836), .A2(n5834), .ZN(n10131) );
  OR2_X1 U5318 ( .A1(n5837), .A2(n5833), .ZN(n5834) );
  OAI22_X1 U5319 ( .A1(n6952), .A2(n8297), .B1(n6990), .B2(n8298), .ZN(n5990)
         );
  INV_X1 U5320 ( .A(n6688), .ZN(n5976) );
  NAND2_X1 U5321 ( .A1(n9132), .A2(n9134), .ZN(n9055) );
  OR2_X1 U5322 ( .A1(n4794), .A2(n4417), .ZN(n4793) );
  NAND2_X1 U5323 ( .A1(n8138), .A2(n9055), .ZN(n9052) );
  NAND2_X1 U5324 ( .A1(n8236), .A2(n8235), .ZN(n9015) );
  NAND2_X1 U5325 ( .A1(n4547), .A2(n4552), .ZN(n4554) );
  INV_X1 U5326 ( .A(n8236), .ZN(n4547) );
  NOR2_X1 U5327 ( .A1(n4552), .A2(n9017), .ZN(n4551) );
  AND2_X1 U5328 ( .A1(n9078), .A2(n4549), .ZN(n4548) );
  OR2_X1 U5329 ( .A1(n8235), .A2(n4550), .ZN(n4549) );
  INV_X1 U5330 ( .A(n7478), .ZN(n4819) );
  NAND2_X1 U5331 ( .A1(n7456), .A2(n7457), .ZN(n7479) );
  NAND2_X1 U5332 ( .A1(n9442), .A2(n9499), .ZN(n6624) );
  AND2_X1 U5333 ( .A1(n8201), .A2(n8200), .ZN(n8395) );
  AND4_X1 U5334 ( .A1(n7287), .A2(n7286), .A3(n7285), .A4(n7284), .ZN(n7804)
         );
  XNOR2_X1 U5335 ( .A(n6251), .B(n5939), .ZN(n6253) );
  AND2_X1 U5336 ( .A1(n5768), .A2(n4562), .ZN(n4910) );
  NOR2_X1 U5337 ( .A1(n6773), .A2(n4472), .ZN(n6774) );
  NOR2_X1 U5338 ( .A1(n6774), .A2(n6775), .ZN(n6883) );
  NOR2_X1 U5339 ( .A1(n9942), .A2(n4780), .ZN(n4779) );
  INV_X1 U5340 ( .A(n9465), .ZN(n4780) );
  NOR2_X1 U5341 ( .A1(n4779), .A2(n4778), .ZN(n9957) );
  INV_X1 U5342 ( .A(n9960), .ZN(n4778) );
  OAI21_X1 U5343 ( .B1(n9983), .B2(n4782), .A(n4781), .ZN(n9992) );
  NAND2_X1 U5344 ( .A1(n4785), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4782) );
  NAND2_X1 U5345 ( .A1(n9469), .A2(n4785), .ZN(n4781) );
  INV_X1 U5346 ( .A(n9993), .ZN(n4785) );
  OR2_X1 U5347 ( .A1(n9983), .A2(n7767), .ZN(n4784) );
  NAND2_X1 U5348 ( .A1(n4935), .A2(n4934), .ZN(n8402) );
  NOR2_X1 U5349 ( .A1(n4936), .A2(n4404), .ZN(n4934) );
  AND4_X1 U5350 ( .A1(n8218), .A2(n8217), .A3(n8216), .A4(n8215), .ZN(n9600)
         );
  OR2_X1 U5351 ( .A1(n9717), .A2(n9634), .ZN(n8397) );
  OR2_X1 U5352 ( .A1(n9264), .A2(n9160), .ZN(n9595) );
  AND2_X1 U5353 ( .A1(n4713), .A2(n9210), .ZN(n9618) );
  AOI21_X1 U5354 ( .B1(n9625), .B2(n9624), .A(n8396), .ZN(n9612) );
  AND2_X1 U5355 ( .A1(n9723), .A2(n9649), .ZN(n8396) );
  NAND2_X1 U5356 ( .A1(n9632), .A2(n9633), .ZN(n9631) );
  AOI21_X1 U5357 ( .B1(n4933), .B2(n8392), .A(n4458), .ZN(n4932) );
  AND2_X1 U5358 ( .A1(n9344), .A2(n9332), .ZN(n9647) );
  AND2_X1 U5359 ( .A1(n9105), .A2(n9665), .ZN(n8392) );
  NOR2_X1 U5360 ( .A1(n4727), .A2(n4726), .ZN(n4725) );
  INV_X1 U5361 ( .A(n9319), .ZN(n4726) );
  OAI21_X1 U5362 ( .B1(n7747), .B2(n7746), .A(n7745), .ZN(n7828) );
  NAND2_X1 U5363 ( .A1(n7753), .A2(n7752), .ZN(n7840) );
  INV_X1 U5364 ( .A(n7754), .ZN(n7753) );
  INV_X1 U5365 ( .A(n9178), .ZN(n4707) );
  NAND2_X1 U5366 ( .A1(n7578), .A2(n4708), .ZN(n4702) );
  AOI21_X1 U5367 ( .B1(n4718), .B2(n4722), .A(n4717), .ZN(n4716) );
  INV_X1 U5368 ( .A(n9162), .ZN(n4717) );
  NAND2_X1 U5369 ( .A1(n7553), .A2(n7552), .ZN(n9876) );
  NAND2_X1 U5370 ( .A1(n9170), .A2(n7079), .ZN(n7080) );
  NAND2_X1 U5371 ( .A1(n7086), .A2(n4427), .ZN(n7179) );
  NAND2_X1 U5372 ( .A1(n4899), .A2(n4898), .ZN(n7069) );
  AND2_X1 U5373 ( .A1(n4435), .A2(n7028), .ZN(n4898) );
  XNOR2_X1 U5374 ( .A(n5778), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U5375 ( .A1(n5792), .A2(n5791), .ZN(n5794) );
  NAND2_X1 U5376 ( .A1(n4561), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U5377 ( .A1(n5149), .A2(n5148), .ZN(n4490) );
  NAND2_X1 U5378 ( .A1(n8449), .A2(n8448), .ZN(n8451) );
  NAND2_X1 U5379 ( .A1(n8451), .A2(n8450), .ZN(n8507) );
  AOI21_X1 U5380 ( .B1(n8497), .B2(n4476), .A(n4748), .ZN(n8387) );
  OAI21_X1 U5381 ( .B1(n4750), .B2(n4749), .A(n4480), .ZN(n4748) );
  NAND2_X1 U5382 ( .A1(n5210), .A2(n4413), .ZN(n4638) );
  AND4_X1 U5383 ( .A1(n5372), .A2(n5371), .A3(n5370), .A4(n5369), .ZN(n7883)
         );
  NAND2_X1 U5384 ( .A1(n5411), .A2(n5410), .ZN(n8956) );
  INV_X1 U5385 ( .A(n6808), .ZN(n4622) );
  NAND2_X1 U5386 ( .A1(n8616), .A2(n8057), .ZN(n8058) );
  OAI21_X1 U5387 ( .B1(n8588), .B2(n4507), .A(n8076), .ZN(n4629) );
  OR2_X1 U5388 ( .A1(n4410), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n4415) );
  OAI21_X1 U5389 ( .B1(n7964), .B2(n7963), .A(n7962), .ZN(n7966) );
  OAI21_X1 U5390 ( .B1(n4810), .B2(n4807), .A(n4805), .ZN(n8348) );
  AND2_X1 U5391 ( .A1(n4806), .A2(n8302), .ZN(n4805) );
  OR2_X1 U5392 ( .A1(n9005), .A2(n8328), .ZN(n8302) );
  OR2_X1 U5393 ( .A1(n4808), .A2(n4807), .ZN(n4806) );
  AND2_X1 U5394 ( .A1(n6104), .A2(n6102), .ZN(n9139) );
  NAND2_X1 U5395 ( .A1(n9433), .A2(n7142), .ZN(n9434) );
  INV_X1 U5396 ( .A(n8395), .ZN(n9649) );
  OAI22_X1 U5397 ( .A1(n8429), .A2(n9601), .B1(n8431), .B2(n8430), .ZN(n4731)
         );
  XNOR2_X1 U5398 ( .A(n4733), .B(n4909), .ZN(n4732) );
  NAND2_X1 U5399 ( .A1(n4497), .A2(n4496), .ZN(n4495) );
  XNOR2_X1 U5400 ( .A(n9528), .B(n9527), .ZN(n4498) );
  NAND2_X1 U5401 ( .A1(n9529), .A2(n9867), .ZN(n4496) );
  NOR2_X1 U5402 ( .A1(n9822), .A2(n4906), .ZN(n4905) );
  NAND2_X1 U5403 ( .A1(n9187), .A2(n4471), .ZN(n4904) );
  AND2_X1 U5404 ( .A1(n7405), .A2(n5655), .ZN(n5170) );
  NAND2_X1 U5405 ( .A1(n9316), .A2(n4566), .ZN(n4567) );
  NOR2_X1 U5406 ( .A1(n9308), .A2(n9161), .ZN(n4566) );
  AND2_X1 U5407 ( .A1(n4607), .A2(n4605), .ZN(n4603) );
  AND2_X1 U5408 ( .A1(n4462), .A2(n4604), .ZN(n4602) );
  OR2_X1 U5409 ( .A1(n5699), .A2(n4609), .ZN(n4604) );
  NAND2_X1 U5410 ( .A1(n4460), .A2(n4610), .ZN(n4606) );
  NOR2_X1 U5411 ( .A1(n9209), .A2(n9373), .ZN(n4588) );
  NAND2_X1 U5412 ( .A1(n9164), .A2(n4477), .ZN(n9169) );
  NOR2_X1 U5413 ( .A1(n7404), .A2(n5683), .ZN(n5684) );
  INV_X1 U5414 ( .A(n8139), .ZN(n4801) );
  MUX2_X1 U5415 ( .A(n5729), .B(n5573), .S(n5637), .Z(n5574) );
  OAI21_X1 U5416 ( .B1(n5538), .B2(n5537), .A(n4599), .ZN(n4598) );
  INV_X1 U5417 ( .A(n4600), .ZN(n4599) );
  OR2_X1 U5418 ( .A1(n5219), .A2(n4434), .ZN(n4636) );
  OR2_X1 U5419 ( .A1(n4397), .A2(n4641), .ZN(n4635) );
  INV_X1 U5420 ( .A(n4576), .ZN(n4575) );
  AND2_X1 U5421 ( .A1(n4684), .A2(n5373), .ZN(n4683) );
  NAND2_X1 U5422 ( .A1(n5000), .A2(n4658), .ZN(n4657) );
  NAND2_X1 U5423 ( .A1(n4660), .A2(n4662), .ZN(n4658) );
  NOR2_X1 U5424 ( .A1(n5250), .A2(n4666), .ZN(n4665) );
  INV_X1 U5425 ( .A(n5193), .ZN(n4666) );
  NAND2_X1 U5426 ( .A1(n4982), .A2(n4669), .ZN(n4668) );
  INV_X1 U5427 ( .A(n4981), .ZN(n4669) );
  NOR2_X1 U5428 ( .A1(n5271), .A2(n4856), .ZN(n4855) );
  INV_X1 U5429 ( .A(n4984), .ZN(n4856) );
  XNOR2_X1 U5430 ( .A(n4637), .B(n5886), .ZN(n5874) );
  OR2_X1 U5431 ( .A1(n7150), .A2(n5860), .ZN(n5920) );
  NAND2_X1 U5432 ( .A1(n8649), .A2(n8647), .ZN(n4486) );
  INV_X1 U5433 ( .A(n4890), .ZN(n4888) );
  NAND2_X1 U5434 ( .A1(n8774), .A2(n5712), .ZN(n8757) );
  AND2_X1 U5435 ( .A1(n4647), .A2(n4646), .ZN(n4645) );
  NOR2_X1 U5436 ( .A1(n8946), .A2(n8953), .ZN(n4647) );
  NOR2_X1 U5437 ( .A1(n4885), .A2(n4883), .ZN(n4882) );
  INV_X1 U5438 ( .A(n5705), .ZN(n4883) );
  INV_X1 U5439 ( .A(n5706), .ZN(n4885) );
  NAND2_X1 U5440 ( .A1(n4836), .A2(n7881), .ZN(n4828) );
  NAND2_X1 U5441 ( .A1(n4862), .A2(n4860), .ZN(n7607) );
  AOI21_X1 U5442 ( .B1(n4863), .B2(n4867), .A(n4861), .ZN(n4860) );
  NAND2_X1 U5443 ( .A1(n5089), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5346) );
  INV_X1 U5444 ( .A(n7358), .ZN(n4859) );
  NAND2_X1 U5445 ( .A1(n4593), .A2(n7664), .ZN(n7405) );
  NAND2_X1 U5446 ( .A1(n5657), .A2(n7320), .ZN(n5678) );
  NAND2_X1 U5447 ( .A1(n4892), .A2(n5691), .ZN(n5823) );
  NOR2_X1 U5448 ( .A1(n7505), .A2(n7504), .ZN(n7660) );
  NAND3_X1 U5449 ( .A1(n4412), .A2(n7314), .A3(n7004), .ZN(n7505) );
  INV_X1 U5450 ( .A(n4896), .ZN(n4895) );
  INV_X1 U5451 ( .A(n9017), .ZN(n4550) );
  OAI21_X1 U5452 ( .B1(n4798), .B2(n4539), .A(n4449), .ZN(n8221) );
  INV_X1 U5453 ( .A(n4540), .ZN(n4539) );
  AOI21_X1 U5454 ( .B1(n4812), .B2(n9088), .A(n4445), .ZN(n4811) );
  NOR2_X1 U5455 ( .A1(n9957), .A2(n4777), .ZN(n9466) );
  AND2_X1 U5456 ( .A1(n9956), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4777) );
  OR2_X1 U5457 ( .A1(n9692), .A2(n4765), .ZN(n4764) );
  AND2_X1 U5458 ( .A1(n8406), .A2(n4429), .ZN(n4925) );
  OR2_X1 U5459 ( .A1(n9698), .A2(n9703), .ZN(n4765) );
  NAND2_X1 U5460 ( .A1(n4770), .A2(n9644), .ZN(n4769) );
  INV_X1 U5461 ( .A(n4771), .ZN(n4770) );
  OR2_X1 U5462 ( .A1(n9732), .A2(n9105), .ZN(n4771) );
  INV_X1 U5463 ( .A(n9322), .ZN(n4727) );
  INV_X1 U5464 ( .A(n4470), .ZN(n4704) );
  INV_X1 U5465 ( .A(n9294), .ZN(n4720) );
  AND2_X1 U5466 ( .A1(n9608), .A2(n9613), .ZN(n9602) );
  AND2_X1 U5467 ( .A1(n5785), .A2(n5931), .ZN(n4729) );
  NOR2_X1 U5468 ( .A1(n4695), .A2(n4690), .ZN(n4689) );
  INV_X1 U5469 ( .A(n5057), .ZN(n4690) );
  INV_X1 U5470 ( .A(n4696), .ZN(n4695) );
  INV_X1 U5471 ( .A(n4698), .ZN(n4694) );
  INV_X1 U5472 ( .A(n5541), .ZN(n4693) );
  AOI21_X1 U5473 ( .B1(n5438), .B2(n4677), .A(n4481), .ZN(n4675) );
  INV_X1 U5474 ( .A(n4677), .ZN(n4676) );
  AND2_X1 U5475 ( .A1(n5027), .A2(n5026), .ZN(n5407) );
  OAI21_X1 U5476 ( .B1(n4960), .B2(n4503), .A(n4502), .ZN(n4959) );
  INV_X1 U5477 ( .A(n8439), .ZN(n4749) );
  NAND2_X1 U5478 ( .A1(n5094), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5504) );
  INV_X1 U5479 ( .A(n5481), .ZN(n5094) );
  INV_X1 U5480 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5182) );
  AND2_X1 U5481 ( .A1(n5895), .A2(n7126), .ZN(n4527) );
  AOI211_X1 U5482 ( .C1(n5594), .C2(n4674), .A(n4673), .B(n5592), .ZN(n4672)
         );
  NOR2_X1 U5483 ( .A1(n8894), .A2(n5294), .ZN(n4674) );
  OAI21_X1 U5484 ( .B1(n4615), .B2(n4450), .A(n4408), .ZN(n4614) );
  NAND2_X1 U5485 ( .A1(n5241), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5204) );
  XNOR2_X1 U5486 ( .A(n9803), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n9800) );
  NOR2_X1 U5487 ( .A1(n9800), .A2(n4626), .ZN(n9799) );
  NAND2_X1 U5488 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n4626) );
  NOR2_X2 U5489 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5220) );
  AOI21_X1 U5490 ( .B1(n6935), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6934), .ZN(
        n8571) );
  NOR2_X1 U5491 ( .A1(n5324), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5342) );
  AOI21_X1 U5492 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7102), .A(n7101), .ZN(
        n7105) );
  INV_X1 U5493 ( .A(n7329), .ZN(n8052) );
  NAND2_X1 U5494 ( .A1(n5126), .A2(n5125), .ZN(n5409) );
  XNOR2_X1 U5495 ( .A(n8056), .B(n8059), .ZN(n8617) );
  NOR2_X1 U5496 ( .A1(n8597), .A2(n4620), .ZN(n8056) );
  AND2_X1 U5497 ( .A1(n8055), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4620) );
  NAND2_X1 U5498 ( .A1(n8617), .A2(n5444), .ZN(n8616) );
  OR2_X1 U5499 ( .A1(n8699), .A2(n4649), .ZN(n8655) );
  NAND2_X1 U5500 ( .A1(n5730), .A2(n5646), .ZN(n8669) );
  AND2_X1 U5501 ( .A1(n4651), .A2(n4650), .ZN(n8665) );
  AOI21_X1 U5502 ( .B1(n4411), .B2(n4826), .A(n4456), .ZN(n4823) );
  INV_X1 U5503 ( .A(n8645), .ZN(n4826) );
  AND2_X1 U5504 ( .A1(n5562), .A2(n5096), .ZN(n8544) );
  NOR2_X1 U5505 ( .A1(n8739), .A2(n8914), .ZN(n8708) );
  AND2_X1 U5506 ( .A1(n8708), .A2(n8712), .ZN(n8698) );
  NAND2_X1 U5507 ( .A1(n4872), .A2(n4488), .ZN(n8724) );
  OR2_X1 U5508 ( .A1(n8749), .A2(n8921), .ZN(n8739) );
  NAND2_X1 U5509 ( .A1(n5719), .A2(n4875), .ZN(n4871) );
  OR2_X1 U5510 ( .A1(n8751), .A2(n8926), .ZN(n8749) );
  AOI21_X1 U5511 ( .B1(n8785), .B2(n8792), .A(n8638), .ZN(n8770) );
  AND2_X1 U5512 ( .A1(n8865), .A2(n4643), .ZN(n8786) );
  NOR2_X1 U5513 ( .A1(n4644), .A2(n8936), .ZN(n4643) );
  INV_X1 U5514 ( .A(n4645), .ZN(n4644) );
  NAND2_X1 U5515 ( .A1(n8841), .A2(n5709), .ZN(n8817) );
  NAND2_X1 U5516 ( .A1(n8865), .A2(n4647), .ZN(n8812) );
  INV_X1 U5517 ( .A(n4849), .ZN(n4848) );
  OAI21_X1 U5518 ( .B1(n4852), .B2(n4850), .A(n8631), .ZN(n4849) );
  OR2_X1 U5519 ( .A1(n5429), .A2(n5092), .ZN(n5445) );
  NAND2_X1 U5520 ( .A1(n8865), .A2(n8834), .ZN(n8831) );
  AND2_X1 U5521 ( .A1(n8864), .A2(n8872), .ZN(n8865) );
  NAND2_X1 U5522 ( .A1(n4884), .A2(n5705), .ZN(n8850) );
  NAND2_X1 U5523 ( .A1(n7863), .A2(n5704), .ZN(n4884) );
  NAND2_X1 U5524 ( .A1(n5091), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5429) );
  INV_X1 U5525 ( .A(n5397), .ZN(n5091) );
  OR2_X1 U5526 ( .A1(n7876), .A2(n8967), .ZN(n4957) );
  NOR2_X1 U5527 ( .A1(n7640), .A2(n10193), .ZN(n7696) );
  NAND2_X1 U5528 ( .A1(n7411), .A2(n4652), .ZN(n7640) );
  NOR2_X1 U5529 ( .A1(n4654), .A2(n7730), .ZN(n4652) );
  NAND2_X1 U5530 ( .A1(n7411), .A2(n4653), .ZN(n8001) );
  NAND2_X1 U5531 ( .A1(n4869), .A2(n5694), .ZN(n7991) );
  NAND2_X1 U5532 ( .A1(n7364), .A2(n5693), .ZN(n4869) );
  NAND2_X1 U5533 ( .A1(n7362), .A2(n7360), .ZN(n4821) );
  NAND2_X1 U5534 ( .A1(n7411), .A2(n4409), .ZN(n7999) );
  AND2_X1 U5535 ( .A1(n7411), .A2(n10179), .ZN(n7369) );
  OR2_X1 U5536 ( .A1(n7659), .A2(n7540), .ZN(n7535) );
  AND2_X1 U5537 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5153) );
  OR2_X1 U5538 ( .A1(n8566), .A2(n7004), .ZN(n7499) );
  NAND2_X1 U5539 ( .A1(n7499), .A2(n5233), .ZN(n6999) );
  INV_X1 U5540 ( .A(n6999), .ZN(n7006) );
  INV_X1 U5541 ( .A(n7425), .ZN(n7434) );
  AND2_X1 U5542 ( .A1(n5678), .A2(n5656), .ZN(n7433) );
  INV_X1 U5543 ( .A(n8759), .ZN(n8863) );
  NAND2_X1 U5544 ( .A1(n5395), .A2(n5394), .ZN(n8962) );
  INV_X1 U5545 ( .A(n5758), .ZN(n5759) );
  OAI21_X1 U5546 ( .B1(n5134), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5751) );
  NOR2_X1 U5547 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(n4407), .ZN(n4755) );
  NOR2_X1 U5548 ( .A1(n5072), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n4876) );
  NOR2_X1 U5549 ( .A1(n5072), .A2(n5146), .ZN(n5273) );
  OAI21_X1 U5550 ( .B1(n7113), .B2(n4535), .A(n4533), .ZN(n4537) );
  INV_X1 U5551 ( .A(n4534), .ZN(n4533) );
  NAND2_X1 U5552 ( .A1(n8283), .A2(n8285), .ZN(n8286) );
  INV_X1 U5553 ( .A(n8228), .ZN(n8229) );
  NOR2_X1 U5554 ( .A1(n6158), .A2(n7460), .ZN(n7189) );
  AND2_X1 U5555 ( .A1(n7914), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8027) );
  INV_X1 U5556 ( .A(n8286), .ZN(n4807) );
  INV_X1 U5557 ( .A(n8258), .ZN(n8259) );
  INV_X1 U5558 ( .A(n8243), .ZN(n8244) );
  NAND2_X1 U5559 ( .A1(n8244), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8258) );
  INV_X1 U5560 ( .A(n6915), .ZN(n4795) );
  NAND2_X1 U5561 ( .A1(n4797), .A2(n6014), .ZN(n4796) );
  INV_X1 U5562 ( .A(n6866), .ZN(n4797) );
  NAND2_X1 U5563 ( .A1(n4798), .A2(n4545), .ZN(n4542) );
  OR2_X1 U5564 ( .A1(n7559), .A2(n7558), .ZN(n7570) );
  NOR2_X1 U5565 ( .A1(n8193), .A2(n9039), .ZN(n8213) );
  AND2_X1 U5566 ( .A1(n8159), .A2(n8158), .ZN(n9108) );
  NOR2_X1 U5567 ( .A1(n6051), .A2(n6111), .ZN(n6105) );
  NAND2_X1 U5568 ( .A1(n6031), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6051) );
  INV_X1 U5569 ( .A(n8274), .ZN(n8275) );
  AND2_X1 U5570 ( .A1(n9121), .A2(n4809), .ZN(n4808) );
  AND2_X1 U5571 ( .A1(n8124), .A2(n8120), .ZN(n4531) );
  NAND2_X1 U5572 ( .A1(n8126), .A2(n8114), .ZN(n4530) );
  OR2_X1 U5573 ( .A1(n9431), .A2(n9189), .ZN(n9191) );
  NOR2_X1 U5574 ( .A1(n6883), .A2(n4473), .ZN(n6884) );
  NAND2_X1 U5575 ( .A1(n6884), .A2(n6885), .ZN(n9464) );
  NOR2_X1 U5576 ( .A1(n10003), .A2(n4792), .ZN(n10022) );
  AND2_X1 U5577 ( .A1(n10008), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4792) );
  NOR2_X1 U5578 ( .A1(n10022), .A2(n10023), .ZN(n10021) );
  XNOR2_X1 U5579 ( .A(n4790), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9498) );
  OR2_X1 U5580 ( .A1(n10021), .A2(n4791), .ZN(n4790) );
  AND2_X1 U5581 ( .A1(n10027), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4791) );
  NAND2_X1 U5582 ( .A1(n9156), .A2(n9155), .ZN(n9513) );
  AND4_X1 U5583 ( .A1(n8318), .A2(n8317), .A3(n8316), .A4(n8315), .ZN(n8429)
         );
  AOI21_X1 U5584 ( .B1(n9541), .B2(n9423), .A(n8419), .ZN(n9528) );
  NAND2_X1 U5585 ( .A1(n9554), .A2(n9865), .ZN(n4497) );
  NAND2_X1 U5586 ( .A1(n4763), .A2(n9526), .ZN(n4762) );
  INV_X1 U5587 ( .A(n4764), .ZN(n4763) );
  INV_X1 U5588 ( .A(n4918), .ZN(n4917) );
  OAI22_X1 U5589 ( .A1(n9423), .A2(n4919), .B1(n9692), .B2(n9554), .ZN(n4918)
         );
  OAI21_X1 U5590 ( .B1(n9553), .B2(n9547), .A(n9422), .ZN(n9541) );
  NOR2_X1 U5591 ( .A1(n9583), .A2(n4764), .ZN(n9534) );
  INV_X1 U5592 ( .A(n4925), .ZN(n4924) );
  NOR2_X1 U5593 ( .A1(n9583), .A2(n4765), .ZN(n9548) );
  NAND2_X1 U5594 ( .A1(n4713), .A2(n9343), .ZN(n4710) );
  NAND2_X1 U5595 ( .A1(n4713), .A2(n4711), .ZN(n4492) );
  NOR2_X1 U5596 ( .A1(n9717), .A2(n9626), .ZN(n9613) );
  AOI21_X1 U5597 ( .B1(n4930), .B2(n4931), .A(n4446), .ZN(n4928) );
  NOR2_X1 U5598 ( .A1(n8034), .A2(n4771), .ZN(n9655) );
  AND2_X1 U5599 ( .A1(n9329), .A2(n9331), .ZN(n9664) );
  NOR2_X1 U5600 ( .A1(n8034), .A2(n9105), .ZN(n9654) );
  AND2_X1 U5601 ( .A1(n9330), .A2(n9202), .ZN(n9181) );
  OR2_X1 U5602 ( .A1(n8016), .A2(n8015), .ZN(n8020) );
  OR2_X1 U5603 ( .A1(n7911), .A2(n9745), .ZN(n8034) );
  NOR2_X1 U5604 ( .A1(n7570), .A2(n7973), .ZN(n7579) );
  NOR2_X1 U5605 ( .A1(n7766), .A2(n9754), .ZN(n7842) );
  NAND2_X1 U5606 ( .A1(n7751), .A2(n9310), .ZN(n7754) );
  AND4_X1 U5607 ( .A1(n7762), .A2(n7761), .A3(n7760), .A4(n7759), .ZN(n8131)
         );
  OR2_X1 U5608 ( .A1(n7589), .A2(n7979), .ZN(n7766) );
  AOI21_X1 U5609 ( .B1(n4913), .B2(n4915), .A(n4479), .ZN(n4911) );
  NOR2_X1 U5610 ( .A1(n9875), .A2(n4775), .ZN(n4773) );
  OR2_X1 U5611 ( .A1(n7282), .A2(n7819), .ZN(n7559) );
  NAND2_X1 U5612 ( .A1(n7200), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7282) );
  OAI21_X1 U5613 ( .B1(n7250), .B2(n4722), .A(n4718), .ZN(n7577) );
  INV_X1 U5614 ( .A(n4776), .ZN(n4774) );
  NAND2_X1 U5615 ( .A1(n4724), .A2(n9292), .ZN(n7281) );
  NAND2_X1 U5616 ( .A1(n7250), .A2(n9294), .ZN(n4724) );
  AOI21_X1 U5617 ( .B1(n7086), .B2(n4439), .A(n4940), .ZN(n7195) );
  NAND2_X1 U5618 ( .A1(n4454), .A2(n4941), .ZN(n4940) );
  NAND2_X1 U5619 ( .A1(n9235), .A2(n4714), .ZN(n4508) );
  NAND2_X1 U5620 ( .A1(n4510), .A2(n9235), .ZN(n4509) );
  INV_X1 U5621 ( .A(n9274), .ZN(n4510) );
  AND4_X1 U5622 ( .A1(n6145), .A2(n6144), .A3(n6143), .A4(n6142), .ZN(n7251)
         );
  AND2_X1 U5623 ( .A1(n7074), .A2(n10094), .ZN(n7092) );
  AOI21_X1 U5624 ( .B1(n7037), .B2(n4584), .A(n4583), .ZN(n4582) );
  INV_X1 U5625 ( .A(n7055), .ZN(n4584) );
  INV_X1 U5626 ( .A(n7057), .ZN(n4583) );
  OR2_X1 U5627 ( .A1(n7056), .A2(n9232), .ZN(n4581) );
  OR2_X1 U5628 ( .A1(n7030), .A2(n7112), .ZN(n7045) );
  NAND2_X1 U5629 ( .A1(n7056), .A2(n7055), .ZN(n7038) );
  AND2_X1 U5630 ( .A1(n9230), .A2(n7057), .ZN(n9166) );
  NOR2_X1 U5631 ( .A1(n6989), .A2(n6959), .ZN(n6972) );
  NAND2_X1 U5632 ( .A1(n6972), .A2(n10072), .ZN(n7030) );
  NAND2_X1 U5633 ( .A1(n9274), .A2(n9406), .ZN(n7056) );
  NAND2_X1 U5634 ( .A1(n4761), .A2(n6990), .ZN(n6989) );
  AND2_X1 U5635 ( .A1(n6617), .A2(n6086), .ZN(n9766) );
  OR2_X1 U5636 ( .A1(n6637), .A2(n9396), .ZN(n10101) );
  XNOR2_X1 U5637 ( .A(n5622), .B(n5621), .ZN(n9148) );
  XNOR2_X1 U5638 ( .A(n5600), .B(n5581), .ZN(n8407) );
  NAND2_X1 U5639 ( .A1(n5805), .A2(n5804), .ZN(n8427) );
  INV_X1 U5640 ( .A(n5803), .ZN(n5804) );
  MUX2_X1 U5641 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5802), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5805) );
  OAI21_X1 U5642 ( .B1(n5783), .B2(n4945), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5802) );
  NAND2_X1 U5643 ( .A1(n4691), .A2(n4696), .ZN(n5542) );
  NAND2_X1 U5644 ( .A1(n5522), .A2(n4698), .ZN(n4691) );
  NAND2_X1 U5645 ( .A1(n4803), .A2(n4802), .ZN(n5799) );
  INV_X1 U5646 ( .A(n5783), .ZN(n4803) );
  AND2_X1 U5647 ( .A1(n5057), .A2(n5056), .ZN(n5135) );
  NAND2_X1 U5648 ( .A1(n4679), .A2(n4677), .ZN(n5471) );
  NAND2_X1 U5649 ( .A1(n4679), .A2(n5036), .ZN(n5457) );
  NAND2_X1 U5650 ( .A1(n4680), .A2(n4684), .ZN(n5374) );
  OR2_X1 U5651 ( .A1(n5341), .A2(n4686), .ZN(n4680) );
  OR2_X1 U5652 ( .A1(n5341), .A2(n5340), .ZN(n5355) );
  OR3_X1 U5653 ( .A1(n6241), .A2(P1_IR_REG_10__SCAN_IN), .A3(
        P1_IR_REG_11__SCAN_IN), .ZN(n6319) );
  OAI21_X1 U5654 ( .B1(n5282), .B2(n4662), .A(n4660), .ZN(n5321) );
  INV_X1 U5655 ( .A(n4659), .ZN(n5299) );
  AOI21_X1 U5656 ( .B1(n5282), .B2(n4951), .A(n4662), .ZN(n4659) );
  NAND2_X1 U5657 ( .A1(n5251), .A2(n4982), .ZN(n4857) );
  XNOR2_X1 U5658 ( .A(n4965), .B(SI_2_), .ZN(n5217) );
  INV_X1 U5659 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4505) );
  AND2_X1 U5660 ( .A1(n7303), .A2(n5901), .ZN(n7230) );
  NAND2_X1 U5661 ( .A1(n4747), .A2(n4750), .ZN(n8440) );
  NAND2_X1 U5662 ( .A1(n8287), .A2(n5623), .ZN(n5549) );
  AND4_X1 U5663 ( .A1(n5293), .A2(n5292), .A3(n5291), .A4(n5290), .ZN(n7993)
         );
  OR2_X1 U5664 ( .A1(n5412), .A2(n5289), .ZN(n5290) );
  OR2_X1 U5665 ( .A1(n8382), .A2(n8381), .ZN(n8383) );
  AND4_X1 U5666 ( .A1(n5334), .A2(n5333), .A3(n5332), .A4(n5331), .ZN(n7992)
         );
  NAND2_X1 U5667 ( .A1(n4528), .A2(n7126), .ZN(n7163) );
  OR2_X1 U5668 ( .A1(n5926), .A2(n5925), .ZN(n8502) );
  NAND2_X1 U5669 ( .A1(n7943), .A2(n4758), .ZN(n8530) );
  NAND2_X1 U5670 ( .A1(n7943), .A2(n7942), .ZN(n7948) );
  INV_X1 U5671 ( .A(n8508), .ZN(n4517) );
  NAND2_X1 U5672 ( .A1(n5885), .A2(n5884), .ZN(n7130) );
  INV_X1 U5673 ( .A(n10146), .ZN(n7314) );
  NAND2_X1 U5674 ( .A1(n8460), .A2(n8087), .ZN(n8519) );
  AOI21_X1 U5675 ( .B1(n4737), .B2(n4522), .A(n4521), .ZN(n4520) );
  INV_X1 U5676 ( .A(n4737), .ZN(n4523) );
  INV_X1 U5677 ( .A(n7673), .ZN(n4521) );
  AND3_X1 U5678 ( .A1(n5509), .A2(n5508), .A3(n5507), .ZN(n8641) );
  AND4_X1 U5679 ( .A1(n5351), .A2(n5350), .A3(n5349), .A4(n5348), .ZN(n7683)
         );
  AND4_X1 U5680 ( .A1(n5311), .A2(n5310), .A3(n5309), .A4(n5308), .ZN(n7397)
         );
  INV_X1 U5681 ( .A(n4742), .ZN(n4739) );
  INV_X1 U5682 ( .A(n8547), .ZN(n8523) );
  NAND2_X1 U5683 ( .A1(n4513), .A2(n4516), .ZN(n4511) );
  NAND2_X1 U5684 ( .A1(n4526), .A2(n4524), .ZN(n7303) );
  NAND2_X1 U5685 ( .A1(n7130), .A2(n4527), .ZN(n4526) );
  AND2_X1 U5686 ( .A1(n5897), .A2(n4525), .ZN(n4524) );
  NAND2_X1 U5687 ( .A1(n4527), .A2(n7127), .ZN(n4525) );
  AND4_X1 U5688 ( .A1(n5385), .A2(n5384), .A3(n5383), .A4(n5382), .ZN(n7898)
         );
  AND4_X1 U5689 ( .A1(n5416), .A2(n5415), .A3(n5414), .A4(n5413), .ZN(n7952)
         );
  OR2_X1 U5690 ( .A1(n8502), .A2(n8853), .ZN(n8548) );
  OR2_X1 U5691 ( .A1(n8502), .A2(n8851), .ZN(n8547) );
  INV_X1 U5692 ( .A(n8551), .ZN(n8541) );
  INV_X1 U5693 ( .A(n8108), .ZN(n6998) );
  NOR2_X1 U5694 ( .A1(n5743), .A2(n5742), .ZN(n5744) );
  NAND2_X1 U5695 ( .A1(n5241), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5270) );
  OR2_X1 U5696 ( .A1(n5412), .A2(n5185), .ZN(n5186) );
  OR2_X1 U5697 ( .A1(n5412), .A2(n5142), .ZN(n5143) );
  NAND2_X1 U5698 ( .A1(n5241), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5214) );
  CLKBUF_X1 U5699 ( .A(n5872), .Z(n7441) );
  NAND2_X1 U5700 ( .A1(n6706), .A2(n10144), .ZN(n8567) );
  NAND2_X1 U5701 ( .A1(n10129), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4627) );
  AOI21_X1 U5702 ( .B1(n9814), .B2(P2_REG2_REG_2__SCAN_IN), .A(n9810), .ZN(
        n6821) );
  NOR2_X1 U5703 ( .A1(n6807), .A2(n4621), .ZN(n6845) );
  AND2_X1 U5704 ( .A1(n6741), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4621) );
  NOR2_X1 U5705 ( .A1(n6843), .A2(n4625), .ZN(n6857) );
  NOR2_X1 U5706 ( .A1(n6852), .A2(n6742), .ZN(n4625) );
  NOR2_X1 U5707 ( .A1(n6857), .A2(n6856), .ZN(n6855) );
  OR2_X1 U5708 ( .A1(n6855), .A2(n4624), .ZN(n6746) );
  NOR2_X1 U5709 ( .A1(n6863), .A2(n5261), .ZN(n4624) );
  AND2_X1 U5710 ( .A1(n6763), .A2(n6764), .ZN(n6934) );
  AND2_X1 U5711 ( .A1(n5074), .A2(n4760), .ZN(n5375) );
  XNOR2_X1 U5712 ( .A(n8622), .B(n8042), .ZN(n8881) );
  INV_X1 U5713 ( .A(n8041), .ZN(n8888) );
  OAI21_X1 U5714 ( .B1(n8654), .B2(n8759), .A(n8653), .ZN(n8891) );
  NAND2_X1 U5715 ( .A1(n4824), .A2(n8645), .ZN(n8677) );
  NAND2_X1 U5716 ( .A1(n5725), .A2(n5724), .ZN(n8693) );
  NAND2_X1 U5717 ( .A1(n8919), .A2(n4947), .ZN(n8720) );
  NAND2_X1 U5718 ( .A1(n8737), .A2(n8736), .ZN(n8919) );
  NOR2_X1 U5719 ( .A1(n8858), .A2(n4854), .ZN(n8829) );
  OR2_X1 U5720 ( .A1(n8858), .A2(n4852), .ZN(n8827) );
  NAND2_X1 U5721 ( .A1(n7682), .A2(n5702), .ZN(n7882) );
  NAND2_X1 U5722 ( .A1(n4839), .A2(n4837), .ZN(n7868) );
  NAND2_X1 U5723 ( .A1(n4839), .A2(n4840), .ZN(n7687) );
  NAND2_X1 U5724 ( .A1(n8846), .A2(n5917), .ZN(n8871) );
  OR2_X1 U5725 ( .A1(n10130), .A2(n7015), .ZN(n8835) );
  INV_X1 U5726 ( .A(n8871), .ZN(n8691) );
  INV_X1 U5727 ( .A(n8656), .ZN(n8876) );
  AND2_X2 U5728 ( .A1(n7019), .A2(n7155), .ZN(n10217) );
  AND2_X2 U5729 ( .A1(n7156), .A2(n7155), .ZN(n10204) );
  INV_X1 U5730 ( .A(n10138), .ZN(n10141) );
  NAND2_X1 U5731 ( .A1(n8998), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5099) );
  NAND2_X1 U5732 ( .A1(n5097), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5083) );
  NAND2_X1 U5733 ( .A1(n4619), .A2(n4618), .ZN(n5097) );
  XNOR2_X1 U5734 ( .A(n5751), .B(n5750), .ZN(n8108) );
  XNOR2_X1 U5735 ( .A(n5133), .B(n5132), .ZN(n7160) );
  NAND2_X1 U5736 ( .A1(n5641), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5643) );
  INV_X1 U5737 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6192) );
  INV_X1 U5738 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6408) );
  INV_X1 U5739 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U5740 ( .A1(n9120), .A2(n8286), .ZN(n9007) );
  INV_X1 U5741 ( .A(n4554), .ZN(n9014) );
  NAND2_X1 U5742 ( .A1(n7479), .A2(n7478), .ZN(n7702) );
  AND4_X1 U5743 ( .A1(n6110), .A2(n6109), .A3(n6108), .A4(n6107), .ZN(n7082)
         );
  NAND2_X1 U5744 ( .A1(n9077), .A2(n8253), .ZN(n9045) );
  NAND2_X1 U5745 ( .A1(n9067), .A2(n9068), .ZN(n9066) );
  NAND2_X1 U5746 ( .A1(n9052), .A2(n8139), .ZN(n9067) );
  NAND2_X1 U5747 ( .A1(n9015), .A2(n9017), .ZN(n4553) );
  NAND2_X1 U5748 ( .A1(n4796), .A2(n4794), .ZN(n6914) );
  AND4_X1 U5749 ( .A1(n7194), .A2(n7193), .A3(n7192), .A4(n7191), .ZN(n7712)
         );
  INV_X1 U5750 ( .A(n4405), .ZN(n4555) );
  NAND2_X1 U5751 ( .A1(n4405), .A2(n4818), .ZN(n4556) );
  NAND2_X1 U5752 ( .A1(n7479), .A2(n4818), .ZN(n7797) );
  NAND2_X1 U5753 ( .A1(n4810), .A2(n4808), .ZN(n9120) );
  AND2_X1 U5754 ( .A1(n6099), .A2(n6098), .ZN(n9142) );
  AND2_X1 U5755 ( .A1(n6690), .A2(n9766), .ZN(n9144) );
  NOR2_X1 U5756 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n4560) );
  INV_X1 U5757 ( .A(n8429), .ZN(n9542) );
  OR2_X1 U5758 ( .A1(n5996), .A2(n5937), .ZN(n5944) );
  OR2_X1 U5759 ( .A1(n8425), .A2(n6587), .ZN(n5945) );
  OR2_X1 U5760 ( .A1(n8332), .A2(n10043), .ZN(n5942) );
  OR2_X1 U5761 ( .A1(n8332), .A2(n5958), .ZN(n5962) );
  XNOR2_X1 U5762 ( .A(n6023), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9907) );
  OAI21_X1 U5763 ( .B1(n9919), .B2(n9920), .A(n4787), .ZN(n6283) );
  OR2_X1 U5764 ( .A1(n9918), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4787) );
  NOR2_X1 U5765 ( .A1(n6283), .A2(n6284), .ZN(n6310) );
  NOR2_X1 U5766 ( .A1(n6310), .A2(n4786), .ZN(n6312) );
  NOR2_X1 U5767 ( .A1(n6286), .A2(n7049), .ZN(n4786) );
  NAND2_X1 U5768 ( .A1(n6312), .A2(n6313), .ZN(n6670) );
  INV_X1 U5769 ( .A(n4779), .ZN(n9959) );
  INV_X1 U5770 ( .A(n4784), .ZN(n9982) );
  INV_X1 U5771 ( .A(n9469), .ZN(n4783) );
  NAND2_X1 U5772 ( .A1(n9559), .A2(n9159), .ZN(n4926) );
  AND2_X1 U5773 ( .A1(n4935), .A2(n4939), .ZN(n9573) );
  NAND2_X1 U5774 ( .A1(n8398), .A2(n8397), .ZN(n9593) );
  NAND2_X1 U5775 ( .A1(n9631), .A2(n9343), .ZN(n9619) );
  NAND2_X1 U5776 ( .A1(n4929), .A2(n4932), .ZN(n9639) );
  NAND2_X1 U5777 ( .A1(n8393), .A2(n4933), .ZN(n4929) );
  NAND2_X1 U5778 ( .A1(n7840), .A2(n9319), .ZN(n7918) );
  NAND2_X1 U5779 ( .A1(n4702), .A2(n4706), .ZN(n4955) );
  NAND2_X1 U5780 ( .A1(n7578), .A2(n9298), .ZN(n7725) );
  NAND2_X1 U5781 ( .A1(n9876), .A2(n7554), .ZN(n7720) );
  NAND2_X1 U5782 ( .A1(n7179), .A2(n7178), .ZN(n7252) );
  NAND2_X1 U5783 ( .A1(n7086), .A2(n7085), .ZN(n7088) );
  NAND2_X1 U5784 ( .A1(n4494), .A2(n9151), .ZN(n4493) );
  INV_X1 U5785 ( .A(n6191), .ZN(n4494) );
  OR2_X1 U5786 ( .A1(n10065), .A2(n6900), .ZN(n10042) );
  INV_X1 U5787 ( .A(n9660), .ZN(n9874) );
  INV_X1 U5788 ( .A(n5940), .ZN(n7923) );
  OR2_X1 U5789 ( .A1(n5803), .A2(n6320), .ZN(n5801) );
  NAND2_X1 U5790 ( .A1(n4431), .A2(n4406), .ZN(n5955) );
  INV_X1 U5791 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6174) );
  OR2_X1 U5792 ( .A1(n6041), .A2(n6040), .ZN(n6276) );
  NAND2_X1 U5793 ( .A1(n5950), .A2(n4788), .ZN(n6251) );
  AOI22_X1 U5794 ( .A1(n4455), .A2(P1_IR_REG_0__SCAN_IN), .B1(n4789), .B2(
        n6320), .ZN(n4788) );
  INV_X1 U5795 ( .A(n4623), .ZN(n6809) );
  OAI211_X1 U5796 ( .C1(n8075), .C2(n5458), .A(n4630), .B(n4628), .ZN(P2_U3264) );
  INV_X1 U5797 ( .A(n4629), .ZN(n4628) );
  NAND2_X1 U5798 ( .A1(n4631), .A2(n5458), .ZN(n4630) );
  NOR2_X1 U5799 ( .A1(n9690), .A2(n4399), .ZN(n9530) );
  OR2_X1 U5800 ( .A1(n10117), .A2(n4908), .ZN(n4907) );
  NAND2_X1 U5801 ( .A1(n4901), .A2(n4905), .ZN(n4900) );
  INV_X1 U5802 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n4908) );
  INV_X1 U5803 ( .A(n4700), .ZN(P1_U3520) );
  NOR2_X1 U5804 ( .A1(n10107), .A2(n8334), .ZN(n4701) );
  AND2_X1 U5805 ( .A1(n9709), .A2(n9567), .ZN(n4404) );
  OR2_X1 U5806 ( .A1(n7795), .A2(n7794), .ZN(n4405) );
  AND2_X1 U5807 ( .A1(n4396), .A2(n4950), .ZN(n4406) );
  INV_X1 U5808 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5274) );
  NAND2_X1 U5809 ( .A1(n5524), .A2(n5523), .ZN(n8914) );
  OR2_X1 U5810 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n4407) );
  OAI211_X1 U5811 ( .C1(n5965), .C2(n6279), .A(n5989), .B(n5988), .ZN(n6991)
         );
  NAND2_X1 U5812 ( .A1(n5693), .A2(n5694), .ZN(n7362) );
  OR2_X1 U5813 ( .A1(n5638), .A2(n5294), .ZN(n4408) );
  AND2_X1 U5814 ( .A1(n7376), .A2(n10179), .ZN(n4409) );
  AND2_X1 U5815 ( .A1(n8683), .A2(n4825), .ZN(n4411) );
  AND3_X1 U5816 ( .A1(n4466), .A2(n4635), .A3(n4636), .ZN(n4412) );
  INV_X1 U5817 ( .A(n9159), .ZN(n4923) );
  NAND3_X1 U5818 ( .A1(n5143), .A2(n4594), .A3(n4441), .ZN(n8564) );
  INV_X1 U5819 ( .A(n8564), .ZN(n4593) );
  AND2_X1 U5820 ( .A1(n5952), .A2(n4436), .ZN(n10045) );
  INV_X1 U5821 ( .A(n10045), .ZN(n4728) );
  AND2_X1 U5822 ( .A1(n4402), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4413) );
  INV_X1 U5823 ( .A(n9088), .ZN(n4816) );
  AND2_X1 U5824 ( .A1(n8188), .A2(n8187), .ZN(n9088) );
  OAI21_X1 U5825 ( .B1(n9633), .B2(n4712), .A(n9210), .ZN(n4711) );
  AND2_X1 U5826 ( .A1(n8888), .A2(n4650), .ZN(n4414) );
  NAND2_X1 U5827 ( .A1(n5644), .A2(n5637), .ZN(n4416) );
  NOR2_X1 U5828 ( .A1(n6029), .A2(n6028), .ZN(n4417) );
  NOR2_X1 U5829 ( .A1(n8914), .A2(n4846), .ZN(n4418) );
  INV_X1 U5830 ( .A(n7043), .ZN(n4580) );
  AND2_X1 U5831 ( .A1(n7796), .A2(n4557), .ZN(n4419) );
  AND2_X1 U5832 ( .A1(n7752), .A2(n4568), .ZN(n4420) );
  NAND2_X1 U5833 ( .A1(n6093), .A2(n6625), .ZN(n7710) );
  XNOR2_X1 U5834 ( .A(n5643), .B(n5642), .ZN(n5741) );
  OR2_X1 U5835 ( .A1(n7256), .A2(n4774), .ZN(n4421) );
  AND2_X1 U5836 ( .A1(n4796), .A2(n6867), .ZN(n4422) );
  NAND4_X1 U5837 ( .A1(n5202), .A2(n5201), .A3(n5200), .A4(n5199), .ZN(n5875)
         );
  OR2_X1 U5838 ( .A1(n8956), .A2(n7952), .ZN(n5706) );
  AND2_X1 U5839 ( .A1(n7703), .A2(n7704), .ZN(n4423) );
  NAND2_X1 U5840 ( .A1(n4989), .A2(n4988), .ZN(n5271) );
  NAND4_X1 U5841 ( .A1(n5945), .A2(n5944), .A3(n5943), .A4(n5942), .ZN(n5973)
         );
  NAND4_X1 U5842 ( .A1(n5963), .A2(n5962), .A3(n5961), .A4(n5960), .ZN(n6229)
         );
  INV_X1 U5843 ( .A(n8184), .ZN(n8322) );
  AND2_X1 U5844 ( .A1(n6100), .A2(n6624), .ZN(n8184) );
  NOR2_X1 U5845 ( .A1(n7686), .A2(n4838), .ZN(n4837) );
  NAND2_X1 U5846 ( .A1(n4798), .A2(n4799), .ZN(n9024) );
  INV_X1 U5847 ( .A(n4571), .ZN(n6630) );
  AND2_X1 U5848 ( .A1(n8757), .A2(n5719), .ZN(n4424) );
  AND2_X1 U5849 ( .A1(n6944), .A2(n6943), .ZN(n4425) );
  INV_X1 U5850 ( .A(n4722), .ZN(n4721) );
  OR2_X1 U5851 ( .A1(n7280), .A2(n4723), .ZN(n4722) );
  OR2_X1 U5852 ( .A1(n4894), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4426) );
  AND2_X1 U5853 ( .A1(n4943), .A2(n7085), .ZN(n4427) );
  XNOR2_X1 U5854 ( .A(n9682), .B(n9529), .ZN(n9187) );
  INV_X1 U5855 ( .A(n9187), .ZN(n4909) );
  AND2_X1 U5856 ( .A1(n8166), .A2(n4954), .ZN(n4428) );
  INV_X1 U5857 ( .A(n9406), .ZN(n4714) );
  OR2_X1 U5858 ( .A1(n9703), .A2(n8403), .ZN(n4429) );
  INV_X1 U5859 ( .A(n4867), .ZN(n4866) );
  OR2_X1 U5860 ( .A1(n5697), .A2(n4868), .ZN(n4867) );
  INV_X1 U5861 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4802) );
  AND2_X1 U5862 ( .A1(n4817), .A2(n4816), .ZN(n4430) );
  INV_X1 U5863 ( .A(n7664), .ZN(n10169) );
  AND2_X1 U5864 ( .A1(n5865), .A2(n5864), .ZN(n8365) );
  INV_X1 U5865 ( .A(n5693), .ZN(n4865) );
  INV_X1 U5866 ( .A(n5694), .ZN(n4868) );
  AND2_X1 U5867 ( .A1(n6123), .A2(n5787), .ZN(n4431) );
  AOI21_X1 U5868 ( .B1(n8679), .B2(n5589), .A(n5552), .ZN(n8697) );
  INV_X1 U5869 ( .A(n5698), .ZN(n4861) );
  NAND2_X1 U5870 ( .A1(n5427), .A2(n5426), .ZN(n8953) );
  XNOR2_X1 U5871 ( .A(n5102), .B(n5101), .ZN(n5103) );
  OR3_X1 U5872 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        n10129), .ZN(n4432) );
  NAND2_X1 U5873 ( .A1(n4542), .A2(n4543), .ZN(n9085) );
  INV_X1 U5874 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5190) );
  AND2_X1 U5875 ( .A1(n9698), .A2(n9568), .ZN(n4433) );
  NAND2_X1 U5876 ( .A1(n5530), .A2(n5721), .ZN(n8736) );
  AND2_X1 U5877 ( .A1(n6189), .A2(n6180), .ZN(n4434) );
  NOR2_X1 U5878 ( .A1(n9166), .A2(n7066), .ZN(n4435) );
  AND2_X1 U5879 ( .A1(n5951), .A2(n4572), .ZN(n4436) );
  AND2_X1 U5880 ( .A1(n4582), .A2(n4580), .ZN(n4437) );
  INV_X1 U5881 ( .A(n9343), .ZN(n4712) );
  AND2_X1 U5882 ( .A1(n5728), .A2(n5727), .ZN(n4438) );
  XNOR2_X1 U5883 ( .A(n4983), .B(SI_7_), .ZN(n5250) );
  NAND2_X1 U5884 ( .A1(n7551), .A2(n7550), .ZN(n9875) );
  NOR2_X1 U5885 ( .A1(n4423), .A2(n4819), .ZN(n4818) );
  NAND2_X2 U5886 ( .A1(n5938), .A2(n7923), .ZN(n5996) );
  INV_X1 U5887 ( .A(n4651), .ZN(n8678) );
  OR2_X1 U5888 ( .A1(n8894), .A2(n8684), .ZN(n5730) );
  AND2_X1 U5889 ( .A1(n4427), .A2(n7184), .ZN(n4439) );
  AND2_X1 U5890 ( .A1(n5703), .A2(n5404), .ZN(n7869) );
  INV_X1 U5891 ( .A(n7869), .ZN(n7881) );
  AND2_X1 U5892 ( .A1(n4944), .A2(n5800), .ZN(n4440) );
  INV_X1 U5893 ( .A(n9161), .ZN(n7752) );
  AND2_X1 U5894 ( .A1(n5145), .A2(n5144), .ZN(n4441) );
  AND2_X1 U5895 ( .A1(n4784), .A2(n4783), .ZN(n4442) );
  INV_X1 U5896 ( .A(n9309), .ZN(n4568) );
  NOR2_X1 U5897 ( .A1(n9583), .A2(n9703), .ZN(n4766) );
  AND2_X1 U5898 ( .A1(n9321), .A2(n9320), .ZN(n4443) );
  OR2_X1 U5899 ( .A1(n9085), .A2(n9086), .ZN(n4817) );
  OR2_X1 U5900 ( .A1(n7492), .A2(n7712), .ZN(n9288) );
  INV_X1 U5901 ( .A(n9288), .ZN(n4719) );
  INV_X1 U5902 ( .A(n6868), .ZN(n6014) );
  AND2_X1 U5903 ( .A1(n4511), .A2(n8528), .ZN(n4444) );
  NOR2_X1 U5904 ( .A1(n8207), .A2(n8206), .ZN(n4445) );
  NOR2_X1 U5905 ( .A1(n9644), .A2(n9032), .ZN(n4446) );
  AND4_X1 U5906 ( .A1(n5777), .A2(n5946), .A3(n5787), .A4(n5791), .ZN(n4447)
         );
  INV_X1 U5907 ( .A(n4546), .ZN(n4545) );
  NAND2_X1 U5908 ( .A1(n4428), .A2(n4799), .ZN(n4546) );
  AND3_X1 U5909 ( .A1(n5124), .A2(n4592), .A3(n5125), .ZN(n4448) );
  INV_X1 U5910 ( .A(n4840), .ZN(n4838) );
  OR2_X1 U5911 ( .A1(n10193), .A2(n8558), .ZN(n4840) );
  INV_X1 U5912 ( .A(n4654), .ZN(n4653) );
  NAND2_X1 U5913 ( .A1(n4409), .A2(n4655), .ZN(n4654) );
  INV_X1 U5914 ( .A(n4813), .ZN(n4812) );
  NAND2_X1 U5915 ( .A1(n4815), .A2(n4814), .ZN(n4813) );
  NAND2_X1 U5916 ( .A1(n5461), .A2(n5460), .ZN(n8942) );
  INV_X1 U5917 ( .A(n8942), .ZN(n4646) );
  AND2_X1 U5918 ( .A1(n4538), .A2(n4811), .ZN(n4449) );
  NAND2_X1 U5919 ( .A1(n5553), .A2(n8681), .ZN(n8694) );
  INV_X1 U5920 ( .A(n8694), .ZN(n4891) );
  INV_X1 U5921 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5946) );
  AND2_X1 U5922 ( .A1(n5737), .A2(n5612), .ZN(n4450) );
  NAND2_X1 U5923 ( .A1(n4804), .A2(n4730), .ZN(n5783) );
  INV_X1 U5924 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5073) );
  AND2_X1 U5925 ( .A1(n5016), .A2(SI_14_), .ZN(n4451) );
  NAND2_X1 U5926 ( .A1(n8972), .A2(n8557), .ZN(n4452) );
  OR2_X1 U5927 ( .A1(n6868), .A2(n4417), .ZN(n4453) );
  NAND2_X1 U5928 ( .A1(n7451), .A2(n9454), .ZN(n4454) );
  AND2_X1 U5929 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4455) );
  AND2_X1 U5930 ( .A1(n4827), .A2(n8697), .ZN(n4456) );
  AND2_X1 U5931 ( .A1(n5798), .A2(n5797), .ZN(n4457) );
  NOR2_X1 U5932 ( .A1(n9661), .A2(n9114), .ZN(n4458) );
  NOR2_X1 U5933 ( .A1(n9728), .A2(n9666), .ZN(n4459) );
  OR2_X1 U5934 ( .A1(n4861), .A2(n4608), .ZN(n4460) );
  INV_X1 U5935 ( .A(n9209), .ZN(n4713) );
  NAND2_X1 U5936 ( .A1(n8152), .A2(n8151), .ZN(n9732) );
  NAND2_X1 U5937 ( .A1(n8290), .A2(n8289), .ZN(n9692) );
  AND2_X1 U5938 ( .A1(n4926), .A2(n4429), .ZN(n4461) );
  AND2_X1 U5939 ( .A1(n7686), .A2(n4606), .ZN(n4462) );
  AND2_X1 U5940 ( .A1(n5704), .A2(n5707), .ZN(n4463) );
  NAND2_X1 U5941 ( .A1(n8273), .A2(n8272), .ZN(n9698) );
  INV_X1 U5942 ( .A(n9698), .ZN(n8405) );
  XNOR2_X1 U5943 ( .A(n5015), .B(SI_14_), .ZN(n5373) );
  AND2_X1 U5944 ( .A1(n8919), .A2(n4844), .ZN(n4464) );
  AND2_X1 U5945 ( .A1(n9316), .A2(n4420), .ZN(n4465) );
  AND2_X1 U5946 ( .A1(n5222), .A2(n5211), .ZN(n4466) );
  INV_X1 U5947 ( .A(n5712), .ZN(n4875) );
  NAND2_X1 U5948 ( .A1(n4707), .A2(n9216), .ZN(n4706) );
  AND2_X1 U5949 ( .A1(n4553), .A2(n4554), .ZN(n4467) );
  AND2_X1 U5950 ( .A1(n4567), .A2(n4443), .ZN(n4468) );
  OR2_X1 U5951 ( .A1(n9504), .A2(n9503), .ZN(P1_U3260) );
  AND2_X1 U5952 ( .A1(n9310), .A2(n9312), .ZN(n4470) );
  AND2_X1 U5953 ( .A1(n5706), .A2(n5707), .ZN(n8855) );
  INV_X1 U5954 ( .A(n8855), .ZN(n4850) );
  AOI21_X1 U5955 ( .B1(n8721), .B2(n5589), .A(n5529), .ZN(n8642) );
  INV_X1 U5956 ( .A(n8642), .ZN(n4846) );
  NAND2_X1 U5957 ( .A1(n4512), .A2(n4444), .ZN(n8459) );
  NAND2_X1 U5958 ( .A1(n4876), .A2(n4879), .ZN(n5276) );
  NOR2_X1 U5959 ( .A1(n4426), .A2(n5324), .ZN(n5758) );
  NAND2_X1 U5960 ( .A1(n9688), .A2(n9542), .ZN(n4471) );
  NAND2_X1 U5961 ( .A1(n5560), .A2(n5559), .ZN(n8894) );
  INV_X1 U5962 ( .A(n8894), .ZN(n4650) );
  AND2_X1 U5963 ( .A1(n7181), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4472) );
  AND2_X1 U5964 ( .A1(n7186), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4473) );
  XNOR2_X1 U5965 ( .A(n7930), .B(n7928), .ZN(n7927) );
  NOR2_X1 U5966 ( .A1(n8393), .A2(n8392), .ZN(n4474) );
  INV_X1 U5967 ( .A(n8496), .ZN(n4754) );
  AND2_X1 U5968 ( .A1(n6739), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4475) );
  NAND2_X1 U5969 ( .A1(n5074), .A2(n5073), .ZN(n5324) );
  AND2_X1 U5970 ( .A1(n4753), .A2(n8439), .ZN(n4476) );
  NAND2_X1 U5971 ( .A1(n5701), .A2(n5700), .ZN(n7681) );
  AND3_X1 U5972 ( .A1(n9163), .A2(n9165), .A3(n4571), .ZN(n4477) );
  NOR3_X1 U5973 ( .A1(n8034), .A2(n9723), .A3(n4769), .ZN(n4767) );
  NAND2_X1 U5974 ( .A1(n5549), .A2(n5548), .ZN(n8899) );
  INV_X1 U5975 ( .A(n5074), .ZN(n5300) );
  OR2_X1 U5976 ( .A1(n5324), .A2(n4894), .ZN(n4478) );
  AND2_X1 U5977 ( .A1(n9759), .A2(n9868), .ZN(n4479) );
  NAND2_X1 U5978 ( .A1(n8865), .A2(n4645), .ZN(n4648) );
  INV_X1 U5979 ( .A(n4768), .ZN(n9640) );
  NOR2_X1 U5980 ( .A1(n8034), .A2(n4769), .ZN(n4768) );
  NAND2_X1 U5981 ( .A1(n8375), .A2(n8374), .ZN(n4480) );
  AND2_X1 U5982 ( .A1(n8240), .A2(n8239), .ZN(n9590) );
  NAND2_X1 U5983 ( .A1(n5470), .A2(n5473), .ZN(n4481) );
  AND2_X1 U5984 ( .A1(n6179), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4482) );
  INV_X1 U5985 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8997) );
  INV_X1 U5986 ( .A(n4939), .ZN(n4936) );
  NAND2_X1 U5987 ( .A1(n9714), .A2(n8399), .ZN(n4939) );
  INV_X1 U5988 ( .A(n10117), .ZN(n4906) );
  AND2_X1 U5989 ( .A1(n5794), .A2(n5793), .ZN(n5948) );
  NAND2_X1 U5990 ( .A1(n7674), .A2(n7675), .ZN(n7857) );
  NAND2_X1 U5991 ( .A1(n4528), .A2(n4527), .ZN(n7161) );
  NAND2_X1 U5992 ( .A1(n9393), .A2(n10039), .ZN(n9373) );
  NAND2_X1 U5993 ( .A1(n4899), .A2(n7028), .ZN(n7062) );
  NAND2_X1 U5994 ( .A1(n7303), .A2(n4756), .ZN(n7267) );
  OAI21_X1 U5995 ( .B1(n6866), .B2(n4453), .A(n4793), .ZN(n7113) );
  NAND2_X1 U5996 ( .A1(n5825), .A2(n5692), .ZN(n7364) );
  OAI21_X1 U5997 ( .B1(n7396), .B2(n7395), .A(n4739), .ZN(n7624) );
  NAND2_X1 U5998 ( .A1(n4870), .A2(n5678), .ZN(n7432) );
  AND2_X1 U5999 ( .A1(n4581), .A2(n4582), .ZN(n4483) );
  NAND2_X1 U6000 ( .A1(n4804), .A2(n6123), .ZN(n4484) );
  NOR2_X1 U6001 ( .A1(n7256), .A2(n7451), .ZN(n4485) );
  OAI211_X1 U6002 ( .C1(n5219), .C2(n6189), .A(n5222), .B(n4640), .ZN(n4639)
         );
  INV_X1 U6003 ( .A(n6625), .ZN(n6100) );
  XNOR2_X1 U6004 ( .A(n5083), .B(n5082), .ZN(n5763) );
  NAND4_X1 U6005 ( .A1(n5189), .A2(n5188), .A3(n5187), .A4(n5186), .ZN(n8563)
         );
  INV_X1 U6006 ( .A(n8563), .ZN(n4487) );
  NAND2_X1 U6007 ( .A1(n5303), .A2(n5302), .ZN(n10185) );
  INV_X1 U6008 ( .A(n10185), .ZN(n4655) );
  INV_X1 U6009 ( .A(n6988), .ZN(n4761) );
  INV_X1 U6010 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n4503) );
  INV_X1 U6011 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4504) );
  INV_X1 U6012 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4562) );
  INV_X1 U6013 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4789) );
  INV_X1 U6014 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5642) );
  INV_X1 U6015 ( .A(n5105), .ZN(n8435) );
  XNOR2_X1 U6016 ( .A(n5099), .B(n5098), .ZN(n5105) );
  INV_X1 U6017 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4506) );
  INV_X1 U6018 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4507) );
  NOR2_X2 U6019 ( .A1(n6902), .A2(n10039), .ZN(n9884) );
  AOI21_X2 U6020 ( .B1(n8670), .B2(n8663), .A(n5731), .ZN(n8649) );
  INV_X2 U6021 ( .A(n7540), .ZN(n10172) );
  INV_X1 U6022 ( .A(n7407), .ZN(n5683) );
  NAND2_X1 U6023 ( .A1(n4487), .A2(n7540), .ZN(n7407) );
  NAND3_X1 U6024 ( .A1(n8774), .A2(n5720), .A3(n5712), .ZN(n4488) );
  OAI21_X1 U6025 ( .B1(n4402), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n4489), .ZN(
        n4965) );
  NAND2_X1 U6026 ( .A1(n4402), .A2(n6178), .ZN(n4489) );
  XNOR2_X2 U6027 ( .A(n5194), .B(n5193), .ZN(n6191) );
  NAND2_X2 U6028 ( .A1(n4490), .A2(n4978), .ZN(n5194) );
  AND2_X1 U6029 ( .A1(n5691), .A2(n5317), .ZN(n4491) );
  OR2_X2 U6030 ( .A1(n5690), .A2(n5689), .ZN(n5691) );
  NAND2_X2 U6031 ( .A1(n9645), .A2(n9332), .ZN(n9632) );
  NAND3_X1 U6032 ( .A1(n9863), .A2(n9214), .A3(n4706), .ZN(n4499) );
  NAND2_X1 U6033 ( .A1(n4960), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4502) );
  NAND3_X1 U6034 ( .A1(n4504), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4500) );
  NAND3_X1 U6035 ( .A1(n4507), .A2(n4506), .A3(n4505), .ZN(n4501) );
  NAND3_X1 U6036 ( .A1(n4509), .A2(n9408), .A3(n4508), .ZN(n7079) );
  AND2_X1 U6037 ( .A1(n9229), .A2(n9275), .ZN(n9235) );
  NAND2_X1 U6038 ( .A1(n7938), .A2(n4513), .ZN(n4512) );
  AND3_X2 U6039 ( .A1(n4879), .A2(n4877), .A3(n4878), .ZN(n5074) );
  OAI21_X2 U6040 ( .B1(n7396), .B2(n4523), .A(n4520), .ZN(n7674) );
  NAND2_X2 U6041 ( .A1(n5763), .A2(n8044), .ZN(n5210) );
  XNOR2_X2 U6042 ( .A(n5085), .B(n5081), .ZN(n8044) );
  NAND2_X1 U6043 ( .A1(n8113), .A2(n8112), .ZN(n8126) );
  NAND2_X1 U6044 ( .A1(n8116), .A2(n8115), .ZN(n8124) );
  NAND2_X1 U6045 ( .A1(n7113), .A2(n6047), .ZN(n4532) );
  NAND2_X1 U6046 ( .A1(n4532), .A2(n6050), .ZN(n6119) );
  NAND2_X1 U6047 ( .A1(n6120), .A2(n4537), .ZN(n7345) );
  NOR2_X1 U6048 ( .A1(n8221), .A2(n8220), .ZN(n9095) );
  OAI22_X1 U6049 ( .A1(n7456), .A2(n4556), .B1(n4555), .B2(n4419), .ZN(n7964)
         );
  NAND2_X1 U6050 ( .A1(n5947), .A2(n5946), .ZN(n4561) );
  NAND2_X1 U6051 ( .A1(n4559), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U6052 ( .A1(n5947), .A2(n4560), .ZN(n4559) );
  XNOR2_X1 U6053 ( .A(n5957), .B(n8184), .ZN(n5972) );
  NAND4_X1 U6054 ( .A1(n4406), .A2(n6123), .A3(n5788), .A4(n5787), .ZN(n5789)
         );
  NAND2_X1 U6055 ( .A1(n5949), .A2(n4562), .ZN(n5986) );
  NAND2_X1 U6056 ( .A1(n4468), .A2(n4563), .ZN(n9326) );
  NAND3_X1 U6057 ( .A1(n4565), .A2(n4564), .A3(n4465), .ZN(n4563) );
  NAND2_X1 U6058 ( .A1(n9301), .A2(n9379), .ZN(n4564) );
  NAND2_X1 U6059 ( .A1(n9300), .A2(n9373), .ZN(n4565) );
  NAND2_X1 U6060 ( .A1(n4571), .A2(n6631), .ZN(n6950) );
  NAND2_X1 U6061 ( .A1(n6950), .A2(n4569), .ZN(n6634) );
  NAND2_X1 U6062 ( .A1(n4570), .A2(n6630), .ZN(n4569) );
  INV_X1 U6063 ( .A(n6631), .ZN(n4570) );
  NAND2_X1 U6064 ( .A1(n5965), .A2(n4482), .ZN(n4572) );
  NAND2_X4 U6065 ( .A1(n6102), .A2(n8427), .ZN(n5965) );
  NAND2_X2 U6066 ( .A1(n5965), .A2(n4398), .ZN(n9154) );
  OR2_X1 U6067 ( .A1(n9360), .A2(n4578), .ZN(n4573) );
  OR2_X1 U6068 ( .A1(n9350), .A2(n4579), .ZN(n4574) );
  AND3_X2 U6069 ( .A1(n4574), .A2(n4573), .A3(n4575), .ZN(n9372) );
  NAND2_X1 U6070 ( .A1(n4581), .A2(n4437), .ZN(n9284) );
  NAND3_X1 U6071 ( .A1(n4587), .A2(n4586), .A3(n9348), .ZN(n4585) );
  NAND2_X1 U6072 ( .A1(n9342), .A2(n9373), .ZN(n4586) );
  OAI21_X1 U6073 ( .B1(n9347), .B2(n9346), .A(n4588), .ZN(n4587) );
  INV_X1 U6074 ( .A(n5772), .ZN(n4589) );
  NAND2_X1 U6075 ( .A1(n4589), .A2(n5785), .ZN(n4590) );
  NAND2_X1 U6076 ( .A1(n4591), .A2(n4895), .ZN(n4894) );
  NAND2_X1 U6077 ( .A1(n5241), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4594) );
  NAND3_X1 U6078 ( .A1(n4598), .A2(n5554), .A3(n5555), .ZN(n4597) );
  OR2_X1 U6079 ( .A1(n5353), .A2(n4603), .ZN(n4601) );
  NAND2_X1 U6080 ( .A1(n4601), .A2(n4602), .ZN(n5389) );
  INV_X1 U6081 ( .A(n4610), .ZN(n4607) );
  NAND2_X1 U6082 ( .A1(n5700), .A2(n5294), .ZN(n4609) );
  NAND2_X1 U6083 ( .A1(n5613), .A2(n4613), .ZN(n4612) );
  NOR2_X1 U6084 ( .A1(n5324), .A2(n4410), .ZN(n4616) );
  NOR2_X1 U6085 ( .A1(n5324), .A2(n4403), .ZN(n4618) );
  NAND2_X1 U6086 ( .A1(n4619), .A2(n4617), .ZN(n8998) );
  NOR2_X1 U6087 ( .A1(n5324), .A2(n4415), .ZN(n4617) );
  AND2_X1 U6088 ( .A1(n5079), .A2(n5078), .ZN(n4634) );
  NAND2_X1 U6089 ( .A1(n5758), .A2(n5080), .ZN(n5084) );
  NAND2_X1 U6090 ( .A1(n4412), .A2(n7314), .ZN(n7428) );
  INV_X1 U6091 ( .A(n7004), .ZN(n7518) );
  INV_X1 U6092 ( .A(n4648), .ZN(n8799) );
  NOR2_X1 U6093 ( .A1(n8699), .A2(n8899), .ZN(n4651) );
  MUX2_X1 U6094 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n4398), .Z(n5208) );
  MUX2_X1 U6095 ( .A(n6175), .B(n6187), .S(n6179), .Z(n4973) );
  MUX2_X1 U6096 ( .A(n6173), .B(n6195), .S(n6179), .Z(n4969) );
  MUX2_X1 U6097 ( .A(n6174), .B(n6408), .S(n6179), .Z(n4976) );
  MUX2_X1 U6098 ( .A(n6411), .B(n6444), .S(n6179), .Z(n4986) );
  MUX2_X1 U6099 ( .A(n6177), .B(n6192), .S(n6179), .Z(n4979) );
  MUX2_X1 U6100 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6179), .Z(n4983) );
  MUX2_X1 U6101 ( .A(n6227), .B(n6219), .S(n6179), .Z(n4992) );
  MUX2_X1 U6102 ( .A(n6233), .B(n6231), .S(n6179), .Z(n4997) );
  AOI21_X1 U6103 ( .B1(n5282), .B2(n4660), .A(n4657), .ZN(n4656) );
  INV_X1 U6104 ( .A(n4656), .ZN(n5004) );
  NAND2_X1 U6105 ( .A1(n5194), .A2(n4665), .ZN(n4664) );
  NAND2_X1 U6106 ( .A1(n4664), .A2(n4667), .ZN(n4990) );
  NAND2_X1 U6107 ( .A1(n4672), .A2(n4671), .ZN(n5613) );
  OAI21_X1 U6108 ( .B1(n5594), .B2(n5294), .A(n5593), .ZN(n4671) );
  NOR2_X1 U6109 ( .A1(n5646), .A2(n5637), .ZN(n4673) );
  OAI21_X1 U6110 ( .B1(n5439), .B2(n4676), .A(n4675), .ZN(n5043) );
  NAND2_X1 U6111 ( .A1(n5341), .A2(n4683), .ZN(n4682) );
  NAND2_X1 U6112 ( .A1(n5058), .A2(n5057), .ZN(n5522) );
  NAND2_X1 U6113 ( .A1(n5058), .A2(n4689), .ZN(n4688) );
  NOR2_X1 U6114 ( .A1(n4709), .A2(n9213), .ZN(n4708) );
  NAND2_X1 U6115 ( .A1(n7250), .A2(n4718), .ZN(n4715) );
  NAND2_X1 U6116 ( .A1(n4715), .A2(n4716), .ZN(n9863) );
  NAND2_X1 U6117 ( .A1(n7840), .A2(n4725), .ZN(n7919) );
  NAND2_X1 U6118 ( .A1(n6950), .A2(n6949), .ZN(n9405) );
  NAND4_X1 U6119 ( .A1(n4804), .A2(n4440), .A3(n6123), .A4(n4729), .ZN(n5933)
         );
  NAND2_X1 U6120 ( .A1(n6951), .A2(n9402), .ZN(n9236) );
  AOI22_X2 U6121 ( .A1(n8416), .A2(n9270), .B1(n9201), .B2(n9202), .ZN(n9663)
         );
  NAND2_X1 U6122 ( .A1(n7919), .A2(n9323), .ZN(n8416) );
  NAND2_X1 U6123 ( .A1(n9663), .A2(n9664), .ZN(n9662) );
  NAND2_X1 U6124 ( .A1(n5177), .A2(n5176), .ZN(n5163) );
  NAND2_X1 U6125 ( .A1(n5028), .A2(n5027), .ZN(n5421) );
  AOI21_X2 U6126 ( .B1(n9576), .B2(n8418), .A(n9354), .ZN(n9553) );
  NAND2_X1 U6127 ( .A1(n7197), .A2(n9291), .ZN(n7250) );
  OAI21_X1 U6128 ( .B1(n9686), .B2(n9822), .A(n9685), .ZN(n9773) );
  NAND2_X1 U6129 ( .A1(n5874), .A2(n5873), .ZN(n4734) );
  OAI21_X1 U6130 ( .B1(n7396), .B2(n4743), .A(n4740), .ZN(n7672) );
  NAND2_X1 U6131 ( .A1(n7623), .A2(n4744), .ZN(n4743) );
  OAI21_X1 U6132 ( .B1(n8497), .B2(n8492), .A(n8496), .ZN(n8543) );
  OAI211_X2 U6133 ( .C1(n8450), .C2(n8361), .A(n8360), .B(n8359), .ZN(n8497)
         );
  NAND2_X1 U6134 ( .A1(n8497), .A2(n4753), .ZN(n4747) );
  NAND2_X1 U6135 ( .A1(n5126), .A2(n4755), .ZN(n5440) );
  INV_X1 U6136 ( .A(n5440), .ZN(n5131) );
  NAND2_X1 U6137 ( .A1(n7267), .A2(n7266), .ZN(n7269) );
  AND2_X1 U6138 ( .A1(n5907), .A2(n5901), .ZN(n4756) );
  NAND2_X1 U6139 ( .A1(n8460), .A2(n4757), .ZN(n8517) );
  NAND2_X1 U6140 ( .A1(n8517), .A2(n8093), .ZN(n8094) );
  NAND2_X1 U6141 ( .A1(n5074), .A2(n4759), .ZN(n5392) );
  INV_X1 U6142 ( .A(n4766), .ZN(n9560) );
  INV_X1 U6143 ( .A(n4767), .ZN(n9626) );
  INV_X1 U6144 ( .A(n7256), .ZN(n4772) );
  NAND2_X1 U6145 ( .A1(n4772), .A2(n4773), .ZN(n9880) );
  NOR2_X1 U6146 ( .A1(n7256), .A2(n4775), .ZN(n9882) );
  XNOR2_X1 U6147 ( .A(n9468), .B(n9485), .ZN(n9983) );
  NAND3_X1 U6148 ( .A1(n8138), .A2(n9055), .A3(n9068), .ZN(n4798) );
  NAND2_X1 U6149 ( .A1(n9045), .A2(n9046), .ZN(n4810) );
  AND2_X1 U6150 ( .A1(n4810), .A2(n4809), .ZN(n9122) );
  NAND2_X1 U6151 ( .A1(n8269), .A2(n8268), .ZN(n4809) );
  INV_X1 U6152 ( .A(n9038), .ZN(n4815) );
  AND2_X1 U6153 ( .A1(n7986), .A2(n4821), .ZN(n7361) );
  NAND2_X1 U6154 ( .A1(n8690), .A2(n4411), .ZN(n4822) );
  NAND2_X1 U6155 ( .A1(n8690), .A2(n8694), .ZN(n4824) );
  NAND2_X1 U6156 ( .A1(n4822), .A2(n4823), .ZN(n8664) );
  INV_X1 U6157 ( .A(n8899), .ZN(n4827) );
  NAND2_X1 U6158 ( .A1(n7684), .A2(n4840), .ZN(n4830) );
  NAND2_X1 U6159 ( .A1(n4831), .A2(n4836), .ZN(n7874) );
  NAND2_X1 U6160 ( .A1(n7685), .A2(n4837), .ZN(n4831) );
  AOI21_X1 U6161 ( .B1(n4834), .B2(n4836), .A(n4833), .ZN(n4832) );
  NOR2_X1 U6162 ( .A1(n4837), .A2(n7869), .ZN(n4834) );
  INV_X1 U6163 ( .A(n4843), .ZN(n8707) );
  NAND2_X1 U6164 ( .A1(n8856), .A2(n4851), .ZN(n4847) );
  NAND2_X1 U6165 ( .A1(n4847), .A2(n4848), .ZN(n8811) );
  AND2_X1 U6166 ( .A1(n8956), .A2(n8630), .ZN(n4854) );
  NAND2_X1 U6167 ( .A1(n4857), .A2(n4984), .ZN(n5272) );
  NAND2_X1 U6168 ( .A1(n7601), .A2(n4858), .ZN(n7596) );
  NAND2_X1 U6169 ( .A1(n4859), .A2(n7362), .ZN(n7982) );
  OAI21_X1 U6170 ( .B1(n7364), .B2(n4867), .A(n4863), .ZN(n7637) );
  NAND2_X1 U6171 ( .A1(n7364), .A2(n4863), .ZN(n4862) );
  OAI211_X1 U6172 ( .C1(n8774), .C2(n4874), .A(n4871), .B(n5720), .ZN(n8733)
         );
  AOI21_X1 U6173 ( .B1(n4874), .B2(n5720), .A(n4873), .ZN(n4872) );
  INV_X1 U6174 ( .A(n5721), .ZN(n4873) );
  INV_X1 U6175 ( .A(n5719), .ZN(n4874) );
  INV_X1 U6176 ( .A(n5072), .ZN(n4877) );
  NAND2_X1 U6177 ( .A1(n7863), .A2(n4463), .ZN(n4880) );
  NAND2_X1 U6178 ( .A1(n4880), .A2(n4881), .ZN(n8843) );
  OAI21_X2 U6179 ( .B1(n4889), .B2(n5725), .A(n4886), .ZN(n8670) );
  AOI21_X1 U6180 ( .B1(n5727), .B2(n4888), .A(n4887), .ZN(n4886) );
  INV_X1 U6181 ( .A(n5727), .ZN(n4889) );
  NAND2_X1 U6182 ( .A1(n5725), .A2(n4890), .ZN(n5728) );
  NAND2_X1 U6183 ( .A1(n7026), .A2(n9167), .ZN(n4899) );
  NAND2_X1 U6184 ( .A1(n9517), .A2(n4909), .ZN(n4902) );
  OAI211_X1 U6185 ( .C1(n9685), .C2(n4906), .A(n4900), .B(n4907), .ZN(P1_U3552) );
  NAND2_X1 U6186 ( .A1(n5949), .A2(n4910), .ZN(n6022) );
  NAND2_X1 U6187 ( .A1(n7553), .A2(n4913), .ZN(n4912) );
  NAND2_X1 U6188 ( .A1(n9559), .A2(n4920), .ZN(n4916) );
  NAND2_X1 U6189 ( .A1(n4916), .A2(n4917), .ZN(n9518) );
  NAND2_X1 U6190 ( .A1(n8393), .A2(n4930), .ZN(n4927) );
  NAND2_X1 U6191 ( .A1(n4927), .A2(n4928), .ZN(n9625) );
  INV_X1 U6192 ( .A(n8394), .ZN(n4933) );
  NAND2_X1 U6193 ( .A1(n8398), .A2(n4937), .ZN(n4935) );
  MUX2_X1 U6194 ( .A(n9367), .B(n9366), .S(n9373), .Z(n9368) );
  INV_X1 U6195 ( .A(n5864), .ZN(n5742) );
  INV_X1 U6196 ( .A(n5741), .ZN(n5855) );
  OR2_X1 U6197 ( .A1(n8353), .A2(n8352), .ZN(n8354) );
  NAND2_X1 U6198 ( .A1(n6149), .A2(n6148), .ZN(n7454) );
  INV_X1 U6199 ( .A(n5392), .ZN(n5126) );
  INV_X1 U6200 ( .A(n6151), .ZN(n6149) );
  OAI21_X2 U6201 ( .B1(n5489), .B2(n5047), .A(n5046), .ZN(n5499) );
  NAND2_X1 U6202 ( .A1(n8018), .A2(n8017), .ZN(n8393) );
  OR2_X1 U6203 ( .A1(n5100), .A2(n8997), .ZN(n5102) );
  NAND2_X1 U6204 ( .A1(n5131), .A2(n5130), .ZN(n5134) );
  NOR2_X2 U6205 ( .A1(n7045), .A2(n7051), .ZN(n7074) );
  NAND2_X2 U6206 ( .A1(n7605), .A2(n7604), .ZN(n7685) );
  INV_X1 U6207 ( .A(n9582), .ZN(n8403) );
  AND4_X1 U6208 ( .A1(n8248), .A2(n8247), .A3(n8246), .A4(n8245), .ZN(n9598)
         );
  AND4_X1 U6209 ( .A1(n8233), .A2(n8232), .A3(n8231), .A4(n8230), .ZN(n9581)
         );
  INV_X1 U6210 ( .A(n9581), .ZN(n8399) );
  AND2_X1 U6211 ( .A1(n6629), .A2(n9438), .ZN(n9865) );
  AND2_X1 U6212 ( .A1(n5320), .A2(n4999), .ZN(n4946) );
  NOR2_X1 U6213 ( .A1(n4974), .A2(n5164), .ZN(n4949) );
  AND4_X1 U6214 ( .A1(n6908), .A2(n6236), .A3(n5776), .A4(n5775), .ZN(n4950)
         );
  NAND2_X1 U6215 ( .A1(n5553), .A2(n5724), .ZN(n4952) );
  INV_X1 U6216 ( .A(n9703), .ZN(n9564) );
  AND4_X1 U6217 ( .A1(n5495), .A2(n5494), .A3(n5493), .A4(n5492), .ZN(n8762)
         );
  AOI21_X1 U6218 ( .B1(n6229), .B2(n8324), .A(n5970), .ZN(n6604) );
  AND3_X1 U6219 ( .A1(n5515), .A2(n5650), .A3(n5649), .ZN(n4953) );
  OR2_X1 U6220 ( .A1(n8165), .A2(n9028), .ZN(n4954) );
  INV_X1 U6221 ( .A(n8946), .ZN(n8816) );
  NAND2_X1 U6222 ( .A1(n8777), .A2(n8776), .ZN(n4956) );
  INV_X1 U6223 ( .A(n8906), .ZN(n8366) );
  OR2_X1 U6224 ( .A1(n8773), .A2(n8762), .ZN(n4958) );
  NOR2_X1 U6225 ( .A1(n5295), .A2(n5294), .ZN(n5296) );
  NOR2_X1 U6226 ( .A1(n4868), .A2(n5296), .ZN(n5297) );
  OAI21_X1 U6227 ( .B1(n5298), .B2(n5637), .A(n5297), .ZN(n5315) );
  AND2_X1 U6228 ( .A1(n7869), .A2(n5387), .ZN(n5388) );
  AND2_X1 U6229 ( .A1(n5650), .A2(n5714), .ZN(n5496) );
  NAND2_X1 U6230 ( .A1(n4953), .A2(n5294), .ZN(n5517) );
  OAI211_X1 U6231 ( .C1(n5518), .C2(n5294), .A(n5517), .B(n5516), .ZN(n5519)
         );
  NAND2_X1 U6232 ( .A1(n4952), .A2(n5294), .ZN(n5539) );
  INV_X1 U6233 ( .A(n5645), .ZN(n5592) );
  NOR2_X1 U6234 ( .A1(n5645), .A2(n5637), .ZN(n5608) );
  NOR2_X1 U6235 ( .A1(n5609), .A2(n5608), .ZN(n5611) );
  OAI211_X1 U6236 ( .C1(n5733), .C2(n8623), .A(n5762), .B(n6611), .ZN(n5734)
         );
  AND2_X1 U6237 ( .A1(n5611), .A2(n5636), .ZN(n5612) );
  INV_X1 U6238 ( .A(n8643), .ZN(n8644) );
  NAND2_X1 U6239 ( .A1(n7344), .A2(n7348), .ZN(n6151) );
  INV_X1 U6240 ( .A(n5380), .ZN(n5090) );
  INV_X1 U6241 ( .A(n5329), .ZN(n5089) );
  INV_X1 U6242 ( .A(n5445), .ZN(n5093) );
  NAND2_X1 U6243 ( .A1(n8366), .A2(n8644), .ZN(n8645) );
  INV_X1 U6244 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5125) );
  INV_X1 U6245 ( .A(n6150), .ZN(n6148) );
  NAND2_X1 U6246 ( .A1(n5965), .A2(n4402), .ZN(n6003) );
  INV_X1 U6247 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5787) );
  AND2_X1 U6248 ( .A1(n5354), .A2(n5357), .ZN(n5012) );
  AND2_X1 U6249 ( .A1(n5322), .A2(n5320), .ZN(n5000) );
  INV_X1 U6250 ( .A(n5250), .ZN(n4982) );
  NAND2_X1 U6251 ( .A1(n5090), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5397) );
  OR2_X1 U6252 ( .A1(n5346), .A2(n5345), .ZN(n5367) );
  INV_X1 U6253 ( .A(n5287), .ZN(n5088) );
  INV_X1 U6254 ( .A(n8520), .ZN(n8092) );
  OR2_X1 U6255 ( .A1(n5367), .A2(n7107), .ZN(n5380) );
  OR2_X1 U6256 ( .A1(n5116), .A2(n8545), .ZN(n5562) );
  OR2_X1 U6257 ( .A1(n5463), .A2(n8464), .ZN(n5481) );
  NOR2_X1 U6258 ( .A1(n5183), .A2(n5182), .ZN(n5243) );
  NAND2_X1 U6259 ( .A1(n8229), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8243) );
  INV_X1 U6260 ( .A(n8284), .ZN(n8285) );
  NAND2_X1 U6261 ( .A1(n8259), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8274) );
  AND2_X1 U6262 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6031) );
  INV_X1 U6263 ( .A(n6867), .ZN(n6013) );
  NAND2_X1 U6264 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n8275), .ZN(n8310) );
  OR2_X1 U6265 ( .A1(n7757), .A2(n9058), .ZN(n7833) );
  NOR2_X1 U6266 ( .A1(n9714), .A2(n8399), .ZN(n8400) );
  INV_X1 U6267 ( .A(n9163), .ZN(n6945) );
  NAND2_X1 U6268 ( .A1(n5018), .A2(n5017), .ZN(n5021) );
  NAND2_X1 U6269 ( .A1(n5007), .A2(n5006), .ZN(n5354) );
  NAND2_X1 U6270 ( .A1(n5153), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5183) );
  INV_X1 U6271 ( .A(n7949), .ZN(n7950) );
  NAND2_X1 U6272 ( .A1(n5088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5305) );
  INV_X1 U6273 ( .A(n7160), .ZN(n5762) );
  INV_X1 U6274 ( .A(n5265), .ZN(n5589) );
  AND2_X1 U6275 ( .A1(n8936), .A2(n8806), .ZN(n8638) );
  NOR2_X1 U6276 ( .A1(n8946), .A2(n8805), .ZN(n8633) );
  NAND2_X1 U6277 ( .A1(n7985), .A2(n7600), .ZN(n7983) );
  OR2_X1 U6278 ( .A1(n5263), .A2(n5262), .ZN(n5287) );
  OR2_X1 U6279 ( .A1(n5849), .A2(n10130), .ZN(n5853) );
  AND2_X1 U6280 ( .A1(n5826), .A2(n5864), .ZN(n8759) );
  OR3_X1 U6281 ( .A1(n7381), .A2(n7742), .A3(n7647), .ZN(n5922) );
  NAND2_X1 U6282 ( .A1(n7966), .A2(n7965), .ZN(n8116) );
  NOR2_X1 U6283 ( .A1(n8329), .A2(n9146), .ZN(n8330) );
  OR2_X1 U6284 ( .A1(n6140), .A2(n6166), .ZN(n6158) );
  NAND2_X1 U6285 ( .A1(n8252), .A2(n8251), .ZN(n8253) );
  OR2_X1 U6286 ( .A1(n8173), .A2(n8172), .ZN(n8193) );
  OR2_X1 U6287 ( .A1(n8332), .A2(n9536), .ZN(n8294) );
  NAND2_X1 U6288 ( .A1(n8027), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8173) );
  NOR2_X1 U6289 ( .A1(n7833), .A2(n7832), .ZN(n7914) );
  OR2_X1 U6290 ( .A1(n5996), .A2(n5979), .ZN(n5983) );
  INV_X1 U6291 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U6292 ( .A1(n9590), .A2(n9598), .ZN(n8401) );
  INV_X1 U6293 ( .A(n9450), .ZN(n9060) );
  AND2_X1 U6294 ( .A1(n9302), .A2(n9298), .ZN(n9879) );
  AND2_X1 U6295 ( .A1(n9218), .A2(n9291), .ZN(n9171) );
  INV_X1 U6296 ( .A(n6976), .ZN(n10072) );
  NAND2_X1 U6297 ( .A1(n5354), .A2(n5009), .ZN(n5340) );
  NAND2_X1 U6298 ( .A1(n4990), .A2(n4989), .ZN(n5282) );
  INV_X1 U6299 ( .A(n7468), .ZN(n7412) );
  NAND2_X1 U6300 ( .A1(n7269), .A2(n7268), .ZN(n7396) );
  NAND2_X1 U6301 ( .A1(n8094), .A2(n8480), .ZN(n8483) );
  NAND2_X1 U6302 ( .A1(n7145), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8546) );
  INV_X1 U6303 ( .A(n8553), .ZN(n8476) );
  NAND2_X1 U6304 ( .A1(n5919), .A2(n8835), .ZN(n8551) );
  AND2_X1 U6305 ( .A1(n5571), .A2(n5570), .ZN(n8684) );
  AND4_X1 U6306 ( .A1(n5435), .A2(n5434), .A3(n5433), .A4(n5432), .ZN(n8852)
         );
  AND2_X1 U6307 ( .A1(n6727), .A2(n6726), .ZN(n10119) );
  INV_X1 U6308 ( .A(n8879), .ZN(n8042) );
  INV_X1 U6309 ( .A(n8669), .ZN(n8663) );
  NAND2_X1 U6310 ( .A1(n5649), .A2(n5648), .ZN(n8761) );
  INV_X1 U6311 ( .A(n8851), .ZN(n8821) );
  NAND2_X1 U6312 ( .A1(n5853), .A2(n8835), .ZN(n8846) );
  OR2_X1 U6313 ( .A1(n5862), .A2(n5861), .ZN(n10186) );
  INV_X1 U6314 ( .A(n10177), .ZN(n10199) );
  NAND2_X1 U6315 ( .A1(n8859), .A2(n8977), .ZN(n10177) );
  NAND2_X1 U6316 ( .A1(n5922), .A2(n10144), .ZN(n10130) );
  AND4_X1 U6317 ( .A1(n8264), .A2(n8263), .A3(n8262), .A4(n8261), .ZN(n9582)
         );
  INV_X1 U6318 ( .A(n6276), .ZN(n9918) );
  INV_X1 U6319 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6166) );
  AND2_X1 U6320 ( .A1(n8415), .A2(n8414), .ZN(n9325) );
  AND2_X1 U6321 ( .A1(n9220), .A2(n9216), .ZN(n9178) );
  INV_X1 U6322 ( .A(n9599), .ZN(n9867) );
  MUX2_X1 U6323 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9798), .S(n5965), .Z(n6904) );
  AND2_X1 U6324 ( .A1(n6083), .A2(n6200), .ZN(n6897) );
  AND2_X1 U6325 ( .A1(n9680), .A2(n10065), .ZN(n9822) );
  OR2_X1 U6326 ( .A1(n9373), .A2(n9396), .ZN(n10065) );
  AND2_X1 U6327 ( .A1(n6125), .A2(n6124), .ZN(n6671) );
  XNOR2_X1 U6328 ( .A(n4969), .B(SI_3_), .ZN(n5176) );
  INV_X1 U6329 ( .A(n8588), .ZN(n10124) );
  INV_X1 U6330 ( .A(n8914), .ZN(n8723) );
  OR3_X1 U6331 ( .A1(n5926), .A2(n6708), .A3(n10194), .ZN(n8553) );
  INV_X1 U6332 ( .A(n9815), .ZN(n10121) );
  INV_X1 U6333 ( .A(n10217), .ZN(n10215) );
  INV_X1 U6334 ( .A(n10204), .ZN(n10202) );
  AND2_X1 U6335 ( .A1(n5921), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10144) );
  XNOR2_X1 U6336 ( .A(n5757), .B(n5756), .ZN(n7381) );
  INV_X1 U6337 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6444) );
  INV_X1 U6338 ( .A(n9728), .ZN(n9644) );
  INV_X1 U6339 ( .A(n9598), .ZN(n9567) );
  INV_X1 U6340 ( .A(n6952), .ZN(n9461) );
  INV_X1 U6341 ( .A(n9513), .ZN(n9679) );
  INV_X1 U6342 ( .A(n10107), .ZN(n10105) );
  AND2_X1 U6343 ( .A1(n6093), .A2(n6085), .ZN(n9439) );
  INV_X1 U6344 ( .A(n9442), .ZN(n9393) );
  INV_X1 U6345 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6411) );
  INV_X1 U6346 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6175) );
  INV_X1 U6347 ( .A(n8567), .ZN(P2_U3966) );
  NAND2_X1 U6348 ( .A1(n4959), .A2(SI_0_), .ZN(n4961) );
  XNOR2_X1 U6349 ( .A(n4961), .B(SI_1_), .ZN(n5209) );
  NAND2_X1 U6350 ( .A1(n5209), .A2(n5208), .ZN(n4964) );
  INV_X1 U6351 ( .A(n4961), .ZN(n4962) );
  NAND2_X1 U6352 ( .A1(n4962), .A2(SI_1_), .ZN(n4963) );
  NAND2_X1 U6353 ( .A1(n4964), .A2(n4963), .ZN(n5218) );
  INV_X1 U6354 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6190) );
  INV_X1 U6355 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U6356 ( .A1(n5218), .A2(n5217), .ZN(n4968) );
  INV_X1 U6357 ( .A(n4965), .ZN(n4966) );
  NAND2_X1 U6358 ( .A1(n4966), .A2(SI_2_), .ZN(n4967) );
  NAND2_X1 U6359 ( .A1(n4968), .A2(n4967), .ZN(n5177) );
  INV_X1 U6360 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6195) );
  INV_X1 U6361 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6173) );
  INV_X1 U6362 ( .A(n4969), .ZN(n4970) );
  NAND2_X1 U6363 ( .A1(n4970), .A2(SI_3_), .ZN(n5162) );
  INV_X1 U6364 ( .A(n4973), .ZN(n4971) );
  NAND2_X1 U6365 ( .A1(n4971), .A2(SI_4_), .ZN(n4972) );
  AND2_X1 U6366 ( .A1(n5162), .A2(n4972), .ZN(n4975) );
  INV_X1 U6367 ( .A(n4972), .ZN(n4974) );
  INV_X1 U6368 ( .A(n4976), .ZN(n4977) );
  NAND2_X1 U6369 ( .A1(n4977), .A2(SI_5_), .ZN(n4978) );
  INV_X1 U6370 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6177) );
  INV_X1 U6371 ( .A(n4979), .ZN(n4980) );
  NAND2_X1 U6372 ( .A1(n4980), .A2(SI_6_), .ZN(n4981) );
  NAND2_X1 U6373 ( .A1(n4983), .A2(SI_7_), .ZN(n4984) );
  INV_X1 U6374 ( .A(SI_8_), .ZN(n4985) );
  INV_X1 U6375 ( .A(n4986), .ZN(n4987) );
  NAND2_X1 U6376 ( .A1(n4987), .A2(SI_8_), .ZN(n4988) );
  INV_X1 U6377 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6219) );
  INV_X1 U6378 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6227) );
  INV_X1 U6379 ( .A(SI_9_), .ZN(n4991) );
  INV_X1 U6380 ( .A(n4992), .ZN(n4993) );
  NAND2_X1 U6381 ( .A1(n4993), .A2(SI_9_), .ZN(n4994) );
  INV_X1 U6382 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6231) );
  INV_X1 U6383 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6233) );
  INV_X1 U6384 ( .A(SI_10_), .ZN(n4996) );
  INV_X1 U6385 ( .A(n4997), .ZN(n4998) );
  NAND2_X1 U6386 ( .A1(n4998), .A2(SI_10_), .ZN(n4999) );
  INV_X1 U6387 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6457) );
  INV_X1 U6388 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6551) );
  MUX2_X1 U6389 ( .A(n6457), .B(n6551), .S(n4402), .Z(n5001) );
  INV_X1 U6390 ( .A(n5001), .ZN(n5002) );
  NAND2_X1 U6391 ( .A1(n5002), .A2(SI_11_), .ZN(n5003) );
  NAND2_X1 U6392 ( .A1(n5004), .A2(n5003), .ZN(n5341) );
  INV_X1 U6393 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6549) );
  INV_X1 U6394 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5005) );
  MUX2_X1 U6395 ( .A(n6549), .B(n5005), .S(n4402), .Z(n5007) );
  INV_X1 U6396 ( .A(SI_12_), .ZN(n5006) );
  INV_X1 U6397 ( .A(n5007), .ZN(n5008) );
  NAND2_X1 U6398 ( .A1(n5008), .A2(SI_12_), .ZN(n5009) );
  INV_X1 U6399 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6323) );
  INV_X1 U6400 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5010) );
  MUX2_X1 U6401 ( .A(n6323), .B(n5010), .S(n4402), .Z(n5013) );
  INV_X1 U6402 ( .A(SI_13_), .ZN(n5011) );
  NAND2_X1 U6403 ( .A1(n5013), .A2(n5011), .ZN(n5357) );
  INV_X1 U6404 ( .A(n5013), .ZN(n5014) );
  NAND2_X1 U6405 ( .A1(n5014), .A2(SI_13_), .ZN(n5356) );
  INV_X1 U6406 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6596) );
  INV_X1 U6407 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6601) );
  MUX2_X1 U6408 ( .A(n6596), .B(n6601), .S(n4402), .Z(n5015) );
  INV_X1 U6409 ( .A(n5015), .ZN(n5016) );
  INV_X1 U6410 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6696) );
  INV_X1 U6411 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6699) );
  MUX2_X1 U6412 ( .A(n6696), .B(n6699), .S(n4402), .Z(n5018) );
  INV_X1 U6413 ( .A(SI_15_), .ZN(n5017) );
  INV_X1 U6414 ( .A(n5018), .ZN(n5019) );
  NAND2_X1 U6415 ( .A1(n5019), .A2(SI_15_), .ZN(n5020) );
  OAI21_X1 U6416 ( .B1(n5391), .B2(n5390), .A(n5021), .ZN(n5408) );
  INV_X1 U6417 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6701) );
  INV_X1 U6418 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5022) );
  MUX2_X1 U6419 ( .A(n6701), .B(n5022), .S(n4402), .Z(n5024) );
  INV_X1 U6420 ( .A(SI_16_), .ZN(n5023) );
  NAND2_X1 U6421 ( .A1(n5024), .A2(n5023), .ZN(n5027) );
  INV_X1 U6422 ( .A(n5024), .ZN(n5025) );
  NAND2_X1 U6423 ( .A1(n5025), .A2(SI_16_), .ZN(n5026) );
  NAND2_X1 U6424 ( .A1(n5408), .A2(n5407), .ZN(n5028) );
  INV_X1 U6425 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6784) );
  INV_X1 U6426 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5029) );
  MUX2_X1 U6427 ( .A(n6784), .B(n5029), .S(n4402), .Z(n5030) );
  XNOR2_X1 U6428 ( .A(n5030), .B(SI_17_), .ZN(n5420) );
  INV_X1 U6429 ( .A(n5420), .ZN(n5033) );
  INV_X1 U6430 ( .A(n5030), .ZN(n5031) );
  NAND2_X1 U6431 ( .A1(n5031), .A2(SI_17_), .ZN(n5032) );
  OAI21_X2 U6432 ( .B1(n5421), .B2(n5033), .A(n5032), .ZN(n5439) );
  MUX2_X1 U6433 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4402), .Z(n5035) );
  XNOR2_X1 U6434 ( .A(n5035), .B(SI_18_), .ZN(n5438) );
  INV_X1 U6435 ( .A(n5438), .ZN(n5034) );
  NAND2_X1 U6436 ( .A1(n5035), .A2(SI_18_), .ZN(n5036) );
  INV_X1 U6437 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6982) );
  INV_X1 U6438 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6979) );
  MUX2_X1 U6439 ( .A(n6982), .B(n6979), .S(n4402), .Z(n5037) );
  INV_X1 U6440 ( .A(SI_19_), .ZN(n6524) );
  NAND2_X1 U6441 ( .A1(n5037), .A2(n6524), .ZN(n5470) );
  INV_X1 U6442 ( .A(n5037), .ZN(n5038) );
  NAND2_X1 U6443 ( .A1(n5038), .A2(SI_19_), .ZN(n5039) );
  NAND2_X1 U6444 ( .A1(n5470), .A2(n5039), .ZN(n5456) );
  INV_X1 U6445 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7960) );
  INV_X1 U6446 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8169) );
  MUX2_X1 U6447 ( .A(n7960), .B(n8169), .S(n4402), .Z(n5041) );
  INV_X1 U6448 ( .A(SI_20_), .ZN(n5040) );
  NAND2_X1 U6449 ( .A1(n5041), .A2(n5040), .ZN(n5473) );
  INV_X1 U6450 ( .A(n5041), .ZN(n5042) );
  NAND2_X1 U6451 ( .A1(n5042), .A2(SI_20_), .ZN(n5472) );
  INV_X1 U6452 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7159) );
  INV_X1 U6453 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8190) );
  MUX2_X1 U6454 ( .A(n7159), .B(n8190), .S(n4402), .Z(n5044) );
  XNOR2_X1 U6455 ( .A(n5044), .B(SI_21_), .ZN(n5488) );
  INV_X1 U6456 ( .A(n5488), .ZN(n5047) );
  INV_X1 U6457 ( .A(n5044), .ZN(n5045) );
  NAND2_X1 U6458 ( .A1(n5045), .A2(SI_21_), .ZN(n5046) );
  INV_X1 U6459 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8111) );
  INV_X1 U6460 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8209) );
  MUX2_X1 U6461 ( .A(n8111), .B(n8209), .S(n4402), .Z(n5049) );
  INV_X1 U6462 ( .A(SI_22_), .ZN(n5048) );
  NAND2_X1 U6463 ( .A1(n5049), .A2(n5048), .ZN(n5052) );
  INV_X1 U6464 ( .A(n5049), .ZN(n5050) );
  NAND2_X1 U6465 ( .A1(n5050), .A2(SI_22_), .ZN(n5051) );
  NAND2_X1 U6466 ( .A1(n5052), .A2(n5051), .ZN(n5498) );
  INV_X1 U6467 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7302) );
  INV_X1 U6468 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8223) );
  MUX2_X1 U6469 ( .A(n7302), .B(n8223), .S(n4402), .Z(n5054) );
  INV_X1 U6470 ( .A(SI_23_), .ZN(n5053) );
  NAND2_X1 U6471 ( .A1(n5054), .A2(n5053), .ZN(n5057) );
  INV_X1 U6472 ( .A(n5054), .ZN(n5055) );
  NAND2_X1 U6473 ( .A1(n5055), .A2(SI_23_), .ZN(n5056) );
  NAND2_X1 U6474 ( .A1(n5136), .A2(n5135), .ZN(n5058) );
  INV_X1 U6475 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7380) );
  INV_X1 U6476 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8238) );
  MUX2_X1 U6477 ( .A(n7380), .B(n8238), .S(n4402), .Z(n5059) );
  XNOR2_X1 U6478 ( .A(n5059), .B(SI_24_), .ZN(n5521) );
  INV_X1 U6479 ( .A(n5521), .ZN(n5062) );
  INV_X1 U6480 ( .A(n5059), .ZN(n5060) );
  NAND2_X1 U6481 ( .A1(n5060), .A2(SI_24_), .ZN(n5061) );
  INV_X1 U6482 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7649) );
  INV_X1 U6483 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8255) );
  MUX2_X1 U6484 ( .A(n7649), .B(n8255), .S(n4402), .Z(n5063) );
  INV_X1 U6485 ( .A(SI_25_), .ZN(n6493) );
  NAND2_X1 U6486 ( .A1(n5063), .A2(n6493), .ZN(n5066) );
  INV_X1 U6487 ( .A(n5063), .ZN(n5064) );
  NAND2_X1 U6488 ( .A1(n5064), .A2(SI_25_), .ZN(n5065) );
  NAND2_X1 U6489 ( .A1(n5066), .A2(n5065), .ZN(n5111) );
  INV_X1 U6490 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7741) );
  INV_X1 U6491 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8271) );
  MUX2_X1 U6492 ( .A(n7741), .B(n8271), .S(n4402), .Z(n5068) );
  INV_X1 U6493 ( .A(SI_26_), .ZN(n5067) );
  NAND2_X1 U6494 ( .A1(n5068), .A2(n5067), .ZN(n5543) );
  INV_X1 U6495 ( .A(n5068), .ZN(n5069) );
  NAND2_X1 U6496 ( .A1(n5069), .A2(SI_26_), .ZN(n5070) );
  AND2_X1 U6497 ( .A1(n5543), .A2(n5070), .ZN(n5541) );
  NAND2_X1 U6498 ( .A1(n5220), .A2(n5071), .ZN(n5146) );
  NOR2_X1 U6499 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5075) );
  INV_X1 U6500 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U6501 ( .A1(n5642), .A2(n5639), .ZN(n5129) );
  INV_X1 U6502 ( .A(n5129), .ZN(n5076) );
  NOR2_X1 U6503 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5079) );
  NOR2_X1 U6504 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5078) );
  NOR2_X1 U6505 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5077) );
  INV_X1 U6506 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5080) );
  INV_X1 U6507 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5081) );
  INV_X1 U6508 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5082) );
  NAND2_X1 U6509 ( .A1(n5084), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5085) );
  NAND2_X1 U6510 ( .A1(n8270), .A2(n5623), .ZN(n5087) );
  OR2_X1 U6511 ( .A1(n4397), .A2(n7741), .ZN(n5086) );
  NAND2_X1 U6512 ( .A1(n5243), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5263) );
  INV_X1 U6513 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5262) );
  INV_X1 U6514 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5304) );
  INV_X1 U6515 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5345) );
  INV_X1 U6516 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7107) );
  NAND2_X1 U6517 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_17__SCAN_IN), 
        .ZN(n5092) );
  INV_X1 U6518 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8464) );
  NAND2_X1 U6519 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n5095) );
  INV_X1 U6520 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8453) );
  OR2_X2 U6521 ( .A1(n5505), .A2(n8453), .ZN(n5525) );
  INV_X1 U6522 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8501) );
  INV_X1 U6523 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8512) );
  OR3_X2 U6524 ( .A1(n5525), .A2(n8501), .A3(n8512), .ZN(n5116) );
  INV_X1 U6525 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U6526 ( .A1(n5116), .A2(n8545), .ZN(n5096) );
  INV_X1 U6527 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5101) );
  INV_X1 U6528 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5098) );
  INV_X1 U6529 ( .A(n5103), .ZN(n5104) );
  NAND2_X2 U6530 ( .A1(n8435), .A2(n5104), .ZN(n5265) );
  NAND2_X1 U6531 ( .A1(n8544), .A2(n5589), .ZN(n5110) );
  INV_X1 U6532 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n6491) );
  NAND2_X1 U6533 ( .A1(n5603), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5107) );
  NAND2_X1 U6534 ( .A1(n5604), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5106) );
  OAI211_X1 U6535 ( .C1(n5629), .C2(n6491), .A(n5107), .B(n5106), .ZN(n5108)
         );
  INV_X1 U6536 ( .A(n5108), .ZN(n5109) );
  NAND2_X1 U6537 ( .A1(n5110), .A2(n5109), .ZN(n8643) );
  NAND2_X1 U6538 ( .A1(n8366), .A2(n8643), .ZN(n5553) );
  NAND2_X1 U6539 ( .A1(n8906), .A2(n8644), .ZN(n8681) );
  NAND2_X1 U6540 ( .A1(n8254), .A2(n5623), .ZN(n5114) );
  OR2_X1 U6541 ( .A1(n4397), .A2(n7649), .ZN(n5113) );
  OAI21_X1 U6542 ( .B1(n5525), .B2(n8512), .A(n8501), .ZN(n5115) );
  AND2_X1 U6543 ( .A1(n5116), .A2(n5115), .ZN(n8710) );
  NAND2_X1 U6544 ( .A1(n8710), .A2(n5589), .ZN(n5122) );
  INV_X1 U6545 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n5119) );
  NAND2_X1 U6546 ( .A1(n5604), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5118) );
  NAND2_X1 U6547 ( .A1(n5241), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5117) );
  OAI211_X1 U6548 ( .C1(n5628), .C2(n5119), .A(n5118), .B(n5117), .ZN(n5120)
         );
  INV_X1 U6549 ( .A(n5120), .ZN(n5121) );
  NAND2_X1 U6550 ( .A1(n8910), .A2(n8696), .ZN(n5534) );
  INV_X1 U6551 ( .A(n5534), .ZN(n5123) );
  NOR2_X1 U6552 ( .A1(n8694), .A2(n5123), .ZN(n5540) );
  INV_X1 U6553 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5127) );
  NAND2_X1 U6554 ( .A1(n5131), .A2(n5127), .ZN(n5128) );
  XNOR2_X1 U6555 ( .A(n5640), .B(P2_IR_REG_19__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U6556 ( .A1(n5134), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5133) );
  INV_X1 U6557 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5132) );
  NOR2_X1 U6558 ( .A1(n6980), .A2(n7160), .ZN(n5850) );
  INV_X1 U6559 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U6560 ( .A1(n5850), .A2(n8108), .ZN(n5637) );
  XNOR2_X1 U6561 ( .A(n5136), .B(n5135), .ZN(n8222) );
  NAND2_X1 U6562 ( .A1(n8222), .A2(n5623), .ZN(n5138) );
  OR2_X1 U6563 ( .A1(n4397), .A2(n7302), .ZN(n5137) );
  NAND2_X1 U6564 ( .A1(n5505), .A2(n8453), .ZN(n5139) );
  NAND2_X1 U6565 ( .A1(n5525), .A2(n5139), .ZN(n8741) );
  AOI22_X1 U6566 ( .A1(n5603), .A2(P2_REG1_REG_23__SCAN_IN), .B1(n5241), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6567 ( .A1(n5604), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5140) );
  OAI211_X1 U6568 ( .C1(n8741), .C2(n5265), .A(n5141), .B(n5140), .ZN(n8728)
         );
  INV_X1 U6569 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6714) );
  OR2_X1 U6570 ( .A1(n5628), .A2(n6714), .ZN(n5145) );
  OAI21_X1 U6571 ( .B1(n5153), .B2(P2_REG3_REG_5__SCAN_IN), .A(n5183), .ZN(
        n7657) );
  OR2_X1 U6572 ( .A1(n5265), .A2(n7657), .ZN(n5144) );
  INV_X1 U6573 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5142) );
  NOR2_X1 U6574 ( .A1(n5146), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5191) );
  OR2_X1 U6575 ( .A1(n5191), .A2(n8997), .ZN(n5147) );
  XNOR2_X1 U6576 ( .A(n5147), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6739) );
  INV_X1 U6577 ( .A(n6739), .ZN(n6840) );
  XNOR2_X1 U6578 ( .A(n5149), .B(n5148), .ZN(n6193) );
  OR2_X1 U6579 ( .A1(n5219), .A2(n6193), .ZN(n5151) );
  OR2_X1 U6580 ( .A1(n4397), .A2(n6408), .ZN(n5150) );
  OAI211_X1 U6581 ( .C1(n5210), .C2(n6840), .A(n5151), .B(n5150), .ZN(n7664)
         );
  NAND2_X1 U6582 ( .A1(n5241), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5161) );
  INV_X1 U6583 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6715) );
  OR2_X1 U6584 ( .A1(n5628), .A2(n6715), .ZN(n5160) );
  INV_X1 U6585 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5152) );
  OR2_X1 U6586 ( .A1(n5412), .A2(n5152), .ZN(n5159) );
  INV_X1 U6587 ( .A(n5153), .ZN(n5157) );
  INV_X1 U6588 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5155) );
  INV_X1 U6589 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U6590 ( .A1(n5155), .A2(n5154), .ZN(n5156) );
  NAND2_X1 U6591 ( .A1(n5157), .A2(n5156), .ZN(n7507) );
  OR2_X1 U6592 ( .A1(n5265), .A2(n7507), .ZN(n5158) );
  NAND4_X1 U6593 ( .A1(n5161), .A2(n5160), .A3(n5159), .A4(n5158), .ZN(n8565)
         );
  NAND2_X1 U6594 ( .A1(n5163), .A2(n5162), .ZN(n5165) );
  XNOR2_X1 U6595 ( .A(n5165), .B(n5164), .ZN(n6186) );
  OR2_X1 U6596 ( .A1(n5219), .A2(n6186), .ZN(n5169) );
  OR2_X1 U6597 ( .A1(n4397), .A2(n6187), .ZN(n5168) );
  NAND2_X1 U6598 ( .A1(n5146), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5166) );
  XNOR2_X1 U6599 ( .A(n5166), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6737) );
  INV_X1 U6600 ( .A(n6737), .ZN(n6804) );
  OR2_X1 U6601 ( .A1(n5210), .A2(n6804), .ZN(n5167) );
  AND3_X2 U6602 ( .A1(n5169), .A2(n5168), .A3(n5167), .ZN(n10162) );
  OR2_X1 U6603 ( .A1(n8565), .A2(n10162), .ZN(n5655) );
  NAND2_X1 U6604 ( .A1(n8565), .A2(n10162), .ZN(n7650) );
  NAND2_X1 U6605 ( .A1(n8564), .A2(n10169), .ZN(n5660) );
  AND2_X1 U6606 ( .A1(n7650), .A2(n5660), .ZN(n5682) );
  MUX2_X1 U6607 ( .A(n5170), .B(n5682), .S(n5637), .Z(n5236) );
  NAND2_X1 U6608 ( .A1(n5241), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5175) );
  INV_X1 U6609 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6716) );
  OR2_X1 U6610 ( .A1(n5628), .A2(n6716), .ZN(n5174) );
  INV_X1 U6611 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5171) );
  OR2_X1 U6612 ( .A1(n5412), .A2(n5171), .ZN(n5173) );
  OR2_X1 U6613 ( .A1(n5265), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5172) );
  XNOR2_X1 U6614 ( .A(n5177), .B(n5176), .ZN(n6194) );
  OR2_X1 U6615 ( .A1(n5219), .A2(n6194), .ZN(n5181) );
  INV_X1 U6616 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5179) );
  NAND2_X1 U6617 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4432), .ZN(n5178) );
  XNOR2_X1 U6618 ( .A(n5179), .B(n5178), .ZN(n6828) );
  OR2_X1 U6619 ( .A1(n5210), .A2(n6828), .ZN(n5180) );
  NAND2_X1 U6620 ( .A1(n7499), .A2(n5655), .ZN(n5197) );
  INV_X1 U6621 ( .A(n7405), .ZN(n7527) );
  NAND2_X1 U6622 ( .A1(n5241), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5189) );
  INV_X1 U6623 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6713) );
  OR2_X1 U6624 ( .A1(n5628), .A2(n6713), .ZN(n5188) );
  AND2_X1 U6625 ( .A1(n5183), .A2(n5182), .ZN(n5184) );
  OR2_X1 U6626 ( .A1(n5184), .A2(n5243), .ZN(n7537) );
  OR2_X1 U6627 ( .A1(n5265), .A2(n7537), .ZN(n5187) );
  INV_X1 U6628 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6629 ( .A1(n5191), .A2(n5190), .ZN(n5252) );
  NAND2_X1 U6630 ( .A1(n5252), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5192) );
  XNOR2_X1 U6631 ( .A(n5192), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6741) );
  INV_X1 U6632 ( .A(n6741), .ZN(n6816) );
  OR2_X1 U6633 ( .A1(n4397), .A2(n6192), .ZN(n5195) );
  OAI211_X1 U6634 ( .C1(n5210), .C2(n6816), .A(n5196), .B(n5195), .ZN(n7540)
         );
  AOI211_X1 U6635 ( .C1(n5236), .C2(n5197), .A(n7527), .B(n5683), .ZN(n5231)
         );
  NAND2_X1 U6636 ( .A1(n5241), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5202) );
  INV_X1 U6637 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10205) );
  OR2_X1 U6638 ( .A1(n5628), .A2(n10205), .ZN(n5201) );
  INV_X1 U6639 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5198) );
  OR2_X1 U6640 ( .A1(n5412), .A2(n5198), .ZN(n5200) );
  INV_X1 U6641 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7442) );
  OR2_X1 U6642 ( .A1(n5265), .A2(n7442), .ZN(n5199) );
  NAND2_X1 U6643 ( .A1(n6179), .A2(SI_0_), .ZN(n5203) );
  XNOR2_X1 U6644 ( .A(n5203), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9003) );
  MUX2_X1 U6645 ( .A(n10129), .B(n9003), .S(n5210), .Z(n10146) );
  OR2_X1 U6646 ( .A1(n5875), .A2(n7314), .ZN(n7320) );
  INV_X1 U6647 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7315) );
  OR2_X1 U6648 ( .A1(n5265), .A2(n7315), .ZN(n5207) );
  INV_X1 U6649 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6718) );
  OR2_X1 U6650 ( .A1(n5628), .A2(n6718), .ZN(n5206) );
  NAND2_X1 U6651 ( .A1(n5604), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5205) );
  INV_X1 U6652 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6467) );
  NAND4_X1 U6653 ( .A1(n5207), .A2(n5206), .A3(n5205), .A4(n5204), .ZN(n5872)
         );
  INV_X1 U6654 ( .A(n5872), .ZN(n5212) );
  INV_X1 U6655 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6182) );
  XNOR2_X1 U6656 ( .A(n5209), .B(n5208), .ZN(n6180) );
  INV_X1 U6657 ( .A(n9803), .ZN(n6181) );
  OR2_X1 U6658 ( .A1(n5210), .A2(n6181), .ZN(n5211) );
  NAND2_X1 U6659 ( .A1(n5212), .A2(n4637), .ZN(n5657) );
  INV_X1 U6660 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7427) );
  OR2_X1 U6661 ( .A1(n5265), .A2(n7427), .ZN(n5216) );
  NAND2_X1 U6662 ( .A1(n5604), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5215) );
  INV_X1 U6663 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6717) );
  OR2_X1 U6664 ( .A1(n5628), .A2(n6717), .ZN(n5213) );
  XNOR2_X1 U6665 ( .A(n5218), .B(n5217), .ZN(n6189) );
  OR2_X1 U6666 ( .A1(n5220), .A2(n8997), .ZN(n5221) );
  XNOR2_X1 U6667 ( .A(n5221), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9814) );
  INV_X1 U6668 ( .A(n9814), .ZN(n6188) );
  OR2_X1 U6669 ( .A1(n5210), .A2(n6188), .ZN(n5222) );
  NAND2_X1 U6670 ( .A1(n8568), .A2(n10156), .ZN(n5654) );
  NAND3_X1 U6671 ( .A1(n5678), .A2(n5656), .A3(n5654), .ZN(n5224) );
  NAND2_X1 U6672 ( .A1(n5875), .A2(n7314), .ZN(n7176) );
  NAND4_X1 U6673 ( .A1(n5654), .A2(n5656), .A3(n7176), .A4(n5762), .ZN(n5223)
         );
  NAND3_X1 U6674 ( .A1(n5224), .A2(n5679), .A3(n5223), .ZN(n5228) );
  NAND2_X1 U6675 ( .A1(n5656), .A2(n7176), .ZN(n5225) );
  NAND3_X1 U6676 ( .A1(n5225), .A2(n5679), .A3(n5657), .ZN(n5226) );
  NAND2_X1 U6677 ( .A1(n5226), .A2(n5654), .ZN(n5227) );
  MUX2_X1 U6678 ( .A(n5228), .B(n5227), .S(n5294), .Z(n5229) );
  NAND2_X1 U6679 ( .A1(n8566), .A2(n7004), .ZN(n5233) );
  NAND3_X1 U6680 ( .A1(n5229), .A2(n7006), .A3(n5236), .ZN(n5230) );
  OAI21_X1 U6681 ( .B1(n5231), .B2(n5294), .A(n5230), .ZN(n5232) );
  NAND2_X1 U6682 ( .A1(n8563), .A2(n10172), .ZN(n5659) );
  NAND2_X1 U6683 ( .A1(n5232), .A2(n5659), .ZN(n5240) );
  INV_X1 U6684 ( .A(n5660), .ZN(n5235) );
  NAND2_X1 U6685 ( .A1(n5682), .A2(n5233), .ZN(n5234) );
  OAI21_X1 U6686 ( .B1(n5236), .B2(n5235), .A(n5234), .ZN(n5237) );
  NAND2_X1 U6687 ( .A1(n5237), .A2(n5659), .ZN(n5238) );
  NAND2_X1 U6688 ( .A1(n5238), .A2(n5294), .ZN(n5239) );
  NAND2_X1 U6689 ( .A1(n5240), .A2(n5239), .ZN(n5260) );
  NOR2_X1 U6690 ( .A1(n7407), .A2(n5637), .ZN(n5258) );
  NAND2_X1 U6691 ( .A1(n5241), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5249) );
  INV_X1 U6692 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6712) );
  OR2_X1 U6693 ( .A1(n5628), .A2(n6712), .ZN(n5248) );
  INV_X1 U6694 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5242) );
  OR2_X1 U6695 ( .A1(n5412), .A2(n5242), .ZN(n5247) );
  INV_X1 U6696 ( .A(n5243), .ZN(n5244) );
  INV_X1 U6697 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7231) );
  NAND2_X1 U6698 ( .A1(n5244), .A2(n7231), .ZN(n5245) );
  NAND2_X1 U6699 ( .A1(n5263), .A2(n5245), .ZN(n7467) );
  OR2_X1 U6700 ( .A1(n5265), .A2(n7467), .ZN(n5246) );
  NAND4_X1 U6701 ( .A1(n5249), .A2(n5248), .A3(n5247), .A4(n5246), .ZN(n5902)
         );
  XNOR2_X1 U6702 ( .A(n5251), .B(n5250), .ZN(n6196) );
  NAND2_X1 U6703 ( .A1(n6196), .A2(n5623), .ZN(n5257) );
  OAI21_X1 U6704 ( .B1(n5252), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5253) );
  XNOR2_X1 U6705 ( .A(n5254), .B(n5253), .ZN(n6852) );
  OR2_X1 U6706 ( .A1(n5210), .A2(n6852), .ZN(n5256) );
  INV_X1 U6707 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6513) );
  OR2_X1 U6708 ( .A1(n4397), .A2(n6513), .ZN(n5255) );
  OR2_X1 U6709 ( .A1(n5902), .A2(n7468), .ZN(n5316) );
  NAND2_X1 U6710 ( .A1(n5902), .A2(n7468), .ZN(n5688) );
  NAND2_X1 U6711 ( .A1(n5316), .A2(n5688), .ZN(n7404) );
  NOR2_X1 U6712 ( .A1(n5258), .A2(n7404), .ZN(n5259) );
  NAND2_X1 U6713 ( .A1(n5260), .A2(n5259), .ZN(n5319) );
  INV_X1 U6714 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n5261) );
  INV_X1 U6715 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6711) );
  OR2_X1 U6716 ( .A1(n5628), .A2(n6711), .ZN(n5269) );
  NAND2_X1 U6717 ( .A1(n5263), .A2(n5262), .ZN(n5264) );
  NAND2_X1 U6718 ( .A1(n5287), .A2(n5264), .ZN(n7244) );
  OR2_X1 U6719 ( .A1(n5265), .A2(n7244), .ZN(n5268) );
  INV_X1 U6720 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5266) );
  OR2_X1 U6721 ( .A1(n5412), .A2(n5266), .ZN(n5267) );
  NAND4_X1 U6722 ( .A1(n5270), .A2(n5269), .A3(n5268), .A4(n5267), .ZN(n8562)
         );
  XNOR2_X1 U6723 ( .A(n5272), .B(n5271), .ZN(n6202) );
  NAND2_X1 U6724 ( .A1(n6202), .A2(n5623), .ZN(n5279) );
  OR2_X1 U6725 ( .A1(n5273), .A2(n8997), .ZN(n5275) );
  MUX2_X1 U6726 ( .A(n5275), .B(P2_IR_REG_31__SCAN_IN), .S(n5274), .Z(n5277)
         );
  NAND2_X1 U6727 ( .A1(n5277), .A2(n5276), .ZN(n6863) );
  INV_X1 U6728 ( .A(n6863), .ZN(n6725) );
  AOI22_X1 U6729 ( .A1(n5459), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6592), .B2(
        n6725), .ZN(n5278) );
  AND2_X2 U6730 ( .A1(n5279), .A2(n5278), .ZN(n10179) );
  OR2_X2 U6731 ( .A1(n8562), .A2(n10179), .ZN(n5692) );
  NAND2_X1 U6732 ( .A1(n8562), .A2(n10179), .ZN(n5295) );
  NAND2_X2 U6733 ( .A1(n5692), .A2(n5295), .ZN(n5822) );
  INV_X1 U6734 ( .A(n5688), .ZN(n5685) );
  NOR2_X1 U6735 ( .A1(n5822), .A2(n5685), .ZN(n5281) );
  INV_X1 U6736 ( .A(n5692), .ZN(n5280) );
  AOI21_X1 U6737 ( .B1(n5319), .B2(n5281), .A(n5280), .ZN(n5298) );
  XNOR2_X1 U6738 ( .A(n5282), .B(n4951), .ZN(n7180) );
  NAND2_X1 U6739 ( .A1(n7180), .A2(n5623), .ZN(n5285) );
  NAND2_X1 U6740 ( .A1(n5276), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5283) );
  XNOR2_X1 U6741 ( .A(n5283), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6759) );
  AOI22_X1 U6742 ( .A1(n5459), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6592), .B2(
        n6759), .ZN(n5284) );
  NAND2_X1 U6743 ( .A1(n5603), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5293) );
  INV_X1 U6744 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6732) );
  OR2_X1 U6745 ( .A1(n5629), .A2(n6732), .ZN(n5292) );
  INV_X1 U6746 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6747 ( .A1(n5287), .A2(n5286), .ZN(n5288) );
  NAND2_X1 U6748 ( .A1(n5305), .A2(n5288), .ZN(n7372) );
  OR2_X1 U6749 ( .A1(n5265), .A2(n7372), .ZN(n5291) );
  INV_X1 U6750 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6751 ( .A1(n7598), .A2(n7993), .ZN(n5694) );
  XNOR2_X1 U6752 ( .A(n5299), .B(n4946), .ZN(n7185) );
  NAND2_X1 U6753 ( .A1(n7185), .A2(n5623), .ZN(n5303) );
  NAND2_X1 U6754 ( .A1(n5300), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5301) );
  XNOR2_X1 U6755 ( .A(n5301), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6935) );
  AOI22_X1 U6756 ( .A1(n5459), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6592), .B2(
        n6935), .ZN(n5302) );
  NAND2_X1 U6757 ( .A1(n5603), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5311) );
  INV_X1 U6758 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7998) );
  OR2_X1 U6759 ( .A1(n5629), .A2(n7998), .ZN(n5310) );
  NAND2_X1 U6760 ( .A1(n5305), .A2(n5304), .ZN(n5306) );
  NAND2_X1 U6761 ( .A1(n5329), .A2(n5306), .ZN(n7997) );
  OR2_X1 U6762 ( .A1(n5265), .A2(n7997), .ZN(n5309) );
  INV_X1 U6763 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5307) );
  OR2_X1 U6764 ( .A1(n5412), .A2(n5307), .ZN(n5308) );
  OR2_X1 U6765 ( .A1(n10185), .A2(n7397), .ZN(n5696) );
  OR2_X1 U6766 ( .A1(n7598), .A2(n7993), .ZN(n5693) );
  AND2_X1 U6767 ( .A1(n5696), .A2(n5693), .ZN(n5314) );
  NAND2_X1 U6768 ( .A1(n10185), .A2(n7397), .ZN(n5695) );
  NAND2_X1 U6769 ( .A1(n5695), .A2(n5694), .ZN(n5312) );
  NAND2_X1 U6770 ( .A1(n5312), .A2(n5637), .ZN(n5313) );
  AND2_X1 U6771 ( .A1(n5314), .A2(n5313), .ZN(n5318) );
  NAND2_X1 U6772 ( .A1(n5315), .A2(n5318), .ZN(n5339) );
  INV_X1 U6773 ( .A(n5822), .ZN(n5317) );
  NAND4_X1 U6774 ( .A1(n5319), .A2(n5318), .A3(n5317), .A4(n5316), .ZN(n5336)
         );
  NAND2_X1 U6775 ( .A1(n5321), .A2(n5320), .ZN(n5323) );
  XNOR2_X1 U6776 ( .A(n5323), .B(n5322), .ZN(n7277) );
  NAND2_X1 U6777 ( .A1(n7277), .A2(n5623), .ZN(n5327) );
  NAND2_X1 U6778 ( .A1(n5324), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5325) );
  XNOR2_X1 U6779 ( .A(n5325), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8575) );
  AOI22_X1 U6780 ( .A1(n5459), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6592), .B2(
        n8575), .ZN(n5326) );
  NAND2_X1 U6781 ( .A1(n5241), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5334) );
  INV_X1 U6782 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5328) );
  OR2_X1 U6783 ( .A1(n5412), .A2(n5328), .ZN(n5333) );
  INV_X1 U6784 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U6785 ( .A1(n5329), .A2(n8573), .ZN(n5330) );
  NAND2_X1 U6786 ( .A1(n5346), .A2(n5330), .ZN(n7731) );
  OR2_X1 U6787 ( .A1(n5265), .A2(n7731), .ZN(n5332) );
  INV_X1 U6788 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6925) );
  OR2_X1 U6789 ( .A1(n5628), .A2(n6925), .ZN(n5331) );
  OR2_X1 U6790 ( .A1(n7730), .A2(n7992), .ZN(n7606) );
  NAND2_X1 U6791 ( .A1(n5695), .A2(n4865), .ZN(n5335) );
  NAND4_X1 U6792 ( .A1(n5336), .A2(n5696), .A3(n7606), .A4(n5335), .ZN(n5337)
         );
  NAND2_X1 U6793 ( .A1(n5337), .A2(n5637), .ZN(n5338) );
  NAND2_X1 U6794 ( .A1(n5339), .A2(n5338), .ZN(n5353) );
  XNOR2_X1 U6795 ( .A(n5341), .B(n5340), .ZN(n7549) );
  NAND2_X1 U6796 ( .A1(n7549), .A2(n5623), .ZN(n5344) );
  OR2_X1 U6797 ( .A1(n5342), .A2(n8997), .ZN(n5361) );
  XNOR2_X1 U6798 ( .A(n5361), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7102) );
  AOI22_X1 U6799 ( .A1(n5459), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6592), .B2(
        n7102), .ZN(n5343) );
  NAND2_X1 U6800 ( .A1(n5604), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5351) );
  INV_X1 U6801 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6924) );
  OR2_X1 U6802 ( .A1(n5628), .A2(n6924), .ZN(n5350) );
  INV_X1 U6803 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7612) );
  OR2_X1 U6804 ( .A1(n5629), .A2(n7612), .ZN(n5349) );
  NAND2_X1 U6805 ( .A1(n5346), .A2(n5345), .ZN(n5347) );
  NAND2_X1 U6806 ( .A1(n5367), .A2(n5347), .ZN(n7631) );
  OR2_X1 U6807 ( .A1(n5265), .A2(n7631), .ZN(n5348) );
  NAND2_X1 U6808 ( .A1(n10193), .A2(n7683), .ZN(n5700) );
  NAND2_X1 U6809 ( .A1(n7730), .A2(n7992), .ZN(n5698) );
  OR2_X1 U6810 ( .A1(n10193), .A2(n7683), .ZN(n5663) );
  NAND2_X1 U6811 ( .A1(n5698), .A2(n5695), .ZN(n5352) );
  AND2_X1 U6812 ( .A1(n5663), .A2(n7606), .ZN(n5699) );
  NAND2_X1 U6813 ( .A1(n5355), .A2(n5354), .ZN(n5359) );
  AND2_X1 U6814 ( .A1(n5357), .A2(n5356), .ZN(n5358) );
  XNOR2_X1 U6815 ( .A(n5359), .B(n5358), .ZN(n7555) );
  NAND2_X1 U6816 ( .A1(n7555), .A2(n5623), .ZN(n5365) );
  INV_X1 U6817 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U6818 ( .A1(n5361), .A2(n5360), .ZN(n5362) );
  NAND2_X1 U6819 ( .A1(n5362), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5363) );
  XNOR2_X1 U6820 ( .A(n5363), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7220) );
  AOI22_X1 U6821 ( .A1(n5459), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6592), .B2(
        n7220), .ZN(n5364) );
  NAND2_X1 U6822 ( .A1(n5604), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5372) );
  INV_X1 U6823 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5366) );
  OR2_X1 U6824 ( .A1(n5628), .A2(n5366), .ZN(n5371) );
  INV_X1 U6825 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7693) );
  OR2_X1 U6826 ( .A1(n5629), .A2(n7693), .ZN(n5370) );
  NAND2_X1 U6827 ( .A1(n5367), .A2(n7107), .ZN(n5368) );
  NAND2_X1 U6828 ( .A1(n5380), .A2(n5368), .ZN(n7692) );
  OR2_X1 U6829 ( .A1(n5265), .A2(n7692), .ZN(n5369) );
  OR2_X1 U6830 ( .A1(n8972), .A2(n7883), .ZN(n5386) );
  NAND2_X1 U6831 ( .A1(n8972), .A2(n7883), .ZN(n5702) );
  XNOR2_X1 U6832 ( .A(n5374), .B(n5373), .ZN(n7567) );
  NAND2_X1 U6833 ( .A1(n7567), .A2(n5623), .ZN(n5378) );
  OR2_X1 U6834 ( .A1(n5375), .A2(n8997), .ZN(n5376) );
  XNOR2_X1 U6835 ( .A(n5376), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7330) );
  AOI22_X1 U6836 ( .A1(n5459), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6592), .B2(
        n7330), .ZN(n5377) );
  NAND2_X1 U6837 ( .A1(n5604), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5385) );
  INV_X1 U6838 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7216) );
  OR2_X1 U6839 ( .A1(n5628), .A2(n7216), .ZN(n5384) );
  INV_X1 U6840 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7328) );
  OR2_X1 U6841 ( .A1(n5629), .A2(n7328), .ZN(n5383) );
  INV_X1 U6842 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6843 ( .A1(n5380), .A2(n5379), .ZN(n5381) );
  NAND2_X1 U6844 ( .A1(n5397), .A2(n5381), .ZN(n7877) );
  OR2_X1 U6845 ( .A1(n5265), .A2(n7877), .ZN(n5382) );
  NAND2_X1 U6846 ( .A1(n8967), .A2(n7898), .ZN(n5404) );
  MUX2_X1 U6847 ( .A(n5702), .B(n5386), .S(n5637), .Z(n5387) );
  NAND2_X1 U6848 ( .A1(n5389), .A2(n5388), .ZN(n5406) );
  XNOR2_X1 U6849 ( .A(n5391), .B(n5390), .ZN(n7748) );
  NAND2_X1 U6850 ( .A1(n7748), .A2(n5623), .ZN(n5395) );
  NAND2_X1 U6851 ( .A1(n5392), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5393) );
  XNOR2_X1 U6852 ( .A(n5393), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8053) );
  AOI22_X1 U6853 ( .A1(n5459), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6592), .B2(
        n8053), .ZN(n5394) );
  NAND2_X1 U6854 ( .A1(n5603), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5403) );
  INV_X1 U6855 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7865) );
  OR2_X1 U6856 ( .A1(n5629), .A2(n7865), .ZN(n5402) );
  INV_X1 U6857 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U6858 ( .A1(n5397), .A2(n5396), .ZN(n5398) );
  NAND2_X1 U6859 ( .A1(n5429), .A2(n5398), .ZN(n7897) );
  OR2_X1 U6860 ( .A1(n5265), .A2(n7897), .ZN(n5401) );
  INV_X1 U6861 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n5399) );
  OR2_X1 U6862 ( .A1(n5412), .A2(n5399), .ZN(n5400) );
  XNOR2_X1 U6863 ( .A(n8962), .B(n8854), .ZN(n7870) );
  INV_X1 U6864 ( .A(n7870), .ZN(n5704) );
  MUX2_X1 U6865 ( .A(n5703), .B(n5404), .S(n5637), .Z(n5405) );
  NAND3_X1 U6866 ( .A1(n5406), .A2(n5704), .A3(n5405), .ZN(n5419) );
  XNOR2_X1 U6867 ( .A(n5408), .B(n5407), .ZN(n7829) );
  NAND2_X1 U6868 ( .A1(n7829), .A2(n5623), .ZN(n5411) );
  NAND2_X1 U6869 ( .A1(n5409), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5423) );
  XNOR2_X1 U6870 ( .A(n5423), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8594) );
  AOI22_X1 U6871 ( .A1(n5459), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6592), .B2(
        n8594), .ZN(n5410) );
  NAND2_X1 U6872 ( .A1(n5241), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5416) );
  INV_X1 U6873 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8066) );
  OR2_X1 U6874 ( .A1(n5628), .A2(n8066), .ZN(n5415) );
  INV_X1 U6875 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5428) );
  XNOR2_X1 U6876 ( .A(n5429), .B(n5428), .ZN(n8867) );
  OR2_X1 U6877 ( .A1(n5265), .A2(n8867), .ZN(n5414) );
  INV_X1 U6878 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n6478) );
  OR2_X1 U6879 ( .A1(n5412), .A2(n6478), .ZN(n5413) );
  NAND2_X1 U6880 ( .A1(n8956), .A2(n7952), .ZN(n5707) );
  INV_X1 U6881 ( .A(n8962), .ZN(n7903) );
  INV_X1 U6882 ( .A(n8854), .ZN(n8627) );
  MUX2_X1 U6883 ( .A(n8962), .B(n8627), .S(n5637), .Z(n5417) );
  OAI21_X1 U6884 ( .B1(n7903), .B2(n8854), .A(n5417), .ZN(n5418) );
  NAND3_X1 U6885 ( .A1(n5419), .A2(n8855), .A3(n5418), .ZN(n5437) );
  XNOR2_X1 U6886 ( .A(n5421), .B(n5420), .ZN(n7904) );
  NAND2_X1 U6887 ( .A1(n7904), .A2(n5623), .ZN(n5427) );
  INV_X1 U6888 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U6889 ( .A1(n5423), .A2(n5422), .ZN(n5424) );
  NAND2_X1 U6890 ( .A1(n5424), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5425) );
  XNOR2_X1 U6891 ( .A(n5425), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8055) );
  AOI22_X1 U6892 ( .A1(n5459), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6592), .B2(
        n8055), .ZN(n5426) );
  NAND2_X1 U6893 ( .A1(n5241), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5435) );
  INV_X1 U6894 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8068) );
  OR2_X1 U6895 ( .A1(n5628), .A2(n8068), .ZN(n5434) );
  INV_X1 U6896 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7955) );
  OAI21_X1 U6897 ( .B1(n5429), .B2(n5428), .A(n7955), .ZN(n5430) );
  NAND2_X1 U6898 ( .A1(n5430), .A2(n5445), .ZN(n8836) );
  OR2_X1 U6899 ( .A1(n5265), .A2(n8836), .ZN(n5433) );
  INV_X1 U6900 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n5431) );
  OR2_X1 U6901 ( .A1(n5412), .A2(n5431), .ZN(n5432) );
  XNOR2_X1 U6902 ( .A(n8953), .B(n8852), .ZN(n8828) );
  INV_X1 U6903 ( .A(n8828), .ZN(n8842) );
  MUX2_X1 U6904 ( .A(n5706), .B(n5707), .S(n5637), .Z(n5436) );
  NAND3_X1 U6905 ( .A1(n5437), .A2(n8842), .A3(n5436), .ZN(n5455) );
  OR2_X1 U6906 ( .A1(n8953), .A2(n8852), .ZN(n5709) );
  INV_X1 U6907 ( .A(n5709), .ZN(n5452) );
  INV_X1 U6908 ( .A(n8953), .ZN(n8834) );
  INV_X1 U6909 ( .A(n8852), .ZN(n8820) );
  XNOR2_X1 U6910 ( .A(n5439), .B(n5438), .ZN(n8006) );
  NAND2_X1 U6911 ( .A1(n8006), .A2(n5623), .ZN(n5443) );
  NAND2_X1 U6912 ( .A1(n5440), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5441) );
  XNOR2_X1 U6913 ( .A(n5441), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8059) );
  AOI22_X1 U6914 ( .A1(n5459), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6592), .B2(
        n8059), .ZN(n5442) );
  NAND2_X1 U6915 ( .A1(n5603), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5450) );
  INV_X1 U6916 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5444) );
  OR2_X1 U6917 ( .A1(n5629), .A2(n5444), .ZN(n5449) );
  INV_X1 U6918 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8536) );
  NAND2_X1 U6919 ( .A1(n5445), .A2(n8536), .ZN(n5446) );
  NAND2_X1 U6920 ( .A1(n5463), .A2(n5446), .ZN(n8535) );
  OR2_X1 U6921 ( .A1(n5265), .A2(n8535), .ZN(n5448) );
  INV_X1 U6922 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n6510) );
  OR2_X1 U6923 ( .A1(n5412), .A2(n6510), .ZN(n5447) );
  NAND4_X1 U6924 ( .A1(n5450), .A2(n5449), .A3(n5448), .A4(n5447), .ZN(n8805)
         );
  INV_X1 U6925 ( .A(n8805), .ZN(n8632) );
  NAND2_X1 U6926 ( .A1(n8946), .A2(n8632), .ZN(n5710) );
  OAI21_X1 U6927 ( .B1(n8834), .B2(n8820), .A(n5710), .ZN(n5451) );
  MUX2_X1 U6928 ( .A(n5452), .B(n5451), .S(n5294), .Z(n5453) );
  NOR2_X1 U6929 ( .A1(n5453), .A2(n5711), .ZN(n5454) );
  NAND2_X1 U6930 ( .A1(n5455), .A2(n5454), .ZN(n5512) );
  NAND2_X1 U6931 ( .A1(n5512), .A2(n5710), .ZN(n5469) );
  XNOR2_X1 U6932 ( .A(n5457), .B(n5456), .ZN(n8148) );
  NAND2_X1 U6933 ( .A1(n8148), .A2(n5623), .ZN(n5461) );
  AOI22_X1 U6934 ( .A1(n5459), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5458), .B2(
        n6592), .ZN(n5460) );
  NAND2_X1 U6935 ( .A1(n5604), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5468) );
  INV_X1 U6936 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8070) );
  OR2_X1 U6937 ( .A1(n5628), .A2(n8070), .ZN(n5467) );
  INV_X1 U6938 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5462) );
  OR2_X1 U6939 ( .A1(n5629), .A2(n5462), .ZN(n5466) );
  NAND2_X1 U6940 ( .A1(n5463), .A2(n8464), .ZN(n5464) );
  NAND2_X1 U6941 ( .A1(n5481), .A2(n5464), .ZN(n8800) );
  OR2_X1 U6942 ( .A1(n5265), .A2(n8800), .ZN(n5465) );
  NAND4_X1 U6943 ( .A1(n5468), .A2(n5467), .A3(n5466), .A4(n5465), .ZN(n8822)
         );
  INV_X1 U6944 ( .A(n8822), .ZN(n8636) );
  OR2_X1 U6945 ( .A1(n8942), .A2(n8636), .ZN(n5652) );
  NAND2_X1 U6946 ( .A1(n5469), .A2(n5652), .ZN(n5487) );
  NAND2_X1 U6947 ( .A1(n5471), .A2(n5470), .ZN(n5475) );
  AND2_X1 U6948 ( .A1(n5473), .A2(n5472), .ZN(n5474) );
  NAND2_X1 U6949 ( .A1(n8168), .A2(n5623), .ZN(n5477) );
  OR2_X1 U6950 ( .A1(n4397), .A2(n7960), .ZN(n5476) );
  NAND2_X2 U6951 ( .A1(n5477), .A2(n5476), .ZN(n8936) );
  NAND2_X1 U6952 ( .A1(n5604), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5486) );
  INV_X1 U6953 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n5478) );
  OR2_X1 U6954 ( .A1(n5628), .A2(n5478), .ZN(n5485) );
  INV_X1 U6955 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5479) );
  OR2_X1 U6956 ( .A1(n5629), .A2(n5479), .ZN(n5484) );
  INV_X1 U6957 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U6958 ( .A1(n5481), .A2(n5480), .ZN(n5482) );
  NAND2_X1 U6959 ( .A1(n5504), .A2(n5482), .ZN(n8521) );
  OR2_X1 U6960 ( .A1(n5265), .A2(n8521), .ZN(n5483) );
  NAND2_X1 U6961 ( .A1(n8936), .A2(n8487), .ZN(n5651) );
  NAND2_X1 U6962 ( .A1(n8942), .A2(n8636), .ZN(n8790) );
  NAND3_X1 U6963 ( .A1(n5487), .A2(n5651), .A3(n8790), .ZN(n5497) );
  XNOR2_X1 U6964 ( .A(n5489), .B(n5488), .ZN(n8189) );
  NAND2_X1 U6965 ( .A1(n8189), .A2(n5623), .ZN(n5491) );
  OR2_X1 U6966 ( .A1(n4397), .A2(n7159), .ZN(n5490) );
  XNOR2_X1 U6967 ( .A(n5504), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n8771) );
  NAND2_X1 U6968 ( .A1(n8771), .A2(n5589), .ZN(n5495) );
  NAND2_X1 U6969 ( .A1(n5603), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U6970 ( .A1(n5241), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U6971 ( .A1(n5604), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5492) );
  OR2_X1 U6972 ( .A1(n8931), .A2(n8762), .ZN(n5650) );
  OR2_X2 U6973 ( .A1(n8936), .A2(n8487), .ZN(n5714) );
  NAND2_X1 U6974 ( .A1(n5497), .A2(n5496), .ZN(n5510) );
  NAND2_X1 U6975 ( .A1(n8931), .A2(n8762), .ZN(n8758) );
  XNOR2_X1 U6976 ( .A(n5499), .B(n5498), .ZN(n8208) );
  NAND2_X1 U6977 ( .A1(n8208), .A2(n5623), .ZN(n5501) );
  OR2_X1 U6978 ( .A1(n4397), .A2(n8111), .ZN(n5500) );
  NAND2_X1 U6979 ( .A1(n5603), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U6980 ( .A1(n5241), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5502) );
  AND2_X1 U6981 ( .A1(n5503), .A2(n5502), .ZN(n5509) );
  INV_X1 U6982 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8486) );
  INV_X1 U6983 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8100) );
  OAI21_X1 U6984 ( .B1(n5504), .B2(n8486), .A(n8100), .ZN(n5506) );
  NAND2_X1 U6985 ( .A1(n5506), .A2(n5505), .ZN(n8752) );
  OR2_X1 U6986 ( .A1(n8752), .A2(n5265), .ZN(n5508) );
  NAND2_X1 U6987 ( .A1(n5604), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U6988 ( .A1(n8926), .A2(n8641), .ZN(n5648) );
  NAND3_X1 U6989 ( .A1(n5510), .A2(n8758), .A3(n5648), .ZN(n5518) );
  INV_X1 U6990 ( .A(n5711), .ZN(n5511) );
  INV_X1 U6991 ( .A(n8790), .ZN(n5715) );
  AOI21_X1 U6992 ( .B1(n5512), .B2(n5511), .A(n5715), .ZN(n5514) );
  NAND2_X1 U6993 ( .A1(n5714), .A2(n5652), .ZN(n5513) );
  OAI211_X1 U6994 ( .C1(n5514), .C2(n5513), .A(n5651), .B(n8758), .ZN(n5515)
         );
  OR2_X1 U6995 ( .A1(n8921), .A2(n8763), .ZN(n5530) );
  INV_X1 U6996 ( .A(n8736), .ZN(n5516) );
  OAI21_X1 U6997 ( .B1(n5294), .B2(n5721), .A(n5519), .ZN(n5533) );
  INV_X1 U6998 ( .A(n5649), .ZN(n8732) );
  NAND2_X1 U6999 ( .A1(n5721), .A2(n8732), .ZN(n5520) );
  MUX2_X1 U7000 ( .A(n5648), .B(n5520), .S(n5637), .Z(n5532) );
  XNOR2_X1 U7001 ( .A(n5522), .B(n5521), .ZN(n8237) );
  NAND2_X1 U7002 ( .A1(n8237), .A2(n5623), .ZN(n5524) );
  OR2_X1 U7003 ( .A1(n4397), .A2(n7380), .ZN(n5523) );
  XNOR2_X1 U7004 ( .A(n5525), .B(P2_REG3_REG_24__SCAN_IN), .ZN(n8721) );
  INV_X1 U7005 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n5528) );
  NAND2_X1 U7006 ( .A1(n5603), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U7007 ( .A1(n5604), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5526) );
  OAI211_X1 U7008 ( .C1(n5629), .C2(n5528), .A(n5527), .B(n5526), .ZN(n5529)
         );
  NAND2_X1 U7009 ( .A1(n8914), .A2(n8642), .ZN(n5535) );
  NAND2_X1 U7010 ( .A1(n8725), .A2(n5530), .ZN(n5647) );
  NAND2_X1 U7011 ( .A1(n5535), .A2(n5637), .ZN(n5531) );
  AOI22_X1 U7012 ( .A1(n5533), .A2(n5532), .B1(n5647), .B2(n5531), .ZN(n5538)
         );
  MUX2_X1 U7013 ( .A(n5535), .B(n5722), .S(n5637), .Z(n5536) );
  NAND2_X1 U7014 ( .A1(n8714), .A2(n5536), .ZN(n5537) );
  INV_X1 U7015 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7776) );
  INV_X1 U7016 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8288) );
  MUX2_X1 U7017 ( .A(n7776), .B(n8288), .S(n4402), .Z(n5545) );
  INV_X1 U7018 ( .A(SI_27_), .ZN(n6522) );
  NAND2_X1 U7019 ( .A1(n5545), .A2(n6522), .ZN(n5558) );
  INV_X1 U7020 ( .A(n5545), .ZN(n5546) );
  NAND2_X1 U7021 ( .A1(n5546), .A2(SI_27_), .ZN(n5547) );
  AND2_X1 U7022 ( .A1(n5558), .A2(n5547), .ZN(n5557) );
  OR2_X1 U7023 ( .A1(n4397), .A2(n7776), .ZN(n5548) );
  XNOR2_X1 U7024 ( .A(n5562), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8679) );
  INV_X1 U7025 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6571) );
  NAND2_X1 U7026 ( .A1(n5241), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U7027 ( .A1(n5603), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5550) );
  OAI211_X1 U7028 ( .C1(n6571), .C2(n5412), .A(n5551), .B(n5550), .ZN(n5552)
         );
  NAND2_X1 U7029 ( .A1(n8899), .A2(n8697), .ZN(n5572) );
  INV_X1 U7030 ( .A(n8683), .ZN(n5555) );
  MUX2_X1 U7031 ( .A(n8681), .B(n5553), .S(n5637), .Z(n5554) );
  INV_X1 U7032 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8106) );
  INV_X1 U7033 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8304) );
  MUX2_X1 U7034 ( .A(n8106), .B(n8304), .S(n4402), .Z(n5578) );
  XNOR2_X1 U7035 ( .A(n5578), .B(SI_28_), .ZN(n5575) );
  OR2_X1 U7036 ( .A1(n4397), .A2(n8106), .ZN(n5559) );
  INV_X1 U7037 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8441) );
  INV_X1 U7038 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5561) );
  OAI21_X1 U7039 ( .B1(n5562), .B2(n8441), .A(n5561), .ZN(n5565) );
  INV_X1 U7040 ( .A(n5562), .ZN(n5564) );
  AND2_X1 U7041 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n5563) );
  NAND2_X1 U7042 ( .A1(n5564), .A2(n5563), .ZN(n5584) );
  NAND2_X1 U7043 ( .A1(n5565), .A2(n5584), .ZN(n8666) );
  OR2_X1 U7044 ( .A1(n8666), .A2(n5265), .ZN(n5571) );
  INV_X1 U7045 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U7046 ( .A1(n5604), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5567) );
  NAND2_X1 U7047 ( .A1(n5241), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5566) );
  OAI211_X1 U7048 ( .C1(n5628), .C2(n5568), .A(n5567), .B(n5566), .ZN(n5569)
         );
  INV_X1 U7049 ( .A(n5569), .ZN(n5570) );
  NAND2_X1 U7050 ( .A1(n8894), .A2(n8684), .ZN(n5646) );
  AND2_X1 U7051 ( .A1(n5646), .A2(n5572), .ZN(n5573) );
  INV_X1 U7052 ( .A(SI_28_), .ZN(n5577) );
  NAND2_X1 U7053 ( .A1(n5578), .A2(n5577), .ZN(n5579) );
  INV_X1 U7054 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8349) );
  INV_X1 U7055 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8408) );
  MUX2_X1 U7056 ( .A(n8349), .B(n8408), .S(n4402), .Z(n5596) );
  XNOR2_X1 U7057 ( .A(n5596), .B(SI_29_), .ZN(n5581) );
  NAND2_X1 U7058 ( .A1(n8407), .A2(n5623), .ZN(n5583) );
  OR2_X1 U7059 ( .A1(n4397), .A2(n8349), .ZN(n5582) );
  INV_X1 U7060 ( .A(n5584), .ZN(n8657) );
  INV_X1 U7061 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7062 ( .A1(n5241), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U7063 ( .A1(n5604), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5585) );
  OAI211_X1 U7064 ( .C1(n5628), .C2(n5587), .A(n5586), .B(n5585), .ZN(n5588)
         );
  AOI21_X1 U7065 ( .B1(n8657), .B2(n5589), .A(n5588), .ZN(n8555) );
  NAND2_X1 U7066 ( .A1(n8041), .A2(n8555), .ZN(n5732) );
  INV_X1 U7067 ( .A(n5732), .ZN(n5590) );
  NAND2_X1 U7068 ( .A1(n5591), .A2(n5732), .ZN(n5593) );
  INV_X1 U7069 ( .A(SI_29_), .ZN(n5595) );
  AND2_X1 U7070 ( .A1(n5596), .A2(n5595), .ZN(n5599) );
  INV_X1 U7071 ( .A(n5596), .ZN(n5597) );
  NAND2_X1 U7072 ( .A1(n5597), .A2(SI_29_), .ZN(n5598) );
  MUX2_X1 U7073 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n4402), .Z(n5616) );
  NAND2_X1 U7074 ( .A1(n9152), .A2(n5623), .ZN(n5602) );
  INV_X1 U7075 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8437) );
  OR2_X1 U7076 ( .A1(n4397), .A2(n8437), .ZN(n5601) );
  INV_X1 U7077 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U7078 ( .A1(n5603), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7079 ( .A1(n5604), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5605) );
  OAI211_X1 U7080 ( .C1(n5629), .C2(n5607), .A(n5606), .B(n5605), .ZN(n8650)
         );
  INV_X1 U7081 ( .A(n8650), .ZN(n5610) );
  NAND2_X1 U7082 ( .A1(n8623), .A2(n5610), .ZN(n5633) );
  NOR2_X1 U7083 ( .A1(n8623), .A2(n5610), .ZN(n5736) );
  INV_X1 U7084 ( .A(n5736), .ZN(n5636) );
  INV_X1 U7085 ( .A(n5614), .ZN(n5615) );
  NAND2_X1 U7086 ( .A1(n5615), .A2(SI_30_), .ZN(n5619) );
  NAND2_X1 U7087 ( .A1(n5617), .A2(n5616), .ZN(n5618) );
  NAND2_X1 U7088 ( .A1(n5619), .A2(n5618), .ZN(n5622) );
  MUX2_X1 U7089 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n4402), .Z(n5620) );
  XNOR2_X1 U7090 ( .A(n5620), .B(SI_31_), .ZN(n5621) );
  NAND2_X1 U7091 ( .A1(n9148), .A2(n5623), .ZN(n5627) );
  INV_X1 U7092 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5624) );
  OR2_X1 U7093 ( .A1(n4397), .A2(n5624), .ZN(n5626) );
  NAND2_X1 U7094 ( .A1(n5604), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5632) );
  INV_X1 U7095 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6429) );
  OR2_X1 U7096 ( .A1(n5628), .A2(n6429), .ZN(n5631) );
  INV_X1 U7097 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8043) );
  OR2_X1 U7098 ( .A1(n5629), .A2(n8043), .ZN(n5630) );
  AND3_X1 U7099 ( .A1(n5632), .A2(n5631), .A3(n5630), .ZN(n6611) );
  NAND2_X1 U7100 ( .A1(n5638), .A2(n5633), .ZN(n5738) );
  NAND2_X1 U7101 ( .A1(n5738), .A2(n5294), .ZN(n5635) );
  NAND2_X1 U7102 ( .A1(n8879), .A2(n6611), .ZN(n5737) );
  INV_X1 U7103 ( .A(n5737), .ZN(n5634) );
  NAND2_X1 U7104 ( .A1(n5737), .A2(n5636), .ZN(n5644) );
  NAND2_X1 U7105 ( .A1(n5640), .A2(n5639), .ZN(n5641) );
  INV_X1 U7106 ( .A(n5738), .ZN(n5674) );
  INV_X1 U7107 ( .A(n5644), .ZN(n5673) );
  INV_X1 U7108 ( .A(n5647), .ZN(n5670) );
  NAND2_X1 U7109 ( .A1(n5650), .A2(n8758), .ZN(n8769) );
  NAND2_X2 U7110 ( .A1(n5714), .A2(n5651), .ZN(n8792) );
  INV_X1 U7111 ( .A(n5710), .ZN(n5653) );
  NOR2_X1 U7112 ( .A1(n5711), .A2(n5653), .ZN(n8818) );
  NAND2_X1 U7113 ( .A1(n7320), .A2(n7176), .ZN(n10147) );
  INV_X1 U7114 ( .A(n10147), .ZN(n7446) );
  NAND3_X1 U7115 ( .A1(n7434), .A2(n7446), .A3(n5855), .ZN(n5658) );
  NAND2_X1 U7116 ( .A1(n5655), .A2(n7650), .ZN(n7497) );
  NOR4_X1 U7117 ( .A1(n5658), .A2(n7497), .A3(n5806), .A4(n6999), .ZN(n5661)
         );
  INV_X1 U7118 ( .A(n7404), .ZN(n7408) );
  NAND2_X1 U7119 ( .A1(n7407), .A2(n5659), .ZN(n7525) );
  INV_X1 U7120 ( .A(n7525), .ZN(n7528) );
  AND2_X1 U7121 ( .A1(n7405), .A2(n5660), .ZN(n7655) );
  NAND4_X1 U7122 ( .A1(n5661), .A2(n7408), .A3(n7528), .A4(n7655), .ZN(n5662)
         );
  AND2_X1 U7123 ( .A1(n5696), .A2(n5695), .ZN(n7990) );
  INV_X1 U7124 ( .A(n7990), .ZN(n7600) );
  NOR4_X1 U7125 ( .A1(n5662), .A2(n7600), .A3(n5822), .A4(n7362), .ZN(n5665)
         );
  NAND2_X1 U7126 ( .A1(n7606), .A2(n5698), .ZN(n7638) );
  INV_X1 U7127 ( .A(n7638), .ZN(n5664) );
  NAND4_X1 U7128 ( .A1(n7686), .A2(n5665), .A3(n7684), .A4(n5664), .ZN(n5666)
         );
  NOR4_X1 U7129 ( .A1(n4850), .A2(n7870), .A3(n7881), .A4(n5666), .ZN(n5667)
         );
  NAND4_X1 U7130 ( .A1(n8804), .A2(n8818), .A3(n5667), .A4(n8842), .ZN(n5668)
         );
  NOR4_X1 U7131 ( .A1(n8761), .A2(n8769), .A3(n8792), .A4(n5668), .ZN(n5669)
         );
  NAND4_X1 U7132 ( .A1(n8714), .A2(n5670), .A3(n5669), .A4(n5721), .ZN(n5671)
         );
  NOR4_X1 U7133 ( .A1(n8669), .A2(n8683), .A3(n8694), .A4(n5671), .ZN(n5672)
         );
  NAND4_X1 U7134 ( .A1(n5674), .A2(n5673), .A3(n8647), .A4(n5672), .ZN(n5675)
         );
  XNOR2_X1 U7135 ( .A(n5675), .B(n6980), .ZN(n5676) );
  NAND2_X1 U7136 ( .A1(n6998), .A2(n5458), .ZN(n5826) );
  OAI22_X1 U7137 ( .A1(n5676), .A2(n5762), .B1(n5855), .B2(n5826), .ZN(n5748)
         );
  INV_X1 U7138 ( .A(n5826), .ZN(n5677) );
  NAND2_X1 U7139 ( .A1(n7005), .A2(n7006), .ZN(n7500) );
  INV_X1 U7140 ( .A(n7499), .ZN(n5680) );
  NOR2_X1 U7141 ( .A1(n5680), .A2(n7497), .ZN(n5681) );
  NAND2_X1 U7142 ( .A1(n7500), .A2(n5681), .ZN(n7651) );
  NAND2_X1 U7143 ( .A1(n7651), .A2(n5682), .ZN(n7531) );
  OR2_X1 U7144 ( .A1(n5685), .A2(n5684), .ZN(n5687) );
  AND2_X1 U7145 ( .A1(n7405), .A2(n5687), .ZN(n5686) );
  INV_X1 U7146 ( .A(n5687), .ZN(n5690) );
  AND2_X1 U7147 ( .A1(n7528), .A2(n5688), .ZN(n5689) );
  INV_X1 U7148 ( .A(n5695), .ZN(n5697) );
  NAND2_X1 U7149 ( .A1(n7607), .A2(n5699), .ZN(n5701) );
  OR2_X1 U7150 ( .A1(n8962), .A2(n8854), .ZN(n5705) );
  INV_X1 U7151 ( .A(n5707), .ZN(n5708) );
  NAND2_X1 U7152 ( .A1(n8843), .A2(n8842), .ZN(n8841) );
  AND2_X1 U7153 ( .A1(n8804), .A2(n5714), .ZN(n8775) );
  INV_X1 U7154 ( .A(n8769), .ZN(n8779) );
  AND2_X1 U7155 ( .A1(n8775), .A2(n8779), .ZN(n5712) );
  INV_X1 U7156 ( .A(n8758), .ZN(n5713) );
  NOR2_X1 U7157 ( .A1(n8761), .A2(n5713), .ZN(n5718) );
  INV_X1 U7158 ( .A(n5714), .ZN(n5717) );
  NOR2_X1 U7159 ( .A1(n8792), .A2(n5715), .ZN(n5716) );
  OR2_X1 U7160 ( .A1(n5717), .A2(n5716), .ZN(n8776) );
  OR2_X1 U7161 ( .A1(n8769), .A2(n8776), .ZN(n8756) );
  AND2_X1 U7162 ( .A1(n5718), .A2(n8756), .ZN(n5719) );
  NOR2_X1 U7163 ( .A1(n8736), .A2(n8732), .ZN(n5720) );
  INV_X1 U7164 ( .A(n8725), .ZN(n5723) );
  INV_X1 U7165 ( .A(n8681), .ZN(n5726) );
  NOR2_X1 U7166 ( .A1(n8683), .A2(n5726), .ZN(n5727) );
  INV_X1 U7167 ( .A(n5730), .ZN(n5731) );
  OAI21_X1 U7168 ( .B1(n5736), .B2(n5735), .A(n5734), .ZN(n5739) );
  OAI21_X1 U7169 ( .B1(n5739), .B2(n5738), .A(n5737), .ZN(n5740) );
  XNOR2_X1 U7170 ( .A(n5740), .B(n6980), .ZN(n5745) );
  NOR2_X1 U7171 ( .A1(n5745), .A2(n5744), .ZN(n5746) );
  NAND2_X1 U7172 ( .A1(n5751), .A2(n5750), .ZN(n5752) );
  NAND2_X1 U7173 ( .A1(n5752), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5754) );
  INV_X1 U7174 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5753) );
  XNOR2_X1 U7175 ( .A(n5754), .B(n5753), .ZN(n5921) );
  OR2_X1 U7176 ( .A1(n5921), .A2(n7777), .ZN(n7300) );
  NAND2_X1 U7177 ( .A1(n5754), .A2(n5753), .ZN(n5755) );
  NAND2_X1 U7178 ( .A1(n5755), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5757) );
  INV_X1 U7179 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U7180 ( .A1(n5759), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5760) );
  XNOR2_X1 U7181 ( .A(n5760), .B(P2_IR_REG_26__SCAN_IN), .ZN(n5836) );
  INV_X1 U7182 ( .A(n5836), .ZN(n7742) );
  NAND2_X1 U7183 ( .A1(n4478), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5761) );
  XNOR2_X1 U7184 ( .A(n5761), .B(P2_IR_REG_25__SCAN_IN), .ZN(n5837) );
  INV_X1 U7185 ( .A(n5837), .ZN(n7647) );
  NAND2_X1 U7186 ( .A1(n6998), .A2(n5762), .ZN(n6591) );
  INV_X1 U7187 ( .A(n6591), .ZN(n6708) );
  INV_X1 U7188 ( .A(n5763), .ZN(n5827) );
  INV_X1 U7189 ( .A(n5861), .ZN(n5925) );
  NOR4_X1 U7190 ( .A1(n10130), .A2(n8853), .A3(n8044), .A4(n5925), .ZN(n5765)
         );
  OAI21_X1 U7191 ( .B1(n7300), .B2(n6998), .A(P2_B_REG_SCAN_IN), .ZN(n5764) );
  OR2_X1 U7192 ( .A1(n5765), .A2(n5764), .ZN(n5766) );
  OAI21_X1 U7193 ( .B1(n5767), .B2(n7300), .A(n5766), .ZN(P2_U3244) );
  NAND4_X1 U7194 ( .A1(n6038), .A2(n5771), .A3(n5770), .A4(n5769), .ZN(n5772)
         );
  NOR2_X1 U7195 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5774) );
  INV_X1 U7196 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5776) );
  INV_X1 U7197 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5775) );
  NOR2_X1 U7198 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5777) );
  NAND2_X1 U7199 ( .A1(n5799), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5779) );
  INV_X1 U7200 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U7201 ( .A1(n5779), .A2(n5798), .ZN(n5781) );
  NAND2_X1 U7202 ( .A1(n5781), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5778) );
  INV_X1 U7203 ( .A(n5779), .ZN(n5780) );
  NAND2_X1 U7204 ( .A1(n5780), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n5782) );
  NAND2_X1 U7205 ( .A1(n5782), .A2(n5781), .ZN(n7646) );
  NAND2_X1 U7206 ( .A1(n5783), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5784) );
  XNOR2_X1 U7207 ( .A(n5784), .B(n4802), .ZN(n7403) );
  NAND2_X1 U7208 ( .A1(n4484), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5786) );
  XNOR2_X1 U7209 ( .A(n5786), .B(n5785), .ZN(n7297) );
  INV_X1 U7210 ( .A(n7297), .ZN(n5795) );
  OR2_X1 U7211 ( .A1(n6093), .A2(n5795), .ZN(n6204) );
  OR2_X2 U7212 ( .A1(n6204), .A2(P1_U3084), .ZN(n9462) );
  INV_X1 U7213 ( .A(n9462), .ZN(P1_U4006) );
  INV_X1 U7214 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U7215 ( .A1(n5789), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5947) );
  XNOR2_X1 U7216 ( .A(n5790), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9442) );
  OR2_X1 U7217 ( .A1(n5792), .A2(n5791), .ZN(n5793) );
  NAND2_X1 U7218 ( .A1(n9442), .A2(n5948), .ZN(n9390) );
  OR2_X1 U7219 ( .A1(n9390), .A2(n5795), .ZN(n5796) );
  AND2_X1 U7220 ( .A1(n5796), .A2(n6204), .ZN(n6249) );
  INV_X1 U7221 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5797) );
  INV_X1 U7222 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5800) );
  INV_X1 U7223 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5931) );
  XNOR2_X2 U7224 ( .A(n5801), .B(n5931), .ZN(n6102) );
  NAND2_X1 U7225 ( .A1(n6249), .A2(n5965), .ZN(n6212) );
  NAND2_X1 U7226 ( .A1(n6212), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NAND2_X1 U7227 ( .A1(n5875), .A2(n10146), .ZN(n7319) );
  NAND2_X1 U7228 ( .A1(n5806), .A2(n7319), .ZN(n7318) );
  NAND2_X1 U7229 ( .A1(n5212), .A2(n10150), .ZN(n5807) );
  NAND2_X1 U7230 ( .A1(n7318), .A2(n5807), .ZN(n7426) );
  NAND2_X1 U7231 ( .A1(n7426), .A2(n7425), .ZN(n7424) );
  INV_X1 U7232 ( .A(n8568), .ZN(n7008) );
  NAND2_X1 U7233 ( .A1(n7008), .A2(n10156), .ZN(n5808) );
  NAND2_X1 U7234 ( .A1(n7424), .A2(n5808), .ZN(n7000) );
  NAND2_X1 U7235 ( .A1(n7000), .A2(n6999), .ZN(n7002) );
  INV_X1 U7236 ( .A(n8566), .ZN(n5809) );
  NAND2_X1 U7237 ( .A1(n5809), .A2(n7004), .ZN(n5810) );
  NAND2_X1 U7238 ( .A1(n7002), .A2(n5810), .ZN(n7496) );
  NAND2_X1 U7239 ( .A1(n7496), .A2(n7497), .ZN(n7495) );
  INV_X1 U7240 ( .A(n8565), .ZN(n7007) );
  NAND2_X1 U7241 ( .A1(n7007), .A2(n10162), .ZN(n5811) );
  NAND2_X1 U7242 ( .A1(n7495), .A2(n5811), .ZN(n7656) );
  NAND2_X1 U7243 ( .A1(n8564), .A2(n7664), .ZN(n5812) );
  NAND2_X1 U7244 ( .A1(n7656), .A2(n5812), .ZN(n5814) );
  NAND2_X1 U7245 ( .A1(n4593), .A2(n10169), .ZN(n5813) );
  NOR2_X1 U7246 ( .A1(n8563), .A2(n7540), .ZN(n5816) );
  NAND2_X1 U7247 ( .A1(n8563), .A2(n7540), .ZN(n5815) );
  OR2_X1 U7248 ( .A1(n7597), .A2(n7408), .ZN(n5818) );
  INV_X1 U7249 ( .A(n5902), .ZN(n7534) );
  NAND2_X1 U7250 ( .A1(n7534), .A2(n7468), .ZN(n5817) );
  AND2_X1 U7251 ( .A1(n5818), .A2(n5817), .ZN(n5820) );
  AND2_X1 U7252 ( .A1(n5822), .A2(n5817), .ZN(n7355) );
  NAND2_X1 U7253 ( .A1(n5818), .A2(n7355), .ZN(n5819) );
  OAI21_X1 U7254 ( .B1(n5820), .B2(n5822), .A(n5819), .ZN(n10178) );
  NAND2_X1 U7255 ( .A1(n5863), .A2(n5925), .ZN(n5821) );
  INV_X1 U7256 ( .A(n10145), .ZN(n5862) );
  NAND3_X1 U7257 ( .A1(n5821), .A2(n6591), .A3(n5862), .ZN(n8859) );
  OR2_X1 U7258 ( .A1(n10178), .A2(n8859), .ZN(n5832) );
  NAND2_X1 U7259 ( .A1(n5823), .A2(n5822), .ZN(n5824) );
  NAND2_X1 U7260 ( .A1(n5825), .A2(n5824), .ZN(n5830) );
  NAND2_X1 U7261 ( .A1(n5902), .A2(n8819), .ZN(n5828) );
  OAI21_X1 U7262 ( .B1(n7993), .B2(n8851), .A(n5828), .ZN(n5829) );
  AOI21_X1 U7263 ( .B1(n5830), .B2(n8863), .A(n5829), .ZN(n5831) );
  NAND2_X1 U7264 ( .A1(n5832), .A2(n5831), .ZN(n10181) );
  AND2_X1 U7265 ( .A1(n7381), .A2(n7742), .ZN(n10139) );
  XOR2_X1 U7266 ( .A(n7381), .B(P2_B_REG_SCAN_IN), .Z(n5833) );
  INV_X1 U7267 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10140) );
  AND2_X1 U7268 ( .A1(n10131), .A2(n10140), .ZN(n5835) );
  INV_X1 U7269 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10142) );
  NOR2_X1 U7270 ( .A1(n5837), .A2(n5836), .ZN(n10143) );
  AOI21_X1 U7271 ( .B1(n10131), .B2(n10142), .A(n10143), .ZN(n7018) );
  NOR4_X1 U7272 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5841) );
  NOR4_X1 U7273 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n5840) );
  NOR4_X1 U7274 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5839) );
  NOR4_X1 U7275 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5838) );
  NAND4_X1 U7276 ( .A1(n5841), .A2(n5840), .A3(n5839), .A4(n5838), .ZN(n5847)
         );
  NOR2_X1 U7277 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .ZN(
        n5845) );
  NOR4_X1 U7278 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5844) );
  NOR4_X1 U7279 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n5843) );
  NOR4_X1 U7280 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n5842) );
  NAND4_X1 U7281 ( .A1(n5845), .A2(n5844), .A3(n5843), .A4(n5842), .ZN(n5846)
         );
  OAI21_X1 U7282 ( .B1(n5847), .B2(n5846), .A(n10131), .ZN(n7154) );
  NAND2_X1 U7283 ( .A1(n7018), .A2(n7154), .ZN(n5860) );
  INV_X1 U7284 ( .A(n5860), .ZN(n5848) );
  OR2_X1 U7285 ( .A1(n6591), .A2(n5861), .ZN(n7014) );
  NAND3_X1 U7286 ( .A1(n7150), .A2(n5848), .A3(n7014), .ZN(n5849) );
  NAND2_X1 U7287 ( .A1(n10195), .A2(n5458), .ZN(n7015) );
  INV_X2 U7288 ( .A(n8846), .ZN(n8878) );
  MUX2_X1 U7289 ( .A(n10181), .B(P2_REG2_REG_8__SCAN_IN), .S(n8878), .Z(n5859)
         );
  NAND2_X1 U7290 ( .A1(n5850), .A2(n5741), .ZN(n5851) );
  NOR2_X1 U7291 ( .A1(n5853), .A2(n5851), .ZN(n7378) );
  INV_X1 U7292 ( .A(n7378), .ZN(n8873) );
  NOR2_X1 U7293 ( .A1(n10178), .A2(n8873), .ZN(n5858) );
  INV_X1 U7294 ( .A(n10162), .ZN(n7504) );
  NAND2_X1 U7295 ( .A1(n7660), .A2(n10169), .ZN(n7659) );
  NOR2_X1 U7296 ( .A1(n7411), .A2(n10179), .ZN(n5852) );
  OR2_X1 U7297 ( .A1(n7369), .A2(n5852), .ZN(n10180) );
  INV_X1 U7298 ( .A(n5853), .ZN(n5854) );
  NAND2_X1 U7299 ( .A1(n5854), .A2(n5743), .ZN(n8656) );
  NOR2_X1 U7300 ( .A1(n10180), .A2(n8656), .ZN(n5857) );
  AND2_X1 U7301 ( .A1(n10145), .A2(n5855), .ZN(n5917) );
  OAI22_X1 U7302 ( .A1(n8871), .A2(n10179), .B1(n8835), .B2(n7244), .ZN(n5856)
         );
  OR4_X1 U7303 ( .A1(n5859), .A2(n5858), .A3(n5857), .A4(n5856), .ZN(P2_U3288)
         );
  INV_X1 U7304 ( .A(n5922), .ZN(n6706) );
  NOR2_X1 U7305 ( .A1(n5920), .A2(n10130), .ZN(n5918) );
  INV_X1 U7306 ( .A(n5918), .ZN(n5926) );
  NAND2_X1 U7307 ( .A1(n5863), .A2(n7160), .ZN(n5865) );
  XNOR2_X1 U7308 ( .A(n7598), .B(n8365), .ZN(n5870) );
  INV_X1 U7309 ( .A(n5870), .ZN(n5867) );
  NOR2_X1 U7310 ( .A1(n7993), .A2(n5743), .ZN(n5868) );
  INV_X1 U7311 ( .A(n5868), .ZN(n5866) );
  NAND2_X1 U7312 ( .A1(n5867), .A2(n5866), .ZN(n7268) );
  INV_X1 U7313 ( .A(n7268), .ZN(n5869) );
  AND2_X1 U7314 ( .A1(n5870), .A2(n5868), .ZN(n7263) );
  NOR3_X1 U7315 ( .A1(n8553), .A2(n5869), .A3(n7263), .ZN(n5916) );
  NAND2_X1 U7316 ( .A1(n8476), .A2(n8367), .ZN(n8531) );
  INV_X1 U7317 ( .A(n8531), .ZN(n8493) );
  INV_X1 U7318 ( .A(n7993), .ZN(n8561) );
  NAND3_X1 U7319 ( .A1(n8493), .A2(n5870), .A3(n8561), .ZN(n5871) );
  OAI21_X1 U7320 ( .B1(n8553), .B2(n7268), .A(n5871), .ZN(n5915) );
  NAND2_X1 U7321 ( .A1(n5872), .A2(n8367), .ZN(n5873) );
  NAND2_X1 U7322 ( .A1(n5875), .A2(n8367), .ZN(n5876) );
  MUX2_X1 U7323 ( .A(n5876), .B(n8365), .S(n7314), .Z(n8474) );
  AND2_X1 U7324 ( .A1(n8568), .A2(n8367), .ZN(n5878) );
  XNOR2_X1 U7325 ( .A(n5886), .B(n10156), .ZN(n5877) );
  XNOR2_X1 U7326 ( .A(n5878), .B(n5877), .ZN(n7144) );
  INV_X1 U7327 ( .A(n5877), .ZN(n5880) );
  INV_X1 U7328 ( .A(n5878), .ZN(n5879) );
  OAI22_X1 U7329 ( .A1(n7143), .A2(n7144), .B1(n5880), .B2(n5879), .ZN(n7136)
         );
  XNOR2_X1 U7330 ( .A(n5886), .B(n7004), .ZN(n5882) );
  NAND2_X1 U7331 ( .A1(n8566), .A2(n8367), .ZN(n5881) );
  XNOR2_X1 U7332 ( .A(n5882), .B(n5881), .ZN(n7137) );
  NAND2_X1 U7333 ( .A1(n7136), .A2(n7137), .ZN(n5885) );
  INV_X1 U7334 ( .A(n5881), .ZN(n5883) );
  NAND2_X1 U7335 ( .A1(n5883), .A2(n5882), .ZN(n5884) );
  AND2_X1 U7336 ( .A1(n8565), .A2(n8367), .ZN(n5888) );
  XNOR2_X1 U7337 ( .A(n8376), .B(n10162), .ZN(n5887) );
  AND2_X1 U7338 ( .A1(n5888), .A2(n5887), .ZN(n7127) );
  INV_X1 U7339 ( .A(n5887), .ZN(n5890) );
  INV_X1 U7340 ( .A(n5888), .ZN(n5889) );
  NAND2_X1 U7341 ( .A1(n5890), .A2(n5889), .ZN(n7126) );
  AND2_X1 U7342 ( .A1(n8564), .A2(n8367), .ZN(n5891) );
  XNOR2_X1 U7343 ( .A(n8376), .B(n10169), .ZN(n7306) );
  NAND2_X1 U7344 ( .A1(n5891), .A2(n7306), .ZN(n5896) );
  INV_X1 U7345 ( .A(n7306), .ZN(n5893) );
  INV_X1 U7346 ( .A(n5891), .ZN(n5892) );
  NAND2_X1 U7347 ( .A1(n5893), .A2(n5892), .ZN(n5894) );
  NAND2_X1 U7348 ( .A1(n5896), .A2(n5894), .ZN(n7164) );
  INV_X1 U7349 ( .A(n7164), .ZN(n5895) );
  XNOR2_X1 U7350 ( .A(n8376), .B(n10172), .ZN(n5898) );
  NAND2_X1 U7351 ( .A1(n8563), .A2(n8367), .ZN(n5900) );
  XNOR2_X1 U7352 ( .A(n5898), .B(n5900), .ZN(n7304) );
  AND2_X1 U7353 ( .A1(n7304), .A2(n5896), .ZN(n5897) );
  INV_X1 U7354 ( .A(n5898), .ZN(n5899) );
  NAND2_X1 U7355 ( .A1(n5900), .A2(n5899), .ZN(n5901) );
  AND2_X1 U7356 ( .A1(n5902), .A2(n8367), .ZN(n5904) );
  XNOR2_X1 U7357 ( .A(n7468), .B(n8376), .ZN(n5903) );
  NAND2_X1 U7358 ( .A1(n5904), .A2(n5903), .ZN(n5912) );
  INV_X1 U7359 ( .A(n5903), .ZN(n7239) );
  INV_X1 U7360 ( .A(n5904), .ZN(n5905) );
  NAND2_X1 U7361 ( .A1(n7239), .A2(n5905), .ZN(n5906) );
  AND2_X1 U7362 ( .A1(n5912), .A2(n5906), .ZN(n7229) );
  XNOR2_X1 U7363 ( .A(n10179), .B(n8376), .ZN(n5910) );
  NAND2_X1 U7364 ( .A1(n8562), .A2(n8367), .ZN(n5908) );
  XNOR2_X1 U7365 ( .A(n5910), .B(n5908), .ZN(n5911) );
  AND2_X1 U7366 ( .A1(n7229), .A2(n5911), .ZN(n5907) );
  INV_X1 U7367 ( .A(n5908), .ZN(n5909) );
  NAND2_X1 U7368 ( .A1(n5910), .A2(n5909), .ZN(n5913) );
  INV_X1 U7369 ( .A(n5911), .ZN(n7237) );
  OR2_X1 U7370 ( .A1(n7237), .A2(n5912), .ZN(n7240) );
  AND2_X1 U7371 ( .A1(n5913), .A2(n7240), .ZN(n7264) );
  NAND2_X1 U7372 ( .A1(n7267), .A2(n7264), .ZN(n5914) );
  MUX2_X1 U7373 ( .A(n5916), .B(n5915), .S(n5914), .Z(n5930) );
  NAND2_X1 U7374 ( .A1(n5918), .A2(n5917), .ZN(n5919) );
  INV_X1 U7375 ( .A(n7598), .ZN(n7376) );
  NOR2_X1 U7376 ( .A1(n8541), .A2(n7376), .ZN(n5929) );
  NAND2_X1 U7377 ( .A1(n5920), .A2(n7015), .ZN(n5924) );
  AND3_X1 U7378 ( .A1(n5922), .A2(n5921), .A3(n7014), .ZN(n5923) );
  NAND2_X1 U7379 ( .A1(n5924), .A2(n5923), .ZN(n7145) );
  NAND2_X1 U7380 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(n7777), .ZN(n6710) );
  OAI21_X1 U7381 ( .B1(n8546), .B2(n7372), .A(n6710), .ZN(n5928) );
  INV_X1 U7382 ( .A(n8562), .ZN(n7232) );
  OAI22_X1 U7383 ( .A1(n7232), .A2(n8548), .B1(n8547), .B2(n7397), .ZN(n5927)
         );
  OR4_X1 U7384 ( .A1(n5930), .A2(n5929), .A3(n5928), .A4(n5927), .ZN(P2_U3233)
         );
  INV_X1 U7385 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9790) );
  NAND2_X1 U7386 ( .A1(n5933), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5934) );
  INV_X1 U7387 ( .A(n5935), .ZN(n9793) );
  AND2_X2 U7388 ( .A1(n5936), .A2(n9793), .ZN(n5940) );
  NAND2_X2 U7389 ( .A1(n5938), .A2(n5940), .ZN(n8425) );
  INV_X1 U7390 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6587) );
  INV_X1 U7391 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5937) );
  NAND2_X2 U7393 ( .A1(n5941), .A2(n7923), .ZN(n8333) );
  INV_X1 U7394 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5939) );
  OR2_X1 U7395 ( .A1(n8333), .A2(n5939), .ZN(n5943) );
  NAND2_X4 U7396 ( .A1(n5941), .A2(n5940), .ZN(n8332) );
  INV_X1 U7397 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10043) );
  XNOR2_X1 U7398 ( .A(n5947), .B(n5946), .ZN(n7142) );
  NAND2_X1 U7399 ( .A1(n4400), .A2(n7480), .ZN(n5954) );
  OR2_X1 U7400 ( .A1(n6003), .A2(n6180), .ZN(n5952) );
  INV_X1 U7401 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6172) );
  INV_X1 U7402 ( .A(n5949), .ZN(n5950) );
  OR2_X1 U7403 ( .A1(n5965), .A2(n6251), .ZN(n5951) );
  NAND2_X1 U7404 ( .A1(n5954), .A2(n5953), .ZN(n5957) );
  NAND2_X1 U7405 ( .A1(n5955), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5956) );
  XNOR2_X1 U7406 ( .A(n5956), .B(n5788), .ZN(n9499) );
  NAND2_X1 U7407 ( .A1(n6030), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5963) );
  INV_X1 U7408 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U7409 ( .A1(n8421), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5961) );
  INV_X1 U7410 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5959) );
  OR2_X1 U7411 ( .A1(n8333), .A2(n5959), .ZN(n5960) );
  INV_X2 U7412 ( .A(n7710), .ZN(n7480) );
  NAND2_X1 U7413 ( .A1(n6229), .A2(n7480), .ZN(n5968) );
  NAND2_X1 U7414 ( .A1(n4402), .A2(SI_0_), .ZN(n5964) );
  XNOR2_X1 U7415 ( .A(n5964), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9798) );
  INV_X1 U7416 ( .A(n6093), .ZN(n5966) );
  AOI22_X1 U7417 ( .A1(n6904), .A2(n8307), .B1(n5966), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U7418 ( .A1(n5968), .A2(n5967), .ZN(n6606) );
  AND2_X1 U7419 ( .A1(n7142), .A2(n9499), .ZN(n6091) );
  NAND2_X1 U7420 ( .A1(n9393), .A2(n6091), .ZN(n6626) );
  INV_X1 U7421 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6207) );
  INV_X2 U7422 ( .A(n7710), .ZN(n8319) );
  NAND2_X1 U7423 ( .A1(n6904), .A2(n8319), .ZN(n5969) );
  OAI21_X1 U7424 ( .B1(n6207), .B2(n6093), .A(n5969), .ZN(n5970) );
  NAND2_X1 U7425 ( .A1(n6606), .A2(n6604), .ZN(n6605) );
  OAI21_X1 U7426 ( .B1(n6606), .B2(n8184), .A(n6605), .ZN(n5971) );
  NAND2_X1 U7427 ( .A1(n5971), .A2(n5972), .ZN(n5978) );
  OAI21_X1 U7428 ( .B1(n5972), .B2(n5971), .A(n5978), .ZN(n6687) );
  INV_X1 U7429 ( .A(n6687), .ZN(n5977) );
  NAND2_X1 U7430 ( .A1(n4400), .A2(n8324), .ZN(n5975) );
  OR2_X1 U7431 ( .A1(n10045), .A2(n8297), .ZN(n5974) );
  NAND2_X1 U7432 ( .A1(n5975), .A2(n5974), .ZN(n6688) );
  NAND2_X1 U7433 ( .A1(n5977), .A2(n5976), .ZN(n6685) );
  NAND2_X1 U7434 ( .A1(n6685), .A2(n5978), .ZN(n6787) );
  INV_X1 U7435 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5979) );
  INV_X1 U7436 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6789) );
  OR2_X1 U7437 ( .A1(n8332), .A2(n6789), .ZN(n5982) );
  INV_X1 U7438 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6260) );
  OR2_X1 U7439 ( .A1(n8425), .A2(n6260), .ZN(n5981) );
  NAND2_X1 U7440 ( .A1(n5995), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5980) );
  AND4_X2 U7441 ( .A1(n5983), .A2(n5982), .A3(n5981), .A4(n5980), .ZN(n6952)
         );
  NOR2_X1 U7442 ( .A1(n5949), .A2(n6320), .ZN(n5984) );
  MUX2_X1 U7443 ( .A(n6320), .B(n5984), .S(P1_IR_REG_2__SCAN_IN), .Z(n5985) );
  INV_X1 U7444 ( .A(n5985), .ZN(n5987) );
  NAND2_X1 U7445 ( .A1(n5987), .A2(n5986), .ZN(n6279) );
  OR2_X1 U7446 ( .A1(n9154), .A2(n6178), .ZN(n5989) );
  OR2_X1 U7447 ( .A1(n6003), .A2(n6189), .ZN(n5988) );
  INV_X1 U7448 ( .A(n6991), .ZN(n6990) );
  XNOR2_X1 U7449 ( .A(n5990), .B(n8184), .ZN(n5991) );
  OAI22_X1 U7450 ( .A1(n6952), .A2(n8300), .B1(n6990), .B2(n8297), .ZN(n5992)
         );
  XNOR2_X1 U7451 ( .A(n5991), .B(n5992), .ZN(n6786) );
  INV_X1 U7452 ( .A(n5991), .ZN(n5993) );
  OR2_X1 U7453 ( .A1(n5993), .A2(n5992), .ZN(n5994) );
  NAND2_X1 U7454 ( .A1(n6788), .A2(n5994), .ZN(n6866) );
  NAND2_X1 U7455 ( .A1(n5995), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6001) );
  OR2_X1 U7456 ( .A1(n8332), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6000) );
  INV_X1 U7457 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6261) );
  OR2_X1 U7458 ( .A1(n8425), .A2(n6261), .ZN(n5999) );
  INV_X1 U7459 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5997) );
  OR2_X1 U7460 ( .A1(n5996), .A2(n5997), .ZN(n5998) );
  NAND2_X1 U7461 ( .A1(n5986), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6002) );
  XNOR2_X1 U7462 ( .A(n6002), .B(n5768), .ZN(n6290) );
  OR2_X1 U7463 ( .A1(n9154), .A2(n6173), .ZN(n6005) );
  OR2_X1 U7464 ( .A1(n6003), .A2(n6194), .ZN(n6004) );
  OAI211_X1 U7465 ( .C1(n5965), .C2(n6290), .A(n6005), .B(n6004), .ZN(n6959)
         );
  INV_X1 U7466 ( .A(n6959), .ZN(n10066) );
  OAI22_X1 U7467 ( .A1(n6966), .A2(n8297), .B1(n10066), .B2(n8298), .ZN(n6006)
         );
  XNOR2_X1 U7468 ( .A(n6006), .B(n8184), .ZN(n6010) );
  OR2_X1 U7469 ( .A1(n6966), .A2(n8300), .ZN(n6008) );
  NAND2_X1 U7470 ( .A1(n6959), .A2(n7480), .ZN(n6007) );
  NAND2_X1 U7471 ( .A1(n6008), .A2(n6007), .ZN(n6011) );
  INV_X1 U7472 ( .A(n6011), .ZN(n6009) );
  AND2_X1 U7473 ( .A1(n6010), .A2(n6009), .ZN(n6868) );
  INV_X1 U7474 ( .A(n6010), .ZN(n6012) );
  NAND2_X1 U7475 ( .A1(n6012), .A2(n6011), .ZN(n6867) );
  NAND2_X1 U7476 ( .A1(n5995), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6021) );
  INV_X1 U7477 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6015) );
  OR2_X1 U7478 ( .A1(n5996), .A2(n6015), .ZN(n6020) );
  INV_X1 U7479 ( .A(n6031), .ZN(n6017) );
  INV_X1 U7480 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6295) );
  INV_X1 U7481 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6916) );
  NAND2_X1 U7482 ( .A1(n6295), .A2(n6916), .ZN(n6016) );
  NAND2_X1 U7483 ( .A1(n6017), .A2(n6016), .ZN(n6970) );
  OR2_X1 U7484 ( .A1(n8332), .A2(n6970), .ZN(n6019) );
  INV_X1 U7485 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9908) );
  OR2_X1 U7486 ( .A1(n8425), .A2(n9908), .ZN(n6018) );
  NAND2_X1 U7487 ( .A1(n6022), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6023) );
  INV_X1 U7488 ( .A(n9907), .ZN(n6176) );
  OR2_X1 U7489 ( .A1(n6003), .A2(n6186), .ZN(n6025) );
  OR2_X1 U7490 ( .A1(n9154), .A2(n6175), .ZN(n6024) );
  OAI211_X1 U7491 ( .C1(n5965), .C2(n6176), .A(n6025), .B(n6024), .ZN(n6976)
         );
  OAI22_X1 U7492 ( .A1(n7027), .A2(n8297), .B1(n10072), .B2(n8298), .ZN(n6026)
         );
  XNOR2_X1 U7493 ( .A(n6026), .B(n8184), .ZN(n6027) );
  OAI22_X1 U7494 ( .A1(n7027), .A2(n8300), .B1(n10072), .B2(n8297), .ZN(n6028)
         );
  XNOR2_X1 U7495 ( .A(n6027), .B(n6028), .ZN(n6915) );
  INV_X1 U7496 ( .A(n6027), .ZN(n6029) );
  NAND2_X1 U7497 ( .A1(n6030), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6036) );
  INV_X1 U7498 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6275) );
  OR2_X1 U7499 ( .A1(n8333), .A2(n6275), .ZN(n6035) );
  OAI21_X1 U7500 ( .B1(n6031), .B2(P1_REG3_REG_5__SCAN_IN), .A(n6051), .ZN(
        n7121) );
  OR2_X1 U7501 ( .A1(n8332), .A2(n7121), .ZN(n6034) );
  INV_X1 U7502 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6032) );
  OR2_X1 U7503 ( .A1(n5996), .A2(n6032), .ZN(n6033) );
  NOR2_X1 U7504 ( .A1(n6022), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6039) );
  NOR2_X1 U7505 ( .A1(n6039), .A2(n6320), .ZN(n6037) );
  MUX2_X1 U7506 ( .A(n6320), .B(n6037), .S(P1_IR_REG_5__SCAN_IN), .Z(n6041) );
  NAND2_X1 U7507 ( .A1(n6039), .A2(n6038), .ZN(n6121) );
  INV_X1 U7508 ( .A(n6121), .ZN(n6040) );
  AOI22_X1 U7509 ( .A1(n8150), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8149), .B2(
        n9918), .ZN(n6043) );
  OR2_X1 U7510 ( .A1(n6193), .A2(n6003), .ZN(n6042) );
  NAND2_X1 U7511 ( .A1(n6043), .A2(n6042), .ZN(n7112) );
  INV_X1 U7512 ( .A(n7112), .ZN(n7022) );
  OAI22_X1 U7513 ( .A1(n7021), .A2(n8297), .B1(n7022), .B2(n8298), .ZN(n6044)
         );
  XNOR2_X1 U7514 ( .A(n6044), .B(n8184), .ZN(n7115) );
  OR2_X1 U7515 ( .A1(n7021), .A2(n8300), .ZN(n6046) );
  NAND2_X1 U7516 ( .A1(n7112), .A2(n7480), .ZN(n6045) );
  NAND2_X1 U7517 ( .A1(n6046), .A2(n6045), .ZN(n6048) );
  INV_X1 U7518 ( .A(n6048), .ZN(n7114) );
  NAND2_X1 U7519 ( .A1(n7115), .A2(n7114), .ZN(n6047) );
  INV_X1 U7520 ( .A(n7115), .ZN(n6049) );
  NAND2_X1 U7521 ( .A1(n6049), .A2(n6048), .ZN(n6050) );
  NAND2_X1 U7522 ( .A1(n8421), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6057) );
  INV_X1 U7523 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7049) );
  OR2_X1 U7524 ( .A1(n8333), .A2(n7049), .ZN(n6056) );
  AND2_X1 U7525 ( .A1(n6051), .A2(n6111), .ZN(n6052) );
  OR2_X1 U7526 ( .A1(n6052), .A2(n6105), .ZN(n7048) );
  OR2_X1 U7527 ( .A1(n8332), .A2(n7048), .ZN(n6055) );
  INV_X1 U7528 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6053) );
  OR2_X1 U7529 ( .A1(n8425), .A2(n6053), .ZN(n6054) );
  OR2_X1 U7530 ( .A1(n7064), .A2(n8300), .ZN(n6061) );
  NAND2_X1 U7531 ( .A1(n6121), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6058) );
  XNOR2_X1 U7532 ( .A(n6058), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6311) );
  AOI22_X1 U7533 ( .A1(n8150), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8149), .B2(
        n6311), .ZN(n6059) );
  NAND2_X1 U7534 ( .A1(n7051), .A2(n7480), .ZN(n6060) );
  NAND2_X1 U7535 ( .A1(n6061), .A2(n6060), .ZN(n6118) );
  NAND2_X1 U7536 ( .A1(n7051), .A2(n8307), .ZN(n6062) );
  OAI21_X1 U7537 ( .B1(n7064), .B2(n8297), .A(n6062), .ZN(n6063) );
  XNOR2_X1 U7538 ( .A(n6063), .B(n8322), .ZN(n6117) );
  XOR2_X1 U7539 ( .A(n6118), .B(n6117), .Z(n6064) );
  XNOR2_X1 U7540 ( .A(n6119), .B(n6064), .ZN(n6088) );
  NAND2_X1 U7541 ( .A1(n7646), .A2(P1_B_REG_SCAN_IN), .ZN(n6066) );
  INV_X1 U7542 ( .A(n7403), .ZN(n6065) );
  MUX2_X1 U7543 ( .A(n6066), .B(P1_B_REG_SCAN_IN), .S(n6065), .Z(n6067) );
  NAND2_X1 U7544 ( .A1(n6067), .A2(n6068), .ZN(n6199) );
  INV_X1 U7545 ( .A(n6199), .ZN(n6082) );
  INV_X1 U7546 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U7547 ( .A1(n6082), .A2(n6185), .ZN(n6070) );
  INV_X1 U7548 ( .A(n6068), .ZN(n7744) );
  NAND2_X1 U7549 ( .A1(n7744), .A2(n7646), .ZN(n6069) );
  NAND2_X1 U7550 ( .A1(n6070), .A2(n6069), .ZN(n6896) );
  INV_X1 U7551 ( .A(n6896), .ZN(n6183) );
  NOR2_X1 U7552 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .ZN(
        n6074) );
  NOR4_X1 U7553 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n6073) );
  NOR4_X1 U7554 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6072) );
  NOR4_X1 U7555 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6071) );
  NAND4_X1 U7556 ( .A1(n6074), .A2(n6073), .A3(n6072), .A4(n6071), .ZN(n6080)
         );
  NOR4_X1 U7557 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6078) );
  NOR4_X1 U7558 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n6077) );
  NOR4_X1 U7559 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6076) );
  NOR4_X1 U7560 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6075) );
  NAND4_X1 U7561 ( .A1(n6078), .A2(n6077), .A3(n6076), .A4(n6075), .ZN(n6079)
         );
  NOR2_X1 U7562 ( .A1(n6080), .A2(n6079), .ZN(n6081) );
  NOR2_X1 U7563 ( .A1(n6199), .A2(n6081), .ZN(n6614) );
  INV_X1 U7564 ( .A(n6614), .ZN(n6084) );
  INV_X1 U7565 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6421) );
  NAND2_X1 U7566 ( .A1(n6082), .A2(n6421), .ZN(n6083) );
  NAND2_X1 U7567 ( .A1(n7744), .A2(n7403), .ZN(n6200) );
  NAND3_X1 U7568 ( .A1(n6183), .A2(n6084), .A3(n6897), .ZN(n6095) );
  AND2_X1 U7569 ( .A1(n7297), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6085) );
  INV_X1 U7570 ( .A(n9439), .ZN(n6089) );
  NOR2_X1 U7571 ( .A1(n6095), .A2(n6089), .ZN(n6101) );
  INV_X1 U7572 ( .A(n5948), .ZN(n9190) );
  NAND2_X1 U7573 ( .A1(n9393), .A2(n9190), .ZN(n6637) );
  INV_X1 U7574 ( .A(n6637), .ZN(n6617) );
  INV_X1 U7575 ( .A(n6091), .ZN(n6086) );
  INV_X1 U7576 ( .A(n9390), .ZN(n6629) );
  NOR2_X1 U7577 ( .A1(n9766), .A2(n6629), .ZN(n6087) );
  NAND2_X1 U7578 ( .A1(n6101), .A2(n6087), .ZN(n9146) );
  NOR2_X1 U7579 ( .A1(n6088), .A2(n9146), .ZN(n6116) );
  AND2_X1 U7580 ( .A1(n7051), .A2(n9766), .ZN(n10084) );
  OR2_X1 U7581 ( .A1(n6637), .A2(n7142), .ZN(n10044) );
  NOR2_X1 U7582 ( .A1(n10044), .A2(n6089), .ZN(n6090) );
  NAND2_X1 U7583 ( .A1(n6095), .A2(n6090), .ZN(n6098) );
  OR2_X1 U7584 ( .A1(n9390), .A2(n6091), .ZN(n6094) );
  NAND2_X1 U7585 ( .A1(n6094), .A2(n9439), .ZN(n6615) );
  INV_X1 U7586 ( .A(n6615), .ZN(n6092) );
  AND2_X1 U7587 ( .A1(n6098), .A2(n6092), .ZN(n6690) );
  AND2_X1 U7588 ( .A1(n10084), .A2(n6690), .ZN(n6115) );
  AND3_X1 U7589 ( .A1(n6094), .A2(n6093), .A3(n7297), .ZN(n6096) );
  INV_X1 U7590 ( .A(n9766), .ZN(n10093) );
  NAND2_X1 U7591 ( .A1(n6095), .A2(n10093), .ZN(n6603) );
  NAND2_X1 U7592 ( .A1(n6096), .A2(n6603), .ZN(n6097) );
  NAND2_X1 U7593 ( .A1(n6097), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6099) );
  NOR2_X1 U7594 ( .A1(n9142), .A2(n7048), .ZN(n6114) );
  OR2_X1 U7595 ( .A1(n6100), .A2(n6624), .ZN(n9441) );
  INV_X1 U7596 ( .A(n9441), .ZN(n6618) );
  NAND2_X1 U7597 ( .A1(n6101), .A2(n6618), .ZN(n6103) );
  OR2_X1 U7598 ( .A1(n6103), .A2(n6102), .ZN(n9137) );
  INV_X1 U7599 ( .A(n6103), .ZN(n6104) );
  NAND2_X1 U7600 ( .A1(n8421), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6110) );
  INV_X1 U7601 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7072) );
  OR2_X1 U7602 ( .A1(n8333), .A2(n7072), .ZN(n6109) );
  NAND2_X1 U7603 ( .A1(n6105), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6140) );
  OR2_X1 U7604 ( .A1(n6105), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U7605 ( .A1(n6140), .A2(n6106), .ZN(n7343) );
  OR2_X1 U7606 ( .A1(n8332), .A2(n7343), .ZN(n6108) );
  OR2_X1 U7607 ( .A1(n8425), .A2(n10114), .ZN(n6107) );
  INV_X1 U7608 ( .A(n7082), .ZN(n9456) );
  NAND2_X1 U7609 ( .A1(n9139), .A2(n9456), .ZN(n6112) );
  OR2_X1 U7610 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6111), .ZN(n6285) );
  OAI211_X1 U7611 ( .C1(n7021), .C2(n9137), .A(n6112), .B(n6285), .ZN(n6113)
         );
  OR4_X1 U7612 ( .A1(n6116), .A2(n6115), .A3(n6114), .A4(n6113), .ZN(P1_U3237)
         );
  NAND2_X1 U7613 ( .A1(n6119), .A2(n6118), .ZN(n6120) );
  NAND2_X1 U7614 ( .A1(n6196), .A2(n9151), .ZN(n6127) );
  OAI21_X1 U7615 ( .B1(n6121), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6122) );
  MUX2_X1 U7616 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6122), .S(
        P1_IR_REG_7__SCAN_IN), .Z(n6125) );
  INV_X1 U7617 ( .A(n6123), .ZN(n6124) );
  AOI22_X1 U7618 ( .A1(n8150), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8149), .B2(
        n6671), .ZN(n6126) );
  NAND2_X1 U7619 ( .A1(n6127), .A2(n6126), .ZN(n7352) );
  NAND2_X1 U7620 ( .A1(n7352), .A2(n8307), .ZN(n6129) );
  OR2_X1 U7621 ( .A1(n7082), .A2(n8297), .ZN(n6128) );
  NAND2_X1 U7622 ( .A1(n6129), .A2(n6128), .ZN(n6130) );
  XNOR2_X1 U7623 ( .A(n6130), .B(n8184), .ZN(n6133) );
  NAND2_X1 U7624 ( .A1(n9456), .A2(n8324), .ZN(n6132) );
  NAND2_X1 U7625 ( .A1(n7352), .A2(n7480), .ZN(n6131) );
  AND2_X1 U7626 ( .A1(n6132), .A2(n6131), .ZN(n6134) );
  NAND2_X1 U7627 ( .A1(n6133), .A2(n6134), .ZN(n7346) );
  NAND2_X1 U7628 ( .A1(n7345), .A2(n7346), .ZN(n7344) );
  INV_X1 U7629 ( .A(n6133), .ZN(n6136) );
  INV_X1 U7630 ( .A(n6134), .ZN(n6135) );
  NAND2_X1 U7631 ( .A1(n6136), .A2(n6135), .ZN(n7348) );
  NAND2_X1 U7632 ( .A1(n6202), .A2(n9151), .ZN(n6139) );
  OR2_X1 U7633 ( .A1(n6123), .A2(n6320), .ZN(n6137) );
  XNOR2_X1 U7634 ( .A(n6137), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9929) );
  AOI22_X1 U7635 ( .A1(n8150), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8149), .B2(
        n9929), .ZN(n6138) );
  NAND2_X1 U7636 ( .A1(n6139), .A2(n6138), .ZN(n7177) );
  NAND2_X1 U7637 ( .A1(n7177), .A2(n7480), .ZN(n6147) );
  NAND2_X1 U7638 ( .A1(n8421), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6145) );
  INV_X1 U7639 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7090) );
  OR2_X1 U7640 ( .A1(n8333), .A2(n7090), .ZN(n6144) );
  NAND2_X1 U7641 ( .A1(n6140), .A2(n6166), .ZN(n6141) );
  NAND2_X1 U7642 ( .A1(n6158), .A2(n6141), .ZN(n7089) );
  OR2_X1 U7643 ( .A1(n8332), .A2(n7089), .ZN(n6143) );
  INV_X1 U7644 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6662) );
  OR2_X1 U7645 ( .A1(n8425), .A2(n6662), .ZN(n6142) );
  INV_X1 U7646 ( .A(n7251), .ZN(n9455) );
  NAND2_X1 U7647 ( .A1(n9455), .A2(n8324), .ZN(n6146) );
  NAND2_X1 U7648 ( .A1(n6147), .A2(n6146), .ZN(n6150) );
  NAND2_X1 U7649 ( .A1(n6151), .A2(n6150), .ZN(n7453) );
  NAND2_X1 U7650 ( .A1(n7454), .A2(n7453), .ZN(n6155) );
  NAND2_X1 U7651 ( .A1(n7177), .A2(n8307), .ZN(n6153) );
  NAND2_X1 U7652 ( .A1(n9455), .A2(n7480), .ZN(n6152) );
  NAND2_X1 U7653 ( .A1(n6153), .A2(n6152), .ZN(n6154) );
  XNOR2_X1 U7654 ( .A(n6154), .B(n8184), .ZN(n7452) );
  XNOR2_X1 U7655 ( .A(n6155), .B(n7452), .ZN(n6156) );
  NOR2_X1 U7656 ( .A1(n6156), .A2(n9146), .ZN(n6171) );
  NAND2_X1 U7657 ( .A1(n7177), .A2(n9766), .ZN(n10098) );
  INV_X1 U7658 ( .A(n6690), .ZN(n7125) );
  NOR2_X1 U7659 ( .A1(n10098), .A2(n7125), .ZN(n6170) );
  NOR2_X1 U7660 ( .A1(n9142), .A2(n7089), .ZN(n6169) );
  INV_X1 U7661 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6157) );
  OR2_X1 U7662 ( .A1(n8425), .A2(n6157), .ZN(n6165) );
  INV_X1 U7663 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7460) );
  AND2_X1 U7664 ( .A1(n6158), .A2(n7460), .ZN(n6159) );
  OR2_X1 U7665 ( .A1(n6159), .A2(n7189), .ZN(n7459) );
  OR2_X1 U7666 ( .A1(n8332), .A2(n7459), .ZN(n6164) );
  INV_X1 U7667 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6160) );
  OR2_X1 U7668 ( .A1(n8333), .A2(n6160), .ZN(n6163) );
  INV_X1 U7669 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n6161) );
  OR2_X1 U7670 ( .A1(n5996), .A2(n6161), .ZN(n6162) );
  NAND4_X1 U7671 ( .A1(n6165), .A2(n6164), .A3(n6163), .A4(n6162), .ZN(n9454)
         );
  NAND2_X1 U7672 ( .A1(n9139), .A2(n9454), .ZN(n6167) );
  OR2_X1 U7673 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6166), .ZN(n9940) );
  OAI211_X1 U7674 ( .C1(n7082), .C2(n9137), .A(n6167), .B(n9940), .ZN(n6168)
         );
  OR4_X1 U7675 ( .A1(n6171), .A2(n6170), .A3(n6169), .A4(n6168), .ZN(P1_U3219)
         );
  NAND2_X2 U7676 ( .A1(n6179), .A2(P1_U3084), .ZN(n9791) );
  NAND2_X1 U7677 ( .A1(n4402), .A2(P1_U3084), .ZN(n9796) );
  OAI222_X1 U7678 ( .A1(n9791), .A2(n6172), .B1(n9796), .B2(n6180), .C1(
        P1_U3084), .C2(n6251), .ZN(P1_U3352) );
  OAI222_X1 U7679 ( .A1(n9791), .A2(n6173), .B1(n9796), .B2(n6194), .C1(n6290), 
        .C2(P1_U3084), .ZN(P1_U3350) );
  OAI222_X1 U7680 ( .A1(n9791), .A2(n6174), .B1(n9796), .B2(n6193), .C1(n6276), 
        .C2(P1_U3084), .ZN(P1_U3348) );
  INV_X1 U7681 ( .A(n9796), .ZN(n7773) );
  INV_X1 U7682 ( .A(n7773), .ZN(n7925) );
  OAI222_X1 U7683 ( .A1(n6176), .A2(P1_U3084), .B1(n7925), .B2(n6186), .C1(
        n6175), .C2(n9791), .ZN(P1_U3349) );
  INV_X1 U7684 ( .A(n6311), .ZN(n6286) );
  OAI222_X1 U7685 ( .A1(n6286), .A2(P1_U3084), .B1(n7925), .B2(n6191), .C1(
        n6177), .C2(n9791), .ZN(P1_U3347) );
  OAI222_X1 U7686 ( .A1(n9791), .A2(n6178), .B1(n7925), .B2(n6189), .C1(n6279), 
        .C2(P1_U3084), .ZN(P1_U3351) );
  AND2_X1 U7687 ( .A1(n4402), .A2(P2_U3152), .ZN(n9000) );
  NAND2_X1 U7688 ( .A1(n6179), .A2(P2_U3152), .ZN(n8110) );
  OAI222_X1 U7689 ( .A1(n8438), .A2(n6182), .B1(n6181), .B2(P2_U3152), .C1(
        n8110), .C2(n6180), .ZN(P2_U3357) );
  NAND2_X1 U7690 ( .A1(n6183), .A2(n9439), .ZN(n6184) );
  OAI21_X1 U7691 ( .B1(n9439), .B2(n6185), .A(n6184), .ZN(P1_U3441) );
  INV_X1 U7692 ( .A(n8110), .ZN(n7299) );
  INV_X1 U7693 ( .A(n7299), .ZN(n9002) );
  OAI222_X1 U7694 ( .A1(n8438), .A2(n6187), .B1(n9002), .B2(n6186), .C1(
        P2_U3152), .C2(n6804), .ZN(P2_U3354) );
  OAI222_X1 U7695 ( .A1(n8438), .A2(n6190), .B1(n9002), .B2(n6189), .C1(n7777), 
        .C2(n6188), .ZN(P2_U3356) );
  OAI222_X1 U7696 ( .A1(n8438), .A2(n6192), .B1(n9002), .B2(n6191), .C1(
        P2_U3152), .C2(n6816), .ZN(P2_U3352) );
  OAI222_X1 U7697 ( .A1(n8438), .A2(n6408), .B1(n9002), .B2(n6193), .C1(n7777), 
        .C2(n6840), .ZN(P2_U3353) );
  OAI222_X1 U7698 ( .A1(n8438), .A2(n6195), .B1(n9002), .B2(n6194), .C1(
        P2_U3152), .C2(n6828), .ZN(P2_U3355) );
  INV_X1 U7699 ( .A(n6671), .ZN(n6309) );
  INV_X1 U7700 ( .A(n6196), .ZN(n6198) );
  INV_X1 U7701 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6197) );
  OAI222_X1 U7702 ( .A1(n6309), .A2(P1_U3084), .B1(n9796), .B2(n6198), .C1(
        n6197), .C2(n9791), .ZN(P1_U3346) );
  OAI222_X1 U7703 ( .A1(n8438), .A2(n6513), .B1(n9002), .B2(n6198), .C1(n7777), 
        .C2(n6852), .ZN(P2_U3351) );
  NAND2_X1 U7704 ( .A1(n9439), .A2(n6199), .ZN(n10058) );
  INV_X1 U7705 ( .A(n10058), .ZN(n10057) );
  OAI21_X1 U7706 ( .B1(n10057), .B2(P1_D_REG_0__SCAN_IN), .A(n6200), .ZN(n6201) );
  OAI21_X1 U7707 ( .B1(n9439), .B2(n6421), .A(n6201), .ZN(P1_U3440) );
  INV_X1 U7708 ( .A(n6202), .ZN(n6203) );
  OAI222_X1 U7709 ( .A1(n8438), .A2(n6444), .B1(n9002), .B2(n6203), .C1(n7777), 
        .C2(n6863), .ZN(P2_U3350) );
  INV_X1 U7710 ( .A(n9929), .ZN(n6669) );
  OAI222_X1 U7711 ( .A1(n6669), .A2(P1_U3084), .B1(n9796), .B2(n6203), .C1(
        n6411), .C2(n9791), .ZN(P1_U3345) );
  INV_X1 U7712 ( .A(n6204), .ZN(n6205) );
  OR2_X1 U7713 ( .A1(P1_U3083), .A2(n6205), .ZN(n10035) );
  INV_X1 U7714 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6218) );
  NOR2_X1 U7715 ( .A1(n8427), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6206) );
  OR2_X1 U7716 ( .A1(n6206), .A2(n6102), .ZN(n6208) );
  NAND2_X1 U7717 ( .A1(n6208), .A2(n6207), .ZN(n6648) );
  INV_X1 U7718 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6622) );
  INV_X1 U7719 ( .A(n6102), .ZN(n9438) );
  INV_X1 U7720 ( .A(n8427), .ZN(n9437) );
  NAND2_X1 U7721 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6647) );
  NAND2_X1 U7722 ( .A1(n9437), .A2(n6647), .ZN(n6209) );
  OAI211_X1 U7723 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n6622), .A(n9438), .B(n6209), .ZN(n6210) );
  NAND3_X1 U7724 ( .A1(n6648), .A2(P1_STATE_REG_SCAN_IN), .A3(n6210), .ZN(
        n6211) );
  NOR2_X1 U7725 ( .A1(n6212), .A2(n6211), .ZN(n6216) );
  NAND2_X1 U7726 ( .A1(n8427), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6213) );
  NOR2_X1 U7727 ( .A1(n6102), .A2(n6213), .ZN(n6214) );
  AND2_X1 U7728 ( .A1(n6249), .A2(n6214), .ZN(n10012) );
  AND3_X1 U7729 ( .A1(n10012), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6622), .ZN(
        n6215) );
  AOI211_X1 U7730 ( .C1(P1_REG3_REG_0__SCAN_IN), .C2(P1_U3084), .A(n6216), .B(
        n6215), .ZN(n6217) );
  OAI21_X1 U7731 ( .B1(n10035), .B2(n6218), .A(n6217), .ZN(P1_U3241) );
  INV_X1 U7732 ( .A(n7180), .ZN(n6228) );
  INV_X1 U7733 ( .A(n6759), .ZN(n6750) );
  OAI222_X1 U7734 ( .A1(n8110), .A2(n6228), .B1(n6750), .B2(n7777), .C1(n6219), 
        .C2(n8438), .ZN(P2_U3349) );
  INV_X1 U7735 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6220) );
  NOR2_X1 U7736 ( .A1(n8425), .A2(n6220), .ZN(n6224) );
  INV_X1 U7737 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9505) );
  NOR2_X1 U7738 ( .A1(n8333), .A2(n9505), .ZN(n6223) );
  INV_X1 U7739 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6221) );
  NOR2_X1 U7740 ( .A1(n5996), .A2(n6221), .ZN(n6222) );
  OR3_X1 U7741 ( .A1(n6224), .A2(n6223), .A3(n6222), .ZN(n9507) );
  NAND2_X1 U7742 ( .A1(n9507), .A2(P1_U4006), .ZN(n6225) );
  OAI21_X1 U7743 ( .B1(P1_U4006), .B2(n5624), .A(n6225), .ZN(P1_U3586) );
  OR2_X1 U7744 ( .A1(n4431), .A2(n6320), .ZN(n6226) );
  XNOR2_X1 U7745 ( .A(n6226), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7181) );
  INV_X1 U7746 ( .A(n7181), .ZN(n6667) );
  OAI222_X1 U7747 ( .A1(P1_U3084), .A2(n6667), .B1(n9796), .B2(n6228), .C1(
        n6227), .C2(n9791), .ZN(P1_U3344) );
  NAND2_X1 U7748 ( .A1(n6229), .A2(P1_U4006), .ZN(n6230) );
  OAI21_X1 U7749 ( .B1(P1_U4006), .B2(n4503), .A(n6230), .ZN(P1_U3555) );
  INV_X1 U7750 ( .A(n7185), .ZN(n6234) );
  INV_X1 U7751 ( .A(n6935), .ZN(n6927) );
  OAI222_X1 U7752 ( .A1(n8110), .A2(n6234), .B1(n6927), .B2(n7777), .C1(n6231), 
        .C2(n8438), .ZN(P2_U3348) );
  NAND2_X1 U7753 ( .A1(n4431), .A2(n6232), .ZN(n6241) );
  NAND2_X1 U7754 ( .A1(n6241), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6237) );
  XNOR2_X1 U7755 ( .A(n6237), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7186) );
  INV_X1 U7756 ( .A(n7186), .ZN(n6877) );
  OAI222_X1 U7757 ( .A1(P1_U3084), .A2(n6877), .B1(n9796), .B2(n6234), .C1(
        n6233), .C2(n9791), .ZN(P1_U3343) );
  INV_X1 U7758 ( .A(n7277), .ZN(n6240) );
  INV_X1 U7759 ( .A(n8575), .ZN(n6235) );
  OAI222_X1 U7760 ( .A1(n8110), .A2(n6240), .B1(n6235), .B2(P2_U3152), .C1(
        n6457), .C2(n8438), .ZN(P2_U3347) );
  NAND2_X1 U7761 ( .A1(n6237), .A2(n6236), .ZN(n6238) );
  NAND2_X1 U7762 ( .A1(n6238), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6239) );
  XNOR2_X1 U7763 ( .A(n6239), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9476) );
  INV_X1 U7764 ( .A(n9476), .ZN(n6878) );
  OAI222_X1 U7765 ( .A1(P1_U3084), .A2(n6878), .B1(n9796), .B2(n6240), .C1(
        n6551), .C2(n9791), .ZN(P1_U3342) );
  INV_X1 U7766 ( .A(n7549), .ZN(n6244) );
  NAND2_X1 U7767 ( .A1(n6319), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6242) );
  XNOR2_X1 U7768 ( .A(n6242), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9947) );
  INV_X1 U7769 ( .A(n9791), .ZN(n6704) );
  AOI22_X1 U7770 ( .A1(n9947), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n6704), .ZN(n6243) );
  OAI21_X1 U7771 ( .B1(n6244), .B2(n9796), .A(n6243), .ZN(P1_U3341) );
  INV_X1 U7772 ( .A(n7102), .ZN(n7098) );
  OAI222_X1 U7773 ( .A1(n8438), .A2(n6549), .B1(n9002), .B2(n6244), .C1(
        P2_U3152), .C2(n7098), .ZN(P2_U3346) );
  INV_X1 U7774 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6257) );
  XNOR2_X1 U7775 ( .A(n6251), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n6246) );
  AND2_X1 U7776 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6245) );
  NAND2_X1 U7777 ( .A1(n6246), .A2(n6245), .ZN(n6259) );
  OAI211_X1 U7778 ( .C1(n6246), .C2(n6245), .A(n10012), .B(n6259), .ZN(n6247)
         );
  OAI21_X1 U7779 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n10043), .A(n6247), .ZN(
        n6248) );
  INV_X1 U7780 ( .A(n6248), .ZN(n6256) );
  INV_X1 U7781 ( .A(n6249), .ZN(n6250) );
  OR2_X1 U7782 ( .A1(n8427), .A2(P1_U3084), .ZN(n7774) );
  NOR2_X1 U7783 ( .A1(n6250), .A2(n7774), .ZN(n9475) );
  AND2_X1 U7784 ( .A1(n9475), .A2(n6102), .ZN(n10026) );
  INV_X1 U7785 ( .A(n6251), .ZN(n6278) );
  NOR2_X1 U7786 ( .A1(n6253), .A2(n6647), .ZN(n6277) );
  INV_X1 U7787 ( .A(n9475), .ZN(n6252) );
  OR2_X1 U7788 ( .A1(n6252), .A2(n6102), .ZN(n10020) );
  AOI211_X1 U7789 ( .C1(n6647), .C2(n6253), .A(n6277), .B(n10020), .ZN(n6254)
         );
  AOI21_X1 U7790 ( .B1(n10026), .B2(n6278), .A(n6254), .ZN(n6255) );
  OAI211_X1 U7791 ( .C1(n10035), .C2(n6257), .A(n6256), .B(n6255), .ZN(
        P1_U3242) );
  NAND2_X1 U7792 ( .A1(n9918), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6269) );
  MUX2_X1 U7793 ( .A(n6260), .B(P1_REG1_REG_2__SCAN_IN), .S(n6279), .Z(n6652)
         );
  NAND2_X1 U7794 ( .A1(n6278), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6258) );
  NAND2_X1 U7795 ( .A1(n6259), .A2(n6258), .ZN(n6651) );
  NAND2_X1 U7796 ( .A1(n6652), .A2(n6651), .ZN(n6650) );
  OR2_X1 U7797 ( .A1(n6279), .A2(n6260), .ZN(n6292) );
  NAND2_X1 U7798 ( .A1(n6650), .A2(n6292), .ZN(n6263) );
  MUX2_X1 U7799 ( .A(n6261), .B(P1_REG1_REG_3__SCAN_IN), .S(n6290), .Z(n6262)
         );
  NAND2_X1 U7800 ( .A1(n6263), .A2(n6262), .ZN(n6294) );
  OR2_X1 U7801 ( .A1(n6290), .A2(n6261), .ZN(n6264) );
  AND2_X1 U7802 ( .A1(n6294), .A2(n6264), .ZN(n9906) );
  MUX2_X1 U7803 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9908), .S(n9907), .Z(n6265)
         );
  NAND2_X1 U7804 ( .A1(n9906), .A2(n6265), .ZN(n9912) );
  INV_X1 U7805 ( .A(n9912), .ZN(n6267) );
  NOR2_X1 U7806 ( .A1(n9907), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6266) );
  NOR2_X1 U7807 ( .A1(n6267), .A2(n6266), .ZN(n9923) );
  INV_X1 U7808 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10111) );
  INV_X1 U7809 ( .A(n6269), .ZN(n6268) );
  AOI21_X1 U7810 ( .B1(n10111), .B2(n6276), .A(n6268), .ZN(n9924) );
  NAND2_X1 U7811 ( .A1(n9923), .A2(n9924), .ZN(n9922) );
  NAND2_X1 U7812 ( .A1(n6269), .A2(n9922), .ZN(n6271) );
  AOI22_X1 U7813 ( .A1(n6311), .A2(n6053), .B1(P1_REG1_REG_6__SCAN_IN), .B2(
        n6286), .ZN(n6270) );
  NOR2_X1 U7814 ( .A1(n6271), .A2(n6270), .ZN(n6305) );
  AOI21_X1 U7815 ( .B1(n6271), .B2(n6270), .A(n6305), .ZN(n6273) );
  INV_X1 U7816 ( .A(n10012), .ZN(n10032) );
  INV_X1 U7817 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6272) );
  OAI22_X1 U7818 ( .A1(n6273), .A2(n10032), .B1(n10035), .B2(n6272), .ZN(n6289) );
  NAND2_X1 U7819 ( .A1(n6311), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6274) );
  OAI21_X1 U7820 ( .B1(n6311), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6274), .ZN(
        n6284) );
  XNOR2_X1 U7821 ( .A(n6276), .B(n6275), .ZN(n9920) );
  INV_X1 U7822 ( .A(n6290), .ZN(n6303) );
  INV_X1 U7823 ( .A(n6279), .ZN(n6659) );
  AOI21_X1 U7824 ( .B1(n6278), .B2(P1_REG2_REG_1__SCAN_IN), .A(n6277), .ZN(
        n6656) );
  XOR2_X1 U7825 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6279), .Z(n6655) );
  NOR2_X1 U7826 ( .A1(n6656), .A2(n6655), .ZN(n6654) );
  AOI21_X1 U7827 ( .B1(n6659), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6654), .ZN(
        n6300) );
  INV_X1 U7828 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6280) );
  MUX2_X1 U7829 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6280), .S(n6290), .Z(n6299)
         );
  NOR2_X1 U7830 ( .A1(n6300), .A2(n6299), .ZN(n6298) );
  AOI21_X1 U7831 ( .B1(n6303), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6298), .ZN(
        n9904) );
  NOR2_X1 U7832 ( .A1(n9907), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6281) );
  AOI21_X1 U7833 ( .B1(n9907), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6281), .ZN(
        n9903) );
  NAND2_X1 U7834 ( .A1(n9904), .A2(n9903), .ZN(n9902) );
  OAI21_X1 U7835 ( .B1(n9907), .B2(P1_REG2_REG_4__SCAN_IN), .A(n9902), .ZN(
        n6282) );
  INV_X1 U7836 ( .A(n6282), .ZN(n9919) );
  AOI211_X1 U7837 ( .C1(n6284), .C2(n6283), .A(n10020), .B(n6310), .ZN(n6288)
         );
  INV_X1 U7838 ( .A(n10026), .ZN(n6668) );
  OAI21_X1 U7839 ( .B1(n6668), .B2(n6286), .A(n6285), .ZN(n6287) );
  OR3_X1 U7840 ( .A1(n6289), .A2(n6288), .A3(n6287), .ZN(P1_U3247) );
  MUX2_X1 U7841 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6261), .S(n6290), .Z(n6291)
         );
  NAND3_X1 U7842 ( .A1(n6650), .A2(n6292), .A3(n6291), .ZN(n6293) );
  NAND3_X1 U7843 ( .A1(n10012), .A2(n6294), .A3(n6293), .ZN(n6297) );
  NOR2_X1 U7844 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6295), .ZN(n6870) );
  INV_X1 U7845 ( .A(n6870), .ZN(n6296) );
  NAND2_X1 U7846 ( .A1(n6297), .A2(n6296), .ZN(n6302) );
  AOI211_X1 U7847 ( .C1(n6300), .C2(n6299), .A(n6298), .B(n10020), .ZN(n6301)
         );
  AOI211_X1 U7848 ( .C1(n10026), .C2(n6303), .A(n6302), .B(n6301), .ZN(n6304)
         );
  OAI21_X1 U7849 ( .B1(n10035), .B2(n6548), .A(n6304), .ZN(P1_U3244) );
  NOR2_X1 U7850 ( .A1(n6311), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6306) );
  NOR2_X1 U7851 ( .A1(n6306), .A2(n6305), .ZN(n6308) );
  INV_X1 U7852 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10114) );
  AOI22_X1 U7853 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6309), .B1(n6671), .B2(
        n10114), .ZN(n6307) );
  NOR2_X1 U7854 ( .A1(n6308), .A2(n6307), .ZN(n6664) );
  AOI21_X1 U7855 ( .B1(n6308), .B2(n6307), .A(n6664), .ZN(n6318) );
  INV_X1 U7856 ( .A(n10020), .ZN(n10007) );
  AOI22_X1 U7857 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6671), .B1(n6309), .B2(
        n7072), .ZN(n6313) );
  OAI21_X1 U7858 ( .B1(n6313), .B2(n6312), .A(n6670), .ZN(n6316) );
  INV_X1 U7859 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6395) );
  NAND2_X1 U7860 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7339) );
  NAND2_X1 U7861 ( .A1(n10026), .A2(n6671), .ZN(n6314) );
  OAI211_X1 U7862 ( .C1(n10035), .C2(n6395), .A(n7339), .B(n6314), .ZN(n6315)
         );
  AOI21_X1 U7863 ( .B1(n10007), .B2(n6316), .A(n6315), .ZN(n6317) );
  OAI21_X1 U7864 ( .B1(n6318), .B2(n10032), .A(n6317), .ZN(P1_U3248) );
  INV_X1 U7865 ( .A(n7555), .ZN(n6324) );
  NOR2_X1 U7866 ( .A1(n6319), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6598) );
  OR2_X1 U7867 ( .A1(n6598), .A2(n6320), .ZN(n6321) );
  XNOR2_X1 U7868 ( .A(n6321), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9956) );
  AOI22_X1 U7869 ( .A1(n9956), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n6704), .ZN(n6322) );
  OAI21_X1 U7870 ( .B1(n6324), .B2(n9796), .A(n6322), .ZN(P1_U3340) );
  INV_X1 U7871 ( .A(n7220), .ZN(n7215) );
  OAI222_X1 U7872 ( .A1(n8110), .A2(n6324), .B1(n7215), .B2(P2_U3152), .C1(
        n6323), .C2(n8438), .ZN(P2_U3345) );
  MUX2_X1 U7873 ( .A(n7441), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8567), .Z(n6590)
         );
  NAND2_X1 U7874 ( .A1(keyinput76), .A2(keyinput23), .ZN(n6325) );
  NOR3_X1 U7875 ( .A1(keyinput70), .A2(keyinput6), .A3(n6325), .ZN(n6392) );
  NAND3_X1 U7876 ( .A1(keyinput38), .A2(keyinput69), .A3(keyinput109), .ZN(
        n6326) );
  NOR2_X1 U7877 ( .A1(keyinput77), .A2(n6326), .ZN(n6391) );
  NAND2_X1 U7878 ( .A1(keyinput30), .A2(keyinput27), .ZN(n6327) );
  NOR3_X1 U7879 ( .A1(keyinput106), .A2(keyinput17), .A3(n6327), .ZN(n6328) );
  NAND3_X1 U7880 ( .A1(keyinput35), .A2(keyinput81), .A3(n6328), .ZN(n6338) );
  INV_X1 U7881 ( .A(keyinput94), .ZN(n6329) );
  NOR4_X1 U7882 ( .A1(keyinput114), .A2(keyinput37), .A3(keyinput40), .A4(
        n6329), .ZN(n6336) );
  NAND2_X1 U7883 ( .A1(keyinput127), .A2(keyinput63), .ZN(n6330) );
  NOR3_X1 U7884 ( .A1(keyinput36), .A2(keyinput123), .A3(n6330), .ZN(n6335) );
  INV_X1 U7885 ( .A(keyinput47), .ZN(n6331) );
  NOR4_X1 U7886 ( .A1(keyinput121), .A2(keyinput15), .A3(keyinput25), .A4(
        n6331), .ZN(n6334) );
  NAND2_X1 U7887 ( .A1(keyinput78), .A2(keyinput24), .ZN(n6332) );
  NOR3_X1 U7888 ( .A1(keyinput56), .A2(keyinput72), .A3(n6332), .ZN(n6333) );
  NAND4_X1 U7889 ( .A1(n6336), .A2(n6335), .A3(n6334), .A4(n6333), .ZN(n6337)
         );
  NOR4_X1 U7890 ( .A1(keyinput73), .A2(keyinput115), .A3(n6338), .A4(n6337), 
        .ZN(n6390) );
  INV_X1 U7891 ( .A(keyinput119), .ZN(n6341) );
  INV_X1 U7892 ( .A(keyinput28), .ZN(n6339) );
  NAND4_X1 U7893 ( .A1(keyinput46), .A2(keyinput80), .A3(keyinput29), .A4(
        n6339), .ZN(n6340) );
  NOR4_X1 U7894 ( .A1(keyinput89), .A2(keyinput42), .A3(n6341), .A4(n6340), 
        .ZN(n6354) );
  NAND2_X1 U7895 ( .A1(keyinput51), .A2(keyinput107), .ZN(n6342) );
  NOR3_X1 U7896 ( .A1(keyinput86), .A2(keyinput9), .A3(n6342), .ZN(n6353) );
  INV_X1 U7897 ( .A(keyinput118), .ZN(n6343) );
  NOR4_X1 U7898 ( .A1(keyinput93), .A2(keyinput64), .A3(keyinput79), .A4(n6343), .ZN(n6352) );
  NAND4_X1 U7899 ( .A1(keyinput33), .A2(keyinput90), .A3(keyinput57), .A4(
        keyinput125), .ZN(n6350) );
  NOR2_X1 U7900 ( .A1(keyinput97), .A2(keyinput122), .ZN(n6344) );
  NAND3_X1 U7901 ( .A1(keyinput8), .A2(keyinput53), .A3(n6344), .ZN(n6349) );
  INV_X1 U7902 ( .A(keyinput3), .ZN(n6345) );
  NAND4_X1 U7903 ( .A1(keyinput7), .A2(keyinput85), .A3(keyinput74), .A4(n6345), .ZN(n6348) );
  NOR2_X1 U7904 ( .A1(keyinput75), .A2(keyinput55), .ZN(n6346) );
  NAND3_X1 U7905 ( .A1(keyinput45), .A2(keyinput41), .A3(n6346), .ZN(n6347) );
  NOR4_X1 U7906 ( .A1(n6350), .A2(n6349), .A3(n6348), .A4(n6347), .ZN(n6351)
         );
  NAND4_X1 U7907 ( .A1(n6354), .A2(n6353), .A3(n6352), .A4(n6351), .ZN(n6388)
         );
  NOR4_X1 U7908 ( .A1(keyinput34), .A2(keyinput10), .A3(keyinput88), .A4(
        keyinput16), .ZN(n6368) );
  NAND2_X1 U7909 ( .A1(keyinput60), .A2(keyinput105), .ZN(n6355) );
  NOR3_X1 U7910 ( .A1(keyinput65), .A2(keyinput20), .A3(n6355), .ZN(n6367) );
  NAND2_X1 U7911 ( .A1(keyinput68), .A2(keyinput83), .ZN(n6356) );
  NOR3_X1 U7912 ( .A1(keyinput58), .A2(keyinput71), .A3(n6356), .ZN(n6357) );
  NAND3_X1 U7913 ( .A1(keyinput26), .A2(keyinput120), .A3(n6357), .ZN(n6358)
         );
  NOR3_X1 U7914 ( .A1(keyinput111), .A2(keyinput126), .A3(n6358), .ZN(n6366)
         );
  NAND4_X1 U7915 ( .A1(keyinput31), .A2(keyinput96), .A3(keyinput2), .A4(
        keyinput44), .ZN(n6364) );
  NOR2_X1 U7916 ( .A1(keyinput5), .A2(keyinput84), .ZN(n6359) );
  NAND3_X1 U7917 ( .A1(keyinput117), .A2(keyinput87), .A3(n6359), .ZN(n6363)
         );
  NAND4_X1 U7918 ( .A1(keyinput110), .A2(keyinput32), .A3(keyinput112), .A4(
        keyinput82), .ZN(n6362) );
  NOR2_X1 U7919 ( .A1(keyinput14), .A2(keyinput54), .ZN(n6360) );
  NAND3_X1 U7920 ( .A1(keyinput18), .A2(keyinput124), .A3(n6360), .ZN(n6361)
         );
  NOR4_X1 U7921 ( .A1(n6364), .A2(n6363), .A3(n6362), .A4(n6361), .ZN(n6365)
         );
  NAND4_X1 U7922 ( .A1(n6368), .A2(n6367), .A3(n6366), .A4(n6365), .ZN(n6387)
         );
  NAND3_X1 U7923 ( .A1(keyinput91), .A2(keyinput19), .A3(keyinput104), .ZN(
        n6369) );
  NOR2_X1 U7924 ( .A1(keyinput61), .A2(n6369), .ZN(n6376) );
  NAND2_X1 U7925 ( .A1(keyinput100), .A2(keyinput103), .ZN(n6370) );
  NOR3_X1 U7926 ( .A1(keyinput21), .A2(keyinput50), .A3(n6370), .ZN(n6375) );
  INV_X1 U7927 ( .A(keyinput59), .ZN(n6371) );
  NOR4_X1 U7928 ( .A1(keyinput0), .A2(keyinput22), .A3(keyinput12), .A4(n6371), 
        .ZN(n6374) );
  NAND2_X1 U7929 ( .A1(keyinput66), .A2(keyinput43), .ZN(n6372) );
  NOR3_X1 U7930 ( .A1(keyinput67), .A2(keyinput113), .A3(n6372), .ZN(n6373) );
  NAND4_X1 U7931 ( .A1(n6376), .A2(n6375), .A3(n6374), .A4(n6373), .ZN(n6386)
         );
  NAND2_X1 U7932 ( .A1(keyinput52), .A2(keyinput99), .ZN(n6377) );
  NOR3_X1 U7933 ( .A1(keyinput4), .A2(keyinput62), .A3(n6377), .ZN(n6384) );
  INV_X1 U7934 ( .A(keyinput48), .ZN(n6378) );
  NOR4_X1 U7935 ( .A1(keyinput116), .A2(keyinput39), .A3(keyinput1), .A4(n6378), .ZN(n6383) );
  INV_X1 U7936 ( .A(keyinput49), .ZN(n6379) );
  NOR4_X1 U7937 ( .A1(keyinput92), .A2(keyinput102), .A3(keyinput95), .A4(
        n6379), .ZN(n6382) );
  NAND2_X1 U7938 ( .A1(keyinput98), .A2(keyinput108), .ZN(n6380) );
  NOR3_X1 U7939 ( .A1(keyinput101), .A2(keyinput11), .A3(n6380), .ZN(n6381) );
  NAND4_X1 U7940 ( .A1(n6384), .A2(n6383), .A3(n6382), .A4(n6381), .ZN(n6385)
         );
  NOR4_X1 U7941 ( .A1(n6388), .A2(n6387), .A3(n6386), .A4(n6385), .ZN(n6389)
         );
  NAND4_X1 U7942 ( .A1(n6392), .A2(n6391), .A3(n6390), .A4(n6389), .ZN(n6393)
         );
  AND2_X1 U7943 ( .A1(n6393), .A2(keyinput13), .ZN(n6588) );
  INV_X1 U7944 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7581) );
  AOI22_X1 U7945 ( .A1(n7581), .A2(keyinput16), .B1(keyinput5), .B2(n6395), 
        .ZN(n6394) );
  OAI221_X1 U7946 ( .B1(n7581), .B2(keyinput16), .C1(n6395), .C2(keyinput5), 
        .A(n6394), .ZN(n6405) );
  INV_X1 U7947 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6889) );
  INV_X1 U7948 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6397) );
  AOI22_X1 U7949 ( .A1(n6889), .A2(keyinput20), .B1(keyinput34), .B2(n6397), 
        .ZN(n6396) );
  OAI221_X1 U7950 ( .B1(n6889), .B2(keyinput20), .C1(n6397), .C2(keyinput34), 
        .A(n6396), .ZN(n6404) );
  INV_X1 U7951 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n6399) );
  AOI22_X1 U7952 ( .A1(n6032), .A2(keyinput10), .B1(n6399), .B2(keyinput88), 
        .ZN(n6398) );
  OAI221_X1 U7953 ( .B1(n6032), .B2(keyinput10), .C1(n6399), .C2(keyinput88), 
        .A(n6398), .ZN(n6403) );
  XNOR2_X1 U7954 ( .A(P1_STATE_REG_SCAN_IN), .B(keyinput105), .ZN(n6401) );
  XNOR2_X1 U7955 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput60), .ZN(n6400) );
  NAND2_X1 U7956 ( .A1(n6401), .A2(n6400), .ZN(n6402) );
  NOR4_X1 U7957 ( .A1(n6405), .A2(n6404), .A3(n6403), .A4(n6402), .ZN(n6439)
         );
  AOI22_X1 U7958 ( .A1(n6924), .A2(keyinput117), .B1(n5098), .B2(keyinput31), 
        .ZN(n6406) );
  OAI221_X1 U7959 ( .B1(n6924), .B2(keyinput117), .C1(n5098), .C2(keyinput31), 
        .A(n6406), .ZN(n6415) );
  INV_X1 U7960 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10136) );
  AOI22_X1 U7961 ( .A1(n6408), .A2(keyinput96), .B1(keyinput84), .B2(n10136), 
        .ZN(n6407) );
  OAI221_X1 U7962 ( .B1(n6408), .B2(keyinput96), .C1(n10136), .C2(keyinput84), 
        .A(n6407), .ZN(n6414) );
  INV_X1 U7963 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n8291) );
  INV_X1 U7964 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9981) );
  AOI22_X1 U7965 ( .A1(n8291), .A2(keyinput87), .B1(keyinput2), .B2(n9981), 
        .ZN(n6409) );
  OAI221_X1 U7966 ( .B1(n8291), .B2(keyinput87), .C1(n9981), .C2(keyinput2), 
        .A(n6409), .ZN(n6413) );
  INV_X1 U7967 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10052) );
  AOI22_X1 U7968 ( .A1(n10052), .A2(keyinput44), .B1(keyinput111), .B2(n6411), 
        .ZN(n6410) );
  OAI221_X1 U7969 ( .B1(n10052), .B2(keyinput44), .C1(n6411), .C2(keyinput111), 
        .A(n6410), .ZN(n6412) );
  NOR4_X1 U7970 ( .A1(n6415), .A2(n6414), .A3(n6413), .A4(n6412), .ZN(n6438)
         );
  INV_X1 U7971 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n6417) );
  AOI22_X1 U7972 ( .A1(n6699), .A2(keyinput126), .B1(keyinput26), .B2(n6417), 
        .ZN(n6416) );
  OAI221_X1 U7973 ( .B1(n6699), .B2(keyinput126), .C1(n6417), .C2(keyinput26), 
        .A(n6416), .ZN(n6425) );
  INV_X1 U7974 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7224) );
  AOI22_X1 U7975 ( .A1(n7224), .A2(keyinput120), .B1(n6979), .B2(keyinput83), 
        .ZN(n6418) );
  OAI221_X1 U7976 ( .B1(n7224), .B2(keyinput120), .C1(n6979), .C2(keyinput83), 
        .A(n6418), .ZN(n6424) );
  INV_X1 U7977 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n8227) );
  AOI22_X1 U7978 ( .A1(n8068), .A2(keyinput71), .B1(n8227), .B2(keyinput58), 
        .ZN(n6419) );
  OAI221_X1 U7979 ( .B1(n8068), .B2(keyinput71), .C1(n8227), .C2(keyinput58), 
        .A(n6419), .ZN(n6423) );
  AOI22_X1 U7980 ( .A1(n6421), .A2(keyinput68), .B1(keyinput18), .B2(n5185), 
        .ZN(n6420) );
  OAI221_X1 U7981 ( .B1(n6421), .B2(keyinput68), .C1(n5185), .C2(keyinput18), 
        .A(n6420), .ZN(n6422) );
  NOR4_X1 U7982 ( .A1(n6425), .A2(n6424), .A3(n6423), .A4(n6422), .ZN(n6437)
         );
  INV_X1 U7983 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10018) );
  AOI22_X1 U7984 ( .A1(n10018), .A2(keyinput82), .B1(n7315), .B2(keyinput116), 
        .ZN(n6426) );
  OAI221_X1 U7985 ( .B1(n10018), .B2(keyinput82), .C1(n7315), .C2(keyinput116), 
        .A(n6426), .ZN(n6435) );
  INV_X1 U7986 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10133) );
  AOI22_X1 U7987 ( .A1(n4504), .A2(keyinput54), .B1(keyinput110), .B2(n10133), 
        .ZN(n6427) );
  OAI221_X1 U7988 ( .B1(n4504), .B2(keyinput54), .C1(n10133), .C2(keyinput110), 
        .A(n6427), .ZN(n6434) );
  AOI22_X1 U7989 ( .A1(n4562), .A2(keyinput14), .B1(keyinput124), .B2(n6429), 
        .ZN(n6428) );
  OAI221_X1 U7990 ( .B1(n4562), .B2(keyinput14), .C1(n6429), .C2(keyinput124), 
        .A(n6428), .ZN(n6433) );
  XNOR2_X1 U7991 ( .A(P2_REG2_REG_24__SCAN_IN), .B(keyinput32), .ZN(n6431) );
  XNOR2_X1 U7992 ( .A(P1_REG2_REG_2__SCAN_IN), .B(keyinput112), .ZN(n6430) );
  NAND2_X1 U7993 ( .A1(n6431), .A2(n6430), .ZN(n6432) );
  NOR4_X1 U7994 ( .A1(n6435), .A2(n6434), .A3(n6433), .A4(n6432), .ZN(n6436)
         );
  NAND4_X1 U7995 ( .A1(n6439), .A2(n6438), .A3(n6437), .A4(n6436), .ZN(n6585)
         );
  INV_X1 U7996 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6441) );
  INV_X1 U7997 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7819) );
  AOI22_X1 U7998 ( .A1(n6441), .A2(keyinput52), .B1(n7819), .B2(keyinput101), 
        .ZN(n6440) );
  OAI221_X1 U7999 ( .B1(n6441), .B2(keyinput52), .C1(n7819), .C2(keyinput101), 
        .A(n6440), .ZN(n6451) );
  INV_X1 U8000 ( .A(P2_B_REG_SCAN_IN), .ZN(n6443) );
  AOI22_X1 U8001 ( .A1(n6444), .A2(keyinput48), .B1(keyinput99), .B2(n6443), 
        .ZN(n6442) );
  OAI221_X1 U8002 ( .B1(n6444), .B2(keyinput48), .C1(n6443), .C2(keyinput99), 
        .A(n6442), .ZN(n6450) );
  INV_X1 U8003 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n8226) );
  INV_X1 U8004 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n8242) );
  AOI22_X1 U8005 ( .A1(n8226), .A2(keyinput62), .B1(n8242), .B2(keyinput4), 
        .ZN(n6445) );
  OAI221_X1 U8006 ( .B1(n8226), .B2(keyinput62), .C1(n8242), .C2(keyinput4), 
        .A(n6445), .ZN(n6449) );
  XNOR2_X1 U8007 ( .A(P2_REG1_REG_20__SCAN_IN), .B(keyinput39), .ZN(n6447) );
  XNOR2_X1 U8008 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput1), .ZN(n6446) );
  NAND2_X1 U8009 ( .A1(n6447), .A2(n6446), .ZN(n6448) );
  NOR4_X1 U8010 ( .A1(n6451), .A2(n6450), .A3(n6449), .A4(n6448), .ZN(n6488)
         );
  INV_X1 U8011 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n6453) );
  AOI22_X1 U8012 ( .A1(n6453), .A2(keyinput102), .B1(n4789), .B2(keyinput49), 
        .ZN(n6452) );
  OAI221_X1 U8013 ( .B1(n6453), .B2(keyinput102), .C1(n4789), .C2(keyinput49), 
        .A(n6452), .ZN(n6463) );
  INV_X1 U8014 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9058) );
  INV_X1 U8015 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6455) );
  AOI22_X1 U8016 ( .A1(n9058), .A2(keyinput108), .B1(n6455), .B2(keyinput98), 
        .ZN(n6454) );
  OAI221_X1 U8017 ( .B1(n9058), .B2(keyinput108), .C1(n6455), .C2(keyinput98), 
        .A(n6454), .ZN(n6462) );
  INV_X1 U8018 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6879) );
  AOI22_X1 U8019 ( .A1(n6879), .A2(keyinput11), .B1(n6457), .B2(keyinput92), 
        .ZN(n6456) );
  OAI221_X1 U8020 ( .B1(n6879), .B2(keyinput11), .C1(n6457), .C2(keyinput92), 
        .A(n6456), .ZN(n6461) );
  XOR2_X1 U8021 ( .A(n5266), .B(keyinput95), .Z(n6459) );
  XNOR2_X1 U8022 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput103), .ZN(n6458) );
  NAND2_X1 U8023 ( .A1(n6459), .A2(n6458), .ZN(n6460) );
  NOR4_X1 U8024 ( .A1(n6463), .A2(n6462), .A3(n6461), .A4(n6460), .ZN(n6487)
         );
  AOI22_X1 U8025 ( .A1(n6701), .A2(keyinput21), .B1(keyinput100), .B2(n6260), 
        .ZN(n6464) );
  OAI221_X1 U8026 ( .B1(n6701), .B2(keyinput21), .C1(n6260), .C2(keyinput100), 
        .A(n6464), .ZN(n6474) );
  AOI22_X1 U8027 ( .A1(n8453), .A2(keyinput50), .B1(n8441), .B2(keyinput19), 
        .ZN(n6465) );
  OAI221_X1 U8028 ( .B1(n8453), .B2(keyinput50), .C1(n8441), .C2(keyinput19), 
        .A(n6465), .ZN(n6473) );
  INV_X1 U8029 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10222) );
  AOI22_X1 U8030 ( .A1(n6467), .A2(keyinput104), .B1(keyinput61), .B2(n10222), 
        .ZN(n6466) );
  OAI221_X1 U8031 ( .B1(n6467), .B2(keyinput104), .C1(n10222), .C2(keyinput61), 
        .A(n6466), .ZN(n6472) );
  INV_X1 U8032 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6470) );
  INV_X1 U8033 ( .A(SI_6_), .ZN(n6469) );
  AOI22_X1 U8034 ( .A1(n6470), .A2(keyinput91), .B1(n6469), .B2(keyinput43), 
        .ZN(n6468) );
  OAI221_X1 U8035 ( .B1(n6470), .B2(keyinput91), .C1(n6469), .C2(keyinput43), 
        .A(n6468), .ZN(n6471) );
  NOR4_X1 U8036 ( .A1(n6474), .A2(n6473), .A3(n6472), .A4(n6471), .ZN(n6486)
         );
  INV_X1 U8037 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9493) );
  INV_X1 U8038 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n8198) );
  AOI22_X1 U8039 ( .A1(n9493), .A2(keyinput113), .B1(n8198), .B2(keyinput67), 
        .ZN(n6475) );
  OAI221_X1 U8040 ( .B1(n9493), .B2(keyinput113), .C1(n8198), .C2(keyinput67), 
        .A(n6475), .ZN(n6484) );
  INV_X1 U8041 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9829) );
  AOI22_X1 U8042 ( .A1(n9829), .A2(keyinput66), .B1(keyinput59), .B2(n8066), 
        .ZN(n6476) );
  OAI221_X1 U8043 ( .B1(n9829), .B2(keyinput66), .C1(n8066), .C2(keyinput59), 
        .A(n6476), .ZN(n6483) );
  INV_X1 U8044 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9893) );
  AOI22_X1 U8045 ( .A1(n9893), .A2(keyinput22), .B1(keyinput0), .B2(n6478), 
        .ZN(n6477) );
  OAI221_X1 U8046 ( .B1(n9893), .B2(keyinput22), .C1(n6478), .C2(keyinput0), 
        .A(n6477), .ZN(n6482) );
  INV_X1 U8047 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10056) );
  INV_X1 U8048 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n6480) );
  AOI22_X1 U8049 ( .A1(n10056), .A2(keyinput89), .B1(keyinput12), .B2(n6480), 
        .ZN(n6479) );
  OAI221_X1 U8050 ( .B1(n10056), .B2(keyinput89), .C1(n6480), .C2(keyinput12), 
        .A(n6479), .ZN(n6481) );
  NOR4_X1 U8051 ( .A1(n6484), .A2(n6483), .A3(n6482), .A4(n6481), .ZN(n6485)
         );
  NAND4_X1 U8052 ( .A1(n6488), .A2(n6487), .A3(n6486), .A4(n6485), .ZN(n6584)
         );
  INV_X1 U8053 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10053) );
  AOI22_X1 U8054 ( .A1(n5607), .A2(keyinput6), .B1(n10053), .B2(keyinput63), 
        .ZN(n6489) );
  OAI221_X1 U8055 ( .B1(n5607), .B2(keyinput6), .C1(n10053), .C2(keyinput63), 
        .A(n6489), .ZN(n6499) );
  AOI22_X1 U8056 ( .A1(n4503), .A2(keyinput77), .B1(keyinput69), .B2(n6491), 
        .ZN(n6490) );
  OAI221_X1 U8057 ( .B1(n4503), .B2(keyinput77), .C1(n6491), .C2(keyinput69), 
        .A(n6490), .ZN(n6498) );
  INV_X1 U8058 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8214) );
  AOI22_X1 U8059 ( .A1(n8214), .A2(keyinput70), .B1(n6493), .B2(keyinput76), 
        .ZN(n6492) );
  OAI221_X1 U8060 ( .B1(n8214), .B2(keyinput70), .C1(n6493), .C2(keyinput76), 
        .A(n6492), .ZN(n6497) );
  XNOR2_X1 U8061 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput38), .ZN(n6495) );
  XNOR2_X1 U8062 ( .A(P1_REG1_REG_21__SCAN_IN), .B(keyinput23), .ZN(n6494) );
  NAND2_X1 U8063 ( .A1(n6495), .A2(n6494), .ZN(n6496) );
  NOR4_X1 U8064 ( .A1(n6499), .A2(n6498), .A3(n6497), .A4(n6496), .ZN(n6534)
         );
  INV_X1 U8065 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6886) );
  AOI22_X1 U8066 ( .A1(n6886), .A2(keyinput27), .B1(n8190), .B2(keyinput73), 
        .ZN(n6500) );
  OAI221_X1 U8067 ( .B1(n6886), .B2(keyinput27), .C1(n8190), .C2(keyinput73), 
        .A(n6500), .ZN(n6508) );
  INV_X1 U8068 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8424) );
  AOI22_X1 U8069 ( .A1(n8424), .A2(keyinput81), .B1(n5642), .B2(keyinput106), 
        .ZN(n6501) );
  OAI221_X1 U8070 ( .B1(n8424), .B2(keyinput81), .C1(n5642), .C2(keyinput106), 
        .A(n6501), .ZN(n6507) );
  INV_X1 U8071 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8178) );
  AOI22_X1 U8072 ( .A1(n5479), .A2(keyinput17), .B1(n8178), .B2(keyinput109), 
        .ZN(n6502) );
  OAI221_X1 U8073 ( .B1(n5479), .B2(keyinput17), .C1(n8178), .C2(keyinput109), 
        .A(n6502), .ZN(n6506) );
  INV_X1 U8074 ( .A(SI_18_), .ZN(n6504) );
  AOI22_X1 U8075 ( .A1(n6504), .A2(keyinput115), .B1(n8209), .B2(keyinput30), 
        .ZN(n6503) );
  OAI221_X1 U8076 ( .B1(n6504), .B2(keyinput115), .C1(n8209), .C2(keyinput30), 
        .A(n6503), .ZN(n6505) );
  NOR4_X1 U8077 ( .A1(n6508), .A2(n6507), .A3(n6506), .A4(n6505), .ZN(n6533)
         );
  AOI22_X1 U8078 ( .A1(n5959), .A2(keyinput78), .B1(keyinput121), .B2(n6510), 
        .ZN(n6509) );
  OAI221_X1 U8079 ( .B1(n5959), .B2(keyinput78), .C1(n6510), .C2(keyinput121), 
        .A(n6509), .ZN(n6519) );
  INV_X1 U8080 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n6512) );
  AOI22_X1 U8081 ( .A1(n6513), .A2(keyinput72), .B1(keyinput56), .B2(n6512), 
        .ZN(n6511) );
  OAI221_X1 U8082 ( .B1(n6513), .B2(keyinput72), .C1(n6512), .C2(keyinput56), 
        .A(n6511), .ZN(n6518) );
  INV_X1 U8083 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10054) );
  AOI22_X1 U8084 ( .A1(n10054), .A2(keyinput47), .B1(keyinput65), .B2(n6784), 
        .ZN(n6514) );
  OAI221_X1 U8085 ( .B1(n10054), .B2(keyinput47), .C1(n6784), .C2(keyinput65), 
        .A(n6514), .ZN(n6517) );
  INV_X1 U8086 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10036) );
  AOI22_X1 U8087 ( .A1(n10036), .A2(keyinput15), .B1(n6601), .B2(keyinput25), 
        .ZN(n6515) );
  OAI221_X1 U8088 ( .B1(n10036), .B2(keyinput15), .C1(n6601), .C2(keyinput25), 
        .A(n6515), .ZN(n6516) );
  NOR4_X1 U8089 ( .A1(n6519), .A2(n6518), .A3(n6517), .A4(n6516), .ZN(n6532)
         );
  INV_X1 U8090 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10137) );
  INV_X1 U8091 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9123) );
  AOI22_X1 U8092 ( .A1(n10137), .A2(keyinput36), .B1(n9123), .B2(keyinput127), 
        .ZN(n6520) );
  OAI221_X1 U8093 ( .B1(n10137), .B2(keyinput36), .C1(n9123), .C2(keyinput127), 
        .A(n6520), .ZN(n6530) );
  INV_X1 U8094 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10055) );
  AOI22_X1 U8095 ( .A1(n6522), .A2(keyinput37), .B1(n10055), .B2(keyinput94), 
        .ZN(n6521) );
  OAI221_X1 U8096 ( .B1(n6522), .B2(keyinput37), .C1(n10055), .C2(keyinput94), 
        .A(n6521), .ZN(n6529) );
  INV_X1 U8097 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10134) );
  AOI22_X1 U8098 ( .A1(n10134), .A2(keyinput123), .B1(n6524), .B2(keyinput114), 
        .ZN(n6523) );
  OAI221_X1 U8099 ( .B1(n10134), .B2(keyinput123), .C1(n6524), .C2(keyinput114), .A(n6523), .ZN(n6528) );
  XOR2_X1 U8100 ( .A(n5756), .B(keyinput24), .Z(n6526) );
  XNOR2_X1 U8101 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput40), .ZN(n6525) );
  NAND2_X1 U8102 ( .A1(n6526), .A2(n6525), .ZN(n6527) );
  NOR4_X1 U8103 ( .A1(n6530), .A2(n6529), .A3(n6528), .A4(n6527), .ZN(n6531)
         );
  NAND4_X1 U8104 ( .A1(n6534), .A2(n6533), .A3(n6532), .A4(n6531), .ZN(n6583)
         );
  AOI22_X1 U8105 ( .A1(n8169), .A2(keyinput125), .B1(keyinput97), .B2(n6716), 
        .ZN(n6535) );
  OAI221_X1 U8106 ( .B1(n8169), .B2(keyinput125), .C1(n6716), .C2(keyinput97), 
        .A(n6535), .ZN(n6544) );
  INV_X1 U8107 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n10135) );
  AOI22_X1 U8108 ( .A1(n5152), .A2(keyinput122), .B1(n10135), .B2(keyinput33), 
        .ZN(n6536) );
  OAI221_X1 U8109 ( .B1(n5152), .B2(keyinput122), .C1(n10135), .C2(keyinput33), 
        .A(n6536), .ZN(n6543) );
  INV_X1 U8110 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n7835) );
  AOI22_X1 U8111 ( .A1(n7835), .A2(keyinput90), .B1(keyinput57), .B2(n8536), 
        .ZN(n6537) );
  OAI221_X1 U8112 ( .B1(n7835), .B2(keyinput90), .C1(n8536), .C2(keyinput57), 
        .A(n6537), .ZN(n6542) );
  INV_X1 U8113 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n6538) );
  XOR2_X1 U8114 ( .A(n6538), .B(keyinput53), .Z(n6540) );
  XNOR2_X1 U8115 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput93), .ZN(n6539) );
  NAND2_X1 U8116 ( .A1(n6540), .A2(n6539), .ZN(n6541) );
  NOR4_X1 U8117 ( .A1(n6544), .A2(n6543), .A3(n6542), .A4(n6541), .ZN(n6581)
         );
  INV_X1 U8118 ( .A(keyinput13), .ZN(n6546) );
  XNOR2_X1 U8119 ( .A(P1_REG0_REG_20__SCAN_IN), .B(keyinput80), .ZN(n6545) );
  OAI21_X1 U8120 ( .B1(P1_REG1_REG_1__SCAN_IN), .B2(n6546), .A(n6545), .ZN(
        n6556) );
  INV_X1 U8121 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6548) );
  AOI22_X1 U8122 ( .A1(n6549), .A2(keyinput42), .B1(keyinput119), .B2(n6548), 
        .ZN(n6547) );
  OAI221_X1 U8123 ( .B1(n6549), .B2(keyinput42), .C1(n6548), .C2(keyinput119), 
        .A(n6547), .ZN(n6555) );
  AOI22_X1 U8124 ( .A1(n7998), .A2(keyinput28), .B1(n6551), .B2(keyinput8), 
        .ZN(n6550) );
  OAI221_X1 U8125 ( .B1(n7998), .B2(keyinput28), .C1(n6551), .C2(keyinput8), 
        .A(n6550), .ZN(n6554) );
  INV_X1 U8126 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10051) );
  INV_X1 U8127 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6613) );
  AOI22_X1 U8128 ( .A1(n10051), .A2(keyinput46), .B1(keyinput29), .B2(n6613), 
        .ZN(n6552) );
  OAI221_X1 U8129 ( .B1(n10051), .B2(keyinput46), .C1(n6613), .C2(keyinput29), 
        .A(n6552), .ZN(n6553) );
  NOR4_X1 U8130 ( .A1(n6556), .A2(n6555), .A3(n6554), .A4(n6553), .ZN(n6580)
         );
  INV_X1 U8131 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n8241) );
  INV_X1 U8132 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10161) );
  AOI22_X1 U8133 ( .A1(n8241), .A2(keyinput55), .B1(keyinput75), .B2(n10161), 
        .ZN(n6557) );
  OAI221_X1 U8134 ( .B1(n8241), .B2(keyinput55), .C1(n10161), .C2(keyinput75), 
        .A(n6557), .ZN(n6565) );
  AOI22_X1 U8135 ( .A1(n6712), .A2(keyinput41), .B1(n7231), .B2(keyinput85), 
        .ZN(n6558) );
  OAI221_X1 U8136 ( .B1(n6712), .B2(keyinput41), .C1(n7231), .C2(keyinput85), 
        .A(n6558), .ZN(n6564) );
  INV_X1 U8137 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10097) );
  XOR2_X1 U8138 ( .A(n10097), .B(keyinput35), .Z(n6561) );
  XNOR2_X1 U8139 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput3), .ZN(n6560) );
  XNOR2_X1 U8140 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput7), .ZN(n6559) );
  NAND3_X1 U8141 ( .A1(n6561), .A2(n6560), .A3(n6559), .ZN(n6563) );
  INV_X1 U8142 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10050) );
  XNOR2_X1 U8143 ( .A(n10050), .B(keyinput74), .ZN(n6562) );
  NOR4_X1 U8144 ( .A1(n6565), .A2(n6564), .A3(n6563), .A4(n6562), .ZN(n6579)
         );
  INV_X1 U8145 ( .A(SI_21_), .ZN(n6567) );
  INV_X1 U8146 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10132) );
  AOI22_X1 U8147 ( .A1(n6567), .A2(keyinput9), .B1(keyinput86), .B2(n10132), 
        .ZN(n6566) );
  OAI221_X1 U8148 ( .B1(n6567), .B2(keyinput9), .C1(n10132), .C2(keyinput86), 
        .A(n6566), .ZN(n6577) );
  INV_X1 U8149 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9135) );
  INV_X1 U8150 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6569) );
  AOI22_X1 U8151 ( .A1(n9135), .A2(keyinput51), .B1(keyinput45), .B2(n6569), 
        .ZN(n6568) );
  OAI221_X1 U8152 ( .B1(n9135), .B2(keyinput51), .C1(n6569), .C2(keyinput45), 
        .A(n6568), .ZN(n6576) );
  AOI22_X1 U8153 ( .A1(n6925), .A2(keyinput64), .B1(n6571), .B2(keyinput118), 
        .ZN(n6570) );
  OAI221_X1 U8154 ( .B1(n6925), .B2(keyinput64), .C1(n6571), .C2(keyinput118), 
        .A(n6570), .ZN(n6575) );
  XNOR2_X1 U8155 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput107), .ZN(n6573) );
  XNOR2_X1 U8156 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput79), .ZN(n6572) );
  NAND2_X1 U8157 ( .A1(n6573), .A2(n6572), .ZN(n6574) );
  NOR4_X1 U8158 ( .A1(n6577), .A2(n6576), .A3(n6575), .A4(n6574), .ZN(n6578)
         );
  NAND4_X1 U8159 ( .A1(n6581), .A2(n6580), .A3(n6579), .A4(n6578), .ZN(n6582)
         );
  NOR4_X1 U8160 ( .A1(n6585), .A2(n6584), .A3(n6583), .A4(n6582), .ZN(n6586)
         );
  OAI21_X1 U8161 ( .B1(n6588), .B2(n6587), .A(n6586), .ZN(n6589) );
  XNOR2_X1 U8162 ( .A(n6590), .B(n6589), .ZN(P2_U3553) );
  OR2_X1 U8163 ( .A1(n10130), .A2(n6591), .ZN(n6595) );
  NAND2_X1 U8164 ( .A1(n10130), .A2(n7300), .ZN(n6593) );
  NAND2_X1 U8165 ( .A1(n6593), .A2(n6592), .ZN(n6594) );
  AND2_X1 U8166 ( .A1(n6595), .A2(n6594), .ZN(n8588) );
  NOR2_X1 U8167 ( .A1(n10124), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8168 ( .A(n7567), .ZN(n6602) );
  INV_X1 U8169 ( .A(n7330), .ZN(n7327) );
  OAI222_X1 U8170 ( .A1(n8110), .A2(n6602), .B1(n7327), .B2(n7777), .C1(n6596), 
        .C2(n8438), .ZN(P2_U3344) );
  INV_X1 U8171 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6597) );
  NAND2_X1 U8172 ( .A1(n6598), .A2(n6597), .ZN(n6682) );
  NAND2_X1 U8173 ( .A1(n6682), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U8174 ( .A1(n6599), .A2(n6680), .ZN(n6697) );
  OR2_X1 U8175 ( .A1(n6599), .A2(n6680), .ZN(n6600) );
  NAND2_X1 U8176 ( .A1(n6697), .A2(n6600), .ZN(n9483) );
  OAI222_X1 U8177 ( .A1(P1_U3084), .A2(n9483), .B1(n9796), .B2(n6602), .C1(
        n6601), .C2(n9791), .ZN(P1_U3339) );
  INV_X1 U8178 ( .A(n9144), .ZN(n9131) );
  INV_X1 U8179 ( .A(n6904), .ZN(n6638) );
  AND2_X1 U8180 ( .A1(n6690), .A2(n6603), .ZN(n6790) );
  INV_X1 U8181 ( .A(n6790), .ZN(n6692) );
  AOI22_X1 U8182 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n6692), .B1(n9139), .B2(
        n4400), .ZN(n6608) );
  OAI21_X1 U8183 ( .B1(n6604), .B2(n6606), .A(n6605), .ZN(n6646) );
  INV_X1 U8184 ( .A(n9146), .ZN(n9119) );
  NAND2_X1 U8185 ( .A1(n6646), .A2(n9119), .ZN(n6607) );
  OAI211_X1 U8186 ( .C1(n9131), .C2(n6638), .A(n6608), .B(n6607), .ZN(P1_U3230) );
  INV_X1 U8187 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6610) );
  NAND2_X1 U8188 ( .A1(n5875), .A2(P2_U3966), .ZN(n6609) );
  OAI21_X1 U8189 ( .B1(n6610), .B2(P2_U3966), .A(n6609), .ZN(P2_U3552) );
  INV_X1 U8190 ( .A(n6611), .ZN(n8047) );
  NAND2_X1 U8191 ( .A1(n8047), .A2(P2_U3966), .ZN(n6612) );
  OAI21_X1 U8192 ( .B1(n6613), .B2(P2_U3966), .A(n6612), .ZN(P2_U3583) );
  OR2_X1 U8193 ( .A1(n6615), .A2(n6614), .ZN(n6895) );
  INV_X1 U8194 ( .A(n9499), .ZN(n10039) );
  INV_X1 U8195 ( .A(n7142), .ZN(n9396) );
  OAI21_X1 U8196 ( .B1(n10065), .B2(n5948), .A(n6896), .ZN(n6616) );
  NOR2_X1 U8197 ( .A1(n6895), .A2(n6616), .ZN(n6642) );
  AND2_X2 U8198 ( .A1(n6642), .A2(n6897), .ZN(n10117) );
  NOR2_X1 U8199 ( .A1(n6229), .A2(n6638), .ZN(n6631) );
  AND2_X1 U8200 ( .A1(n6229), .A2(n6638), .ZN(n9398) );
  NOR2_X1 U8201 ( .A1(n6631), .A2(n9398), .ZN(n9165) );
  OR3_X1 U8202 ( .A1(n9165), .A2(n6618), .A3(n6617), .ZN(n6620) );
  OR2_X1 U8203 ( .A1(n9390), .A2(n9438), .ZN(n9599) );
  NAND2_X1 U8204 ( .A1(n4400), .A2(n9867), .ZN(n6619) );
  AND2_X1 U8205 ( .A1(n6620), .A2(n6619), .ZN(n6907) );
  OAI21_X1 U8206 ( .B1(n6638), .B2(n6637), .A(n6907), .ZN(n6643) );
  NAND2_X1 U8207 ( .A1(n6643), .A2(n10117), .ZN(n6621) );
  OAI21_X1 U8208 ( .B1(n10117), .B2(n6622), .A(n6621), .ZN(P1_U3523) );
  AND2_X1 U8209 ( .A1(n6229), .A2(n6904), .ZN(n6623) );
  NAND2_X1 U8210 ( .A1(n6630), .A2(n6623), .ZN(n6944) );
  OAI21_X1 U8211 ( .B1(n6630), .B2(n6623), .A(n6944), .ZN(n10038) );
  OR2_X1 U8212 ( .A1(n6625), .A2(n6624), .ZN(n6628) );
  OR2_X1 U8213 ( .A1(n6626), .A2(n9190), .ZN(n6627) );
  AND2_X1 U8214 ( .A1(n6628), .A2(n6627), .ZN(n9680) );
  AOI22_X1 U8215 ( .A1(n9461), .A2(n9867), .B1(n9865), .B2(n6229), .ZN(n6636)
         );
  NAND2_X1 U8216 ( .A1(n9442), .A2(n10039), .ZN(n6633) );
  NAND2_X1 U8217 ( .A1(n5948), .A2(n9396), .ZN(n6632) );
  NAND2_X1 U8218 ( .A1(n6633), .A2(n6632), .ZN(n9870) );
  NAND2_X1 U8219 ( .A1(n6634), .A2(n9870), .ZN(n6635) );
  OAI211_X1 U8220 ( .C1(n10038), .C2(n9680), .A(n6636), .B(n6635), .ZN(n10047)
         );
  INV_X1 U8221 ( .A(n10101), .ZN(n9881) );
  NAND2_X1 U8222 ( .A1(n10045), .A2(n6638), .ZN(n6988) );
  OAI211_X1 U8223 ( .C1(n6638), .C2(n10045), .A(n9881), .B(n6988), .ZN(n10037)
         );
  OR2_X1 U8224 ( .A1(n10045), .A2(n10093), .ZN(n6689) );
  OAI211_X1 U8225 ( .C1(n10038), .C2(n10065), .A(n10037), .B(n6689), .ZN(n6639) );
  NOR2_X1 U8226 ( .A1(n10047), .A2(n6639), .ZN(n10059) );
  NAND2_X1 U8227 ( .A1(n4906), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6640) );
  OAI21_X1 U8228 ( .B1(n10059), .B2(n4906), .A(n6640), .ZN(P1_U3524) );
  INV_X1 U8229 ( .A(n6897), .ZN(n6641) );
  AND2_X2 U8230 ( .A1(n6642), .A2(n6641), .ZN(n10107) );
  INV_X1 U8231 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6645) );
  NAND2_X1 U8232 ( .A1(n6643), .A2(n10107), .ZN(n6644) );
  OAI21_X1 U8233 ( .B1(n10107), .B2(n6645), .A(n6644), .ZN(P1_U3454) );
  INV_X1 U8234 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6661) );
  MUX2_X1 U8235 ( .A(n6647), .B(n6646), .S(n8427), .Z(n6649) );
  OAI211_X1 U8236 ( .C1(n6649), .C2(n6102), .A(P1_U4006), .B(n6648), .ZN(n9915) );
  OAI211_X1 U8237 ( .C1(n6652), .C2(n6651), .A(n10012), .B(n6650), .ZN(n6653)
         );
  OAI21_X1 U8238 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6789), .A(n6653), .ZN(n6658) );
  AOI211_X1 U8239 ( .C1(n6656), .C2(n6655), .A(n6654), .B(n10020), .ZN(n6657)
         );
  AOI211_X1 U8240 ( .C1(n10026), .C2(n6659), .A(n6658), .B(n6657), .ZN(n6660)
         );
  OAI211_X1 U8241 ( .C1(n6661), .C2(n10035), .A(n9915), .B(n6660), .ZN(
        P1_U3243) );
  MUX2_X1 U8242 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6662), .S(n9929), .Z(n9936)
         );
  NOR2_X1 U8243 ( .A1(n6671), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6663) );
  NOR2_X1 U8244 ( .A1(n6664), .A2(n6663), .ZN(n9937) );
  NAND2_X1 U8245 ( .A1(n9936), .A2(n9937), .ZN(n9935) );
  OAI21_X1 U8246 ( .B1(n6662), .B2(n6669), .A(n9935), .ZN(n6666) );
  AOI22_X1 U8247 ( .A1(n7181), .A2(n6157), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6667), .ZN(n6665) );
  NOR2_X1 U8248 ( .A1(n6666), .A2(n6665), .ZN(n6767) );
  AOI21_X1 U8249 ( .B1(n6666), .B2(n6665), .A(n6767), .ZN(n6678) );
  INV_X1 U8250 ( .A(n10035), .ZN(n9930) );
  OAI22_X1 U8251 ( .A1(n6668), .A2(n6667), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7460), .ZN(n6676) );
  AOI22_X1 U8252 ( .A1(n9929), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7090), .B2(
        n6669), .ZN(n9932) );
  OAI21_X1 U8253 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6671), .A(n6670), .ZN(
        n9933) );
  NAND2_X1 U8254 ( .A1(n9932), .A2(n9933), .ZN(n9931) );
  OAI21_X1 U8255 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9929), .A(n9931), .ZN(
        n6674) );
  NAND2_X1 U8256 ( .A1(n7181), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6672) );
  OAI21_X1 U8257 ( .B1(n7181), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6672), .ZN(
        n6673) );
  NOR2_X1 U8258 ( .A1(n6673), .A2(n6674), .ZN(n6773) );
  AOI211_X1 U8259 ( .C1(n6674), .C2(n6673), .A(n6773), .B(n10020), .ZN(n6675)
         );
  AOI211_X1 U8260 ( .C1(n9930), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n6676), .B(
        n6675), .ZN(n6677) );
  OAI21_X1 U8261 ( .B1(n6678), .B2(n10032), .A(n6677), .ZN(P1_U3250) );
  INV_X1 U8262 ( .A(n7829), .ZN(n6702) );
  INV_X1 U8263 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6679) );
  NAND2_X1 U8264 ( .A1(n6680), .A2(n6679), .ZN(n6681) );
  OR2_X1 U8265 ( .A1(n6682), .A2(n6681), .ZN(n6703) );
  NAND2_X1 U8266 ( .A1(n6703), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6683) );
  XNOR2_X1 U8267 ( .A(n6683), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9996) );
  AOI22_X1 U8268 ( .A1(n9996), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n6704), .ZN(n6684) );
  OAI21_X1 U8269 ( .B1(n6702), .B2(n9796), .A(n6684), .ZN(P1_U3337) );
  INV_X1 U8270 ( .A(n6685), .ZN(n6686) );
  AOI21_X1 U8271 ( .B1(n6688), .B2(n6687), .A(n6686), .ZN(n6695) );
  INV_X1 U8272 ( .A(n6689), .ZN(n6691) );
  AOI22_X1 U8273 ( .A1(n9139), .A2(n9461), .B1(n6691), .B2(n6690), .ZN(n6694)
         );
  INV_X1 U8274 ( .A(n9137), .ZN(n9128) );
  AOI22_X1 U8275 ( .A1(n9128), .A2(n6229), .B1(n6692), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6693) );
  OAI211_X1 U8276 ( .C1(n6695), .C2(n9146), .A(n6694), .B(n6693), .ZN(P1_U3220) );
  INV_X1 U8277 ( .A(n7748), .ZN(n6700) );
  INV_X1 U8278 ( .A(n8053), .ZN(n8063) );
  OAI222_X1 U8279 ( .A1(n8438), .A2(n6696), .B1(n9002), .B2(n6700), .C1(n7777), 
        .C2(n8063), .ZN(P2_U3343) );
  NAND2_X1 U8280 ( .A1(n6697), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6698) );
  XNOR2_X1 U8281 ( .A(n6698), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9986) );
  INV_X1 U8282 ( .A(n9986), .ZN(n9485) );
  OAI222_X1 U8283 ( .A1(n9485), .A2(P1_U3084), .B1(n7925), .B2(n6700), .C1(
        n6699), .C2(n9791), .ZN(P1_U3338) );
  INV_X1 U8284 ( .A(n8594), .ZN(n8067) );
  OAI222_X1 U8285 ( .A1(n8110), .A2(n6702), .B1(n8067), .B2(P2_U3152), .C1(
        n6701), .C2(n8438), .ZN(P2_U3342) );
  INV_X1 U8286 ( .A(n7904), .ZN(n6785) );
  OAI21_X1 U8287 ( .B1(n6703), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6909) );
  XNOR2_X1 U8288 ( .A(n6909), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10008) );
  AOI22_X1 U8289 ( .A1(n10008), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n6704), .ZN(n6705) );
  OAI21_X1 U8290 ( .B1(n6785), .B2(n9796), .A(n6705), .ZN(P1_U3336) );
  NAND2_X1 U8291 ( .A1(n6706), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6707) );
  OAI211_X1 U8292 ( .C1(n10130), .C2(n6708), .A(n7300), .B(n6707), .ZN(n6727)
         );
  NAND2_X1 U8293 ( .A1(n6727), .A2(n5210), .ZN(n6709) );
  NAND2_X1 U8294 ( .A1(n6709), .A2(n8567), .ZN(n6745) );
  AND2_X1 U8295 ( .A1(n6745), .A2(n5763), .ZN(n9815) );
  INV_X1 U8296 ( .A(n6710), .ZN(n6731) );
  MUX2_X1 U8297 ( .A(n6711), .B(P2_REG1_REG_8__SCAN_IN), .S(n6863), .Z(n6859)
         );
  MUX2_X1 U8298 ( .A(n6712), .B(P2_REG1_REG_7__SCAN_IN), .S(n6852), .Z(n6848)
         );
  NAND2_X1 U8299 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(n6741), .ZN(n6723) );
  MUX2_X1 U8300 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6713), .S(n6741), .Z(n6812)
         );
  NAND2_X1 U8301 ( .A1(n6739), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6722) );
  MUX2_X1 U8302 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6714), .S(n6739), .Z(n6836)
         );
  NAND2_X1 U8303 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(n6737), .ZN(n6721) );
  MUX2_X1 U8304 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6715), .S(n6737), .Z(n6801)
         );
  MUX2_X1 U8305 ( .A(n6716), .B(P2_REG1_REG_3__SCAN_IN), .S(n6828), .Z(n6824)
         );
  NAND2_X1 U8306 ( .A1(n9814), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6720) );
  MUX2_X1 U8307 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6717), .S(n9814), .Z(n9817)
         );
  NAND2_X1 U8308 ( .A1(P2_REG1_REG_1__SCAN_IN), .A2(n9803), .ZN(n6719) );
  MUX2_X1 U8309 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6718), .S(n9803), .Z(n9805)
         );
  NAND3_X1 U8310 ( .A1(n10129), .A2(P2_REG1_REG_0__SCAN_IN), .A3(n9805), .ZN(
        n9804) );
  NAND2_X1 U8311 ( .A1(n6719), .A2(n9804), .ZN(n9818) );
  NAND2_X1 U8312 ( .A1(n9817), .A2(n9818), .ZN(n9816) );
  NAND2_X1 U8313 ( .A1(n6720), .A2(n9816), .ZN(n6825) );
  NAND2_X1 U8314 ( .A1(n6824), .A2(n6825), .ZN(n6823) );
  OAI21_X1 U8315 ( .B1(n6828), .B2(n6716), .A(n6823), .ZN(n6800) );
  NAND2_X1 U8316 ( .A1(n6801), .A2(n6800), .ZN(n6799) );
  NAND2_X1 U8317 ( .A1(n6721), .A2(n6799), .ZN(n6837) );
  NAND2_X1 U8318 ( .A1(n6836), .A2(n6837), .ZN(n6835) );
  NAND2_X1 U8319 ( .A1(n6722), .A2(n6835), .ZN(n6813) );
  NAND2_X1 U8320 ( .A1(n6812), .A2(n6813), .ZN(n6811) );
  NAND2_X1 U8321 ( .A1(n6723), .A2(n6811), .ZN(n6849) );
  NAND2_X1 U8322 ( .A1(n6848), .A2(n6849), .ZN(n6847) );
  OAI21_X1 U8323 ( .B1(n6852), .B2(n6712), .A(n6847), .ZN(n6860) );
  NAND2_X1 U8324 ( .A1(n6859), .A2(n6860), .ZN(n6858) );
  INV_X1 U8325 ( .A(n6858), .ZN(n6724) );
  AOI21_X1 U8326 ( .B1(n6725), .B2(P2_REG1_REG_8__SCAN_IN), .A(n6724), .ZN(
        n6729) );
  INV_X1 U8327 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7388) );
  MUX2_X1 U8328 ( .A(n7388), .B(P2_REG1_REG_9__SCAN_IN), .S(n6759), .Z(n6728)
         );
  NOR2_X1 U8329 ( .A1(n6728), .A2(n6729), .ZN(n6751) );
  AND2_X1 U8330 ( .A1(n5210), .A2(n8044), .ZN(n6726) );
  INV_X1 U8331 ( .A(n10119), .ZN(n8611) );
  AOI211_X1 U8332 ( .C1(n6729), .C2(n6728), .A(n6751), .B(n8611), .ZN(n6730)
         );
  AOI211_X1 U8333 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n10124), .A(n6731), .B(
        n6730), .ZN(n6749) );
  XNOR2_X1 U8334 ( .A(n6759), .B(n6732), .ZN(n6747) );
  INV_X1 U8335 ( .A(n6828), .ZN(n6735) );
  INV_X1 U8336 ( .A(n10129), .ZN(n10127) );
  AOI21_X1 U8337 ( .B1(n9803), .B2(P2_REG2_REG_1__SCAN_IN), .A(n9799), .ZN(
        n9812) );
  NAND2_X1 U8338 ( .A1(n9814), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6733) );
  OAI21_X1 U8339 ( .B1(n9814), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6733), .ZN(
        n9811) );
  NOR2_X1 U8340 ( .A1(n9812), .A2(n9811), .ZN(n9810) );
  INV_X1 U8341 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6734) );
  MUX2_X1 U8342 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6734), .S(n6828), .Z(n6820)
         );
  NOR2_X1 U8343 ( .A1(n6821), .A2(n6820), .ZN(n6819) );
  AOI21_X1 U8344 ( .B1(n6735), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6819), .ZN(
        n6797) );
  NAND2_X1 U8345 ( .A1(P2_REG2_REG_4__SCAN_IN), .A2(n6737), .ZN(n6736) );
  OAI21_X1 U8346 ( .B1(n6737), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6736), .ZN(
        n6796) );
  NOR2_X1 U8347 ( .A1(n6797), .A2(n6796), .ZN(n6795) );
  AOI21_X1 U8348 ( .B1(n6737), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6795), .ZN(
        n6833) );
  NAND2_X1 U8349 ( .A1(n6739), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6738) );
  OAI21_X1 U8350 ( .B1(n6739), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6738), .ZN(
        n6832) );
  NAND2_X1 U8351 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(n6741), .ZN(n6740) );
  OAI21_X1 U8352 ( .B1(n6741), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6740), .ZN(
        n6808) );
  INV_X1 U8353 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6742) );
  MUX2_X1 U8354 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6742), .S(n6852), .Z(n6844)
         );
  NOR2_X1 U8355 ( .A1(n6845), .A2(n6844), .ZN(n6843) );
  MUX2_X1 U8356 ( .A(n5261), .B(P2_REG2_REG_8__SCAN_IN), .S(n6863), .Z(n6743)
         );
  INV_X1 U8357 ( .A(n6743), .ZN(n6856) );
  NOR2_X1 U8358 ( .A1(n5763), .A2(n8044), .ZN(n6744) );
  NAND2_X1 U8359 ( .A1(n6745), .A2(n6744), .ZN(n10122) );
  INV_X1 U8360 ( .A(n10122), .ZN(n10118) );
  NAND2_X1 U8361 ( .A1(n6747), .A2(n6746), .ZN(n6761) );
  OAI211_X1 U8362 ( .C1(n6747), .C2(n6746), .A(n10118), .B(n6761), .ZN(n6748)
         );
  OAI211_X1 U8363 ( .C1(n10121), .C2(n6750), .A(n6749), .B(n6748), .ZN(
        P2_U3254) );
  NAND2_X1 U8364 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(n7777), .ZN(n7270) );
  INV_X1 U8365 ( .A(n7270), .ZN(n6756) );
  AOI21_X1 U8366 ( .B1(n6759), .B2(P2_REG1_REG_9__SCAN_IN), .A(n6751), .ZN(
        n6754) );
  INV_X1 U8367 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10213) );
  MUX2_X1 U8368 ( .A(n10213), .B(P2_REG1_REG_10__SCAN_IN), .S(n6935), .Z(n6753) );
  OR2_X1 U8369 ( .A1(n6754), .A2(n6753), .ZN(n6926) );
  INV_X1 U8370 ( .A(n6926), .ZN(n6752) );
  AOI211_X1 U8371 ( .C1(n6754), .C2(n6753), .A(n6752), .B(n8611), .ZN(n6755)
         );
  AOI211_X1 U8372 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n10124), .A(n6756), .B(
        n6755), .ZN(n6766) );
  OR2_X1 U8373 ( .A1(n6935), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6758) );
  NAND2_X1 U8374 ( .A1(n6935), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6757) );
  AND2_X1 U8375 ( .A1(n6758), .A2(n6757), .ZN(n6764) );
  NAND2_X1 U8376 ( .A1(n6759), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6760) );
  NAND2_X1 U8377 ( .A1(n6761), .A2(n6760), .ZN(n6763) );
  INV_X1 U8378 ( .A(n6934), .ZN(n6762) );
  OAI211_X1 U8379 ( .C1(n6764), .C2(n6763), .A(n10118), .B(n6762), .ZN(n6765)
         );
  OAI211_X1 U8380 ( .C1(n10121), .C2(n6927), .A(n6766), .B(n6765), .ZN(
        P2_U3255) );
  NOR2_X1 U8381 ( .A1(n7181), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6768) );
  NOR2_X1 U8382 ( .A1(n6768), .A2(n6767), .ZN(n6770) );
  AOI22_X1 U8383 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6877), .B1(n7186), .B2(
        n9829), .ZN(n6769) );
  NOR2_X1 U8384 ( .A1(n6770), .A2(n6769), .ZN(n6876) );
  AOI21_X1 U8385 ( .B1(n6770), .B2(n6769), .A(n6876), .ZN(n6783) );
  OR2_X1 U8386 ( .A1(n7186), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6772) );
  NAND2_X1 U8387 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n7186), .ZN(n6771) );
  NAND2_X1 U8388 ( .A1(n6772), .A2(n6771), .ZN(n6775) );
  AOI21_X1 U8389 ( .B1(n6775), .B2(n6774), .A(n6883), .ZN(n6776) );
  NAND2_X1 U8390 ( .A1(n10007), .A2(n6776), .ZN(n6780) );
  NAND2_X1 U8391 ( .A1(n10026), .A2(n7186), .ZN(n6779) );
  INV_X1 U8392 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6777) );
  NOR2_X1 U8393 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6777), .ZN(n7488) );
  INV_X1 U8394 ( .A(n7488), .ZN(n6778) );
  NAND3_X1 U8395 ( .A1(n6780), .A2(n6779), .A3(n6778), .ZN(n6781) );
  AOI21_X1 U8396 ( .B1(n9930), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n6781), .ZN(
        n6782) );
  OAI21_X1 U8397 ( .B1(n6783), .B2(n10032), .A(n6782), .ZN(P1_U3251) );
  INV_X1 U8398 ( .A(n8055), .ZN(n8606) );
  OAI222_X1 U8399 ( .A1(n8110), .A2(n6785), .B1(n8606), .B2(n7777), .C1(n6784), 
        .C2(n8438), .ZN(P2_U3341) );
  OAI21_X1 U8400 ( .B1(n6786), .B2(n6787), .A(n6788), .ZN(n6793) );
  INV_X1 U8401 ( .A(n9139), .ZN(n9125) );
  NAND2_X1 U8402 ( .A1(n6991), .A2(n9766), .ZN(n10060) );
  OAI22_X1 U8403 ( .A1(n9125), .A2(n6966), .B1(n10060), .B2(n7125), .ZN(n6792)
         );
  INV_X1 U8404 ( .A(n4400), .ZN(n6948) );
  OAI22_X1 U8405 ( .A1(n6948), .A2(n9137), .B1(n6790), .B2(n6789), .ZN(n6791)
         );
  AOI211_X1 U8406 ( .C1(n6793), .C2(n9119), .A(n6792), .B(n6791), .ZN(n6794)
         );
  INV_X1 U8407 ( .A(n6794), .ZN(P1_U3235) );
  AOI211_X1 U8408 ( .C1(n6797), .C2(n6796), .A(n6795), .B(n10122), .ZN(n6806)
         );
  NAND2_X1 U8409 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7131) );
  INV_X1 U8410 ( .A(n7131), .ZN(n6798) );
  AOI21_X1 U8411 ( .B1(n10124), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6798), .ZN(
        n6803) );
  OAI211_X1 U8412 ( .C1(n6801), .C2(n6800), .A(n10119), .B(n6799), .ZN(n6802)
         );
  OAI211_X1 U8413 ( .C1(n10121), .C2(n6804), .A(n6803), .B(n6802), .ZN(n6805)
         );
  OR2_X1 U8414 ( .A1(n6806), .A2(n6805), .ZN(P2_U3249) );
  AOI211_X1 U8415 ( .C1(n6809), .C2(n6808), .A(n6807), .B(n10122), .ZN(n6818)
         );
  NAND2_X1 U8416 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(n7777), .ZN(n7308) );
  INV_X1 U8417 ( .A(n7308), .ZN(n6810) );
  AOI21_X1 U8418 ( .B1(n10124), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6810), .ZN(
        n6815) );
  OAI211_X1 U8419 ( .C1(n6813), .C2(n6812), .A(n10119), .B(n6811), .ZN(n6814)
         );
  OAI211_X1 U8420 ( .C1(n10121), .C2(n6816), .A(n6815), .B(n6814), .ZN(n6817)
         );
  OR2_X1 U8421 ( .A1(n6818), .A2(n6817), .ZN(P2_U3251) );
  AOI211_X1 U8422 ( .C1(n6821), .C2(n6820), .A(n6819), .B(n10122), .ZN(n6830)
         );
  NOR2_X1 U8423 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5155), .ZN(n6822) );
  AOI21_X1 U8424 ( .B1(n10124), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6822), .ZN(
        n6827) );
  OAI211_X1 U8425 ( .C1(n6825), .C2(n6824), .A(n10119), .B(n6823), .ZN(n6826)
         );
  OAI211_X1 U8426 ( .C1(n10121), .C2(n6828), .A(n6827), .B(n6826), .ZN(n6829)
         );
  OR2_X1 U8427 ( .A1(n6830), .A2(n6829), .ZN(P2_U3248) );
  AOI211_X1 U8428 ( .C1(n6833), .C2(n6832), .A(n6831), .B(n10122), .ZN(n6842)
         );
  INV_X1 U8429 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7167) );
  NOR2_X1 U8430 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7167), .ZN(n6834) );
  AOI21_X1 U8431 ( .B1(n10124), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6834), .ZN(
        n6839) );
  OAI211_X1 U8432 ( .C1(n6837), .C2(n6836), .A(n10119), .B(n6835), .ZN(n6838)
         );
  OAI211_X1 U8433 ( .C1(n10121), .C2(n6840), .A(n6839), .B(n6838), .ZN(n6841)
         );
  OR2_X1 U8434 ( .A1(n6842), .A2(n6841), .ZN(P2_U3250) );
  AOI211_X1 U8435 ( .C1(n6845), .C2(n6844), .A(n6843), .B(n10122), .ZN(n6854)
         );
  NOR2_X1 U8436 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7231), .ZN(n6846) );
  AOI21_X1 U8437 ( .B1(n10124), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6846), .ZN(
        n6851) );
  OAI211_X1 U8438 ( .C1(n6849), .C2(n6848), .A(n10119), .B(n6847), .ZN(n6850)
         );
  OAI211_X1 U8439 ( .C1(n10121), .C2(n6852), .A(n6851), .B(n6850), .ZN(n6853)
         );
  OR2_X1 U8440 ( .A1(n6854), .A2(n6853), .ZN(P2_U3252) );
  AOI211_X1 U8441 ( .C1(n6857), .C2(n6856), .A(n6855), .B(n10122), .ZN(n6865)
         );
  AND2_X1 U8442 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7246) );
  AOI21_X1 U8443 ( .B1(n10124), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7246), .ZN(
        n6862) );
  OAI211_X1 U8444 ( .C1(n6860), .C2(n6859), .A(n10119), .B(n6858), .ZN(n6861)
         );
  OAI211_X1 U8445 ( .C1(n10121), .C2(n6863), .A(n6862), .B(n6861), .ZN(n6864)
         );
  OR2_X1 U8446 ( .A1(n6865), .A2(n6864), .ZN(P2_U3253) );
  NOR2_X1 U8447 ( .A1(n6013), .A2(n6868), .ZN(n6869) );
  XNOR2_X1 U8448 ( .A(n6866), .B(n6869), .ZN(n6874) );
  AOI22_X1 U8449 ( .A1(n9128), .A2(n9461), .B1(n9144), .B2(n6959), .ZN(n6872)
         );
  INV_X1 U8450 ( .A(n7027), .ZN(n9459) );
  AOI21_X1 U8451 ( .B1(n9139), .B2(n9459), .A(n6870), .ZN(n6871) );
  OAI211_X1 U8452 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9142), .A(n6872), .B(
        n6871), .ZN(n6873) );
  AOI21_X1 U8453 ( .B1(n6874), .B2(n9119), .A(n6873), .ZN(n6875) );
  INV_X1 U8454 ( .A(n6875), .ZN(P1_U3216) );
  AOI21_X1 U8455 ( .B1(n9829), .B2(n6877), .A(n6876), .ZN(n6881) );
  AOI22_X1 U8456 ( .A1(n9476), .A2(n6879), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n6878), .ZN(n6880) );
  NOR2_X1 U8457 ( .A1(n6881), .A2(n6880), .ZN(n9478) );
  AOI21_X1 U8458 ( .B1(n6881), .B2(n6880), .A(n9478), .ZN(n6893) );
  NOR2_X1 U8459 ( .A1(n9476), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6882) );
  AOI21_X1 U8460 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9476), .A(n6882), .ZN(
        n6885) );
  OAI21_X1 U8461 ( .B1(n6885), .B2(n6884), .A(n9464), .ZN(n6891) );
  NOR2_X1 U8462 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6886), .ZN(n7714) );
  INV_X1 U8463 ( .A(n7714), .ZN(n6888) );
  NAND2_X1 U8464 ( .A1(n10026), .A2(n9476), .ZN(n6887) );
  OAI211_X1 U8465 ( .C1(n10035), .C2(n6889), .A(n6888), .B(n6887), .ZN(n6890)
         );
  AOI21_X1 U8466 ( .B1(n6891), .B2(n10007), .A(n6890), .ZN(n6892) );
  OAI21_X1 U8467 ( .B1(n6893), .B2(n10032), .A(n6892), .ZN(P1_U3252) );
  INV_X1 U8468 ( .A(n8006), .ZN(n6913) );
  AOI22_X1 U8469 ( .A1(n8059), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n9000), .ZN(n6894) );
  OAI21_X1 U8470 ( .B1(n6913), .B2(n9002), .A(n6894), .ZN(P2_U3340) );
  INV_X1 U8471 ( .A(n6895), .ZN(n6899) );
  NOR2_X1 U8472 ( .A1(n6897), .A2(n6896), .ZN(n6898) );
  NAND2_X1 U8473 ( .A1(n6899), .A2(n6898), .ZN(n6902) );
  NAND2_X1 U8474 ( .A1(n9439), .A2(n9190), .ZN(n6900) );
  OAI22_X1 U8475 ( .A1(n9610), .A2(n5959), .B1(n5958), .B2(n10042), .ZN(n6901)
         );
  INV_X1 U8476 ( .A(n6901), .ZN(n6906) );
  AND2_X1 U8477 ( .A1(n9884), .A2(n9881), .ZN(n9670) );
  INV_X1 U8478 ( .A(n10044), .ZN(n6903) );
  NAND2_X1 U8479 ( .A1(n9610), .A2(n6903), .ZN(n9660) );
  OAI21_X1 U8480 ( .B1(n9670), .B2(n9874), .A(n6904), .ZN(n6905) );
  OAI211_X1 U8481 ( .C1(n6907), .C2(n4399), .A(n6906), .B(n6905), .ZN(P1_U3291) );
  NAND2_X1 U8482 ( .A1(n6909), .A2(n6908), .ZN(n6910) );
  NAND2_X1 U8483 ( .A1(n6910), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6911) );
  XNOR2_X1 U8484 ( .A(n6911), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10027) );
  INV_X1 U8485 ( .A(n10027), .ZN(n9491) );
  INV_X1 U8486 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6912) );
  OAI222_X1 U8487 ( .A1(n9491), .A2(P1_U3084), .B1(n7925), .B2(n6913), .C1(
        n6912), .C2(n9791), .ZN(P1_U3335) );
  OAI21_X1 U8488 ( .B1(n6915), .B2(n4422), .A(n6914), .ZN(n6922) );
  INV_X1 U8489 ( .A(n7021), .ZN(n9458) );
  NOR2_X1 U8490 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6916), .ZN(n9914) );
  AOI21_X1 U8491 ( .B1(n9139), .B2(n9458), .A(n9914), .ZN(n6920) );
  NAND2_X1 U8492 ( .A1(n9144), .A2(n6976), .ZN(n6919) );
  OR2_X1 U8493 ( .A1(n9142), .A2(n6970), .ZN(n6918) );
  INV_X1 U8494 ( .A(n6966), .ZN(n9460) );
  NAND2_X1 U8495 ( .A1(n9128), .A2(n9460), .ZN(n6917) );
  NAND4_X1 U8496 ( .A1(n6920), .A2(n6919), .A3(n6918), .A4(n6917), .ZN(n6921)
         );
  AOI21_X1 U8497 ( .B1(n6922), .B2(n9119), .A(n6921), .ZN(n6923) );
  INV_X1 U8498 ( .A(n6923), .ZN(P1_U3228) );
  MUX2_X1 U8499 ( .A(n6924), .B(P2_REG1_REG_12__SCAN_IN), .S(n7102), .Z(n6930)
         );
  NAND2_X1 U8500 ( .A1(n8575), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6928) );
  MUX2_X1 U8501 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n6925), .S(n8575), .Z(n8577)
         );
  OAI21_X1 U8502 ( .B1(n10213), .B2(n6927), .A(n6926), .ZN(n8578) );
  NAND2_X1 U8503 ( .A1(n8577), .A2(n8578), .ZN(n8576) );
  NAND2_X1 U8504 ( .A1(n6928), .A2(n8576), .ZN(n6929) );
  NOR2_X1 U8505 ( .A1(n6929), .A2(n6930), .ZN(n7097) );
  AOI21_X1 U8506 ( .B1(n6930), .B2(n6929), .A(n7097), .ZN(n6933) );
  NAND2_X1 U8507 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7630) );
  INV_X1 U8508 ( .A(n7630), .ZN(n6931) );
  AOI21_X1 U8509 ( .B1(n10124), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n6931), .ZN(
        n6932) );
  OAI21_X1 U8510 ( .B1(n8611), .B2(n6933), .A(n6932), .ZN(n6941) );
  NOR2_X1 U8511 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(n8575), .ZN(n6936) );
  AOI21_X1 U8512 ( .B1(n8575), .B2(P2_REG2_REG_11__SCAN_IN), .A(n6936), .ZN(
        n8570) );
  NAND2_X1 U8513 ( .A1(n8571), .A2(n8570), .ZN(n8569) );
  OAI21_X1 U8514 ( .B1(n8575), .B2(P2_REG2_REG_11__SCAN_IN), .A(n8569), .ZN(
        n6939) );
  NAND2_X1 U8515 ( .A1(n7102), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6937) );
  OAI21_X1 U8516 ( .B1(n7102), .B2(P2_REG2_REG_12__SCAN_IN), .A(n6937), .ZN(
        n6938) );
  NOR2_X1 U8517 ( .A1(n6938), .A2(n6939), .ZN(n7101) );
  AOI211_X1 U8518 ( .C1(n6939), .C2(n6938), .A(n7101), .B(n10122), .ZN(n6940)
         );
  AOI211_X1 U8519 ( .C1(n9815), .C2(n7102), .A(n6941), .B(n6940), .ZN(n6942)
         );
  INV_X1 U8520 ( .A(n6942), .ZN(P2_U3257) );
  NAND2_X1 U8521 ( .A1(n4400), .A2(n4728), .ZN(n6943) );
  NAND2_X1 U8522 ( .A1(n9461), .A2(n6990), .ZN(n9403) );
  NAND2_X1 U8523 ( .A1(n6952), .A2(n6991), .ZN(n9402) );
  NAND2_X1 U8524 ( .A1(n4425), .A2(n6945), .ZN(n6987) );
  NAND2_X1 U8525 ( .A1(n6952), .A2(n6990), .ZN(n6946) );
  NAND2_X1 U8526 ( .A1(n6987), .A2(n6946), .ZN(n6947) );
  NAND2_X1 U8527 ( .A1(n6966), .A2(n6959), .ZN(n9406) );
  NAND2_X1 U8528 ( .A1(n9460), .A2(n10066), .ZN(n9234) );
  NAND2_X1 U8529 ( .A1(n9406), .A2(n9234), .ZN(n6965) );
  NAND2_X1 U8530 ( .A1(n6947), .A2(n6965), .ZN(n6964) );
  OAI21_X1 U8531 ( .B1(n6947), .B2(n6965), .A(n6964), .ZN(n10070) );
  INV_X1 U8532 ( .A(n10070), .ZN(n6962) );
  NOR3_X1 U8533 ( .A1(n4399), .A2(n9499), .A3(n6100), .ZN(n7770) );
  INV_X1 U8534 ( .A(n7770), .ZN(n7259) );
  INV_X1 U8535 ( .A(n9870), .ZN(n9596) );
  NAND2_X1 U8536 ( .A1(n6948), .A2(n4728), .ZN(n6949) );
  NAND2_X1 U8537 ( .A1(n9405), .A2(n9163), .ZN(n6951) );
  XNOR2_X1 U8538 ( .A(n9236), .B(n6965), .ZN(n6955) );
  INV_X1 U8539 ( .A(n9680), .ZN(n7765) );
  INV_X1 U8540 ( .A(n9865), .ZN(n9601) );
  OAI22_X1 U8541 ( .A1(n6952), .A2(n9601), .B1(n7027), .B2(n9599), .ZN(n6953)
         );
  AOI21_X1 U8542 ( .B1(n10070), .B2(n7765), .A(n6953), .ZN(n6954) );
  OAI21_X1 U8543 ( .B1(n9596), .B2(n6955), .A(n6954), .ZN(n10068) );
  NAND2_X1 U8544 ( .A1(n10068), .A2(n9610), .ZN(n6961) );
  OAI22_X1 U8545 ( .A1(n9610), .A2(n6280), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10042), .ZN(n6958) );
  INV_X1 U8546 ( .A(n9670), .ZN(n9510) );
  AND2_X1 U8547 ( .A1(n6989), .A2(n6959), .ZN(n6956) );
  OR2_X1 U8548 ( .A1(n6956), .A2(n6972), .ZN(n10067) );
  NOR2_X1 U8549 ( .A1(n9510), .A2(n10067), .ZN(n6957) );
  AOI211_X1 U8550 ( .C1(n9874), .C2(n6959), .A(n6958), .B(n6957), .ZN(n6960)
         );
  OAI211_X1 U8551 ( .C1(n6962), .C2(n7259), .A(n6961), .B(n6960), .ZN(P1_U3288) );
  NAND2_X1 U8552 ( .A1(n6966), .A2(n10066), .ZN(n6963) );
  NAND2_X1 U8553 ( .A1(n6964), .A2(n6963), .ZN(n7026) );
  NAND2_X1 U8554 ( .A1(n7027), .A2(n6976), .ZN(n7036) );
  NAND2_X1 U8555 ( .A1(n9459), .A2(n10072), .ZN(n7055) );
  NAND2_X1 U8556 ( .A1(n7036), .A2(n7055), .ZN(n9167) );
  XOR2_X1 U8557 ( .A(n7026), .B(n9167), .Z(n10071) );
  INV_X1 U8558 ( .A(n6965), .ZN(n9164) );
  NAND2_X1 U8559 ( .A1(n9236), .A2(n9164), .ZN(n9274) );
  XOR2_X1 U8560 ( .A(n7056), .B(n9167), .Z(n6968) );
  OAI22_X1 U8561 ( .A1(n6966), .A2(n9601), .B1(n7021), .B2(n9599), .ZN(n6967)
         );
  AOI21_X1 U8562 ( .B1(n6968), .B2(n9870), .A(n6967), .ZN(n6969) );
  OAI21_X1 U8563 ( .B1(n10071), .B2(n9680), .A(n6969), .ZN(n10074) );
  NAND2_X1 U8564 ( .A1(n10074), .A2(n9610), .ZN(n6978) );
  INV_X1 U8565 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6971) );
  OAI22_X1 U8566 ( .A1(n9610), .A2(n6971), .B1(n6970), .B2(n10042), .ZN(n6975)
         );
  OR2_X1 U8567 ( .A1(n6972), .A2(n10072), .ZN(n6973) );
  NAND2_X1 U8568 ( .A1(n7030), .A2(n6973), .ZN(n10073) );
  NOR2_X1 U8569 ( .A1(n9510), .A2(n10073), .ZN(n6974) );
  AOI211_X1 U8570 ( .C1(n9874), .C2(n6976), .A(n6975), .B(n6974), .ZN(n6977)
         );
  OAI211_X1 U8571 ( .C1(n10071), .C2(n7259), .A(n6978), .B(n6977), .ZN(
        P1_U3287) );
  INV_X1 U8572 ( .A(n8148), .ZN(n6981) );
  OAI222_X1 U8573 ( .A1(P1_U3084), .A2(n9499), .B1(n7925), .B2(n6981), .C1(
        n6979), .C2(n9791), .ZN(P1_U3334) );
  OAI222_X1 U8574 ( .A1(n8438), .A2(n6982), .B1(n9002), .B2(n6981), .C1(
        P2_U3152), .C2(n6980), .ZN(P2_U3339) );
  XNOR2_X1 U8575 ( .A(n9405), .B(n9163), .ZN(n6983) );
  NAND2_X1 U8576 ( .A1(n6983), .A2(n9870), .ZN(n6985) );
  AOI22_X1 U8577 ( .A1(n9460), .A2(n9867), .B1(n9865), .B2(n4400), .ZN(n6984)
         );
  NAND2_X1 U8578 ( .A1(n6985), .A2(n6984), .ZN(n10062) );
  INV_X1 U8579 ( .A(n10062), .ZN(n6996) );
  AND2_X1 U8580 ( .A1(n9441), .A2(n8322), .ZN(n6986) );
  NAND2_X1 U8581 ( .A1(n9610), .A2(n6986), .ZN(n9672) );
  INV_X1 U8582 ( .A(n9672), .ZN(n9885) );
  OAI21_X1 U8583 ( .B1(n4425), .B2(n6945), .A(n6987), .ZN(n10064) );
  OAI21_X1 U8584 ( .B1(n4761), .B2(n6990), .A(n6989), .ZN(n10061) );
  INV_X1 U8585 ( .A(n10042), .ZN(n9872) );
  AOI22_X1 U8586 ( .A1(n4399), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9872), .ZN(n6993) );
  NAND2_X1 U8587 ( .A1(n9874), .A2(n6991), .ZN(n6992) );
  OAI211_X1 U8588 ( .C1(n9510), .C2(n10061), .A(n6993), .B(n6992), .ZN(n6994)
         );
  AOI21_X1 U8589 ( .B1(n9885), .B2(n10064), .A(n6994), .ZN(n6995) );
  OAI21_X1 U8590 ( .B1(n6996), .B2(n4399), .A(n6995), .ZN(P1_U3289) );
  NAND2_X1 U8591 ( .A1(n5741), .A2(n5458), .ZN(n6997) );
  OR2_X1 U8592 ( .A1(n6998), .A2(n6997), .ZN(n8977) );
  INV_X1 U8593 ( .A(n8977), .ZN(n10192) );
  OR2_X1 U8594 ( .A1(n7000), .A2(n6999), .ZN(n7001) );
  AND2_X1 U8595 ( .A1(n7002), .A2(n7001), .ZN(n7521) );
  INV_X1 U8596 ( .A(n7521), .ZN(n7013) );
  NAND2_X1 U8597 ( .A1(n7428), .A2(n7518), .ZN(n7003) );
  NAND2_X1 U8598 ( .A1(n7505), .A2(n7003), .ZN(n7515) );
  INV_X1 U8599 ( .A(n10195), .ZN(n10187) );
  OAI22_X1 U8600 ( .A1(n7515), .A2(n10187), .B1(n7004), .B2(n10186), .ZN(n7012) );
  OAI21_X1 U8601 ( .B1(n7006), .B2(n7005), .A(n7500), .ZN(n7010) );
  OAI22_X1 U8602 ( .A1(n7008), .A2(n8853), .B1(n7007), .B2(n8851), .ZN(n7009)
         );
  AOI21_X1 U8603 ( .B1(n7010), .B2(n8863), .A(n7009), .ZN(n7011) );
  OAI21_X1 U8604 ( .B1(n7521), .B2(n8859), .A(n7011), .ZN(n7523) );
  AOI211_X1 U8605 ( .C1(n10192), .C2(n7013), .A(n7012), .B(n7523), .ZN(n7157)
         );
  NAND2_X1 U8606 ( .A1(n7015), .A2(n7014), .ZN(n7016) );
  OR2_X1 U8607 ( .A1(n10130), .A2(n7016), .ZN(n7151) );
  NOR2_X1 U8608 ( .A1(n7151), .A2(n7150), .ZN(n7017) );
  AND2_X1 U8609 ( .A1(n7154), .A2(n7017), .ZN(n7019) );
  INV_X1 U8610 ( .A(n7018), .ZN(n7155) );
  NAND2_X1 U8611 ( .A1(n10215), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7020) );
  OAI21_X1 U8612 ( .B1(n7157), .B2(n10215), .A(n7020), .ZN(P2_U3523) );
  NAND2_X1 U8613 ( .A1(n7038), .A2(n7036), .ZN(n7023) );
  NAND2_X1 U8614 ( .A1(n7021), .A2(n7112), .ZN(n9230) );
  NAND2_X1 U8615 ( .A1(n9458), .A2(n7022), .ZN(n7057) );
  XNOR2_X1 U8616 ( .A(n7023), .B(n9166), .ZN(n7025) );
  OAI22_X1 U8617 ( .A1(n7027), .A2(n9601), .B1(n7064), .B2(n9599), .ZN(n7024)
         );
  AOI21_X1 U8618 ( .B1(n7025), .B2(n9870), .A(n7024), .ZN(n10082) );
  NAND2_X1 U8619 ( .A1(n7027), .A2(n10072), .ZN(n7028) );
  OR2_X1 U8620 ( .A1(n7062), .A2(n9166), .ZN(n7041) );
  NAND2_X1 U8621 ( .A1(n7062), .A2(n9166), .ZN(n7029) );
  AND2_X1 U8622 ( .A1(n7041), .A2(n7029), .ZN(n10081) );
  AOI21_X1 U8623 ( .B1(n7030), .B2(n7112), .A(n10101), .ZN(n7031) );
  NAND2_X1 U8624 ( .A1(n7031), .A2(n7045), .ZN(n10079) );
  INV_X1 U8625 ( .A(n9884), .ZN(n8038) );
  OAI22_X1 U8626 ( .A1(n9610), .A2(n6275), .B1(n7121), .B2(n10042), .ZN(n7032)
         );
  AOI21_X1 U8627 ( .B1(n9874), .B2(n7112), .A(n7032), .ZN(n7033) );
  OAI21_X1 U8628 ( .B1(n10079), .B2(n8038), .A(n7033), .ZN(n7034) );
  AOI21_X1 U8629 ( .B1(n10081), .B2(n9885), .A(n7034), .ZN(n7035) );
  OAI21_X1 U8630 ( .B1(n10082), .B2(n4399), .A(n7035), .ZN(P1_U3286) );
  NAND2_X1 U8631 ( .A1(n9230), .A2(n7036), .ZN(n9232) );
  INV_X1 U8632 ( .A(n9232), .ZN(n7037) );
  NAND2_X1 U8633 ( .A1(n7064), .A2(n7051), .ZN(n9279) );
  INV_X1 U8634 ( .A(n7051), .ZN(n7063) );
  INV_X1 U8635 ( .A(n7064), .ZN(n9457) );
  NAND2_X1 U8636 ( .A1(n7063), .A2(n9457), .ZN(n9275) );
  NAND2_X1 U8637 ( .A1(n9279), .A2(n9275), .ZN(n7043) );
  OAI21_X1 U8638 ( .B1(n4483), .B2(n4580), .A(n9284), .ZN(n7039) );
  AOI222_X1 U8639 ( .A1(n9870), .A2(n7039), .B1(n9458), .B2(n9865), .C1(n9456), 
        .C2(n9867), .ZN(n10086) );
  NAND2_X1 U8640 ( .A1(n9458), .A2(n7112), .ZN(n7040) );
  AND2_X1 U8641 ( .A1(n7041), .A2(n7040), .ZN(n7044) );
  AND2_X1 U8642 ( .A1(n7043), .A2(n7040), .ZN(n7065) );
  NAND2_X1 U8643 ( .A1(n7041), .A2(n7065), .ZN(n7042) );
  OAI21_X1 U8644 ( .B1(n7044), .B2(n7043), .A(n7042), .ZN(n10089) );
  INV_X1 U8645 ( .A(n7045), .ZN(n7047) );
  INV_X1 U8646 ( .A(n7074), .ZN(n7046) );
  OAI21_X1 U8647 ( .B1(n7063), .B2(n7047), .A(n7046), .ZN(n10087) );
  OAI22_X1 U8648 ( .A1(n9610), .A2(n7049), .B1(n7048), .B2(n10042), .ZN(n7050)
         );
  AOI21_X1 U8649 ( .B1(n9874), .B2(n7051), .A(n7050), .ZN(n7052) );
  OAI21_X1 U8650 ( .B1(n10087), .B2(n9510), .A(n7052), .ZN(n7053) );
  AOI21_X1 U8651 ( .B1(n10089), .B2(n9885), .A(n7053), .ZN(n7054) );
  OAI21_X1 U8652 ( .B1(n10086), .B2(n4399), .A(n7054), .ZN(P1_U3285) );
  AND2_X1 U8653 ( .A1(n7057), .A2(n7055), .ZN(n9229) );
  NAND2_X1 U8654 ( .A1(n9232), .A2(n7057), .ZN(n7058) );
  NAND2_X1 U8655 ( .A1(n7058), .A2(n9279), .ZN(n7059) );
  NAND2_X1 U8656 ( .A1(n7059), .A2(n9275), .ZN(n9408) );
  OR2_X1 U8657 ( .A1(n7352), .A2(n7082), .ZN(n9281) );
  NAND2_X1 U8658 ( .A1(n7352), .A2(n7082), .ZN(n9280) );
  NAND2_X1 U8659 ( .A1(n9281), .A2(n9280), .ZN(n7070) );
  INV_X1 U8660 ( .A(n7070), .ZN(n9170) );
  XNOR2_X1 U8661 ( .A(n7079), .B(n9170), .ZN(n7061) );
  OAI22_X1 U8662 ( .A1(n7251), .A2(n9599), .B1(n7064), .B2(n9601), .ZN(n7060)
         );
  AOI21_X1 U8663 ( .B1(n7061), .B2(n9870), .A(n7060), .ZN(n10092) );
  AND2_X1 U8664 ( .A1(n7064), .A2(n7063), .ZN(n7066) );
  OR2_X1 U8665 ( .A1(n7066), .A2(n7065), .ZN(n7067) );
  AND2_X1 U8666 ( .A1(n7069), .A2(n7067), .ZN(n7071) );
  AND2_X1 U8667 ( .A1(n7067), .A2(n7070), .ZN(n7068) );
  NAND2_X1 U8668 ( .A1(n7069), .A2(n7068), .ZN(n7086) );
  OAI21_X1 U8669 ( .B1(n7071), .B2(n7070), .A(n7086), .ZN(n10096) );
  NAND2_X1 U8670 ( .A1(n10096), .A2(n9885), .ZN(n7078) );
  OAI22_X1 U8671 ( .A1(n9610), .A2(n7072), .B1(n7343), .B2(n10042), .ZN(n7076)
         );
  INV_X1 U8672 ( .A(n7352), .ZN(n10094) );
  INV_X1 U8673 ( .A(n7092), .ZN(n7073) );
  OAI211_X1 U8674 ( .C1(n10094), .C2(n7074), .A(n7073), .B(n9881), .ZN(n10091)
         );
  NOR2_X1 U8675 ( .A1(n10091), .A2(n8038), .ZN(n7075) );
  AOI211_X1 U8676 ( .C1(n9874), .C2(n7352), .A(n7076), .B(n7075), .ZN(n7077)
         );
  OAI211_X1 U8677 ( .C1(n4399), .C2(n10092), .A(n7078), .B(n7077), .ZN(
        P1_U3284) );
  NAND2_X1 U8678 ( .A1(n7080), .A2(n9280), .ZN(n7196) );
  OR2_X1 U8679 ( .A1(n7177), .A2(n7251), .ZN(n9218) );
  NAND2_X1 U8680 ( .A1(n7177), .A2(n7251), .ZN(n9291) );
  XNOR2_X1 U8681 ( .A(n7196), .B(n9171), .ZN(n7084) );
  NAND2_X1 U8682 ( .A1(n9454), .A2(n9867), .ZN(n7081) );
  OAI21_X1 U8683 ( .B1(n7082), .B2(n9601), .A(n7081), .ZN(n7083) );
  AOI21_X1 U8684 ( .B1(n7084), .B2(n9870), .A(n7083), .ZN(n10099) );
  OR2_X1 U8685 ( .A1(n7352), .A2(n9456), .ZN(n7085) );
  INV_X1 U8686 ( .A(n7179), .ZN(n7087) );
  AOI21_X1 U8687 ( .B1(n9171), .B2(n7088), .A(n7087), .ZN(n10104) );
  NAND2_X1 U8688 ( .A1(n10104), .A2(n9885), .ZN(n7096) );
  OAI22_X1 U8689 ( .A1(n9610), .A2(n7090), .B1(n7089), .B2(n10042), .ZN(n7094)
         );
  INV_X1 U8690 ( .A(n7177), .ZN(n7091) );
  NAND2_X1 U8691 ( .A1(n7092), .A2(n7091), .ZN(n7256) );
  OAI21_X1 U8692 ( .B1(n7092), .B2(n7091), .A(n7256), .ZN(n10100) );
  NOR2_X1 U8693 ( .A1(n10100), .A2(n9510), .ZN(n7093) );
  AOI211_X1 U8694 ( .C1(n9874), .C2(n7177), .A(n7094), .B(n7093), .ZN(n7095)
         );
  OAI211_X1 U8695 ( .C1(n4399), .C2(n10099), .A(n7096), .B(n7095), .ZN(
        P1_U3283) );
  AOI21_X1 U8696 ( .B1(n7098), .B2(n6924), .A(n7097), .ZN(n7100) );
  AOI22_X1 U8697 ( .A1(n7220), .A2(n5366), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7215), .ZN(n7099) );
  NOR2_X1 U8698 ( .A1(n7100), .A2(n7099), .ZN(n7214) );
  AOI21_X1 U8699 ( .B1(n7100), .B2(n7099), .A(n7214), .ZN(n7111) );
  NOR2_X1 U8700 ( .A1(n7220), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7103) );
  AOI21_X1 U8701 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n7220), .A(n7103), .ZN(
        n7104) );
  NAND2_X1 U8702 ( .A1(n7105), .A2(n7104), .ZN(n7219) );
  OAI21_X1 U8703 ( .B1(n7105), .B2(n7104), .A(n7219), .ZN(n7106) );
  NAND2_X1 U8704 ( .A1(n7106), .A2(n10118), .ZN(n7110) );
  NOR2_X1 U8705 ( .A1(n7107), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7677) );
  NOR2_X1 U8706 ( .A1(n10121), .A2(n7215), .ZN(n7108) );
  AOI211_X1 U8707 ( .C1(P2_ADDR_REG_13__SCAN_IN), .C2(n10124), .A(n7677), .B(
        n7108), .ZN(n7109) );
  OAI211_X1 U8708 ( .C1(n7111), .C2(n8611), .A(n7110), .B(n7109), .ZN(P2_U3258) );
  NAND2_X1 U8709 ( .A1(n7112), .A2(n9766), .ZN(n10078) );
  XNOR2_X1 U8710 ( .A(n7115), .B(n7114), .ZN(n7116) );
  XNOR2_X1 U8711 ( .A(n7113), .B(n7116), .ZN(n7117) );
  NAND2_X1 U8712 ( .A1(n7117), .A2(n9119), .ZN(n7124) );
  NAND2_X1 U8713 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9927) );
  INV_X1 U8714 ( .A(n9927), .ZN(n7118) );
  AOI21_X1 U8715 ( .B1(n9139), .B2(n9457), .A(n7118), .ZN(n7120) );
  NAND2_X1 U8716 ( .A1(n9128), .A2(n9459), .ZN(n7119) );
  OAI211_X1 U8717 ( .C1(n9142), .C2(n7121), .A(n7120), .B(n7119), .ZN(n7122)
         );
  INV_X1 U8718 ( .A(n7122), .ZN(n7123) );
  OAI211_X1 U8719 ( .C1(n7125), .C2(n10078), .A(n7124), .B(n7123), .ZN(
        P1_U3225) );
  INV_X1 U8720 ( .A(n7126), .ZN(n7128) );
  NOR2_X1 U8721 ( .A1(n7128), .A2(n7127), .ZN(n7129) );
  XNOR2_X1 U8722 ( .A(n7130), .B(n7129), .ZN(n7135) );
  INV_X1 U8723 ( .A(n8548), .ZN(n8522) );
  OAI21_X1 U8724 ( .B1(n8546), .B2(n7507), .A(n7131), .ZN(n7133) );
  OAI22_X1 U8725 ( .A1(n8541), .A2(n10162), .B1(n8547), .B2(n4593), .ZN(n7132)
         );
  AOI211_X1 U8726 ( .C1(n8522), .C2(n8566), .A(n7133), .B(n7132), .ZN(n7134)
         );
  OAI21_X1 U8727 ( .B1(n7135), .B2(n8553), .A(n7134), .ZN(P2_U3232) );
  XNOR2_X1 U8728 ( .A(n7136), .B(n7137), .ZN(n7141) );
  AOI22_X1 U8729 ( .A1(n8523), .A2(n8565), .B1(n7518), .B2(n8551), .ZN(n7140)
         );
  OAI22_X1 U8730 ( .A1(n8546), .A2(P2_REG3_REG_3__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n5155), .ZN(n7138) );
  AOI21_X1 U8731 ( .B1(n8522), .B2(n8568), .A(n7138), .ZN(n7139) );
  OAI211_X1 U8732 ( .C1(n7141), .C2(n8553), .A(n7140), .B(n7139), .ZN(P2_U3220) );
  INV_X1 U8733 ( .A(n8168), .ZN(n7961) );
  OAI222_X1 U8734 ( .A1(n7142), .A2(P1_U3084), .B1(n7925), .B2(n7961), .C1(
        n8169), .C2(n9791), .ZN(P1_U3333) );
  XNOR2_X1 U8735 ( .A(n7144), .B(n7143), .ZN(n7149) );
  AOI22_X1 U8736 ( .A1(n8522), .A2(n7441), .B1(n8523), .B2(n8566), .ZN(n7148)
         );
  INV_X1 U8737 ( .A(n7145), .ZN(n7146) );
  NAND2_X1 U8738 ( .A1(n7146), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8471) );
  AOI22_X1 U8739 ( .A1(n4639), .A2(n8551), .B1(n8471), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n7147) );
  OAI211_X1 U8740 ( .C1(n8553), .C2(n7149), .A(n7148), .B(n7147), .ZN(P2_U3239) );
  INV_X1 U8741 ( .A(n7150), .ZN(n7152) );
  NOR2_X1 U8742 ( .A1(n7152), .A2(n7151), .ZN(n7153) );
  AND2_X1 U8743 ( .A1(n7154), .A2(n7153), .ZN(n7156) );
  OR2_X1 U8744 ( .A1(n7157), .A2(n10202), .ZN(n7158) );
  OAI21_X1 U8745 ( .B1(n10204), .B2(n5171), .A(n7158), .ZN(P2_U3460) );
  INV_X1 U8746 ( .A(n8189), .ZN(n7172) );
  OAI222_X1 U8747 ( .A1(n8110), .A2(n7172), .B1(n7160), .B2(P2_U3152), .C1(
        n7159), .C2(n8438), .ZN(P2_U3337) );
  INV_X1 U8748 ( .A(n7161), .ZN(n7162) );
  AOI211_X1 U8749 ( .C1(n7164), .C2(n7163), .A(n8553), .B(n7162), .ZN(n7171)
         );
  NAND2_X1 U8750 ( .A1(n8563), .A2(n8821), .ZN(n7166) );
  NAND2_X1 U8751 ( .A1(n8565), .A2(n8819), .ZN(n7165) );
  NAND2_X1 U8752 ( .A1(n7166), .A2(n7165), .ZN(n7653) );
  INV_X1 U8753 ( .A(n7653), .ZN(n7168) );
  OAI22_X1 U8754 ( .A1(n8502), .A2(n7168), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7167), .ZN(n7170) );
  OAI22_X1 U8755 ( .A1(n8541), .A2(n10169), .B1(n8546), .B2(n7657), .ZN(n7169)
         );
  OR3_X1 U8756 ( .A1(n7171), .A2(n7170), .A3(n7169), .ZN(P2_U3229) );
  OAI222_X1 U8757 ( .A1(n9190), .A2(P1_U3084), .B1(n7925), .B2(n7172), .C1(
        n8190), .C2(n9791), .ZN(P1_U3332) );
  AOI22_X1 U8758 ( .A1(n8523), .A2(n7441), .B1(n10146), .B2(n8551), .ZN(n7175)
         );
  OAI21_X1 U8759 ( .B1(n7314), .B2(n8367), .A(n7320), .ZN(n7173) );
  AOI22_X1 U8760 ( .A1(n8476), .A2(n7173), .B1(n8471), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n7174) );
  OAI211_X1 U8761 ( .C1(n7176), .C2(n8531), .A(n7175), .B(n7174), .ZN(P2_U3234) );
  NAND2_X1 U8762 ( .A1(n7177), .A2(n9455), .ZN(n7178) );
  NAND2_X1 U8763 ( .A1(n7180), .A2(n9151), .ZN(n7183) );
  AOI22_X1 U8764 ( .A1(n8150), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8149), .B2(
        n7181), .ZN(n7182) );
  OR2_X1 U8765 ( .A1(n7451), .A2(n9454), .ZN(n7184) );
  NAND2_X1 U8766 ( .A1(n7185), .A2(n9151), .ZN(n7188) );
  AOI22_X1 U8767 ( .A1(n8150), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8149), .B2(
        n7186), .ZN(n7187) );
  NAND2_X1 U8768 ( .A1(n8421), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7194) );
  AND2_X2 U8769 ( .A1(n7189), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7200) );
  NOR2_X1 U8770 ( .A1(n7189), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7190) );
  OR2_X1 U8771 ( .A1(n7200), .A2(n7190), .ZN(n7490) );
  OR2_X1 U8772 ( .A1(n8332), .A2(n7490), .ZN(n7193) );
  OR2_X1 U8773 ( .A1(n8333), .A2(n6470), .ZN(n7192) );
  OR2_X1 U8774 ( .A1(n8425), .A2(n9829), .ZN(n7191) );
  NAND2_X1 U8775 ( .A1(n7492), .A2(n7712), .ZN(n9297) );
  NAND2_X1 U8776 ( .A1(n9288), .A2(n9297), .ZN(n7198) );
  NAND2_X1 U8777 ( .A1(n7195), .A2(n7198), .ZN(n7276) );
  OAI21_X1 U8778 ( .B1(n7195), .B2(n7198), .A(n7276), .ZN(n9827) );
  INV_X1 U8779 ( .A(n9827), .ZN(n7213) );
  NAND2_X1 U8780 ( .A1(n7196), .A2(n9171), .ZN(n7197) );
  INV_X1 U8781 ( .A(n9454), .ZN(n7486) );
  OR2_X1 U8782 ( .A1(n7451), .A2(n7486), .ZN(n9294) );
  NAND2_X1 U8783 ( .A1(n7451), .A2(n7486), .ZN(n9292) );
  INV_X1 U8784 ( .A(n7198), .ZN(n9176) );
  XNOR2_X1 U8785 ( .A(n7281), .B(n9176), .ZN(n7199) );
  NAND2_X1 U8786 ( .A1(n7199), .A2(n9870), .ZN(n7208) );
  NAND2_X1 U8787 ( .A1(n6030), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7206) );
  OR2_X1 U8788 ( .A1(n7200), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7201) );
  NAND2_X1 U8789 ( .A1(n7282), .A2(n7201), .ZN(n7716) );
  OR2_X1 U8790 ( .A1(n8332), .A2(n7716), .ZN(n7205) );
  INV_X1 U8791 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7202) );
  OR2_X1 U8792 ( .A1(n5996), .A2(n7202), .ZN(n7204) );
  INV_X1 U8793 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7292) );
  OR2_X1 U8794 ( .A1(n8333), .A2(n7292), .ZN(n7203) );
  NAND4_X1 U8795 ( .A1(n7206), .A2(n7205), .A3(n7204), .A4(n7203), .ZN(n9866)
         );
  AOI22_X1 U8796 ( .A1(n9867), .A2(n9866), .B1(n9454), .B2(n9865), .ZN(n7207)
         );
  NAND2_X1 U8797 ( .A1(n7208), .A2(n7207), .ZN(n9826) );
  INV_X1 U8798 ( .A(n7492), .ZN(n9824) );
  OAI211_X1 U8799 ( .C1(n9824), .C2(n4485), .A(n4421), .B(n9881), .ZN(n9823)
         );
  OAI22_X1 U8800 ( .A1(n9610), .A2(n6470), .B1(n7490), .B2(n10042), .ZN(n7209)
         );
  AOI21_X1 U8801 ( .B1(n7492), .B2(n9874), .A(n7209), .ZN(n7210) );
  OAI21_X1 U8802 ( .B1(n9823), .B2(n8038), .A(n7210), .ZN(n7211) );
  AOI21_X1 U8803 ( .B1(n9826), .B2(n9610), .A(n7211), .ZN(n7212) );
  OAI21_X1 U8804 ( .B1(n7213), .B2(n9672), .A(n7212), .ZN(P1_U3281) );
  AOI21_X1 U8805 ( .B1(n7215), .B2(n5366), .A(n7214), .ZN(n7218) );
  AOI22_X1 U8806 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n7327), .B1(n7330), .B2(
        n7216), .ZN(n7217) );
  NOR2_X1 U8807 ( .A1(n7218), .A2(n7217), .ZN(n7332) );
  AOI21_X1 U8808 ( .B1(n7218), .B2(n7217), .A(n7332), .ZN(n7228) );
  AOI22_X1 U8809 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7330), .B1(n7327), .B2(
        n7328), .ZN(n7222) );
  OAI21_X1 U8810 ( .B1(n7220), .B2(P2_REG2_REG_13__SCAN_IN), .A(n7219), .ZN(
        n7221) );
  OAI21_X1 U8811 ( .B1(n7222), .B2(n7221), .A(n7326), .ZN(n7223) );
  NAND2_X1 U8812 ( .A1(n7223), .A2(n10118), .ZN(n7227) );
  NAND2_X1 U8813 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(n7777), .ZN(n7853) );
  OAI21_X1 U8814 ( .B1(n8588), .B2(n7224), .A(n7853), .ZN(n7225) );
  AOI21_X1 U8815 ( .B1(n9815), .B2(n7330), .A(n7225), .ZN(n7226) );
  OAI211_X1 U8816 ( .C1(n7228), .C2(n8611), .A(n7227), .B(n7226), .ZN(P2_U3259) );
  NAND2_X1 U8817 ( .A1(n7230), .A2(n7229), .ZN(n7238) );
  OAI211_X1 U8818 ( .C1(n7230), .C2(n7229), .A(n7238), .B(n8476), .ZN(n7236)
         );
  OAI22_X1 U8819 ( .A1(n8546), .A2(n7467), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7231), .ZN(n7234) );
  OAI22_X1 U8820 ( .A1(n7232), .A2(n8547), .B1(n8548), .B2(n4487), .ZN(n7233)
         );
  AOI211_X1 U8821 ( .C1(n7412), .C2(n8551), .A(n7234), .B(n7233), .ZN(n7235)
         );
  NAND2_X1 U8822 ( .A1(n7236), .A2(n7235), .ZN(P2_U3215) );
  AOI21_X1 U8823 ( .B1(n7238), .B2(n7237), .A(n8553), .ZN(n7243) );
  NOR3_X1 U8824 ( .A1(n8531), .A2(n7534), .A3(n7239), .ZN(n7242) );
  AND2_X1 U8825 ( .A1(n7267), .A2(n7240), .ZN(n7241) );
  OAI21_X1 U8826 ( .B1(n7243), .B2(n7242), .A(n7241), .ZN(n7249) );
  INV_X1 U8827 ( .A(n7244), .ZN(n7247) );
  INV_X1 U8828 ( .A(n8546), .ZN(n8538) );
  OAI22_X1 U8829 ( .A1(n7534), .A2(n8548), .B1(n8547), .B2(n7993), .ZN(n7245)
         );
  AOI211_X1 U8830 ( .C1(n7247), .C2(n8538), .A(n7246), .B(n7245), .ZN(n7248)
         );
  OAI211_X1 U8831 ( .C1(n10179), .C2(n8541), .A(n7249), .B(n7248), .ZN(
        P2_U3223) );
  NAND2_X1 U8832 ( .A1(n9294), .A2(n9292), .ZN(n9173) );
  XOR2_X1 U8833 ( .A(n7250), .B(n9173), .Z(n7255) );
  OAI22_X1 U8834 ( .A1(n7251), .A2(n9601), .B1(n7712), .B2(n9599), .ZN(n7254)
         );
  XNOR2_X1 U8835 ( .A(n7252), .B(n9173), .ZN(n7420) );
  NOR2_X1 U8836 ( .A1(n7420), .A2(n9680), .ZN(n7253) );
  AOI211_X1 U8837 ( .C1(n7255), .C2(n9870), .A(n7254), .B(n7253), .ZN(n7419)
         );
  AOI21_X1 U8838 ( .B1(n7451), .B2(n7256), .A(n4485), .ZN(n7417) );
  INV_X1 U8839 ( .A(n7451), .ZN(n7465) );
  INV_X1 U8840 ( .A(n7459), .ZN(n7257) );
  AOI22_X1 U8841 ( .A1(n4399), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7257), .B2(
        n9872), .ZN(n7258) );
  OAI21_X1 U8842 ( .B1(n7465), .B2(n9660), .A(n7258), .ZN(n7261) );
  NOR2_X1 U8843 ( .A1(n7420), .A2(n7259), .ZN(n7260) );
  AOI211_X1 U8844 ( .C1(n7417), .C2(n9670), .A(n7261), .B(n7260), .ZN(n7262)
         );
  OAI21_X1 U8845 ( .B1(n7419), .B2(n4399), .A(n7262), .ZN(P1_U3282) );
  INV_X1 U8846 ( .A(n7263), .ZN(n7265) );
  AND2_X1 U8847 ( .A1(n7265), .A2(n7264), .ZN(n7266) );
  XNOR2_X1 U8848 ( .A(n10185), .B(n8365), .ZN(n7391) );
  NOR2_X1 U8849 ( .A1(n7397), .A2(n5743), .ZN(n7392) );
  XNOR2_X1 U8850 ( .A(n7391), .B(n7392), .ZN(n7395) );
  XNOR2_X1 U8851 ( .A(n7396), .B(n7395), .ZN(n7274) );
  OAI21_X1 U8852 ( .B1(n8546), .B2(n7997), .A(n7270), .ZN(n7272) );
  OAI22_X1 U8853 ( .A1(n7992), .A2(n8547), .B1(n8548), .B2(n7993), .ZN(n7271)
         );
  AOI211_X1 U8854 ( .C1(n10185), .C2(n8551), .A(n7272), .B(n7271), .ZN(n7273)
         );
  OAI21_X1 U8855 ( .B1(n7274), .B2(n8553), .A(n7273), .ZN(P2_U3219) );
  INV_X1 U8856 ( .A(n8208), .ZN(n8109) );
  OAI222_X1 U8857 ( .A1(P1_U3084), .A2(n9393), .B1(n7925), .B2(n8109), .C1(
        n8209), .C2(n9791), .ZN(P1_U3331) );
  INV_X1 U8858 ( .A(n7712), .ZN(n9453) );
  OR2_X1 U8859 ( .A1(n7492), .A2(n9453), .ZN(n7275) );
  NAND2_X1 U8860 ( .A1(n7276), .A2(n7275), .ZN(n7546) );
  NAND2_X1 U8861 ( .A1(n7277), .A2(n9151), .ZN(n7279) );
  AOI22_X1 U8862 ( .A1(n8150), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8149), .B2(
        n9476), .ZN(n7278) );
  OR2_X1 U8863 ( .A1(n9765), .A2(n9866), .ZN(n7547) );
  NAND2_X1 U8864 ( .A1(n9765), .A2(n9866), .ZN(n7545) );
  AND2_X1 U8865 ( .A1(n7547), .A2(n7545), .ZN(n9309) );
  XNOR2_X1 U8866 ( .A(n7546), .B(n9309), .ZN(n9764) );
  INV_X1 U8867 ( .A(n9297), .ZN(n7280) );
  XOR2_X1 U8868 ( .A(n7577), .B(n9309), .Z(n7289) );
  NAND2_X1 U8869 ( .A1(n8421), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7287) );
  OR2_X1 U8870 ( .A1(n8333), .A2(n6569), .ZN(n7286) );
  NAND2_X1 U8871 ( .A1(n7282), .A2(n7819), .ZN(n7283) );
  NAND2_X1 U8872 ( .A1(n7559), .A2(n7283), .ZN(n9871) );
  OR2_X1 U8873 ( .A1(n8332), .A2(n9871), .ZN(n7285) );
  INV_X1 U8874 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9479) );
  OR2_X1 U8875 ( .A1(n8425), .A2(n9479), .ZN(n7284) );
  INV_X1 U8876 ( .A(n7804), .ZN(n9452) );
  AOI22_X1 U8877 ( .A1(n9867), .A2(n9452), .B1(n9453), .B2(n9865), .ZN(n7288)
         );
  OAI21_X1 U8878 ( .B1(n7289), .B2(n9596), .A(n7288), .ZN(n7290) );
  AOI21_X1 U8879 ( .B1(n9764), .B2(n7765), .A(n7290), .ZN(n9769) );
  INV_X1 U8880 ( .A(n9765), .ZN(n7291) );
  AOI21_X1 U8881 ( .B1(n9765), .B2(n4421), .A(n9882), .ZN(n9767) );
  NOR2_X1 U8882 ( .A1(n7291), .A2(n9660), .ZN(n7294) );
  OAI22_X1 U8883 ( .A1(n9610), .A2(n7292), .B1(n7716), .B2(n10042), .ZN(n7293)
         );
  AOI211_X1 U8884 ( .C1(n9767), .C2(n9670), .A(n7294), .B(n7293), .ZN(n7296)
         );
  NAND2_X1 U8885 ( .A1(n9764), .A2(n7770), .ZN(n7295) );
  OAI211_X1 U8886 ( .C1(n9769), .C2(n4399), .A(n7296), .B(n7295), .ZN(P1_U3280) );
  NAND2_X1 U8887 ( .A1(n8222), .A2(n7773), .ZN(n7298) );
  OR2_X1 U8888 ( .A1(n7297), .A2(P1_U3084), .ZN(n9445) );
  OAI211_X1 U8889 ( .C1(n8223), .C2(n9791), .A(n7298), .B(n9445), .ZN(P1_U3330) );
  NAND2_X1 U8890 ( .A1(n8222), .A2(n7299), .ZN(n7301) );
  OAI211_X1 U8891 ( .C1(n7302), .C2(n8438), .A(n7301), .B(n7300), .ZN(P2_U3335) );
  OAI21_X1 U8892 ( .B1(n7304), .B2(n7161), .A(n7303), .ZN(n7312) );
  INV_X1 U8893 ( .A(n7304), .ZN(n7305) );
  NAND3_X1 U8894 ( .A1(n8493), .A2(n7306), .A3(n7305), .ZN(n7307) );
  AOI21_X1 U8895 ( .B1(n7307), .B2(n8548), .A(n4593), .ZN(n7311) );
  AOI22_X1 U8896 ( .A1(n8523), .A2(n5902), .B1(n7540), .B2(n8551), .ZN(n7309)
         );
  OAI211_X1 U8897 ( .C1(n7537), .C2(n8546), .A(n7309), .B(n7308), .ZN(n7310)
         );
  AOI211_X1 U8898 ( .C1(n7312), .C2(n8476), .A(n7311), .B(n7310), .ZN(n7313)
         );
  INV_X1 U8899 ( .A(n7313), .ZN(P2_U3241) );
  NOR2_X1 U8900 ( .A1(n8871), .A2(n10150), .ZN(n7317) );
  XNOR2_X1 U8901 ( .A(n7314), .B(n10150), .ZN(n10151) );
  OAI22_X1 U8902 ( .A1(n8656), .A2(n10151), .B1(n7315), .B2(n8835), .ZN(n7316)
         );
  AOI211_X1 U8903 ( .C1(n8878), .C2(P2_REG2_REG_1__SCAN_IN), .A(n7317), .B(
        n7316), .ZN(n7325) );
  INV_X1 U8904 ( .A(n8859), .ZN(n7368) );
  INV_X1 U8905 ( .A(n8849), .ZN(n8738) );
  OAI21_X1 U8906 ( .B1(n5806), .B2(n7319), .A(n7318), .ZN(n10154) );
  XNOR2_X1 U8907 ( .A(n5806), .B(n7320), .ZN(n7321) );
  NAND2_X1 U8908 ( .A1(n7321), .A2(n8863), .ZN(n7323) );
  AOI22_X1 U8909 ( .A1(n8821), .A2(n8568), .B1(n5875), .B2(n8819), .ZN(n7322)
         );
  NAND2_X1 U8910 ( .A1(n7323), .A2(n7322), .ZN(n10152) );
  AOI22_X1 U8911 ( .A1(n8738), .A2(n10154), .B1(n8846), .B2(n10152), .ZN(n7324) );
  NAND2_X1 U8912 ( .A1(n7325), .A2(n7324), .ZN(P2_U3295) );
  XNOR2_X1 U8913 ( .A(n7329), .B(n8063), .ZN(n8051) );
  XNOR2_X1 U8914 ( .A(n8051), .B(n7865), .ZN(n7338) );
  NOR2_X1 U8915 ( .A1(n7330), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7331) );
  NOR2_X1 U8916 ( .A1(n7332), .A2(n7331), .ZN(n8061) );
  XNOR2_X1 U8917 ( .A(n8061), .B(n8053), .ZN(n8065) );
  XNOR2_X1 U8918 ( .A(n8065), .B(P2_REG1_REG_15__SCAN_IN), .ZN(n7336) );
  AND2_X1 U8919 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7333) );
  AOI21_X1 U8920 ( .B1(n10124), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7333), .ZN(
        n7334) );
  OAI21_X1 U8921 ( .B1(n10121), .B2(n8063), .A(n7334), .ZN(n7335) );
  AOI21_X1 U8922 ( .B1(n7336), .B2(n10119), .A(n7335), .ZN(n7337) );
  OAI21_X1 U8923 ( .B1(n7338), .B2(n10122), .A(n7337), .ZN(P2_U3260) );
  INV_X1 U8924 ( .A(n7339), .ZN(n7340) );
  AOI21_X1 U8925 ( .B1(n9139), .B2(n9455), .A(n7340), .ZN(n7342) );
  NAND2_X1 U8926 ( .A1(n9128), .A2(n9457), .ZN(n7341) );
  OAI211_X1 U8927 ( .C1(n9142), .C2(n7343), .A(n7342), .B(n7341), .ZN(n7351)
         );
  INV_X1 U8928 ( .A(n7344), .ZN(n7349) );
  AOI21_X1 U8929 ( .B1(n7348), .B2(n7346), .A(n7345), .ZN(n7347) );
  AOI211_X1 U8930 ( .C1(n7349), .C2(n7348), .A(n9146), .B(n7347), .ZN(n7350)
         );
  AOI211_X1 U8931 ( .C1(n9144), .C2(n7352), .A(n7351), .B(n7350), .ZN(n7353)
         );
  INV_X1 U8932 ( .A(n7353), .ZN(P1_U3211) );
  INV_X1 U8933 ( .A(n10179), .ZN(n7354) );
  AND2_X1 U8934 ( .A1(n8562), .A2(n7354), .ZN(n7356) );
  OR2_X1 U8935 ( .A1(n7408), .A2(n7356), .ZN(n7358) );
  OR2_X1 U8936 ( .A1(n7597), .A2(n7358), .ZN(n7357) );
  OR2_X1 U8937 ( .A1(n7356), .A2(n7355), .ZN(n7359) );
  NAND2_X1 U8938 ( .A1(n7357), .A2(n7359), .ZN(n7363) );
  OR2_X1 U8939 ( .A1(n7597), .A2(n7982), .ZN(n7986) );
  INV_X1 U8940 ( .A(n7359), .ZN(n7360) );
  OAI21_X1 U8941 ( .B1(n7363), .B2(n7362), .A(n7361), .ZN(n7382) );
  XNOR2_X1 U8942 ( .A(n7364), .B(n7362), .ZN(n7366) );
  INV_X1 U8943 ( .A(n7397), .ZN(n8560) );
  AOI22_X1 U8944 ( .A1(n8560), .A2(n8821), .B1(n8819), .B2(n8562), .ZN(n7365)
         );
  OAI21_X1 U8945 ( .B1(n7366), .B2(n8759), .A(n7365), .ZN(n7367) );
  AOI21_X1 U8946 ( .B1(n7382), .B2(n7368), .A(n7367), .ZN(n7385) );
  INV_X1 U8947 ( .A(n7369), .ZN(n7371) );
  INV_X1 U8948 ( .A(n7999), .ZN(n7370) );
  AOI21_X1 U8949 ( .B1(n7598), .B2(n7371), .A(n7370), .ZN(n7383) );
  NAND2_X1 U8950 ( .A1(n7383), .A2(n8876), .ZN(n7375) );
  INV_X1 U8951 ( .A(n7372), .ZN(n7373) );
  INV_X1 U8952 ( .A(n8835), .ZN(n8868) );
  AOI22_X1 U8953 ( .A1(n8878), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7373), .B2(
        n8868), .ZN(n7374) );
  OAI211_X1 U8954 ( .C1(n7376), .C2(n8871), .A(n7375), .B(n7374), .ZN(n7377)
         );
  AOI21_X1 U8955 ( .B1(n7382), .B2(n7378), .A(n7377), .ZN(n7379) );
  OAI21_X1 U8956 ( .B1(n7385), .B2(n8878), .A(n7379), .ZN(P2_U3287) );
  INV_X1 U8957 ( .A(n8237), .ZN(n7402) );
  OAI222_X1 U8958 ( .A1(n8110), .A2(n7402), .B1(n7777), .B2(n7381), .C1(n7380), 
        .C2(n8438), .ZN(P2_U3334) );
  INV_X1 U8959 ( .A(n7382), .ZN(n7386) );
  AOI22_X1 U8960 ( .A1(n7383), .A2(n10195), .B1(n10194), .B2(n7598), .ZN(n7384) );
  OAI211_X1 U8961 ( .C1(n7386), .C2(n8977), .A(n7385), .B(n7384), .ZN(n7389)
         );
  NAND2_X1 U8962 ( .A1(n7389), .A2(n10217), .ZN(n7387) );
  OAI21_X1 U8963 ( .B1(n10217), .B2(n7388), .A(n7387), .ZN(P2_U3529) );
  NAND2_X1 U8964 ( .A1(n7389), .A2(n10204), .ZN(n7390) );
  OAI21_X1 U8965 ( .B1(n10204), .B2(n5289), .A(n7390), .ZN(P2_U3478) );
  INV_X1 U8966 ( .A(n7391), .ZN(n7394) );
  INV_X1 U8967 ( .A(n7392), .ZN(n7393) );
  XNOR2_X1 U8968 ( .A(n7730), .B(n8376), .ZN(n7625) );
  NOR2_X1 U8969 ( .A1(n7992), .A2(n5743), .ZN(n7626) );
  XNOR2_X1 U8970 ( .A(n7625), .B(n7626), .ZN(n7623) );
  XNOR2_X1 U8971 ( .A(n7624), .B(n7623), .ZN(n7401) );
  OAI22_X1 U8972 ( .A1(n8546), .A2(n7731), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8573), .ZN(n7399) );
  OAI22_X1 U8973 ( .A1(n7397), .A2(n8548), .B1(n8547), .B2(n7683), .ZN(n7398)
         );
  AOI211_X1 U8974 ( .C1(n7730), .C2(n8551), .A(n7399), .B(n7398), .ZN(n7400)
         );
  OAI21_X1 U8975 ( .B1(n7401), .B2(n8553), .A(n7400), .ZN(P2_U3238) );
  OAI222_X1 U8976 ( .A1(n7403), .A2(P1_U3084), .B1(n7925), .B2(n7402), .C1(
        n8238), .C2(n9791), .ZN(P1_U3329) );
  XNOR2_X1 U8977 ( .A(n7597), .B(n7404), .ZN(n7474) );
  NAND2_X1 U8978 ( .A1(n7531), .A2(n7405), .ZN(n7406) );
  NAND2_X1 U8979 ( .A1(n7406), .A2(n7528), .ZN(n7529) );
  NAND2_X1 U8980 ( .A1(n7529), .A2(n7407), .ZN(n7409) );
  XNOR2_X1 U8981 ( .A(n7409), .B(n7408), .ZN(n7410) );
  AOI222_X1 U8982 ( .A1(n8563), .A2(n8819), .B1(n8562), .B2(n8821), .C1(n8863), 
        .C2(n7410), .ZN(n7466) );
  AOI21_X1 U8983 ( .B1(n7412), .B2(n7535), .A(n7411), .ZN(n7471) );
  AOI22_X1 U8984 ( .A1(n7471), .A2(n10195), .B1(n10194), .B2(n7412), .ZN(n7413) );
  OAI211_X1 U8985 ( .C1(n10199), .C2(n7474), .A(n7466), .B(n7413), .ZN(n7415)
         );
  NAND2_X1 U8986 ( .A1(n7415), .A2(n10204), .ZN(n7414) );
  OAI21_X1 U8987 ( .B1(n10204), .B2(n5242), .A(n7414), .ZN(P2_U3472) );
  NAND2_X1 U8988 ( .A1(n7415), .A2(n10217), .ZN(n7416) );
  OAI21_X1 U8989 ( .B1(n10217), .B2(n6712), .A(n7416), .ZN(P2_U3527) );
  AOI22_X1 U8990 ( .A1(n7417), .A2(n9881), .B1(n9766), .B2(n7451), .ZN(n7418)
         );
  OAI211_X1 U8991 ( .C1(n10065), .C2(n7420), .A(n7419), .B(n7418), .ZN(n7422)
         );
  NAND2_X1 U8992 ( .A1(n7422), .A2(n10117), .ZN(n7421) );
  OAI21_X1 U8993 ( .B1(n10117), .B2(n6157), .A(n7421), .ZN(P1_U3532) );
  NAND2_X1 U8994 ( .A1(n7422), .A2(n10107), .ZN(n7423) );
  OAI21_X1 U8995 ( .B1(n10107), .B2(n6161), .A(n7423), .ZN(P1_U3481) );
  OAI21_X1 U8996 ( .B1(n7426), .B2(n7425), .A(n7424), .ZN(n10160) );
  INV_X1 U8997 ( .A(n10160), .ZN(n7440) );
  NOR2_X1 U8998 ( .A1(n8835), .A2(n7427), .ZN(n7431) );
  OAI21_X1 U8999 ( .B1(n4637), .B2(n10146), .A(n4639), .ZN(n7429) );
  NAND2_X1 U9000 ( .A1(n7429), .A2(n7428), .ZN(n10157) );
  NOR2_X1 U9001 ( .A1(n8656), .A2(n10157), .ZN(n7430) );
  AOI211_X1 U9002 ( .C1(n8878), .C2(P2_REG2_REG_2__SCAN_IN), .A(n7431), .B(
        n7430), .ZN(n7439) );
  OAI21_X1 U9003 ( .B1(n7434), .B2(n7433), .A(n7432), .ZN(n7435) );
  NAND2_X1 U9004 ( .A1(n7435), .A2(n8863), .ZN(n7437) );
  AOI22_X1 U9005 ( .A1(n8819), .A2(n7441), .B1(n8566), .B2(n8821), .ZN(n7436)
         );
  NAND2_X1 U9006 ( .A1(n7437), .A2(n7436), .ZN(n10158) );
  AOI22_X1 U9007 ( .A1(n10158), .A2(n8846), .B1(n8691), .B2(n4639), .ZN(n7438)
         );
  OAI211_X1 U9008 ( .C1(n7440), .C2(n8849), .A(n7439), .B(n7438), .ZN(P2_U3294) );
  AOI22_X1 U9009 ( .A1(n10147), .A2(n8863), .B1(n8821), .B2(n7441), .ZN(n10149) );
  OAI22_X1 U9010 ( .A1(n8878), .A2(n10149), .B1(n7442), .B2(n8835), .ZN(n7443)
         );
  AOI21_X1 U9011 ( .B1(n8878), .B2(P2_REG2_REG_0__SCAN_IN), .A(n7443), .ZN(
        n7445) );
  OAI21_X1 U9012 ( .B1(n8691), .B2(n8876), .A(n10146), .ZN(n7444) );
  OAI211_X1 U9013 ( .C1(n7446), .C2(n8849), .A(n7445), .B(n7444), .ZN(P2_U3296) );
  NAND2_X1 U9014 ( .A1(n7451), .A2(n8307), .ZN(n7448) );
  NAND2_X1 U9015 ( .A1(n9454), .A2(n7480), .ZN(n7447) );
  NAND2_X1 U9016 ( .A1(n7448), .A2(n7447), .ZN(n7449) );
  XNOR2_X1 U9017 ( .A(n7449), .B(n8322), .ZN(n7475) );
  AND2_X1 U9018 ( .A1(n9454), .A2(n8324), .ZN(n7450) );
  AOI21_X1 U9019 ( .B1(n7451), .B2(n8319), .A(n7450), .ZN(n7476) );
  XNOR2_X1 U9020 ( .A(n7475), .B(n7476), .ZN(n7457) );
  NAND2_X1 U9021 ( .A1(n7453), .A2(n7452), .ZN(n7455) );
  NAND2_X1 U9022 ( .A1(n7455), .A2(n7454), .ZN(n7456) );
  OAI21_X1 U9023 ( .B1(n7457), .B2(n7456), .A(n7479), .ZN(n7458) );
  NAND2_X1 U9024 ( .A1(n7458), .A2(n9119), .ZN(n7464) );
  NOR2_X1 U9025 ( .A1(n9142), .A2(n7459), .ZN(n7462) );
  OAI22_X1 U9026 ( .A1(n9125), .A2(n7712), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7460), .ZN(n7461) );
  AOI211_X1 U9027 ( .C1(n9128), .C2(n9455), .A(n7462), .B(n7461), .ZN(n7463)
         );
  OAI211_X1 U9028 ( .C1(n7465), .C2(n9131), .A(n7464), .B(n7463), .ZN(P1_U3229) );
  OR2_X1 U9029 ( .A1(n7466), .A2(n8878), .ZN(n7473) );
  OAI22_X1 U9030 ( .A1(n8835), .A2(n7467), .B1(n6742), .B2(n8846), .ZN(n7470)
         );
  NOR2_X1 U9031 ( .A1(n8871), .A2(n7468), .ZN(n7469) );
  AOI211_X1 U9032 ( .C1(n7471), .C2(n8876), .A(n7470), .B(n7469), .ZN(n7472)
         );
  OAI211_X1 U9033 ( .C1(n7474), .C2(n8849), .A(n7473), .B(n7472), .ZN(P2_U3289) );
  INV_X1 U9034 ( .A(n7475), .ZN(n7477) );
  NAND2_X1 U9035 ( .A1(n7477), .A2(n7476), .ZN(n7478) );
  NAND2_X1 U9036 ( .A1(n7492), .A2(n8307), .ZN(n7482) );
  NAND2_X1 U9037 ( .A1(n9453), .A2(n7480), .ZN(n7481) );
  NAND2_X1 U9038 ( .A1(n7482), .A2(n7481), .ZN(n7483) );
  XNOR2_X1 U9039 ( .A(n7483), .B(n8184), .ZN(n7703) );
  NOR2_X1 U9040 ( .A1(n7712), .A2(n8300), .ZN(n7484) );
  AOI21_X1 U9041 ( .B1(n7492), .B2(n7480), .A(n7484), .ZN(n7704) );
  XNOR2_X1 U9042 ( .A(n7703), .B(n7704), .ZN(n7485) );
  XNOR2_X1 U9043 ( .A(n7702), .B(n7485), .ZN(n7494) );
  NOR2_X1 U9044 ( .A1(n9137), .A2(n7486), .ZN(n7487) );
  AOI211_X1 U9045 ( .C1(n9139), .C2(n9866), .A(n7488), .B(n7487), .ZN(n7489)
         );
  OAI21_X1 U9046 ( .B1(n9142), .B2(n7490), .A(n7489), .ZN(n7491) );
  AOI21_X1 U9047 ( .B1(n9144), .B2(n7492), .A(n7491), .ZN(n7493) );
  OAI21_X1 U9048 ( .B1(n7494), .B2(n9146), .A(n7493), .ZN(P1_U3215) );
  OAI21_X1 U9049 ( .B1(n7496), .B2(n7497), .A(n7495), .ZN(n10166) );
  INV_X1 U9050 ( .A(n10166), .ZN(n7514) );
  NAND2_X1 U9051 ( .A1(n7651), .A2(n8863), .ZN(n7503) );
  INV_X1 U9052 ( .A(n7497), .ZN(n7498) );
  AOI21_X1 U9053 ( .B1(n7500), .B2(n7499), .A(n7498), .ZN(n7502) );
  AOI22_X1 U9054 ( .A1(n8819), .A2(n8566), .B1(n8564), .B2(n8821), .ZN(n7501)
         );
  OAI21_X1 U9055 ( .B1(n7503), .B2(n7502), .A(n7501), .ZN(n10164) );
  AND2_X1 U9056 ( .A1(n7505), .A2(n7504), .ZN(n7506) );
  OR2_X1 U9057 ( .A1(n7506), .A2(n7660), .ZN(n10163) );
  INV_X1 U9058 ( .A(n10163), .ZN(n7509) );
  NOR2_X1 U9059 ( .A1(n8835), .A2(n7507), .ZN(n7508) );
  AOI21_X1 U9060 ( .B1(n8876), .B2(n7509), .A(n7508), .ZN(n7511) );
  NAND2_X1 U9061 ( .A1(n8878), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7510) );
  OAI211_X1 U9062 ( .C1(n10162), .C2(n8871), .A(n7511), .B(n7510), .ZN(n7512)
         );
  AOI21_X1 U9063 ( .B1(n10164), .B2(n8846), .A(n7512), .ZN(n7513) );
  OAI21_X1 U9064 ( .B1(n7514), .B2(n8849), .A(n7513), .ZN(P2_U3292) );
  OAI22_X1 U9065 ( .A1(n8656), .A2(n7515), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8835), .ZN(n7517) );
  NOR2_X1 U9066 ( .A1(n8846), .A2(n6734), .ZN(n7516) );
  NOR2_X1 U9067 ( .A1(n7517), .A2(n7516), .ZN(n7520) );
  NAND2_X1 U9068 ( .A1(n8691), .A2(n7518), .ZN(n7519) );
  OAI211_X1 U9069 ( .C1(n7521), .C2(n8873), .A(n7520), .B(n7519), .ZN(n7522)
         );
  AOI21_X1 U9070 ( .B1(n7523), .B2(n8846), .A(n7522), .ZN(n7524) );
  INV_X1 U9071 ( .A(n7524), .ZN(P2_U3293) );
  XNOR2_X1 U9072 ( .A(n7526), .B(n7525), .ZN(n10176) );
  INV_X1 U9073 ( .A(n10176), .ZN(n7544) );
  NOR2_X1 U9074 ( .A1(n7528), .A2(n7527), .ZN(n7532) );
  INV_X1 U9075 ( .A(n7529), .ZN(n7530) );
  AOI21_X1 U9076 ( .B1(n7532), .B2(n7531), .A(n7530), .ZN(n7533) );
  OAI222_X1 U9077 ( .A1(n8851), .A2(n7534), .B1(n8853), .B2(n4593), .C1(n8759), 
        .C2(n7533), .ZN(n10174) );
  INV_X1 U9078 ( .A(n7659), .ZN(n7536) );
  OAI21_X1 U9079 ( .B1(n7536), .B2(n10172), .A(n7535), .ZN(n10173) );
  INV_X1 U9080 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7538) );
  OAI22_X1 U9081 ( .A1(n8846), .A2(n7538), .B1(n7537), .B2(n8835), .ZN(n7539)
         );
  AOI21_X1 U9082 ( .B1(n8691), .B2(n7540), .A(n7539), .ZN(n7541) );
  OAI21_X1 U9083 ( .B1(n8656), .B2(n10173), .A(n7541), .ZN(n7542) );
  AOI21_X1 U9084 ( .B1(n10174), .B2(n8846), .A(n7542), .ZN(n7543) );
  OAI21_X1 U9085 ( .B1(n7544), .B2(n8849), .A(n7543), .ZN(P2_U3290) );
  NAND2_X1 U9086 ( .A1(n7546), .A2(n7545), .ZN(n7548) );
  NAND2_X1 U9087 ( .A1(n7548), .A2(n7547), .ZN(n9878) );
  INV_X1 U9088 ( .A(n9878), .ZN(n7553) );
  NAND2_X1 U9089 ( .A1(n7549), .A2(n9151), .ZN(n7551) );
  AOI22_X1 U9090 ( .A1(n8150), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8149), .B2(
        n9947), .ZN(n7550) );
  OR2_X1 U9091 ( .A1(n9875), .A2(n7804), .ZN(n9302) );
  NAND2_X1 U9092 ( .A1(n9875), .A2(n7804), .ZN(n9298) );
  INV_X1 U9093 ( .A(n9879), .ZN(n7552) );
  NAND2_X1 U9094 ( .A1(n9875), .A2(n9452), .ZN(n7554) );
  NAND2_X1 U9095 ( .A1(n7555), .A2(n9151), .ZN(n7557) );
  AOI22_X1 U9096 ( .A1(n8150), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n8149), .B2(
        n9956), .ZN(n7556) );
  NAND2_X1 U9097 ( .A1(n6030), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7565) );
  INV_X1 U9098 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7558) );
  NAND2_X1 U9099 ( .A1(n7559), .A2(n7558), .ZN(n7560) );
  NAND2_X1 U9100 ( .A1(n7570), .A2(n7560), .ZN(n7807) );
  OR2_X1 U9101 ( .A1(n8332), .A2(n7807), .ZN(n7564) );
  INV_X1 U9102 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9463) );
  OR2_X1 U9103 ( .A1(n8333), .A2(n9463), .ZN(n7563) );
  INV_X1 U9104 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7561) );
  OR2_X1 U9105 ( .A1(n5996), .A2(n7561), .ZN(n7562) );
  NAND4_X1 U9106 ( .A1(n7565), .A2(n7564), .A3(n7563), .A4(n7562), .ZN(n9868)
         );
  OR2_X1 U9107 ( .A1(n9759), .A2(n9868), .ZN(n7566) );
  NAND2_X1 U9108 ( .A1(n7567), .A2(n9151), .ZN(n7569) );
  INV_X1 U9109 ( .A(n9483), .ZN(n9974) );
  AOI22_X1 U9110 ( .A1(n8150), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n8149), .B2(
        n9974), .ZN(n7568) );
  NAND2_X1 U9111 ( .A1(n6030), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7576) );
  INV_X1 U9112 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7973) );
  AND2_X1 U9113 ( .A1(n7570), .A2(n7973), .ZN(n7571) );
  OR2_X1 U9114 ( .A1(n7571), .A2(n7579), .ZN(n7977) );
  OR2_X1 U9115 ( .A1(n8332), .A2(n7977), .ZN(n7575) );
  INV_X1 U9116 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n7572) );
  OR2_X1 U9117 ( .A1(n5996), .A2(n7572), .ZN(n7574) );
  INV_X1 U9118 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7590) );
  OR2_X1 U9119 ( .A1(n8333), .A2(n7590), .ZN(n7573) );
  NAND4_X1 U9120 ( .A1(n7576), .A2(n7575), .A3(n7574), .A4(n7573), .ZN(n9451)
         );
  INV_X1 U9121 ( .A(n9451), .ZN(n9136) );
  NAND2_X1 U9122 ( .A1(n7979), .A2(n9136), .ZN(n9312) );
  XNOR2_X1 U9123 ( .A(n7747), .B(n4470), .ZN(n9892) );
  INV_X1 U9124 ( .A(n9892), .ZN(n7595) );
  INV_X1 U9125 ( .A(n9866), .ZN(n7820) );
  NAND2_X1 U9126 ( .A1(n9765), .A2(n7820), .ZN(n9162) );
  OR2_X1 U9127 ( .A1(n9765), .A2(n7820), .ZN(n9862) );
  AND2_X1 U9128 ( .A1(n9302), .A2(n9862), .ZN(n9214) );
  INV_X1 U9129 ( .A(n9868), .ZN(n7974) );
  OR2_X1 U9130 ( .A1(n9759), .A2(n7974), .ZN(n9220) );
  NAND2_X1 U9131 ( .A1(n9759), .A2(n7974), .ZN(n9216) );
  OAI211_X1 U9132 ( .C1(n4955), .C2(n4470), .A(n7751), .B(n9870), .ZN(n7588)
         );
  NAND2_X1 U9133 ( .A1(n7579), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7757) );
  OR2_X1 U9134 ( .A1(n7579), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7580) );
  NAND2_X1 U9135 ( .A1(n7757), .A2(n7580), .ZN(n9141) );
  OR2_X1 U9136 ( .A1(n8332), .A2(n9141), .ZN(n7586) );
  OR2_X1 U9137 ( .A1(n8425), .A2(n7581), .ZN(n7585) );
  INV_X1 U9138 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7582) );
  OR2_X1 U9139 ( .A1(n5996), .A2(n7582), .ZN(n7584) );
  INV_X1 U9140 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7767) );
  OR2_X1 U9141 ( .A1(n8333), .A2(n7767), .ZN(n7583) );
  NAND4_X1 U9142 ( .A1(n7586), .A2(n7585), .A3(n7584), .A4(n7583), .ZN(n9450)
         );
  AOI22_X1 U9143 ( .A1(n9865), .A2(n9868), .B1(n9450), .B2(n9867), .ZN(n7587)
         );
  NAND2_X1 U9144 ( .A1(n7588), .A2(n7587), .ZN(n9891) );
  INV_X1 U9145 ( .A(n9875), .ZN(n9896) );
  INV_X1 U9146 ( .A(n7589), .ZN(n7721) );
  INV_X1 U9147 ( .A(n7979), .ZN(n9889) );
  OAI211_X1 U9148 ( .C1(n7721), .C2(n9889), .A(n9881), .B(n7766), .ZN(n9888)
         );
  OAI22_X1 U9149 ( .A1(n9610), .A2(n7590), .B1(n7977), .B2(n10042), .ZN(n7591)
         );
  AOI21_X1 U9150 ( .B1(n7979), .B2(n9874), .A(n7591), .ZN(n7592) );
  OAI21_X1 U9151 ( .B1(n9888), .B2(n8038), .A(n7592), .ZN(n7593) );
  AOI21_X1 U9152 ( .B1(n9891), .B2(n9610), .A(n7593), .ZN(n7594) );
  OAI21_X1 U9153 ( .B1(n7595), .B2(n9672), .A(n7594), .ZN(P1_U3277) );
  NAND2_X1 U9154 ( .A1(n10185), .A2(n8560), .ZN(n7601) );
  NOR2_X1 U9155 ( .A1(n7597), .A2(n7596), .ZN(n7603) );
  OR2_X1 U9156 ( .A1(n7598), .A2(n8561), .ZN(n7599) );
  AND2_X1 U9157 ( .A1(n7601), .A2(n7983), .ZN(n7602) );
  NOR2_X1 U9158 ( .A1(n7603), .A2(n7602), .ZN(n7636) );
  NAND2_X1 U9159 ( .A1(n7636), .A2(n7638), .ZN(n7605) );
  INV_X1 U9160 ( .A(n7992), .ZN(n8559) );
  NAND2_X1 U9161 ( .A1(n7730), .A2(n8559), .ZN(n7604) );
  XOR2_X1 U9162 ( .A(n7685), .B(n7684), .Z(n10200) );
  NAND2_X1 U9163 ( .A1(n7607), .A2(n7606), .ZN(n7609) );
  INV_X1 U9164 ( .A(n7684), .ZN(n7608) );
  XNOR2_X1 U9165 ( .A(n7609), .B(n7608), .ZN(n7611) );
  OAI22_X1 U9166 ( .A1(n7883), .A2(n8851), .B1(n7992), .B2(n8853), .ZN(n7610)
         );
  AOI21_X1 U9167 ( .B1(n7611), .B2(n8863), .A(n7610), .ZN(n10198) );
  OAI22_X1 U9168 ( .A1(n8846), .A2(n7612), .B1(n7631), .B2(n8835), .ZN(n7613)
         );
  AOI21_X1 U9169 ( .B1(n8691), .B2(n10193), .A(n7613), .ZN(n7616) );
  AND2_X1 U9170 ( .A1(n7640), .A2(n10193), .ZN(n7614) );
  NOR2_X1 U9171 ( .A1(n7696), .A2(n7614), .ZN(n10196) );
  NAND2_X1 U9172 ( .A1(n10196), .A2(n8876), .ZN(n7615) );
  OAI211_X1 U9173 ( .C1(n10198), .C2(n8878), .A(n7616), .B(n7615), .ZN(n7617)
         );
  INV_X1 U9174 ( .A(n7617), .ZN(n7618) );
  OAI21_X1 U9175 ( .B1(n10200), .B2(n8849), .A(n7618), .ZN(P2_U3284) );
  XNOR2_X1 U9176 ( .A(n10193), .B(n8376), .ZN(n7622) );
  INV_X1 U9177 ( .A(n7622), .ZN(n7620) );
  OR2_X1 U9178 ( .A1(n7683), .A2(n5743), .ZN(n7621) );
  INV_X1 U9179 ( .A(n7621), .ZN(n7619) );
  NAND2_X1 U9180 ( .A1(n7620), .A2(n7619), .ZN(n7673) );
  NAND2_X1 U9181 ( .A1(n7622), .A2(n7621), .ZN(n7671) );
  NAND2_X1 U9182 ( .A1(n7673), .A2(n7671), .ZN(n7629) );
  INV_X1 U9183 ( .A(n7625), .ZN(n7627) );
  NAND2_X1 U9184 ( .A1(n7627), .A2(n7626), .ZN(n7628) );
  XOR2_X1 U9185 ( .A(n7629), .B(n7672), .Z(n7635) );
  OAI21_X1 U9186 ( .B1(n8546), .B2(n7631), .A(n7630), .ZN(n7633) );
  OAI22_X1 U9187 ( .A1(n7992), .A2(n8548), .B1(n8547), .B2(n7883), .ZN(n7632)
         );
  AOI211_X1 U9188 ( .C1(n10193), .C2(n8551), .A(n7633), .B(n7632), .ZN(n7634)
         );
  OAI21_X1 U9189 ( .B1(n7635), .B2(n8553), .A(n7634), .ZN(P2_U3226) );
  XNOR2_X1 U9190 ( .A(n7636), .B(n7638), .ZN(n7740) );
  XNOR2_X1 U9191 ( .A(n7637), .B(n7638), .ZN(n7639) );
  INV_X1 U9192 ( .A(n7683), .ZN(n8558) );
  AOI222_X1 U9193 ( .A1(n8863), .A2(n7639), .B1(n8558), .B2(n8821), .C1(n8560), 
        .C2(n8819), .ZN(n7735) );
  INV_X1 U9194 ( .A(n7640), .ZN(n7641) );
  AOI21_X1 U9195 ( .B1(n7730), .B2(n8001), .A(n7641), .ZN(n7738) );
  AOI22_X1 U9196 ( .A1(n7738), .A2(n10195), .B1(n10194), .B2(n7730), .ZN(n7642) );
  OAI211_X1 U9197 ( .C1(n7740), .C2(n10199), .A(n7735), .B(n7642), .ZN(n7644)
         );
  NAND2_X1 U9198 ( .A1(n7644), .A2(n10217), .ZN(n7643) );
  OAI21_X1 U9199 ( .B1(n10217), .B2(n6925), .A(n7643), .ZN(P2_U3531) );
  NAND2_X1 U9200 ( .A1(n7644), .A2(n10204), .ZN(n7645) );
  OAI21_X1 U9201 ( .B1(n10204), .B2(n5328), .A(n7645), .ZN(P2_U3484) );
  INV_X1 U9202 ( .A(n8254), .ZN(n7648) );
  OAI222_X1 U9203 ( .A1(P1_U3084), .A2(n7646), .B1(n7925), .B2(n7648), .C1(
        n8255), .C2(n9791), .ZN(P1_U3328) );
  OAI222_X1 U9204 ( .A1(n8438), .A2(n7649), .B1(n8110), .B2(n7648), .C1(n7647), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  NAND2_X1 U9205 ( .A1(n7651), .A2(n7650), .ZN(n7652) );
  XOR2_X1 U9206 ( .A(n7655), .B(n7652), .Z(n7654) );
  AOI21_X1 U9207 ( .B1(n7654), .B2(n8863), .A(n7653), .ZN(n10168) );
  XOR2_X1 U9208 ( .A(n7656), .B(n7655), .Z(n10171) );
  NAND2_X1 U9209 ( .A1(n10171), .A2(n8738), .ZN(n7666) );
  INV_X1 U9210 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7658) );
  OAI22_X1 U9211 ( .A1(n8846), .A2(n7658), .B1(n7657), .B2(n8835), .ZN(n7663)
         );
  NOR2_X1 U9212 ( .A1(n8878), .A2(n5458), .ZN(n8840) );
  INV_X1 U9213 ( .A(n8840), .ZN(n7661) );
  OAI211_X1 U9214 ( .C1(n7660), .C2(n10169), .A(n7659), .B(n10195), .ZN(n10167) );
  NOR2_X1 U9215 ( .A1(n7661), .A2(n10167), .ZN(n7662) );
  AOI211_X1 U9216 ( .C1(n8691), .C2(n7664), .A(n7663), .B(n7662), .ZN(n7665)
         );
  OAI211_X1 U9217 ( .C1(n8878), .C2(n10168), .A(n7666), .B(n7665), .ZN(
        P2_U3291) );
  INV_X1 U9218 ( .A(n8972), .ZN(n7695) );
  XNOR2_X1 U9219 ( .A(n8972), .B(n8365), .ZN(n7667) );
  NOR2_X1 U9220 ( .A1(n7883), .A2(n5743), .ZN(n7668) );
  NAND2_X1 U9221 ( .A1(n7667), .A2(n7668), .ZN(n7855) );
  INV_X1 U9222 ( .A(n7667), .ZN(n7850) );
  INV_X1 U9223 ( .A(n7668), .ZN(n7669) );
  NAND2_X1 U9224 ( .A1(n7850), .A2(n7669), .ZN(n7670) );
  AND2_X1 U9225 ( .A1(n7855), .A2(n7670), .ZN(n7675) );
  OAI211_X1 U9226 ( .C1(n7675), .C2(n7674), .A(n7857), .B(n8476), .ZN(n7680)
         );
  INV_X1 U9227 ( .A(n7692), .ZN(n7678) );
  OAI22_X1 U9228 ( .A1(n7898), .A2(n8547), .B1(n8548), .B2(n7683), .ZN(n7676)
         );
  AOI211_X1 U9229 ( .C1(n8538), .C2(n7678), .A(n7677), .B(n7676), .ZN(n7679)
         );
  OAI211_X1 U9230 ( .C1(n7695), .C2(n8541), .A(n7680), .B(n7679), .ZN(P2_U3236) );
  OAI21_X1 U9231 ( .B1(n7686), .B2(n7681), .A(n7682), .ZN(n7691) );
  OAI22_X1 U9232 ( .A1(n7683), .A2(n8853), .B1(n7898), .B2(n8851), .ZN(n7690)
         );
  NAND2_X1 U9233 ( .A1(n7687), .A2(n7686), .ZN(n7688) );
  NAND2_X1 U9234 ( .A1(n7868), .A2(n7688), .ZN(n8976) );
  NOR2_X1 U9235 ( .A1(n8976), .A2(n8859), .ZN(n7689) );
  AOI211_X1 U9236 ( .C1(n8863), .C2(n7691), .A(n7690), .B(n7689), .ZN(n8975)
         );
  OAI22_X1 U9237 ( .A1(n8846), .A2(n7693), .B1(n7692), .B2(n8835), .ZN(n7694)
         );
  AOI21_X1 U9238 ( .B1(n8972), .B2(n8691), .A(n7694), .ZN(n7699) );
  OR2_X1 U9239 ( .A1(n7696), .A2(n7695), .ZN(n7697) );
  NAND2_X1 U9240 ( .A1(n7696), .A2(n7695), .ZN(n7876) );
  AND2_X1 U9241 ( .A1(n7697), .A2(n7876), .ZN(n8973) );
  NAND2_X1 U9242 ( .A1(n8973), .A2(n8876), .ZN(n7698) );
  OAI211_X1 U9243 ( .C1(n8976), .C2(n8873), .A(n7699), .B(n7698), .ZN(n7700)
         );
  INV_X1 U9244 ( .A(n7700), .ZN(n7701) );
  OAI21_X1 U9245 ( .B1(n8975), .B2(n8878), .A(n7701), .ZN(P2_U3283) );
  INV_X1 U9246 ( .A(n7703), .ZN(n7706) );
  INV_X1 U9247 ( .A(n7704), .ZN(n7705) );
  NAND2_X1 U9248 ( .A1(n7706), .A2(n7705), .ZN(n7792) );
  NAND2_X1 U9249 ( .A1(n7797), .A2(n7792), .ZN(n7814) );
  NAND2_X1 U9250 ( .A1(n9765), .A2(n8307), .ZN(n7708) );
  NAND2_X1 U9251 ( .A1(n9866), .A2(n7480), .ZN(n7707) );
  NAND2_X1 U9252 ( .A1(n7708), .A2(n7707), .ZN(n7709) );
  XNOR2_X1 U9253 ( .A(n7709), .B(n8322), .ZN(n7785) );
  AND2_X1 U9254 ( .A1(n9866), .A2(n8324), .ZN(n7711) );
  AOI21_X1 U9255 ( .B1(n9765), .B2(n7480), .A(n7711), .ZN(n7783) );
  XNOR2_X1 U9256 ( .A(n7785), .B(n7783), .ZN(n7813) );
  XNOR2_X1 U9257 ( .A(n7814), .B(n7813), .ZN(n7719) );
  NOR2_X1 U9258 ( .A1(n9137), .A2(n7712), .ZN(n7713) );
  AOI211_X1 U9259 ( .C1(n9139), .C2(n9452), .A(n7714), .B(n7713), .ZN(n7715)
         );
  OAI21_X1 U9260 ( .B1(n9142), .B2(n7716), .A(n7715), .ZN(n7717) );
  AOI21_X1 U9261 ( .B1(n9144), .B2(n9765), .A(n7717), .ZN(n7718) );
  OAI21_X1 U9262 ( .B1(n7719), .B2(n9146), .A(n7718), .ZN(P1_U3234) );
  XOR2_X1 U9263 ( .A(n7720), .B(n9178), .Z(n9763) );
  AOI21_X1 U9264 ( .B1(n9759), .B2(n9880), .A(n7721), .ZN(n9760) );
  INV_X1 U9265 ( .A(n9759), .ZN(n7724) );
  INV_X1 U9266 ( .A(n7807), .ZN(n7722) );
  AOI22_X1 U9267 ( .A1(n4399), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7722), .B2(
        n9872), .ZN(n7723) );
  OAI21_X1 U9268 ( .B1(n7724), .B2(n9660), .A(n7723), .ZN(n7728) );
  XNOR2_X1 U9269 ( .A(n7725), .B(n9178), .ZN(n7726) );
  AOI222_X1 U9270 ( .A1(n9870), .A2(n7726), .B1(n9451), .B2(n9867), .C1(n9452), 
        .C2(n9865), .ZN(n9762) );
  NOR2_X1 U9271 ( .A1(n9762), .A2(n4399), .ZN(n7727) );
  AOI211_X1 U9272 ( .C1(n9760), .C2(n9670), .A(n7728), .B(n7727), .ZN(n7729)
         );
  OAI21_X1 U9273 ( .B1(n9763), .B2(n9672), .A(n7729), .ZN(P1_U3278) );
  INV_X1 U9274 ( .A(n7730), .ZN(n7734) );
  INV_X1 U9275 ( .A(n7731), .ZN(n7732) );
  AOI22_X1 U9276 ( .A1(n8878), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7732), .B2(
        n8868), .ZN(n7733) );
  OAI21_X1 U9277 ( .B1(n7734), .B2(n8871), .A(n7733), .ZN(n7737) );
  NOR2_X1 U9278 ( .A1(n7735), .A2(n8878), .ZN(n7736) );
  AOI211_X1 U9279 ( .C1(n7738), .C2(n8876), .A(n7737), .B(n7736), .ZN(n7739)
         );
  OAI21_X1 U9280 ( .B1(n8849), .B2(n7740), .A(n7739), .ZN(P2_U3285) );
  INV_X1 U9281 ( .A(n8270), .ZN(n7743) );
  OAI222_X1 U9282 ( .A1(n8110), .A2(n7743), .B1(P2_U3152), .B2(n7742), .C1(
        n7741), .C2(n8438), .ZN(P2_U3332) );
  OAI222_X1 U9283 ( .A1(n7744), .A2(P1_U3084), .B1(n7925), .B2(n7743), .C1(
        n8271), .C2(n9791), .ZN(P1_U3327) );
  AND2_X1 U9284 ( .A1(n7979), .A2(n9451), .ZN(n7746) );
  OR2_X1 U9285 ( .A1(n7979), .A2(n9451), .ZN(n7745) );
  NAND2_X1 U9286 ( .A1(n7748), .A2(n9151), .ZN(n7750) );
  AOI22_X1 U9287 ( .A1(n8150), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9986), .B2(
        n8149), .ZN(n7749) );
  OR2_X1 U9288 ( .A1(n9754), .A2(n9060), .ZN(n9318) );
  NAND2_X1 U9289 ( .A1(n9754), .A2(n9060), .ZN(n9319) );
  NAND2_X1 U9290 ( .A1(n9318), .A2(n9319), .ZN(n9161) );
  XNOR2_X1 U9291 ( .A(n7828), .B(n9161), .ZN(n9753) );
  NAND2_X1 U9292 ( .A1(n7754), .A2(n9161), .ZN(n7755) );
  AOI21_X1 U9293 ( .B1(n7840), .B2(n7755), .A(n9596), .ZN(n7764) );
  NAND2_X1 U9294 ( .A1(n5995), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7762) );
  INV_X1 U9295 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n7756) );
  OR2_X1 U9296 ( .A1(n5996), .A2(n7756), .ZN(n7761) );
  NAND2_X1 U9297 ( .A1(n7757), .A2(n9058), .ZN(n7758) );
  NAND2_X1 U9298 ( .A1(n7833), .A2(n7758), .ZN(n7845) );
  OR2_X1 U9299 ( .A1(n7845), .A2(n8332), .ZN(n7760) );
  INV_X1 U9300 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9487) );
  OR2_X1 U9301 ( .A1(n8425), .A2(n9487), .ZN(n7759) );
  OAI22_X1 U9302 ( .A1(n9136), .A2(n9601), .B1(n8131), .B2(n9599), .ZN(n7763)
         );
  AOI211_X1 U9303 ( .C1(n9753), .C2(n7765), .A(n7764), .B(n7763), .ZN(n9757)
         );
  AOI21_X1 U9304 ( .B1(n9754), .B2(n7766), .A(n7842), .ZN(n9755) );
  INV_X1 U9305 ( .A(n9754), .ZN(n7826) );
  NOR2_X1 U9306 ( .A1(n7826), .A2(n9660), .ZN(n7769) );
  OAI22_X1 U9307 ( .A1(n9610), .A2(n7767), .B1(n9141), .B2(n10042), .ZN(n7768)
         );
  AOI211_X1 U9308 ( .C1(n9755), .C2(n9670), .A(n7769), .B(n7768), .ZN(n7772)
         );
  NAND2_X1 U9309 ( .A1(n9753), .A2(n7770), .ZN(n7771) );
  OAI211_X1 U9310 ( .C1(n9757), .C2(n4399), .A(n7772), .B(n7771), .ZN(P1_U3276) );
  NAND2_X1 U9311 ( .A1(n8287), .A2(n7773), .ZN(n7775) );
  OAI211_X1 U9312 ( .C1(n9791), .C2(n8288), .A(n7775), .B(n7774), .ZN(P1_U3326) );
  INV_X1 U9313 ( .A(n8287), .ZN(n7778) );
  OAI222_X1 U9314 ( .A1(n9002), .A2(n7778), .B1(n8044), .B2(n7777), .C1(n7776), 
        .C2(n8438), .ZN(P2_U3331) );
  NAND2_X1 U9315 ( .A1(n9875), .A2(n8307), .ZN(n7780) );
  NAND2_X1 U9316 ( .A1(n9452), .A2(n7480), .ZN(n7779) );
  NAND2_X1 U9317 ( .A1(n7780), .A2(n7779), .ZN(n7781) );
  XNOR2_X1 U9318 ( .A(n7781), .B(n8184), .ZN(n7786) );
  NOR2_X1 U9319 ( .A1(n7804), .A2(n8300), .ZN(n7782) );
  AOI21_X1 U9320 ( .B1(n9875), .B2(n8319), .A(n7782), .ZN(n7787) );
  NAND2_X1 U9321 ( .A1(n7786), .A2(n7787), .ZN(n7811) );
  INV_X1 U9322 ( .A(n7811), .ZN(n7791) );
  INV_X1 U9323 ( .A(n7783), .ZN(n7784) );
  NAND2_X1 U9324 ( .A1(n7785), .A2(n7784), .ZN(n7815) );
  INV_X1 U9325 ( .A(n7786), .ZN(n7789) );
  INV_X1 U9326 ( .A(n7787), .ZN(n7788) );
  NAND2_X1 U9327 ( .A1(n7789), .A2(n7788), .ZN(n7812) );
  AND2_X1 U9328 ( .A1(n7815), .A2(n7812), .ZN(n7790) );
  AND2_X1 U9329 ( .A1(n7792), .A2(n7793), .ZN(n7796) );
  INV_X1 U9330 ( .A(n7793), .ZN(n7795) );
  AND2_X1 U9331 ( .A1(n7813), .A2(n7811), .ZN(n7794) );
  NAND2_X1 U9332 ( .A1(n9759), .A2(n7480), .ZN(n7799) );
  NAND2_X1 U9333 ( .A1(n9868), .A2(n8324), .ZN(n7798) );
  NAND2_X1 U9334 ( .A1(n7799), .A2(n7798), .ZN(n7962) );
  NAND2_X1 U9335 ( .A1(n9759), .A2(n8307), .ZN(n7801) );
  NAND2_X1 U9336 ( .A1(n9868), .A2(n7480), .ZN(n7800) );
  NAND2_X1 U9337 ( .A1(n7801), .A2(n7800), .ZN(n7802) );
  XNOR2_X1 U9338 ( .A(n7802), .B(n8322), .ZN(n7963) );
  XOR2_X1 U9339 ( .A(n7962), .B(n7963), .Z(n7803) );
  XNOR2_X1 U9340 ( .A(n7964), .B(n7803), .ZN(n7810) );
  AND2_X1 U9341 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9955) );
  NOR2_X1 U9342 ( .A1(n9137), .A2(n7804), .ZN(n7805) );
  AOI211_X1 U9343 ( .C1(n9139), .C2(n9451), .A(n9955), .B(n7805), .ZN(n7806)
         );
  OAI21_X1 U9344 ( .B1(n9142), .B2(n7807), .A(n7806), .ZN(n7808) );
  AOI21_X1 U9345 ( .B1(n9759), .B2(n9144), .A(n7808), .ZN(n7809) );
  OAI21_X1 U9346 ( .B1(n7810), .B2(n9146), .A(n7809), .ZN(P1_U3232) );
  NAND2_X1 U9347 ( .A1(n7812), .A2(n7811), .ZN(n7818) );
  NAND2_X1 U9348 ( .A1(n7814), .A2(n7813), .ZN(n7816) );
  NAND2_X1 U9349 ( .A1(n7816), .A2(n7815), .ZN(n7817) );
  XOR2_X1 U9350 ( .A(n7818), .B(n7817), .Z(n7825) );
  NOR2_X1 U9351 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7819), .ZN(n9946) );
  NOR2_X1 U9352 ( .A1(n9137), .A2(n7820), .ZN(n7821) );
  AOI211_X1 U9353 ( .C1(n9139), .C2(n9868), .A(n9946), .B(n7821), .ZN(n7822)
         );
  OAI21_X1 U9354 ( .B1(n9142), .B2(n9871), .A(n7822), .ZN(n7823) );
  AOI21_X1 U9355 ( .B1(n9875), .B2(n9144), .A(n7823), .ZN(n7824) );
  OAI21_X1 U9356 ( .B1(n7825), .B2(n9146), .A(n7824), .ZN(P1_U3222) );
  NOR2_X1 U9357 ( .A1(n9754), .A2(n9450), .ZN(n7827) );
  OAI22_X1 U9358 ( .A1(n7828), .A2(n7827), .B1(n7826), .B2(n9060), .ZN(n8011)
         );
  NAND2_X1 U9359 ( .A1(n7829), .A2(n9151), .ZN(n7831) );
  AOI22_X1 U9360 ( .A1(n8150), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8149), .B2(
        n9996), .ZN(n7830) );
  NAND2_X1 U9361 ( .A1(n9750), .A2(n8131), .ZN(n9322) );
  NAND2_X1 U9362 ( .A1(n9323), .A2(n9322), .ZN(n9317) );
  XNOR2_X1 U9363 ( .A(n8011), .B(n9317), .ZN(n9752) );
  INV_X1 U9364 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7832) );
  AND2_X1 U9365 ( .A1(n7833), .A2(n7832), .ZN(n7834) );
  OR2_X1 U9366 ( .A1(n7834), .A2(n7914), .ZN(n9070) );
  OR2_X1 U9367 ( .A1(n5996), .A2(n7835), .ZN(n7837) );
  OR2_X1 U9368 ( .A1(n8333), .A2(n6538), .ZN(n7836) );
  AND2_X1 U9369 ( .A1(n7837), .A2(n7836), .ZN(n7839) );
  NAND2_X1 U9370 ( .A1(n6030), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7838) );
  OAI211_X1 U9371 ( .C1(n9070), .C2(n8332), .A(n7839), .B(n7838), .ZN(n9448)
         );
  INV_X1 U9372 ( .A(n9448), .ZN(n7907) );
  XNOR2_X1 U9373 ( .A(n7918), .B(n9317), .ZN(n7841) );
  OAI222_X1 U9374 ( .A1(n9599), .A2(n7907), .B1(n9601), .B2(n9060), .C1(n7841), 
        .C2(n9596), .ZN(n9748) );
  INV_X1 U9375 ( .A(n9750), .ZN(n9065) );
  INV_X1 U9376 ( .A(n7842), .ZN(n7844) );
  NAND2_X1 U9377 ( .A1(n7842), .A2(n9065), .ZN(n7911) );
  INV_X1 U9378 ( .A(n7911), .ZN(n7843) );
  AOI211_X1 U9379 ( .C1(n9750), .C2(n7844), .A(n10101), .B(n7843), .ZN(n9749)
         );
  NAND2_X1 U9380 ( .A1(n9749), .A2(n9884), .ZN(n7847) );
  INV_X1 U9381 ( .A(n7845), .ZN(n9062) );
  AOI22_X1 U9382 ( .A1(n4399), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9062), .B2(
        n9872), .ZN(n7846) );
  OAI211_X1 U9383 ( .C1(n9065), .C2(n9660), .A(n7847), .B(n7846), .ZN(n7848)
         );
  AOI21_X1 U9384 ( .B1(n9748), .B2(n9610), .A(n7848), .ZN(n7849) );
  OAI21_X1 U9385 ( .B1(n9752), .B2(n9672), .A(n7849), .ZN(P1_U3275) );
  XNOR2_X1 U9386 ( .A(n8967), .B(n8376), .ZN(n7892) );
  NOR2_X1 U9387 ( .A1(n7898), .A2(n5743), .ZN(n7890) );
  XNOR2_X1 U9388 ( .A(n7892), .B(n7890), .ZN(n7862) );
  INV_X1 U9389 ( .A(n7857), .ZN(n7852) );
  NOR3_X1 U9390 ( .A1(n7850), .A2(n7883), .A3(n8531), .ZN(n7851) );
  AOI21_X1 U9391 ( .B1(n7852), .B2(n8476), .A(n7851), .ZN(n7861) );
  INV_X1 U9392 ( .A(n7883), .ZN(n8557) );
  AOI22_X1 U9393 ( .A1(n8523), .A2(n8627), .B1(n8522), .B2(n8557), .ZN(n7854)
         );
  OAI211_X1 U9394 ( .C1(n7877), .C2(n8546), .A(n7854), .B(n7853), .ZN(n7859)
         );
  AND2_X1 U9395 ( .A1(n7862), .A2(n7855), .ZN(n7856) );
  NOR2_X1 U9396 ( .A1(n7894), .A2(n8553), .ZN(n7858) );
  AOI211_X1 U9397 ( .C1(n8967), .C2(n8551), .A(n7859), .B(n7858), .ZN(n7860)
         );
  OAI21_X1 U9398 ( .B1(n7862), .B2(n7861), .A(n7860), .ZN(P2_U3217) );
  INV_X1 U9399 ( .A(n7898), .ZN(n8556) );
  INV_X1 U9400 ( .A(n7952), .ZN(n8630) );
  XNOR2_X1 U9401 ( .A(n7863), .B(n7870), .ZN(n7864) );
  AOI222_X1 U9402 ( .A1(n8556), .A2(n8819), .B1(n8630), .B2(n8821), .C1(n8863), 
        .C2(n7864), .ZN(n8965) );
  AOI21_X1 U9403 ( .B1(n8962), .B2(n4957), .A(n8864), .ZN(n8963) );
  NOR2_X1 U9404 ( .A1(n7903), .A2(n8871), .ZN(n7867) );
  OAI22_X1 U9405 ( .A1(n8846), .A2(n7865), .B1(n7897), .B2(n8835), .ZN(n7866)
         );
  AOI211_X1 U9406 ( .C1(n8963), .C2(n8876), .A(n7867), .B(n7866), .ZN(n7873)
         );
  NAND2_X1 U9407 ( .A1(n7871), .A2(n7870), .ZN(n8629) );
  OAI21_X1 U9408 ( .B1(n7871), .B2(n7870), .A(n8629), .ZN(n8961) );
  NAND2_X1 U9409 ( .A1(n8961), .A2(n8738), .ZN(n7872) );
  OAI211_X1 U9410 ( .C1(n8965), .C2(n8878), .A(n7873), .B(n7872), .ZN(P2_U3281) );
  XNOR2_X1 U9411 ( .A(n7874), .B(n7881), .ZN(n8971) );
  INV_X1 U9412 ( .A(n4957), .ZN(n7875) );
  AOI21_X1 U9413 ( .B1(n8967), .B2(n7876), .A(n7875), .ZN(n8968) );
  INV_X1 U9414 ( .A(n8967), .ZN(n7880) );
  INV_X1 U9415 ( .A(n7877), .ZN(n7878) );
  AOI22_X1 U9416 ( .A1(n8878), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7878), .B2(
        n8868), .ZN(n7879) );
  OAI21_X1 U9417 ( .B1(n7880), .B2(n8871), .A(n7879), .ZN(n7888) );
  AOI21_X1 U9418 ( .B1(n7882), .B2(n7881), .A(n8759), .ZN(n7886) );
  OAI22_X1 U9419 ( .A1(n7883), .A2(n8853), .B1(n8854), .B2(n8851), .ZN(n7884)
         );
  AOI21_X1 U9420 ( .B1(n7886), .B2(n7885), .A(n7884), .ZN(n8970) );
  NOR2_X1 U9421 ( .A1(n8970), .A2(n8878), .ZN(n7887) );
  AOI211_X1 U9422 ( .C1(n8968), .C2(n8876), .A(n7888), .B(n7887), .ZN(n7889)
         );
  OAI21_X1 U9423 ( .B1(n8971), .B2(n8849), .A(n7889), .ZN(P2_U3282) );
  NAND2_X1 U9424 ( .A1(n8493), .A2(n8627), .ZN(n7896) );
  OR2_X1 U9425 ( .A1(n8854), .A2(n5743), .ZN(n7926) );
  NAND2_X1 U9426 ( .A1(n8476), .A2(n7926), .ZN(n7895) );
  INV_X1 U9427 ( .A(n7890), .ZN(n7891) );
  NAND2_X1 U9428 ( .A1(n7892), .A2(n7891), .ZN(n7893) );
  XNOR2_X1 U9429 ( .A(n8962), .B(n8365), .ZN(n7928) );
  MUX2_X1 U9430 ( .A(n7896), .B(n7895), .S(n7927), .Z(n7902) );
  NOR2_X1 U9431 ( .A1(n8546), .A2(n7897), .ZN(n7900) );
  OAI22_X1 U9432 ( .A1(n7952), .A2(n8547), .B1(n8548), .B2(n7898), .ZN(n7899)
         );
  AOI211_X1 U9433 ( .C1(P2_REG3_REG_15__SCAN_IN), .C2(n7777), .A(n7900), .B(
        n7899), .ZN(n7901) );
  OAI211_X1 U9434 ( .C1(n7903), .C2(n8541), .A(n7902), .B(n7901), .ZN(P2_U3243) );
  NAND2_X1 U9435 ( .A1(n7904), .A2(n9151), .ZN(n7906) );
  AOI22_X1 U9436 ( .A1(n10008), .A2(n8149), .B1(n8150), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n7905) );
  OR2_X1 U9437 ( .A1(n9745), .A2(n7907), .ZN(n8415) );
  NAND2_X1 U9438 ( .A1(n9745), .A2(n7907), .ZN(n8414) );
  NAND2_X1 U9439 ( .A1(n8011), .A2(n9317), .ZN(n7908) );
  INV_X1 U9440 ( .A(n8131), .ZN(n9449) );
  NAND2_X1 U9441 ( .A1(n9750), .A2(n9449), .ZN(n8013) );
  NAND2_X1 U9442 ( .A1(n7908), .A2(n8013), .ZN(n7909) );
  XOR2_X1 U9443 ( .A(n9325), .B(n7909), .Z(n9747) );
  INV_X1 U9444 ( .A(n8034), .ZN(n7910) );
  AOI211_X1 U9445 ( .C1(n9745), .C2(n7911), .A(n10101), .B(n7910), .ZN(n9744)
         );
  INV_X1 U9446 ( .A(n9745), .ZN(n9076) );
  NOR2_X1 U9447 ( .A1(n9076), .A2(n9660), .ZN(n7913) );
  OAI22_X1 U9448 ( .A1(n9610), .A2(n6538), .B1(n9070), .B2(n10042), .ZN(n7912)
         );
  AOI211_X1 U9449 ( .C1(n9744), .C2(n9884), .A(n7913), .B(n7912), .ZN(n7922)
         );
  NOR2_X1 U9450 ( .A1(n7914), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7915) );
  OR2_X1 U9451 ( .A1(n8027), .A2(n7915), .ZN(n9113) );
  AOI22_X1 U9452 ( .A1(n5995), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n8421), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n7917) );
  INV_X1 U9453 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9492) );
  OR2_X1 U9454 ( .A1(n8425), .A2(n9492), .ZN(n7916) );
  OAI211_X1 U9455 ( .C1(n9113), .C2(n8332), .A(n7917), .B(n7916), .ZN(n9665)
         );
  INV_X1 U9456 ( .A(n9665), .ZN(n9071) );
  XNOR2_X1 U9457 ( .A(n8416), .B(n9325), .ZN(n7920) );
  OAI222_X1 U9458 ( .A1(n9599), .A2(n9071), .B1(n9601), .B2(n8131), .C1(n9596), 
        .C2(n7920), .ZN(n9743) );
  NAND2_X1 U9459 ( .A1(n9743), .A2(n9610), .ZN(n7921) );
  OAI211_X1 U9460 ( .C1(n9747), .C2(n9672), .A(n7922), .B(n7921), .ZN(P1_U3274) );
  INV_X1 U9461 ( .A(n8407), .ZN(n8350) );
  OAI222_X1 U9462 ( .A1(P1_U3084), .A2(n7923), .B1(n7925), .B2(n8350), .C1(
        n8408), .C2(n9791), .ZN(P1_U3324) );
  INV_X1 U9463 ( .A(n8303), .ZN(n8107) );
  OAI222_X1 U9464 ( .A1(P1_U3084), .A2(n6102), .B1(n7925), .B2(n8107), .C1(
        n8304), .C2(n9791), .ZN(P1_U3325) );
  NAND2_X1 U9465 ( .A1(n7927), .A2(n7926), .ZN(n7932) );
  INV_X1 U9466 ( .A(n7928), .ZN(n7929) );
  NAND2_X1 U9467 ( .A1(n7930), .A2(n7929), .ZN(n7931) );
  NAND2_X1 U9468 ( .A1(n7932), .A2(n7931), .ZN(n7938) );
  XNOR2_X1 U9469 ( .A(n8956), .B(n8376), .ZN(n7941) );
  NOR2_X1 U9470 ( .A1(n7952), .A2(n5743), .ZN(n7939) );
  XNOR2_X1 U9471 ( .A(n7941), .B(n7939), .ZN(n7937) );
  XOR2_X1 U9472 ( .A(n7938), .B(n7937), .Z(n7936) );
  AOI22_X1 U9473 ( .A1(n8523), .A2(n8820), .B1(n8522), .B2(n8627), .ZN(n7933)
         );
  NAND2_X1 U9474 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(n7777), .ZN(n8586) );
  OAI211_X1 U9475 ( .C1(n8867), .C2(n8546), .A(n7933), .B(n8586), .ZN(n7934)
         );
  AOI21_X1 U9476 ( .B1(n8956), .B2(n8551), .A(n7934), .ZN(n7935) );
  OAI21_X1 U9477 ( .B1(n7936), .B2(n8553), .A(n7935), .ZN(P2_U3228) );
  INV_X1 U9478 ( .A(n7939), .ZN(n7940) );
  NAND2_X1 U9479 ( .A1(n7941), .A2(n7940), .ZN(n7942) );
  XNOR2_X1 U9480 ( .A(n8953), .B(n8365), .ZN(n7944) );
  NOR2_X1 U9481 ( .A1(n8852), .A2(n5743), .ZN(n7945) );
  NAND2_X1 U9482 ( .A1(n7944), .A2(n7945), .ZN(n8077) );
  INV_X1 U9483 ( .A(n7944), .ZN(n8532) );
  INV_X1 U9484 ( .A(n7945), .ZN(n7946) );
  NAND2_X1 U9485 ( .A1(n8532), .A2(n7946), .ZN(n7947) );
  NAND2_X1 U9486 ( .A1(n8077), .A2(n7947), .ZN(n7949) );
  AOI21_X1 U9487 ( .B1(n7948), .B2(n7949), .A(n8553), .ZN(n7951) );
  NAND2_X1 U9488 ( .A1(n7951), .A2(n8530), .ZN(n7959) );
  INV_X1 U9489 ( .A(n8836), .ZN(n7957) );
  OR2_X1 U9490 ( .A1(n7952), .A2(n8853), .ZN(n7954) );
  NAND2_X1 U9491 ( .A1(n8805), .A2(n8821), .ZN(n7953) );
  AND2_X1 U9492 ( .A1(n7954), .A2(n7953), .ZN(n8844) );
  OAI22_X1 U9493 ( .A1(n8502), .A2(n8844), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7955), .ZN(n7956) );
  AOI21_X1 U9494 ( .B1(n7957), .B2(n8538), .A(n7956), .ZN(n7958) );
  OAI211_X1 U9495 ( .C1(n8834), .C2(n8541), .A(n7959), .B(n7958), .ZN(P2_U3230) );
  OAI222_X1 U9496 ( .A1(n8110), .A2(n7961), .B1(n5741), .B2(n7777), .C1(n7960), 
        .C2(n8438), .ZN(P2_U3338) );
  NAND2_X1 U9497 ( .A1(n7964), .A2(n7963), .ZN(n7965) );
  NAND2_X1 U9498 ( .A1(n7979), .A2(n8307), .ZN(n7968) );
  NAND2_X1 U9499 ( .A1(n9451), .A2(n8319), .ZN(n7967) );
  NAND2_X1 U9500 ( .A1(n7968), .A2(n7967), .ZN(n7969) );
  XNOR2_X1 U9501 ( .A(n7969), .B(n8184), .ZN(n8123) );
  NAND2_X1 U9502 ( .A1(n7979), .A2(n8319), .ZN(n7971) );
  NAND2_X1 U9503 ( .A1(n9451), .A2(n8324), .ZN(n7970) );
  NAND2_X1 U9504 ( .A1(n7971), .A2(n7970), .ZN(n8115) );
  XNOR2_X1 U9505 ( .A(n8123), .B(n8115), .ZN(n7972) );
  XNOR2_X1 U9506 ( .A(n8116), .B(n7972), .ZN(n7981) );
  NOR2_X1 U9507 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7973), .ZN(n9973) );
  NOR2_X1 U9508 ( .A1(n9137), .A2(n7974), .ZN(n7975) );
  AOI211_X1 U9509 ( .C1(n9139), .C2(n9450), .A(n9973), .B(n7975), .ZN(n7976)
         );
  OAI21_X1 U9510 ( .B1(n9142), .B2(n7977), .A(n7976), .ZN(n7978) );
  AOI21_X1 U9511 ( .B1(n7979), .B2(n9144), .A(n7978), .ZN(n7980) );
  OAI21_X1 U9512 ( .B1(n7981), .B2(n9146), .A(n7980), .ZN(P1_U3213) );
  NOR2_X1 U9513 ( .A1(n7597), .A2(n7982), .ZN(n7984) );
  OR2_X1 U9514 ( .A1(n7984), .A2(n7983), .ZN(n7989) );
  NAND2_X1 U9515 ( .A1(n7986), .A2(n7985), .ZN(n7987) );
  NAND2_X1 U9516 ( .A1(n7987), .A2(n7990), .ZN(n7988) );
  NAND2_X1 U9517 ( .A1(n7989), .A2(n7988), .ZN(n10184) );
  XNOR2_X1 U9518 ( .A(n7991), .B(n7990), .ZN(n7995) );
  OAI22_X1 U9519 ( .A1(n7993), .A2(n8853), .B1(n7992), .B2(n8851), .ZN(n7994)
         );
  AOI21_X1 U9520 ( .B1(n7995), .B2(n8863), .A(n7994), .ZN(n7996) );
  OAI21_X1 U9521 ( .B1(n10184), .B2(n8859), .A(n7996), .ZN(n10189) );
  NAND2_X1 U9522 ( .A1(n10189), .A2(n8846), .ZN(n8005) );
  OAI22_X1 U9523 ( .A1(n8846), .A2(n7998), .B1(n7997), .B2(n8835), .ZN(n8003)
         );
  NAND2_X1 U9524 ( .A1(n7999), .A2(n10185), .ZN(n8000) );
  NAND2_X1 U9525 ( .A1(n8001), .A2(n8000), .ZN(n10188) );
  NOR2_X1 U9526 ( .A1(n10188), .A2(n8656), .ZN(n8002) );
  AOI211_X1 U9527 ( .C1(n8691), .C2(n10185), .A(n8003), .B(n8002), .ZN(n8004)
         );
  OAI211_X1 U9528 ( .C1(n10184), .C2(n8873), .A(n8005), .B(n8004), .ZN(
        P2_U3286) );
  OR2_X1 U9529 ( .A1(n9745), .A2(n9448), .ZN(n8012) );
  AND2_X1 U9530 ( .A1(n9317), .A2(n8012), .ZN(n8019) );
  NAND2_X1 U9531 ( .A1(n8006), .A2(n9151), .ZN(n8008) );
  AOI22_X1 U9532 ( .A1(n10027), .A2(n8149), .B1(n8150), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n8007) );
  OR2_X1 U9533 ( .A1(n9105), .A2(n9071), .ZN(n9330) );
  NAND2_X1 U9534 ( .A1(n9105), .A2(n9071), .ZN(n9202) );
  INV_X1 U9535 ( .A(n9181), .ZN(n8009) );
  AND2_X1 U9536 ( .A1(n8019), .A2(n8009), .ZN(n8010) );
  NAND2_X1 U9537 ( .A1(n8011), .A2(n8010), .ZN(n8018) );
  INV_X1 U9538 ( .A(n8012), .ZN(n8016) );
  NAND2_X1 U9539 ( .A1(n9745), .A2(n9448), .ZN(n8014) );
  AND2_X1 U9540 ( .A1(n8014), .A2(n8013), .ZN(n8015) );
  NAND2_X1 U9541 ( .A1(n8011), .A2(n8019), .ZN(n8021) );
  AND2_X1 U9542 ( .A1(n8021), .A2(n8020), .ZN(n8022) );
  AND2_X1 U9543 ( .A1(n8022), .A2(n9181), .ZN(n8023) );
  OR2_X1 U9544 ( .A1(n8393), .A2(n8023), .ZN(n9742) );
  INV_X1 U9545 ( .A(n8415), .ZN(n8024) );
  AOI21_X1 U9546 ( .B1(n8416), .B2(n8414), .A(n8024), .ZN(n8025) );
  XNOR2_X1 U9547 ( .A(n8025), .B(n9181), .ZN(n8026) );
  NAND2_X1 U9548 ( .A1(n8026), .A2(n9870), .ZN(n8032) );
  OR2_X1 U9549 ( .A1(n8027), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8028) );
  NAND2_X1 U9550 ( .A1(n8173), .A2(n8028), .ZN(n9657) );
  AOI22_X1 U9551 ( .A1(n5995), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n8421), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n8030) );
  OR2_X1 U9552 ( .A1(n8425), .A2(n9493), .ZN(n8029) );
  OAI211_X1 U9553 ( .C1(n9657), .C2(n8332), .A(n8030), .B(n8029), .ZN(n9648)
         );
  AOI22_X1 U9554 ( .A1(n9648), .A2(n9867), .B1(n9865), .B2(n9448), .ZN(n8031)
         );
  NAND2_X1 U9555 ( .A1(n8032), .A2(n8031), .ZN(n9740) );
  NAND2_X1 U9556 ( .A1(n8034), .A2(n9105), .ZN(n8033) );
  NAND2_X1 U9557 ( .A1(n8033), .A2(n9881), .ZN(n8035) );
  OR2_X1 U9558 ( .A1(n8035), .A2(n9654), .ZN(n9737) );
  INV_X1 U9559 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9473) );
  OAI22_X1 U9560 ( .A1(n9610), .A2(n9473), .B1(n9113), .B2(n10042), .ZN(n8036)
         );
  AOI21_X1 U9561 ( .B1(n9105), .B2(n9874), .A(n8036), .ZN(n8037) );
  OAI21_X1 U9562 ( .B1(n9737), .B2(n8038), .A(n8037), .ZN(n8039) );
  AOI21_X1 U9563 ( .B1(n9740), .B2(n9610), .A(n8039), .ZN(n8040) );
  OAI21_X1 U9564 ( .B1(n9742), .B2(n9672), .A(n8040), .ZN(P1_U3273) );
  INV_X1 U9565 ( .A(n8956), .ZN(n8872) );
  INV_X1 U9566 ( .A(n8936), .ZN(n8789) );
  NAND2_X1 U9567 ( .A1(n8786), .A2(n8773), .ZN(n8751) );
  INV_X1 U9568 ( .A(n8910), .ZN(n8712) );
  NOR2_X1 U9569 ( .A1(n8846), .A2(n8043), .ZN(n8048) );
  INV_X1 U9570 ( .A(n8044), .ZN(n8045) );
  AND2_X1 U9571 ( .A1(n8045), .A2(P2_B_REG_SCAN_IN), .ZN(n8046) );
  NOR2_X1 U9572 ( .A1(n8851), .A2(n8046), .ZN(n8651) );
  NAND2_X1 U9573 ( .A1(n8047), .A2(n8651), .ZN(n8884) );
  NOR2_X1 U9574 ( .A1(n8878), .A2(n8884), .ZN(n8624) );
  AOI211_X1 U9575 ( .C1(n8879), .C2(n8691), .A(n8048), .B(n8624), .ZN(n8049)
         );
  OAI21_X1 U9576 ( .B1(n8881), .B2(n8656), .A(n8049), .ZN(P2_U3265) );
  NAND2_X1 U9577 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8594), .ZN(n8050) );
  OAI21_X1 U9578 ( .B1(n8594), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8050), .ZN(
        n8590) );
  OAI22_X1 U9579 ( .A1(n8053), .A2(n8052), .B1(n8051), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n8591) );
  NOR2_X1 U9580 ( .A1(n8590), .A2(n8591), .ZN(n8589) );
  AOI21_X1 U9581 ( .B1(n8594), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8589), .ZN(
        n8599) );
  NAND2_X1 U9582 ( .A1(n8055), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8054) );
  OAI21_X1 U9583 ( .B1(n8055), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8054), .ZN(
        n8598) );
  NOR2_X1 U9584 ( .A1(n8599), .A2(n8598), .ZN(n8597) );
  INV_X1 U9585 ( .A(n8059), .ZN(n8621) );
  NAND2_X1 U9586 ( .A1(n8056), .A2(n8621), .ZN(n8057) );
  XNOR2_X1 U9587 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8058), .ZN(n8073) );
  OR2_X1 U9588 ( .A1(n8059), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8069) );
  NAND2_X1 U9589 ( .A1(n8059), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8060) );
  NAND2_X1 U9590 ( .A1(n8069), .A2(n8060), .ZN(n8610) );
  XNOR2_X1 U9591 ( .A(n8606), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8603) );
  XNOR2_X1 U9592 ( .A(n8594), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8584) );
  INV_X1 U9593 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8064) );
  INV_X1 U9594 ( .A(n8061), .ZN(n8062) );
  OAI22_X1 U9595 ( .A1(n8065), .A2(n8064), .B1(n8063), .B2(n8062), .ZN(n8585)
         );
  NOR2_X1 U9596 ( .A1(n8584), .A2(n8585), .ZN(n8583) );
  AOI21_X1 U9597 ( .B1(n8067), .B2(n8066), .A(n8583), .ZN(n8602) );
  NAND2_X1 U9598 ( .A1(n8603), .A2(n8602), .ZN(n8601) );
  OAI21_X1 U9599 ( .B1(n8068), .B2(n8606), .A(n8601), .ZN(n8609) );
  OR2_X1 U9600 ( .A1(n8610), .A2(n8609), .ZN(n8613) );
  NAND2_X1 U9601 ( .A1(n8613), .A2(n8069), .ZN(n8071) );
  XNOR2_X1 U9602 ( .A(n8071), .B(n8070), .ZN(n8074) );
  INV_X1 U9603 ( .A(n8074), .ZN(n8072) );
  AOI22_X1 U9604 ( .A1(n8073), .A2(n10118), .B1(n8072), .B2(n10119), .ZN(n8075) );
  NAND2_X1 U9605 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8076) );
  XNOR2_X1 U9606 ( .A(n8946), .B(n8365), .ZN(n8078) );
  AND2_X1 U9607 ( .A1(n8805), .A2(n8367), .ZN(n8079) );
  NAND2_X1 U9608 ( .A1(n8078), .A2(n8079), .ZN(n8082) );
  INV_X1 U9609 ( .A(n8078), .ZN(n8461) );
  INV_X1 U9610 ( .A(n8079), .ZN(n8080) );
  NAND2_X1 U9611 ( .A1(n8461), .A2(n8080), .ZN(n8081) );
  XNOR2_X1 U9612 ( .A(n8942), .B(n8365), .ZN(n8084) );
  NAND2_X1 U9613 ( .A1(n8822), .A2(n8367), .ZN(n8085) );
  XNOR2_X1 U9614 ( .A(n8084), .B(n8085), .ZN(n8462) );
  AND2_X1 U9615 ( .A1(n8462), .A2(n8082), .ZN(n8083) );
  NAND2_X1 U9616 ( .A1(n8459), .A2(n8083), .ZN(n8460) );
  INV_X1 U9617 ( .A(n8084), .ZN(n8086) );
  NAND2_X1 U9618 ( .A1(n8086), .A2(n8085), .ZN(n8087) );
  XNOR2_X1 U9619 ( .A(n8936), .B(n8365), .ZN(n8088) );
  NOR2_X1 U9620 ( .A1(n8487), .A2(n5743), .ZN(n8089) );
  NAND2_X1 U9621 ( .A1(n8088), .A2(n8089), .ZN(n8093) );
  INV_X1 U9622 ( .A(n8088), .ZN(n8482) );
  INV_X1 U9623 ( .A(n8089), .ZN(n8090) );
  NAND2_X1 U9624 ( .A1(n8482), .A2(n8090), .ZN(n8091) );
  NAND2_X1 U9625 ( .A1(n8093), .A2(n8091), .ZN(n8520) );
  XNOR2_X1 U9626 ( .A(n8773), .B(n8365), .ZN(n8095) );
  NOR2_X1 U9627 ( .A1(n8762), .A2(n5743), .ZN(n8096) );
  XNOR2_X1 U9628 ( .A(n8095), .B(n8096), .ZN(n8480) );
  INV_X1 U9629 ( .A(n8095), .ZN(n8097) );
  NAND2_X1 U9630 ( .A1(n8097), .A2(n8096), .ZN(n8098) );
  NAND2_X1 U9631 ( .A1(n8483), .A2(n8098), .ZN(n8353) );
  XNOR2_X1 U9632 ( .A(n8926), .B(n8376), .ZN(n8351) );
  XNOR2_X1 U9633 ( .A(n8353), .B(n8351), .ZN(n8103) );
  INV_X1 U9634 ( .A(n8641), .ZN(n8780) );
  NAND2_X1 U9635 ( .A1(n8780), .A2(n8367), .ZN(n8099) );
  NAND2_X1 U9636 ( .A1(n8103), .A2(n8099), .ZN(n8355) );
  OAI22_X1 U9637 ( .A1(n8546), .A2(n8752), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8100), .ZN(n8102) );
  OAI22_X1 U9638 ( .A1(n8762), .A2(n8548), .B1(n8547), .B2(n8763), .ZN(n8101)
         );
  AOI211_X1 U9639 ( .C1(n8926), .C2(n8551), .A(n8102), .B(n8101), .ZN(n8105)
         );
  OR3_X1 U9640 ( .A1(n8103), .A2(n8641), .A3(n8531), .ZN(n8104) );
  OAI211_X1 U9641 ( .C1(n8355), .C2(n8553), .A(n8105), .B(n8104), .ZN(P2_U3237) );
  OAI222_X1 U9642 ( .A1(n9002), .A2(n8107), .B1(n5763), .B2(P2_U3152), .C1(
        n8106), .C2(n8438), .ZN(P2_U3330) );
  OAI222_X1 U9643 ( .A1(n8438), .A2(n8111), .B1(n8110), .B2(n8109), .C1(
        P2_U3152), .C2(n8108), .ZN(P2_U3336) );
  INV_X1 U9644 ( .A(n8116), .ZN(n8113) );
  INV_X1 U9645 ( .A(n8115), .ZN(n8112) );
  INV_X1 U9646 ( .A(n8123), .ZN(n8114) );
  NAND2_X1 U9647 ( .A1(n9754), .A2(n8307), .ZN(n8118) );
  NAND2_X1 U9648 ( .A1(n9450), .A2(n7480), .ZN(n8117) );
  NAND2_X1 U9649 ( .A1(n8118), .A2(n8117), .ZN(n8119) );
  XNOR2_X1 U9650 ( .A(n8119), .B(n8322), .ZN(n8125) );
  INV_X1 U9651 ( .A(n8125), .ZN(n8120) );
  NAND2_X1 U9652 ( .A1(n9754), .A2(n8319), .ZN(n8122) );
  NAND2_X1 U9653 ( .A1(n9450), .A2(n8324), .ZN(n8121) );
  NAND2_X1 U9654 ( .A1(n8122), .A2(n8121), .ZN(n9134) );
  NAND2_X1 U9655 ( .A1(n8124), .A2(n8123), .ZN(n8127) );
  NAND3_X1 U9656 ( .A1(n8127), .A2(n8126), .A3(n8125), .ZN(n9053) );
  NAND2_X1 U9657 ( .A1(n9750), .A2(n8307), .ZN(n8129) );
  NAND2_X1 U9658 ( .A1(n9449), .A2(n7480), .ZN(n8128) );
  NAND2_X1 U9659 ( .A1(n8129), .A2(n8128), .ZN(n8130) );
  XNOR2_X1 U9660 ( .A(n8130), .B(n8184), .ZN(n8133) );
  NOR2_X1 U9661 ( .A1(n8131), .A2(n8300), .ZN(n8132) );
  AOI21_X1 U9662 ( .B1(n9750), .B2(n7480), .A(n8132), .ZN(n8134) );
  NAND2_X1 U9663 ( .A1(n8133), .A2(n8134), .ZN(n8139) );
  INV_X1 U9664 ( .A(n8133), .ZN(n8136) );
  INV_X1 U9665 ( .A(n8134), .ZN(n8135) );
  NAND2_X1 U9666 ( .A1(n8136), .A2(n8135), .ZN(n8137) );
  AND2_X1 U9667 ( .A1(n8139), .A2(n8137), .ZN(n9054) );
  AND2_X1 U9668 ( .A1(n9053), .A2(n9054), .ZN(n8138) );
  NAND2_X1 U9669 ( .A1(n9745), .A2(n8307), .ZN(n8141) );
  NAND2_X1 U9670 ( .A1(n9448), .A2(n8319), .ZN(n8140) );
  NAND2_X1 U9671 ( .A1(n8141), .A2(n8140), .ZN(n8142) );
  XNOR2_X1 U9672 ( .A(n8142), .B(n8322), .ZN(n8144) );
  AND2_X1 U9673 ( .A1(n9448), .A2(n8324), .ZN(n8143) );
  AOI21_X1 U9674 ( .B1(n9745), .B2(n8319), .A(n8143), .ZN(n8145) );
  XNOR2_X1 U9675 ( .A(n8144), .B(n8145), .ZN(n9068) );
  INV_X1 U9676 ( .A(n8144), .ZN(n8146) );
  NAND2_X1 U9677 ( .A1(n8146), .A2(n8145), .ZN(n8147) );
  NAND2_X1 U9678 ( .A1(n8148), .A2(n9151), .ZN(n8152) );
  AOI22_X1 U9679 ( .A1(n8150), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10039), 
        .B2(n8149), .ZN(n8151) );
  NAND2_X1 U9680 ( .A1(n9732), .A2(n8307), .ZN(n8154) );
  NAND2_X1 U9681 ( .A1(n9648), .A2(n8319), .ZN(n8153) );
  NAND2_X1 U9682 ( .A1(n8154), .A2(n8153), .ZN(n8155) );
  XNOR2_X1 U9683 ( .A(n8155), .B(n8322), .ZN(n9029) );
  NAND2_X1 U9684 ( .A1(n9732), .A2(n8319), .ZN(n8157) );
  NAND2_X1 U9685 ( .A1(n9648), .A2(n8324), .ZN(n8156) );
  NAND2_X1 U9686 ( .A1(n8157), .A2(n8156), .ZN(n9028) );
  NAND2_X1 U9687 ( .A1(n9105), .A2(n7480), .ZN(n8159) );
  NAND2_X1 U9688 ( .A1(n9665), .A2(n8324), .ZN(n8158) );
  INV_X1 U9689 ( .A(n9108), .ZN(n8163) );
  NAND2_X1 U9690 ( .A1(n9105), .A2(n8307), .ZN(n8161) );
  NAND2_X1 U9691 ( .A1(n9665), .A2(n8319), .ZN(n8160) );
  NAND2_X1 U9692 ( .A1(n8161), .A2(n8160), .ZN(n8162) );
  XNOR2_X1 U9693 ( .A(n8162), .B(n8184), .ZN(n9027) );
  INV_X1 U9694 ( .A(n9027), .ZN(n9025) );
  AOI22_X1 U9695 ( .A1(n9029), .A2(n9028), .B1(n8163), .B2(n9025), .ZN(n8167)
         );
  NAND2_X1 U9696 ( .A1(n9027), .A2(n9108), .ZN(n8165) );
  AOI21_X1 U9697 ( .B1(n9028), .B2(n8165), .A(n9029), .ZN(n8164) );
  INV_X1 U9698 ( .A(n8164), .ZN(n8166) );
  NAND2_X1 U9699 ( .A1(n8168), .A2(n9151), .ZN(n8171) );
  OR2_X1 U9700 ( .A1(n9154), .A2(n8169), .ZN(n8170) );
  NAND2_X1 U9701 ( .A1(n9728), .A2(n8307), .ZN(n8183) );
  INV_X1 U9702 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8172) );
  NAND2_X1 U9703 ( .A1(n8173), .A2(n8172), .ZN(n8174) );
  AND2_X1 U9704 ( .A1(n8193), .A2(n8174), .ZN(n9642) );
  INV_X1 U9705 ( .A(n8332), .ZN(n8175) );
  NAND2_X1 U9706 ( .A1(n9642), .A2(n8175), .ZN(n8181) );
  NAND2_X1 U9707 ( .A1(n5995), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8177) );
  NAND2_X1 U9708 ( .A1(n8421), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8176) );
  OAI211_X1 U9709 ( .C1(n8425), .C2(n8178), .A(n8177), .B(n8176), .ZN(n8179)
         );
  INV_X1 U9710 ( .A(n8179), .ZN(n8180) );
  NAND2_X1 U9711 ( .A1(n8181), .A2(n8180), .ZN(n9666) );
  NAND2_X1 U9712 ( .A1(n9666), .A2(n8319), .ZN(n8182) );
  NAND2_X1 U9713 ( .A1(n8183), .A2(n8182), .ZN(n8185) );
  XNOR2_X1 U9714 ( .A(n8185), .B(n8184), .ZN(n8188) );
  AND2_X1 U9715 ( .A1(n9666), .A2(n8324), .ZN(n8186) );
  AOI21_X1 U9716 ( .B1(n9728), .B2(n8319), .A(n8186), .ZN(n8187) );
  NOR2_X1 U9717 ( .A1(n8188), .A2(n8187), .ZN(n9086) );
  NAND2_X1 U9718 ( .A1(n8189), .A2(n9151), .ZN(n8192) );
  OR2_X1 U9719 ( .A1(n9154), .A2(n8190), .ZN(n8191) );
  INV_X1 U9720 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9039) );
  NAND2_X1 U9721 ( .A1(n8193), .A2(n9039), .ZN(n8195) );
  INV_X1 U9722 ( .A(n8213), .ZN(n8194) );
  NAND2_X1 U9723 ( .A1(n8195), .A2(n8194), .ZN(n9627) );
  OR2_X1 U9724 ( .A1(n9627), .A2(n8332), .ZN(n8201) );
  NAND2_X1 U9725 ( .A1(n5995), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U9726 ( .A1(n6030), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8196) );
  OAI211_X1 U9727 ( .C1(n8198), .C2(n5996), .A(n8197), .B(n8196), .ZN(n8199)
         );
  INV_X1 U9728 ( .A(n8199), .ZN(n8200) );
  AOI22_X1 U9729 ( .A1(n9723), .A2(n7480), .B1(n8324), .B2(n9649), .ZN(n8205)
         );
  NAND2_X1 U9730 ( .A1(n9723), .A2(n8307), .ZN(n8203) );
  NAND2_X1 U9731 ( .A1(n9649), .A2(n8319), .ZN(n8202) );
  NAND2_X1 U9732 ( .A1(n8203), .A2(n8202), .ZN(n8204) );
  XNOR2_X1 U9733 ( .A(n8204), .B(n8322), .ZN(n8207) );
  XOR2_X1 U9734 ( .A(n8205), .B(n8207), .Z(n9038) );
  INV_X1 U9735 ( .A(n8205), .ZN(n8206) );
  NAND2_X1 U9736 ( .A1(n8208), .A2(n9151), .ZN(n8211) );
  OR2_X1 U9737 ( .A1(n9154), .A2(n8209), .ZN(n8210) );
  NAND2_X1 U9738 ( .A1(n8421), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8218) );
  INV_X1 U9739 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n8212) );
  OR2_X1 U9740 ( .A1(n8333), .A2(n8212), .ZN(n8217) );
  NAND2_X1 U9741 ( .A1(n8213), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8228) );
  OAI21_X1 U9742 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n8213), .A(n8228), .ZN(
        n9614) );
  OR2_X1 U9743 ( .A1(n8332), .A2(n9614), .ZN(n8216) );
  OR2_X1 U9744 ( .A1(n8425), .A2(n8214), .ZN(n8215) );
  INV_X1 U9745 ( .A(n9600), .ZN(n9634) );
  AOI22_X1 U9746 ( .A1(n9717), .A2(n8319), .B1(n8324), .B2(n9634), .ZN(n8220)
         );
  NAND2_X1 U9747 ( .A1(n8221), .A2(n8220), .ZN(n9096) );
  OAI22_X1 U9748 ( .A1(n9617), .A2(n8298), .B1(n9600), .B2(n8297), .ZN(n8219)
         );
  XNOR2_X1 U9749 ( .A(n8219), .B(n8322), .ZN(n9098) );
  AOI21_X1 U9750 ( .B1(n9096), .B2(n9098), .A(n9095), .ZN(n8236) );
  NAND2_X1 U9751 ( .A1(n8222), .A2(n9151), .ZN(n8225) );
  OR2_X1 U9752 ( .A1(n9154), .A2(n8223), .ZN(n8224) );
  NAND2_X1 U9753 ( .A1(n6030), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8233) );
  OR2_X1 U9754 ( .A1(n5996), .A2(n8226), .ZN(n8232) );
  OR2_X1 U9755 ( .A1(n8333), .A2(n8227), .ZN(n8231) );
  OAI21_X1 U9756 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n8229), .A(n8243), .ZN(
        n9604) );
  OR2_X1 U9757 ( .A1(n8332), .A2(n9604), .ZN(n8230) );
  OAI22_X1 U9758 ( .A1(n9608), .A2(n8298), .B1(n9581), .B2(n8297), .ZN(n8234)
         );
  XOR2_X1 U9759 ( .A(n8322), .B(n8234), .Z(n8235) );
  OAI22_X1 U9760 ( .A1(n9608), .A2(n8297), .B1(n9581), .B2(n8300), .ZN(n9017)
         );
  NAND2_X1 U9761 ( .A1(n8237), .A2(n9151), .ZN(n8240) );
  OR2_X1 U9762 ( .A1(n9154), .A2(n8238), .ZN(n8239) );
  NAND2_X1 U9763 ( .A1(n8421), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8248) );
  OR2_X1 U9764 ( .A1(n8333), .A2(n8241), .ZN(n8247) );
  OR2_X1 U9765 ( .A1(n8425), .A2(n8242), .ZN(n8246) );
  OAI21_X1 U9766 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n8244), .A(n8258), .ZN(
        n9586) );
  OR2_X1 U9767 ( .A1(n8332), .A2(n9586), .ZN(n8245) );
  OAI22_X1 U9768 ( .A1(n9590), .A2(n8298), .B1(n9598), .B2(n8297), .ZN(n8249)
         );
  XNOR2_X1 U9769 ( .A(n8249), .B(n8322), .ZN(n8250) );
  AOI22_X1 U9770 ( .A1(n9709), .A2(n7480), .B1(n8324), .B2(n9567), .ZN(n8251)
         );
  XNOR2_X1 U9771 ( .A(n8250), .B(n8251), .ZN(n9078) );
  INV_X1 U9772 ( .A(n8250), .ZN(n8252) );
  NAND2_X1 U9773 ( .A1(n8254), .A2(n9151), .ZN(n8257) );
  OR2_X1 U9774 ( .A1(n9154), .A2(n8255), .ZN(n8256) );
  NAND2_X1 U9775 ( .A1(n8421), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8264) );
  OR2_X1 U9776 ( .A1(n8333), .A2(n6399), .ZN(n8263) );
  OAI21_X1 U9777 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n8259), .A(n8274), .ZN(
        n9561) );
  OR2_X1 U9778 ( .A1(n8332), .A2(n9561), .ZN(n8262) );
  INV_X1 U9779 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n8260) );
  OR2_X1 U9780 ( .A1(n8425), .A2(n8260), .ZN(n8261) );
  OAI22_X1 U9781 ( .A1(n9564), .A2(n8298), .B1(n9582), .B2(n8297), .ZN(n8265)
         );
  XNOR2_X1 U9782 ( .A(n8265), .B(n8322), .ZN(n8267) );
  NOR2_X1 U9783 ( .A1(n9582), .A2(n8300), .ZN(n8266) );
  AOI21_X1 U9784 ( .B1(n9703), .B2(n7480), .A(n8266), .ZN(n8268) );
  XNOR2_X1 U9785 ( .A(n8267), .B(n8268), .ZN(n9046) );
  INV_X1 U9786 ( .A(n8267), .ZN(n8269) );
  NAND2_X1 U9787 ( .A1(n8270), .A2(n9151), .ZN(n8273) );
  OR2_X1 U9788 ( .A1(n9154), .A2(n8271), .ZN(n8272) );
  NAND2_X1 U9789 ( .A1(n6030), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8281) );
  OAI21_X1 U9790 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n8275), .A(n8310), .ZN(
        n9549) );
  OR2_X1 U9791 ( .A1(n8332), .A2(n9549), .ZN(n8280) );
  INV_X1 U9792 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8276) );
  OR2_X1 U9793 ( .A1(n5996), .A2(n8276), .ZN(n8279) );
  INV_X1 U9794 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n8277) );
  OR2_X1 U9795 ( .A1(n8333), .A2(n8277), .ZN(n8278) );
  NAND4_X1 U9796 ( .A1(n8281), .A2(n8280), .A3(n8279), .A4(n8278), .ZN(n9568)
         );
  OAI22_X1 U9797 ( .A1(n8405), .A2(n8298), .B1(n8404), .B2(n8297), .ZN(n8282)
         );
  XNOR2_X1 U9798 ( .A(n8282), .B(n8322), .ZN(n8283) );
  AOI22_X1 U9799 ( .A1(n9698), .A2(n8319), .B1(n8324), .B2(n9568), .ZN(n8284)
         );
  XNOR2_X1 U9800 ( .A(n8283), .B(n8284), .ZN(n9121) );
  NAND2_X1 U9801 ( .A1(n8287), .A2(n9151), .ZN(n8290) );
  OR2_X1 U9802 ( .A1(n9154), .A2(n8288), .ZN(n8289) );
  INV_X1 U9803 ( .A(n9692), .ZN(n9539) );
  NAND2_X1 U9804 ( .A1(n5995), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8296) );
  OR2_X1 U9805 ( .A1(n5996), .A2(n8291), .ZN(n8295) );
  INV_X1 U9806 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9008) );
  XNOR2_X1 U9807 ( .A(n8310), .B(n9008), .ZN(n9536) );
  INV_X1 U9808 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8292) );
  OR2_X1 U9809 ( .A1(n8425), .A2(n8292), .ZN(n8293) );
  AND4_X2 U9810 ( .A1(n8296), .A2(n8295), .A3(n8294), .A4(n8293), .ZN(n9124)
         );
  OAI22_X1 U9811 ( .A1(n9539), .A2(n8298), .B1(n9124), .B2(n8297), .ZN(n8299)
         );
  XNOR2_X1 U9812 ( .A(n8299), .B(n8322), .ZN(n9005) );
  NOR2_X1 U9813 ( .A1(n9124), .A2(n8300), .ZN(n8301) );
  AOI21_X1 U9814 ( .B1(n9692), .B2(n8319), .A(n8301), .ZN(n9004) );
  INV_X1 U9815 ( .A(n9004), .ZN(n8328) );
  NAND2_X1 U9816 ( .A1(n8303), .A2(n9151), .ZN(n8306) );
  OR2_X1 U9817 ( .A1(n9154), .A2(n8304), .ZN(n8305) );
  NAND2_X1 U9818 ( .A1(n9688), .A2(n8307), .ZN(n8321) );
  NAND2_X1 U9819 ( .A1(n5995), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8318) );
  INV_X1 U9820 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n8308) );
  OR2_X1 U9821 ( .A1(n5996), .A2(n8308), .ZN(n8317) );
  INV_X1 U9822 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8309) );
  OAI21_X1 U9823 ( .B1(n8310), .B2(n9008), .A(n8309), .ZN(n8313) );
  INV_X1 U9824 ( .A(n8310), .ZN(n8312) );
  AND2_X1 U9825 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n8311) );
  NAND2_X1 U9826 ( .A1(n8312), .A2(n8311), .ZN(n8411) );
  NAND2_X1 U9827 ( .A1(n8313), .A2(n8411), .ZN(n9523) );
  OR2_X1 U9828 ( .A1(n8332), .A2(n9523), .ZN(n8316) );
  INV_X1 U9829 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8314) );
  OR2_X1 U9830 ( .A1(n8425), .A2(n8314), .ZN(n8315) );
  NAND2_X1 U9831 ( .A1(n9542), .A2(n8319), .ZN(n8320) );
  NAND2_X1 U9832 ( .A1(n8321), .A2(n8320), .ZN(n8323) );
  XNOR2_X1 U9833 ( .A(n8323), .B(n8322), .ZN(n8326) );
  AOI22_X1 U9834 ( .A1(n9688), .A2(n7480), .B1(n8324), .B2(n9542), .ZN(n8325)
         );
  XNOR2_X1 U9835 ( .A(n8326), .B(n8325), .ZN(n8342) );
  INV_X1 U9836 ( .A(n8342), .ZN(n8327) );
  NAND2_X1 U9837 ( .A1(n8327), .A2(n9119), .ZN(n8347) );
  NAND2_X1 U9838 ( .A1(n9005), .A2(n8328), .ZN(n8341) );
  INV_X1 U9839 ( .A(n8341), .ZN(n8329) );
  AND2_X1 U9840 ( .A1(n8342), .A2(n8330), .ZN(n8331) );
  NAND2_X1 U9841 ( .A1(n8348), .A2(n8331), .ZN(n8346) );
  NAND2_X1 U9842 ( .A1(n6030), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8338) );
  OR2_X1 U9843 ( .A1(n8332), .A2(n8411), .ZN(n8337) );
  OR2_X1 U9844 ( .A1(n8333), .A2(n6417), .ZN(n8336) );
  INV_X1 U9845 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8334) );
  OR2_X1 U9846 ( .A1(n5996), .A2(n8334), .ZN(n8335) );
  NAND4_X1 U9847 ( .A1(n8338), .A2(n8337), .A3(n8336), .A4(n8335), .ZN(n9529)
         );
  AOI22_X1 U9848 ( .A1(n9139), .A2(n9529), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8340) );
  INV_X1 U9849 ( .A(n9124), .ZN(n9554) );
  NAND2_X1 U9850 ( .A1(n9128), .A2(n9554), .ZN(n8339) );
  OAI211_X1 U9851 ( .C1(n9142), .C2(n9523), .A(n8340), .B(n8339), .ZN(n8344)
         );
  NOR3_X1 U9852 ( .A1(n8342), .A2(n9146), .A3(n8341), .ZN(n8343) );
  AOI211_X1 U9853 ( .C1(n9144), .C2(n9688), .A(n8344), .B(n8343), .ZN(n8345)
         );
  OAI211_X1 U9854 ( .C1(n8348), .C2(n8347), .A(n8346), .B(n8345), .ZN(P1_U3218) );
  OAI222_X1 U9855 ( .A1(n9002), .A2(n8350), .B1(n5103), .B2(n7777), .C1(n8349), 
        .C2(n8438), .ZN(P2_U3329) );
  INV_X1 U9856 ( .A(n8351), .ZN(n8352) );
  NAND2_X1 U9857 ( .A1(n8355), .A2(n8354), .ZN(n8357) );
  XNOR2_X1 U9858 ( .A(n8921), .B(n8376), .ZN(n8356) );
  XNOR2_X1 U9859 ( .A(n8914), .B(n8376), .ZN(n8508) );
  OR2_X1 U9860 ( .A1(n8642), .A2(n5743), .ZN(n8510) );
  AND2_X1 U9861 ( .A1(n8508), .A2(n8510), .ZN(n8361) );
  NAND2_X1 U9862 ( .A1(n8728), .A2(n8367), .ZN(n8447) );
  AOI21_X1 U9863 ( .B1(n8508), .B2(n8642), .A(n8447), .ZN(n8358) );
  NOR2_X1 U9864 ( .A1(n8696), .A2(n5743), .ZN(n8362) );
  XNOR2_X1 U9865 ( .A(n8910), .B(n8365), .ZN(n8494) );
  AND2_X1 U9866 ( .A1(n8362), .A2(n8494), .ZN(n8492) );
  INV_X1 U9867 ( .A(n8494), .ZN(n8364) );
  INV_X1 U9868 ( .A(n8362), .ZN(n8363) );
  NAND2_X1 U9869 ( .A1(n8364), .A2(n8363), .ZN(n8496) );
  XNOR2_X1 U9870 ( .A(n8366), .B(n8365), .ZN(n8368) );
  NAND2_X1 U9871 ( .A1(n8643), .A2(n8367), .ZN(n8369) );
  XNOR2_X1 U9872 ( .A(n8368), .B(n8369), .ZN(n8542) );
  INV_X1 U9873 ( .A(n8368), .ZN(n8371) );
  INV_X1 U9874 ( .A(n8369), .ZN(n8370) );
  NAND2_X1 U9875 ( .A1(n8371), .A2(n8370), .ZN(n8372) );
  XNOR2_X1 U9876 ( .A(n8899), .B(n8376), .ZN(n8373) );
  NOR2_X1 U9877 ( .A1(n8697), .A2(n5743), .ZN(n8374) );
  XNOR2_X1 U9878 ( .A(n8373), .B(n8374), .ZN(n8439) );
  INV_X1 U9879 ( .A(n8373), .ZN(n8375) );
  NOR2_X1 U9880 ( .A1(n8684), .A2(n5743), .ZN(n8377) );
  XNOR2_X1 U9881 ( .A(n8377), .B(n8376), .ZN(n8379) );
  INV_X1 U9882 ( .A(n8379), .ZN(n8380) );
  NOR3_X1 U9883 ( .A1(n4650), .A2(n8380), .A3(n8551), .ZN(n8378) );
  AOI21_X1 U9884 ( .B1(n4650), .B2(n8380), .A(n8378), .ZN(n8386) );
  NOR3_X1 U9885 ( .A1(n4650), .A2(n8379), .A3(n8551), .ZN(n8382) );
  NOR2_X1 U9886 ( .A1(n8894), .A2(n8380), .ZN(n8381) );
  NAND2_X1 U9887 ( .A1(n8387), .A2(n8383), .ZN(n8385) );
  OAI21_X1 U9888 ( .B1(n4650), .B2(n8541), .A(n8553), .ZN(n8384) );
  OAI211_X1 U9889 ( .C1(n8387), .C2(n8386), .A(n8385), .B(n8384), .ZN(n8391)
         );
  NOR2_X1 U9890 ( .A1(n8546), .A2(n8666), .ZN(n8389) );
  OAI22_X1 U9891 ( .A1(n8697), .A2(n8548), .B1(n8547), .B2(n8555), .ZN(n8388)
         );
  AOI211_X1 U9892 ( .C1(P2_REG3_REG_28__SCAN_IN), .C2(n7777), .A(n8389), .B(
        n8388), .ZN(n8390) );
  NAND2_X1 U9893 ( .A1(n8391), .A2(n8390), .ZN(P2_U3222) );
  INV_X1 U9894 ( .A(n9152), .ZN(n8436) );
  INV_X1 U9895 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9153) );
  OAI222_X1 U9896 ( .A1(n5938), .A2(P1_U3084), .B1(n9796), .B2(n8436), .C1(
        n9153), .C2(n9791), .ZN(P1_U3323) );
  NOR2_X1 U9897 ( .A1(n9732), .A2(n9648), .ZN(n8394) );
  INV_X1 U9898 ( .A(n9732), .ZN(n9661) );
  INV_X1 U9899 ( .A(n9648), .ZN(n9114) );
  INV_X1 U9900 ( .A(n9666), .ZN(n9032) );
  OR2_X1 U9901 ( .A1(n9723), .A2(n8395), .ZN(n9206) );
  NAND2_X1 U9902 ( .A1(n9723), .A2(n8395), .ZN(n9343) );
  NAND2_X1 U9903 ( .A1(n9206), .A2(n9343), .ZN(n9624) );
  OAI21_X1 U9904 ( .B1(n9600), .B2(n9617), .A(n9612), .ZN(n8398) );
  NAND2_X1 U9905 ( .A1(n9703), .A2(n9582), .ZN(n9419) );
  NAND2_X1 U9906 ( .A1(n9254), .A2(n9419), .ZN(n9159) );
  NAND2_X1 U9907 ( .A1(n8405), .A2(n8404), .ZN(n8406) );
  OR2_X2 U9908 ( .A1(n9692), .A2(n9124), .ZN(n9362) );
  NAND2_X1 U9909 ( .A1(n9692), .A2(n9124), .ZN(n9361) );
  NAND2_X1 U9910 ( .A1(n9688), .A2(n8429), .ZN(n9364) );
  AND2_X2 U9911 ( .A1(n9365), .A2(n9364), .ZN(n9527) );
  NAND2_X1 U9912 ( .A1(n8407), .A2(n9151), .ZN(n8410) );
  OR2_X1 U9913 ( .A1(n9154), .A2(n8408), .ZN(n8409) );
  NAND2_X1 U9914 ( .A1(n9590), .A2(n9602), .ZN(n9583) );
  INV_X1 U9915 ( .A(n9688), .ZN(n9526) );
  AOI211_X1 U9916 ( .C1(n9682), .C2(n9520), .A(n10101), .B(n9511), .ZN(n9681)
         );
  INV_X1 U9917 ( .A(n9682), .ZN(n9381) );
  INV_X1 U9918 ( .A(n8411), .ZN(n8412) );
  AOI22_X1 U9919 ( .A1(n4399), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8412), .B2(
        n9872), .ZN(n8413) );
  OAI21_X1 U9920 ( .B1(n9381), .B2(n9660), .A(n8413), .ZN(n8433) );
  AND2_X1 U9921 ( .A1(n9202), .A2(n8414), .ZN(n9270) );
  NAND2_X1 U9922 ( .A1(n9330), .A2(n8415), .ZN(n9201) );
  OR2_X1 U9923 ( .A1(n9732), .A2(n9114), .ZN(n9329) );
  NAND2_X1 U9924 ( .A1(n9732), .A2(n9114), .ZN(n9331) );
  NAND2_X1 U9925 ( .A1(n9662), .A2(n9331), .ZN(n9646) );
  OR2_X1 U9926 ( .A1(n9728), .A2(n9032), .ZN(n9344) );
  NAND2_X1 U9927 ( .A1(n9728), .A2(n9032), .ZN(n9332) );
  NAND2_X1 U9928 ( .A1(n9646), .A2(n9647), .ZN(n9645) );
  INV_X1 U9929 ( .A(n9624), .ZN(n9633) );
  OR2_X1 U9930 ( .A1(n9717), .A2(n9600), .ZN(n9210) );
  AND2_X1 U9931 ( .A1(n9717), .A2(n9600), .ZN(n9209) );
  NAND2_X1 U9932 ( .A1(n9714), .A2(n9581), .ZN(n9340) );
  OR2_X1 U9933 ( .A1(n9709), .A2(n9598), .ZN(n9251) );
  NAND2_X1 U9934 ( .A1(n9709), .A2(n9598), .ZN(n9565) );
  NAND2_X1 U9935 ( .A1(n9251), .A2(n9565), .ZN(n9579) );
  NOR2_X1 U9936 ( .A1(n9579), .A2(n9264), .ZN(n9348) );
  INV_X1 U9937 ( .A(n9565), .ZN(n8417) );
  NOR2_X1 U9938 ( .A1(n9159), .A2(n8417), .ZN(n8418) );
  INV_X1 U9939 ( .A(n9254), .ZN(n9354) );
  NAND2_X1 U9940 ( .A1(n9698), .A2(n8404), .ZN(n9351) );
  NAND2_X1 U9941 ( .A1(n9422), .A2(n9351), .ZN(n9547) );
  INV_X1 U9942 ( .A(n9362), .ZN(n8419) );
  INV_X1 U9943 ( .A(n9527), .ZN(n8420) );
  NAND2_X1 U9944 ( .A1(n5995), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8423) );
  NAND2_X1 U9945 ( .A1(n8421), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8422) );
  OAI211_X1 U9946 ( .C1(n8425), .C2(n8424), .A(n8423), .B(n8422), .ZN(n9447)
         );
  INV_X1 U9947 ( .A(n9447), .ZN(n8431) );
  INV_X1 U9948 ( .A(P1_B_REG_SCAN_IN), .ZN(n8426) );
  NOR2_X1 U9949 ( .A1(n8427), .A2(n8426), .ZN(n8428) );
  NOR2_X1 U9950 ( .A1(n9599), .A2(n8428), .ZN(n9506) );
  INV_X1 U9951 ( .A(n9506), .ZN(n8430) );
  NOR2_X1 U9952 ( .A1(n9684), .A2(n4399), .ZN(n8432) );
  OAI21_X1 U9953 ( .B1(n9686), .B2(n9672), .A(n8434), .ZN(P1_U3355) );
  OAI222_X1 U9954 ( .A1(n8438), .A2(n8437), .B1(n9002), .B2(n8436), .C1(n7777), 
        .C2(n5105), .ZN(P2_U3328) );
  XNOR2_X1 U9955 ( .A(n8440), .B(n8439), .ZN(n8446) );
  INV_X1 U9956 ( .A(n8679), .ZN(n8442) );
  OAI22_X1 U9957 ( .A1(n8546), .A2(n8442), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8441), .ZN(n8444) );
  OAI22_X1 U9958 ( .A1(n8644), .A2(n8548), .B1(n8547), .B2(n8684), .ZN(n8443)
         );
  AOI211_X1 U9959 ( .C1(n8899), .C2(n8551), .A(n8444), .B(n8443), .ZN(n8445)
         );
  OAI21_X1 U9960 ( .B1(n8446), .B2(n8553), .A(n8445), .ZN(P2_U3216) );
  NAND2_X1 U9961 ( .A1(n8449), .A2(n8476), .ZN(n8458) );
  INV_X1 U9962 ( .A(n8447), .ZN(n8448) );
  INV_X1 U9963 ( .A(n8450), .ZN(n8452) );
  OAI211_X1 U9964 ( .C1(n8452), .C2(n8451), .A(n8493), .B(n8728), .ZN(n8457)
         );
  OAI22_X1 U9965 ( .A1(n8546), .A2(n8741), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8453), .ZN(n8455) );
  OAI22_X1 U9966 ( .A1(n8642), .A2(n8547), .B1(n8548), .B2(n8641), .ZN(n8454)
         );
  AOI211_X1 U9967 ( .C1(n8921), .C2(n8551), .A(n8455), .B(n8454), .ZN(n8456)
         );
  OAI211_X1 U9968 ( .C1(n8458), .C2(n8507), .A(n8457), .B(n8456), .ZN(P2_U3218) );
  OAI21_X1 U9969 ( .B1(n8462), .B2(n8459), .A(n8460), .ZN(n8469) );
  NOR3_X1 U9970 ( .A1(n8462), .A2(n8461), .A3(n8531), .ZN(n8463) );
  OAI21_X1 U9971 ( .B1(n8463), .B2(n8522), .A(n8805), .ZN(n8467) );
  INV_X1 U9972 ( .A(n8487), .ZN(n8806) );
  OAI22_X1 U9973 ( .A1(n8546), .A2(n8800), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8464), .ZN(n8465) );
  AOI21_X1 U9974 ( .B1(n8523), .B2(n8806), .A(n8465), .ZN(n8466) );
  OAI211_X1 U9975 ( .C1(n4646), .C2(n8541), .A(n8467), .B(n8466), .ZN(n8468)
         );
  AOI21_X1 U9976 ( .B1(n8469), .B2(n8476), .A(n8468), .ZN(n8470) );
  INV_X1 U9977 ( .A(n8470), .ZN(P2_U3221) );
  AOI22_X1 U9978 ( .A1(n8523), .A2(n8568), .B1(n8522), .B2(n5875), .ZN(n8479)
         );
  AOI22_X1 U9979 ( .A1(n4637), .A2(n8551), .B1(n8471), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n8478) );
  OAI21_X1 U9980 ( .B1(n8474), .B2(n8473), .A(n8472), .ZN(n8475) );
  NAND2_X1 U9981 ( .A1(n8476), .A2(n8475), .ZN(n8477) );
  NAND3_X1 U9982 ( .A1(n8479), .A2(n8478), .A3(n8477), .ZN(P2_U3224) );
  INV_X1 U9983 ( .A(n8480), .ZN(n8481) );
  AOI21_X1 U9984 ( .B1(n8517), .B2(n8481), .A(n8553), .ZN(n8485) );
  NOR3_X1 U9985 ( .A1(n8482), .A2(n8487), .A3(n8531), .ZN(n8484) );
  OAI21_X1 U9986 ( .B1(n8485), .B2(n8484), .A(n8483), .ZN(n8491) );
  NOR2_X1 U9987 ( .A1(n8486), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8489) );
  OAI22_X1 U9988 ( .A1(n8641), .A2(n8547), .B1(n8548), .B2(n8487), .ZN(n8488)
         );
  AOI211_X1 U9989 ( .C1(n8538), .C2(n8771), .A(n8489), .B(n8488), .ZN(n8490)
         );
  OAI211_X1 U9990 ( .C1(n8773), .C2(n8541), .A(n8491), .B(n8490), .ZN(P2_U3225) );
  NOR3_X1 U9991 ( .A1(n4754), .A2(n8492), .A3(n8553), .ZN(n8499) );
  INV_X1 U9992 ( .A(n8696), .ZN(n8727) );
  NAND3_X1 U9993 ( .A1(n8494), .A2(n8493), .A3(n8727), .ZN(n8495) );
  OAI21_X1 U9994 ( .B1(n8496), .B2(n8553), .A(n8495), .ZN(n8498) );
  MUX2_X1 U9995 ( .A(n8499), .B(n8498), .S(n8497), .Z(n8500) );
  INV_X1 U9996 ( .A(n8500), .ZN(n8506) );
  OAI22_X1 U9997 ( .A1(n8644), .A2(n8851), .B1(n8642), .B2(n8853), .ZN(n8715)
         );
  INV_X1 U9998 ( .A(n8715), .ZN(n8503) );
  OAI22_X1 U9999 ( .A1(n8503), .A2(n8502), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8501), .ZN(n8504) );
  AOI21_X1 U10000 ( .B1(n8710), .B2(n8538), .A(n8504), .ZN(n8505) );
  OAI211_X1 U10001 ( .C1(n8712), .C2(n8541), .A(n8506), .B(n8505), .ZN(
        P2_U3227) );
  OAI22_X1 U10002 ( .A1(n8511), .A2(n8553), .B1(n8642), .B2(n8531), .ZN(n8509)
         );
  OAI21_X1 U10003 ( .B1(n8511), .B2(n8510), .A(n8509), .ZN(n8516) );
  NOR2_X1 U10004 ( .A1(n8512), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8514) );
  OAI22_X1 U10005 ( .A1(n8763), .A2(n8548), .B1(n8547), .B2(n8696), .ZN(n8513)
         );
  AOI211_X1 U10006 ( .C1(n8538), .C2(n8721), .A(n8514), .B(n8513), .ZN(n8515)
         );
  OAI211_X1 U10007 ( .C1(n8723), .C2(n8541), .A(n8516), .B(n8515), .ZN(
        P2_U3231) );
  INV_X1 U10008 ( .A(n8517), .ZN(n8518) );
  AOI211_X1 U10009 ( .C1(n8520), .C2(n8519), .A(n8553), .B(n8518), .ZN(n8527)
         );
  INV_X1 U10010 ( .A(n8521), .ZN(n8787) );
  AOI22_X1 U10011 ( .A1(n8538), .A2(n8787), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8525) );
  INV_X1 U10012 ( .A(n8762), .ZN(n8794) );
  AOI22_X1 U10013 ( .A1(n8523), .A2(n8794), .B1(n8522), .B2(n8822), .ZN(n8524)
         );
  OAI211_X1 U10014 ( .C1(n8789), .C2(n8541), .A(n8525), .B(n8524), .ZN(n8526)
         );
  OR2_X1 U10015 ( .A1(n8527), .A2(n8526), .ZN(P2_U3235) );
  INV_X1 U10016 ( .A(n8528), .ZN(n8529) );
  AOI21_X1 U10017 ( .B1(n8530), .B2(n8529), .A(n8553), .ZN(n8534) );
  NOR3_X1 U10018 ( .A1(n8532), .A2(n8852), .A3(n8531), .ZN(n8533) );
  OAI21_X1 U10019 ( .B1(n8534), .B2(n8533), .A(n8459), .ZN(n8540) );
  INV_X1 U10020 ( .A(n8535), .ZN(n8814) );
  NOR2_X1 U10021 ( .A1(n8536), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8615) );
  OAI22_X1 U10022 ( .A1(n8852), .A2(n8548), .B1(n8547), .B2(n8636), .ZN(n8537)
         );
  AOI211_X1 U10023 ( .C1(n8538), .C2(n8814), .A(n8615), .B(n8537), .ZN(n8539)
         );
  OAI211_X1 U10024 ( .C1(n8816), .C2(n8541), .A(n8540), .B(n8539), .ZN(
        P2_U3240) );
  XNOR2_X1 U10025 ( .A(n8543), .B(n8542), .ZN(n8554) );
  INV_X1 U10026 ( .A(n8544), .ZN(n8702) );
  OAI22_X1 U10027 ( .A1(n8546), .A2(n8702), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8545), .ZN(n8550) );
  OAI22_X1 U10028 ( .A1(n8696), .A2(n8548), .B1(n8547), .B2(n8697), .ZN(n8549)
         );
  AOI211_X1 U10029 ( .C1(n8906), .C2(n8551), .A(n8550), .B(n8549), .ZN(n8552)
         );
  OAI21_X1 U10030 ( .B1(n8554), .B2(n8553), .A(n8552), .ZN(P2_U3242) );
  MUX2_X1 U10031 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8650), .S(P2_U3966), .Z(
        P2_U3582) );
  INV_X1 U10032 ( .A(n8555), .ZN(n8672) );
  MUX2_X1 U10033 ( .A(n8672), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8567), .Z(
        P2_U3581) );
  INV_X1 U10034 ( .A(n8684), .ZN(n8652) );
  MUX2_X1 U10035 ( .A(n8652), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8567), .Z(
        P2_U3580) );
  INV_X1 U10036 ( .A(n8697), .ZN(n8671) );
  MUX2_X1 U10037 ( .A(n8671), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8567), .Z(
        P2_U3579) );
  MUX2_X1 U10038 ( .A(n8643), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8567), .Z(
        P2_U3578) );
  MUX2_X1 U10039 ( .A(n8727), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8567), .Z(
        P2_U3577) );
  MUX2_X1 U10040 ( .A(n4846), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8567), .Z(
        P2_U3576) );
  MUX2_X1 U10041 ( .A(n8728), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8567), .Z(
        P2_U3575) );
  MUX2_X1 U10042 ( .A(n8780), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8567), .Z(
        P2_U3574) );
  MUX2_X1 U10043 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8794), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10044 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8806), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10045 ( .A(n8822), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8567), .Z(
        P2_U3571) );
  MUX2_X1 U10046 ( .A(n8805), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8567), .Z(
        P2_U3570) );
  MUX2_X1 U10047 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8820), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10048 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8630), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10049 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8627), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10050 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8556), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10051 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8557), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U10052 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8558), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U10053 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8559), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U10054 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8560), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U10055 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8561), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U10056 ( .A(n8562), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8567), .Z(
        P2_U3560) );
  MUX2_X1 U10057 ( .A(n5902), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8567), .Z(
        P2_U3559) );
  MUX2_X1 U10058 ( .A(n8563), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8567), .Z(
        P2_U3558) );
  MUX2_X1 U10059 ( .A(n8564), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8567), .Z(
        P2_U3557) );
  MUX2_X1 U10060 ( .A(n8565), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8567), .Z(
        P2_U3556) );
  MUX2_X1 U10061 ( .A(n8566), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8567), .Z(
        P2_U3555) );
  MUX2_X1 U10062 ( .A(n8568), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8567), .Z(
        P2_U3554) );
  OAI21_X1 U10063 ( .B1(n8571), .B2(n8570), .A(n8569), .ZN(n8572) );
  NAND2_X1 U10064 ( .A1(n10118), .A2(n8572), .ZN(n8582) );
  NOR2_X1 U10065 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8573), .ZN(n8574) );
  AOI21_X1 U10066 ( .B1(n10124), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8574), .ZN(
        n8581) );
  NAND2_X1 U10067 ( .A1(n9815), .A2(n8575), .ZN(n8580) );
  OAI211_X1 U10068 ( .C1(n8578), .C2(n8577), .A(n10119), .B(n8576), .ZN(n8579)
         );
  NAND4_X1 U10069 ( .A1(n8582), .A2(n8581), .A3(n8580), .A4(n8579), .ZN(
        P2_U3256) );
  AOI21_X1 U10070 ( .B1(n8585), .B2(n8584), .A(n8583), .ZN(n8596) );
  INV_X1 U10071 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8587) );
  OAI21_X1 U10072 ( .B1(n8588), .B2(n8587), .A(n8586), .ZN(n8593) );
  AOI211_X1 U10073 ( .C1(n8591), .C2(n8590), .A(n8589), .B(n10122), .ZN(n8592)
         );
  AOI211_X1 U10074 ( .C1(n9815), .C2(n8594), .A(n8593), .B(n8592), .ZN(n8595)
         );
  OAI21_X1 U10075 ( .B1(n8596), .B2(n8611), .A(n8595), .ZN(P2_U3261) );
  AOI211_X1 U10076 ( .C1(n8599), .C2(n8598), .A(n8597), .B(n10122), .ZN(n8608)
         );
  AND2_X1 U10077 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8600) );
  AOI21_X1 U10078 ( .B1(n10124), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8600), .ZN(
        n8605) );
  OAI211_X1 U10079 ( .C1(n8603), .C2(n8602), .A(n10119), .B(n8601), .ZN(n8604)
         );
  OAI211_X1 U10080 ( .C1(n10121), .C2(n8606), .A(n8605), .B(n8604), .ZN(n8607)
         );
  OR2_X1 U10081 ( .A1(n8608), .A2(n8607), .ZN(P2_U3262) );
  NAND2_X1 U10082 ( .A1(n8610), .A2(n8609), .ZN(n8612) );
  AOI21_X1 U10083 ( .B1(n8613), .B2(n8612), .A(n8611), .ZN(n8614) );
  AOI211_X1 U10084 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n10124), .A(n8615), .B(
        n8614), .ZN(n8620) );
  OAI21_X1 U10085 ( .B1(n8617), .B2(n5444), .A(n8616), .ZN(n8618) );
  NAND2_X1 U10086 ( .A1(n10118), .A2(n8618), .ZN(n8619) );
  OAI211_X1 U10087 ( .C1(n10121), .C2(n8621), .A(n8620), .B(n8619), .ZN(
        P2_U3263) );
  INV_X1 U10088 ( .A(n8623), .ZN(n8886) );
  INV_X1 U10089 ( .A(n8622), .ZN(n8883) );
  NAND2_X1 U10090 ( .A1(n8623), .A2(n8655), .ZN(n8882) );
  NAND3_X1 U10091 ( .A1(n8883), .A2(n8876), .A3(n8882), .ZN(n8626) );
  AOI21_X1 U10092 ( .B1(n8878), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8624), .ZN(
        n8625) );
  OAI211_X1 U10093 ( .C1(n8886), .C2(n8871), .A(n8626), .B(n8625), .ZN(
        P2_U3266) );
  OR2_X1 U10094 ( .A1(n8962), .A2(n8627), .ZN(n8628) );
  NAND2_X1 U10095 ( .A1(n8629), .A2(n8628), .ZN(n8856) );
  NAND2_X1 U10096 ( .A1(n8946), .A2(n8805), .ZN(n8634) );
  NAND2_X1 U10097 ( .A1(n8798), .A2(n8635), .ZN(n8637) );
  NAND2_X1 U10098 ( .A1(n8770), .A2(n4958), .ZN(n8640) );
  NAND2_X1 U10099 ( .A1(n8773), .A2(n8762), .ZN(n8639) );
  NAND2_X1 U10100 ( .A1(n8640), .A2(n8639), .ZN(n8748) );
  INV_X1 U10101 ( .A(n8926), .ZN(n8755) );
  INV_X1 U10102 ( .A(n8921), .ZN(n8744) );
  OAI22_X2 U10103 ( .A1(n8707), .A2(n8714), .B1(n8727), .B2(n8910), .ZN(n8690)
         );
  AOI22_X1 U10104 ( .A1(n8664), .A2(n8669), .B1(n8684), .B2(n4650), .ZN(n8646)
         );
  XNOR2_X1 U10105 ( .A(n8646), .B(n8647), .ZN(n8887) );
  INV_X1 U10106 ( .A(n8887), .ZN(n8662) );
  INV_X1 U10107 ( .A(n8647), .ZN(n8648) );
  XNOR2_X1 U10108 ( .A(n8649), .B(n8648), .ZN(n8654) );
  AOI22_X1 U10109 ( .A1(n8652), .A2(n8819), .B1(n8651), .B2(n8650), .ZN(n8653)
         );
  OAI21_X1 U10110 ( .B1(n8665), .B2(n8888), .A(n8655), .ZN(n8889) );
  NOR2_X1 U10111 ( .A1(n8889), .A2(n8656), .ZN(n8660) );
  AOI22_X1 U10112 ( .A1(n8878), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8657), .B2(
        n8868), .ZN(n8658) );
  OAI21_X1 U10113 ( .B1(n8888), .B2(n8871), .A(n8658), .ZN(n8659) );
  AOI211_X1 U10114 ( .C1(n8891), .C2(n8846), .A(n8660), .B(n8659), .ZN(n8661)
         );
  OAI21_X1 U10115 ( .B1(n8662), .B2(n8849), .A(n8661), .ZN(P2_U3267) );
  XNOR2_X1 U10116 ( .A(n8664), .B(n8663), .ZN(n8898) );
  AOI21_X1 U10117 ( .B1(n8894), .B2(n8678), .A(n8665), .ZN(n8895) );
  INV_X1 U10118 ( .A(n8666), .ZN(n8667) );
  AOI22_X1 U10119 ( .A1(n8878), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8667), .B2(
        n8868), .ZN(n8668) );
  OAI21_X1 U10120 ( .B1(n4650), .B2(n8871), .A(n8668), .ZN(n8675) );
  XNOR2_X1 U10121 ( .A(n8670), .B(n8669), .ZN(n8673) );
  AOI222_X1 U10122 ( .A1(n8863), .A2(n8673), .B1(n8672), .B2(n8821), .C1(n8671), .C2(n8819), .ZN(n8897) );
  NOR2_X1 U10123 ( .A1(n8897), .A2(n8878), .ZN(n8674) );
  AOI211_X1 U10124 ( .C1(n8876), .C2(n8895), .A(n8675), .B(n8674), .ZN(n8676)
         );
  OAI21_X1 U10125 ( .B1(n8898), .B2(n8849), .A(n8676), .ZN(P2_U3268) );
  XOR2_X1 U10126 ( .A(n8677), .B(n8683), .Z(n8903) );
  AOI21_X1 U10127 ( .B1(n8899), .B2(n8699), .A(n4651), .ZN(n8900) );
  AOI22_X1 U10128 ( .A1(n8878), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8679), .B2(
        n8868), .ZN(n8680) );
  OAI21_X1 U10129 ( .B1(n4827), .B2(n8871), .A(n8680), .ZN(n8688) );
  NOR2_X1 U10130 ( .A1(n8693), .A2(n8694), .ZN(n8692) );
  NAND2_X1 U10131 ( .A1(n5728), .A2(n8681), .ZN(n8682) );
  AOI211_X1 U10132 ( .C1(n8683), .C2(n8682), .A(n8759), .B(n4438), .ZN(n8686)
         );
  OAI22_X1 U10133 ( .A1(n8684), .A2(n8851), .B1(n8644), .B2(n8853), .ZN(n8685)
         );
  NOR2_X1 U10134 ( .A1(n8686), .A2(n8685), .ZN(n8902) );
  NOR2_X1 U10135 ( .A1(n8902), .A2(n8878), .ZN(n8687) );
  AOI211_X1 U10136 ( .C1(n8876), .C2(n8900), .A(n8688), .B(n8687), .ZN(n8689)
         );
  OAI21_X1 U10137 ( .B1(n8903), .B2(n8849), .A(n8689), .ZN(P2_U3269) );
  XOR2_X1 U10138 ( .A(n8690), .B(n8694), .Z(n8908) );
  AOI22_X1 U10139 ( .A1(n8906), .A2(n8691), .B1(n8878), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8706) );
  AOI21_X1 U10140 ( .B1(n8694), .B2(n8693), .A(n8692), .ZN(n8695) );
  OAI222_X1 U10141 ( .A1(n8851), .A2(n8697), .B1(n8853), .B2(n8696), .C1(n8759), .C2(n8695), .ZN(n8904) );
  INV_X1 U10142 ( .A(n8698), .ZN(n8701) );
  INV_X1 U10143 ( .A(n8699), .ZN(n8700) );
  AOI211_X1 U10144 ( .C1(n8906), .C2(n8701), .A(n10187), .B(n8700), .ZN(n8905)
         );
  INV_X1 U10145 ( .A(n8905), .ZN(n8703) );
  OAI22_X1 U10146 ( .A1(n8703), .A2(n5458), .B1(n8835), .B2(n8702), .ZN(n8704)
         );
  OAI21_X1 U10147 ( .B1(n8904), .B2(n8704), .A(n8846), .ZN(n8705) );
  OAI211_X1 U10148 ( .C1(n8908), .C2(n8849), .A(n8706), .B(n8705), .ZN(
        P2_U3270) );
  XOR2_X1 U10149 ( .A(n8714), .B(n8707), .Z(n8913) );
  INV_X1 U10150 ( .A(n8708), .ZN(n8709) );
  AOI211_X1 U10151 ( .C1(n8910), .C2(n8709), .A(n10187), .B(n8698), .ZN(n8909)
         );
  AOI22_X1 U10152 ( .A1(n8878), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8710), .B2(
        n8868), .ZN(n8711) );
  OAI21_X1 U10153 ( .B1(n8712), .B2(n8871), .A(n8711), .ZN(n8718) );
  XOR2_X1 U10154 ( .A(n8713), .B(n8714), .Z(n8716) );
  AOI21_X1 U10155 ( .B1(n8716), .B2(n8863), .A(n8715), .ZN(n8912) );
  NOR2_X1 U10156 ( .A1(n8912), .A2(n8878), .ZN(n8717) );
  AOI211_X1 U10157 ( .C1(n8909), .C2(n8840), .A(n8718), .B(n8717), .ZN(n8719)
         );
  OAI21_X1 U10158 ( .B1(n8913), .B2(n8849), .A(n8719), .ZN(P2_U3271) );
  AOI21_X1 U10159 ( .B1(n8725), .B2(n8720), .A(n4464), .ZN(n8918) );
  XNOR2_X1 U10160 ( .A(n8723), .B(n8739), .ZN(n8915) );
  AOI22_X1 U10161 ( .A1(n8878), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8721), .B2(
        n8868), .ZN(n8722) );
  OAI21_X1 U10162 ( .B1(n8723), .B2(n8871), .A(n8722), .ZN(n8730) );
  XNOR2_X1 U10163 ( .A(n8724), .B(n8725), .ZN(n8726) );
  AOI222_X1 U10164 ( .A1(n8728), .A2(n8819), .B1(n8727), .B2(n8821), .C1(n8863), .C2(n8726), .ZN(n8917) );
  NOR2_X1 U10165 ( .A1(n8917), .A2(n8878), .ZN(n8729) );
  AOI211_X1 U10166 ( .C1(n8915), .C2(n8876), .A(n8730), .B(n8729), .ZN(n8731)
         );
  OAI21_X1 U10167 ( .B1(n8918), .B2(n8849), .A(n8731), .ZN(P2_U3272) );
  OAI21_X1 U10168 ( .B1(n4424), .B2(n8732), .A(n8736), .ZN(n8734) );
  NAND2_X1 U10169 ( .A1(n8734), .A2(n8733), .ZN(n8735) );
  AOI222_X1 U10170 ( .A1(n8863), .A2(n8735), .B1(n4846), .B2(n8821), .C1(n8780), .C2(n8819), .ZN(n8924) );
  OR2_X1 U10171 ( .A1(n8737), .A2(n8736), .ZN(n8920) );
  NAND3_X1 U10172 ( .A1(n8920), .A2(n8919), .A3(n8738), .ZN(n8747) );
  INV_X1 U10173 ( .A(n8739), .ZN(n8740) );
  AOI21_X1 U10174 ( .B1(n8921), .B2(n8749), .A(n8740), .ZN(n8922) );
  INV_X1 U10175 ( .A(n8741), .ZN(n8742) );
  AOI22_X1 U10176 ( .A1(n8878), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8742), .B2(
        n8868), .ZN(n8743) );
  OAI21_X1 U10177 ( .B1(n8744), .B2(n8871), .A(n8743), .ZN(n8745) );
  AOI21_X1 U10178 ( .B1(n8922), .B2(n8876), .A(n8745), .ZN(n8746) );
  OAI211_X1 U10179 ( .C1(n8878), .C2(n8924), .A(n8747), .B(n8746), .ZN(
        P2_U3273) );
  XOR2_X1 U10180 ( .A(n8748), .B(n8761), .Z(n8930) );
  INV_X1 U10181 ( .A(n8749), .ZN(n8750) );
  AOI21_X1 U10182 ( .B1(n8926), .B2(n8751), .A(n8750), .ZN(n8927) );
  INV_X1 U10183 ( .A(n8752), .ZN(n8753) );
  AOI22_X1 U10184 ( .A1(n8878), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8753), .B2(
        n8868), .ZN(n8754) );
  OAI21_X1 U10185 ( .B1(n8755), .B2(n8871), .A(n8754), .ZN(n8767) );
  AND2_X1 U10186 ( .A1(n8757), .A2(n8756), .ZN(n8778) );
  NAND2_X1 U10187 ( .A1(n8778), .A2(n8758), .ZN(n8760) );
  AOI211_X1 U10188 ( .C1(n8761), .C2(n8760), .A(n8759), .B(n4424), .ZN(n8765)
         );
  OAI22_X1 U10189 ( .A1(n8763), .A2(n8851), .B1(n8762), .B2(n8853), .ZN(n8764)
         );
  NOR2_X1 U10190 ( .A1(n8765), .A2(n8764), .ZN(n8929) );
  NOR2_X1 U10191 ( .A1(n8929), .A2(n8878), .ZN(n8766) );
  AOI211_X1 U10192 ( .C1(n8927), .C2(n8876), .A(n8767), .B(n8766), .ZN(n8768)
         );
  OAI21_X1 U10193 ( .B1(n8930), .B2(n8849), .A(n8768), .ZN(P2_U3274) );
  XOR2_X1 U10194 ( .A(n8770), .B(n8769), .Z(n8935) );
  XNOR2_X1 U10195 ( .A(n8786), .B(n8931), .ZN(n8932) );
  AOI22_X1 U10196 ( .A1(n8878), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8771), .B2(
        n8868), .ZN(n8772) );
  OAI21_X1 U10197 ( .B1(n8773), .B2(n8871), .A(n8772), .ZN(n8783) );
  NAND2_X1 U10198 ( .A1(n8774), .A2(n8775), .ZN(n8777) );
  OAI21_X1 U10199 ( .B1(n4956), .B2(n8779), .A(n8778), .ZN(n8781) );
  AOI222_X1 U10200 ( .A1(n8863), .A2(n8781), .B1(n8780), .B2(n8821), .C1(n8806), .C2(n8819), .ZN(n8934) );
  NOR2_X1 U10201 ( .A1(n8934), .A2(n8878), .ZN(n8782) );
  AOI211_X1 U10202 ( .C1(n8932), .C2(n8876), .A(n8783), .B(n8782), .ZN(n8784)
         );
  OAI21_X1 U10203 ( .B1(n8935), .B2(n8849), .A(n8784), .ZN(P2_U3275) );
  XNOR2_X1 U10204 ( .A(n8785), .B(n8792), .ZN(n8940) );
  AOI21_X1 U10205 ( .B1(n8936), .B2(n4648), .A(n8786), .ZN(n8937) );
  AOI22_X1 U10206 ( .A1(n8878), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8787), .B2(
        n8868), .ZN(n8788) );
  OAI21_X1 U10207 ( .B1(n8789), .B2(n8871), .A(n8788), .ZN(n8796) );
  NAND2_X1 U10208 ( .A1(n8774), .A2(n8804), .ZN(n8803) );
  NAND2_X1 U10209 ( .A1(n8803), .A2(n8790), .ZN(n8791) );
  XOR2_X1 U10210 ( .A(n8792), .B(n8791), .Z(n8793) );
  AOI222_X1 U10211 ( .A1(n8822), .A2(n8819), .B1(n8794), .B2(n8821), .C1(n8863), .C2(n8793), .ZN(n8939) );
  NOR2_X1 U10212 ( .A1(n8939), .A2(n8878), .ZN(n8795) );
  AOI211_X1 U10213 ( .C1(n8937), .C2(n8876), .A(n8796), .B(n8795), .ZN(n8797)
         );
  OAI21_X1 U10214 ( .B1(n8849), .B2(n8940), .A(n8797), .ZN(P2_U3276) );
  XOR2_X1 U10215 ( .A(n8798), .B(n8804), .Z(n8945) );
  AOI211_X1 U10216 ( .C1(n8942), .C2(n8812), .A(n10187), .B(n8799), .ZN(n8941)
         );
  INV_X1 U10217 ( .A(n8800), .ZN(n8801) );
  AOI22_X1 U10218 ( .A1(n8878), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8801), .B2(
        n8868), .ZN(n8802) );
  OAI21_X1 U10219 ( .B1(n4646), .B2(n8871), .A(n8802), .ZN(n8809) );
  OAI21_X1 U10220 ( .B1(n8804), .B2(n8774), .A(n8803), .ZN(n8807) );
  AOI222_X1 U10221 ( .A1(n8863), .A2(n8807), .B1(n8806), .B2(n8821), .C1(n8805), .C2(n8819), .ZN(n8944) );
  NOR2_X1 U10222 ( .A1(n8944), .A2(n8878), .ZN(n8808) );
  AOI211_X1 U10223 ( .C1(n8941), .C2(n8840), .A(n8809), .B(n8808), .ZN(n8810)
         );
  OAI21_X1 U10224 ( .B1(n8945), .B2(n8849), .A(n8810), .ZN(P2_U3277) );
  XNOR2_X1 U10225 ( .A(n8811), .B(n8818), .ZN(n8950) );
  INV_X1 U10226 ( .A(n8812), .ZN(n8813) );
  AOI21_X1 U10227 ( .B1(n8946), .B2(n8831), .A(n8813), .ZN(n8947) );
  AOI22_X1 U10228 ( .A1(n8878), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8814), .B2(
        n8868), .ZN(n8815) );
  OAI21_X1 U10229 ( .B1(n8816), .B2(n8871), .A(n8815), .ZN(n8825) );
  XOR2_X1 U10230 ( .A(n8818), .B(n8817), .Z(n8823) );
  AOI222_X1 U10231 ( .A1(n8863), .A2(n8823), .B1(n8822), .B2(n8821), .C1(n8820), .C2(n8819), .ZN(n8949) );
  NOR2_X1 U10232 ( .A1(n8949), .A2(n8878), .ZN(n8824) );
  AOI211_X1 U10233 ( .C1(n8947), .C2(n8876), .A(n8825), .B(n8824), .ZN(n8826)
         );
  OAI21_X1 U10234 ( .B1(n8950), .B2(n8849), .A(n8826), .ZN(P2_U3278) );
  OAI21_X1 U10235 ( .B1(n8829), .B2(n8828), .A(n8827), .ZN(n8830) );
  INV_X1 U10236 ( .A(n8830), .ZN(n8955) );
  INV_X1 U10237 ( .A(n8865), .ZN(n8833) );
  INV_X1 U10238 ( .A(n8831), .ZN(n8832) );
  AOI211_X1 U10239 ( .C1(n8953), .C2(n8833), .A(n10187), .B(n8832), .ZN(n8952)
         );
  NOR2_X1 U10240 ( .A1(n8834), .A2(n8871), .ZN(n8839) );
  INV_X1 U10241 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8837) );
  OAI22_X1 U10242 ( .A1(n8846), .A2(n8837), .B1(n8836), .B2(n8835), .ZN(n8838)
         );
  AOI211_X1 U10243 ( .C1(n8952), .C2(n8840), .A(n8839), .B(n8838), .ZN(n8848)
         );
  OAI211_X1 U10244 ( .C1(n8843), .C2(n8842), .A(n8841), .B(n8863), .ZN(n8845)
         );
  NAND2_X1 U10245 ( .A1(n8845), .A2(n8844), .ZN(n8951) );
  NAND2_X1 U10246 ( .A1(n8951), .A2(n8846), .ZN(n8847) );
  OAI211_X1 U10247 ( .C1(n8955), .C2(n8849), .A(n8848), .B(n8847), .ZN(
        P2_U3279) );
  XNOR2_X1 U10248 ( .A(n8850), .B(n4850), .ZN(n8862) );
  OAI22_X1 U10249 ( .A1(n8854), .A2(n8853), .B1(n8852), .B2(n8851), .ZN(n8861)
         );
  AND2_X1 U10250 ( .A1(n8856), .A2(n8855), .ZN(n8857) );
  OR2_X1 U10251 ( .A1(n8858), .A2(n8857), .ZN(n8960) );
  NOR2_X1 U10252 ( .A1(n8960), .A2(n8859), .ZN(n8860) );
  AOI211_X1 U10253 ( .C1(n8863), .C2(n8862), .A(n8861), .B(n8860), .ZN(n8959)
         );
  INV_X1 U10254 ( .A(n8864), .ZN(n8866) );
  AOI21_X1 U10255 ( .B1(n8956), .B2(n8866), .A(n8865), .ZN(n8957) );
  INV_X1 U10256 ( .A(n8867), .ZN(n8869) );
  AOI22_X1 U10257 ( .A1(n8878), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8869), .B2(
        n8868), .ZN(n8870) );
  OAI21_X1 U10258 ( .B1(n8872), .B2(n8871), .A(n8870), .ZN(n8875) );
  NOR2_X1 U10259 ( .A1(n8960), .A2(n8873), .ZN(n8874) );
  AOI211_X1 U10260 ( .C1(n8957), .C2(n8876), .A(n8875), .B(n8874), .ZN(n8877)
         );
  OAI21_X1 U10261 ( .B1(n8959), .B2(n8878), .A(n8877), .ZN(P2_U3280) );
  NAND2_X1 U10262 ( .A1(n8879), .A2(n10194), .ZN(n8880) );
  OAI211_X1 U10263 ( .C1(n8881), .C2(n10187), .A(n8880), .B(n8884), .ZN(n8978)
         );
  MUX2_X1 U10264 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8978), .S(n10217), .Z(
        P2_U3551) );
  NAND3_X1 U10265 ( .A1(n8883), .A2(n10195), .A3(n8882), .ZN(n8885) );
  OAI211_X1 U10266 ( .C1(n8886), .C2(n10186), .A(n8885), .B(n8884), .ZN(n8979)
         );
  MUX2_X1 U10267 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8979), .S(n10217), .Z(
        P2_U3550) );
  NAND2_X1 U10268 ( .A1(n8887), .A2(n10177), .ZN(n8893) );
  OAI22_X1 U10269 ( .A1(n8889), .A2(n10187), .B1(n8888), .B2(n10186), .ZN(
        n8890) );
  NOR2_X1 U10270 ( .A1(n8891), .A2(n8890), .ZN(n8892) );
  NAND2_X1 U10271 ( .A1(n8893), .A2(n8892), .ZN(n8980) );
  MUX2_X1 U10272 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8980), .S(n10217), .Z(
        P2_U3549) );
  AOI22_X1 U10273 ( .A1(n8895), .A2(n10195), .B1(n10194), .B2(n8894), .ZN(
        n8896) );
  OAI211_X1 U10274 ( .C1(n8898), .C2(n10199), .A(n8897), .B(n8896), .ZN(n8981)
         );
  MUX2_X1 U10275 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8981), .S(n10217), .Z(
        P2_U3548) );
  AOI22_X1 U10276 ( .A1(n8900), .A2(n10195), .B1(n10194), .B2(n8899), .ZN(
        n8901) );
  OAI211_X1 U10277 ( .C1(n8903), .C2(n10199), .A(n8902), .B(n8901), .ZN(n8982)
         );
  MUX2_X1 U10278 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8982), .S(n10217), .Z(
        P2_U3547) );
  AOI211_X1 U10279 ( .C1(n10194), .C2(n8906), .A(n8905), .B(n8904), .ZN(n8907)
         );
  OAI21_X1 U10280 ( .B1(n8908), .B2(n10199), .A(n8907), .ZN(n8983) );
  MUX2_X1 U10281 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8983), .S(n10217), .Z(
        P2_U3546) );
  AOI21_X1 U10282 ( .B1(n10194), .B2(n8910), .A(n8909), .ZN(n8911) );
  OAI211_X1 U10283 ( .C1(n8913), .C2(n10199), .A(n8912), .B(n8911), .ZN(n8984)
         );
  MUX2_X1 U10284 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8984), .S(n10217), .Z(
        P2_U3545) );
  AOI22_X1 U10285 ( .A1(n8915), .A2(n10195), .B1(n10194), .B2(n8914), .ZN(
        n8916) );
  OAI211_X1 U10286 ( .C1(n8918), .C2(n10199), .A(n8917), .B(n8916), .ZN(n8985)
         );
  MUX2_X1 U10287 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8985), .S(n10217), .Z(
        P2_U3544) );
  NAND3_X1 U10288 ( .A1(n8920), .A2(n8919), .A3(n10177), .ZN(n8925) );
  AOI22_X1 U10289 ( .A1(n8922), .A2(n10195), .B1(n10194), .B2(n8921), .ZN(
        n8923) );
  NAND3_X1 U10290 ( .A1(n8925), .A2(n8924), .A3(n8923), .ZN(n8986) );
  MUX2_X1 U10291 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8986), .S(n10217), .Z(
        P2_U3543) );
  AOI22_X1 U10292 ( .A1(n8927), .A2(n10195), .B1(n10194), .B2(n8926), .ZN(
        n8928) );
  OAI211_X1 U10293 ( .C1(n8930), .C2(n10199), .A(n8929), .B(n8928), .ZN(n8987)
         );
  MUX2_X1 U10294 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8987), .S(n10217), .Z(
        P2_U3542) );
  AOI22_X1 U10295 ( .A1(n8932), .A2(n10195), .B1(n10194), .B2(n8931), .ZN(
        n8933) );
  OAI211_X1 U10296 ( .C1(n8935), .C2(n10199), .A(n8934), .B(n8933), .ZN(n8988)
         );
  MUX2_X1 U10297 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8988), .S(n10217), .Z(
        P2_U3541) );
  AOI22_X1 U10298 ( .A1(n8937), .A2(n10195), .B1(n10194), .B2(n8936), .ZN(
        n8938) );
  OAI211_X1 U10299 ( .C1(n8940), .C2(n10199), .A(n8939), .B(n8938), .ZN(n8989)
         );
  MUX2_X1 U10300 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8989), .S(n10217), .Z(
        P2_U3540) );
  AOI21_X1 U10301 ( .B1(n10194), .B2(n8942), .A(n8941), .ZN(n8943) );
  OAI211_X1 U10302 ( .C1(n8945), .C2(n10199), .A(n8944), .B(n8943), .ZN(n8990)
         );
  MUX2_X1 U10303 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8990), .S(n10217), .Z(
        P2_U3539) );
  AOI22_X1 U10304 ( .A1(n8947), .A2(n10195), .B1(n10194), .B2(n8946), .ZN(
        n8948) );
  OAI211_X1 U10305 ( .C1(n8950), .C2(n10199), .A(n8949), .B(n8948), .ZN(n8991)
         );
  MUX2_X1 U10306 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8991), .S(n10217), .Z(
        P2_U3538) );
  AOI211_X1 U10307 ( .C1(n10194), .C2(n8953), .A(n8952), .B(n8951), .ZN(n8954)
         );
  OAI21_X1 U10308 ( .B1(n8955), .B2(n10199), .A(n8954), .ZN(n8992) );
  MUX2_X1 U10309 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8992), .S(n10217), .Z(
        P2_U3537) );
  AOI22_X1 U10310 ( .A1(n8957), .A2(n10195), .B1(n10194), .B2(n8956), .ZN(
        n8958) );
  OAI211_X1 U10311 ( .C1(n8977), .C2(n8960), .A(n8959), .B(n8958), .ZN(n8993)
         );
  MUX2_X1 U10312 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8993), .S(n10217), .Z(
        P2_U3536) );
  INV_X1 U10313 ( .A(n8961), .ZN(n8966) );
  AOI22_X1 U10314 ( .A1(n8963), .A2(n10195), .B1(n10194), .B2(n8962), .ZN(
        n8964) );
  OAI211_X1 U10315 ( .C1(n8966), .C2(n10199), .A(n8965), .B(n8964), .ZN(n8994)
         );
  MUX2_X1 U10316 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8994), .S(n10217), .Z(
        P2_U3535) );
  AOI22_X1 U10317 ( .A1(n8968), .A2(n10195), .B1(n10194), .B2(n8967), .ZN(
        n8969) );
  OAI211_X1 U10318 ( .C1(n8971), .C2(n10199), .A(n8970), .B(n8969), .ZN(n8995)
         );
  MUX2_X1 U10319 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8995), .S(n10217), .Z(
        P2_U3534) );
  AOI22_X1 U10320 ( .A1(n8973), .A2(n10195), .B1(n10194), .B2(n8972), .ZN(
        n8974) );
  OAI211_X1 U10321 ( .C1(n8977), .C2(n8976), .A(n8975), .B(n8974), .ZN(n8996)
         );
  MUX2_X1 U10322 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8996), .S(n10217), .Z(
        P2_U3533) );
  MUX2_X1 U10323 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8978), .S(n10204), .Z(
        P2_U3519) );
  MUX2_X1 U10324 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8979), .S(n10204), .Z(
        P2_U3518) );
  MUX2_X1 U10325 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8980), .S(n10204), .Z(
        P2_U3517) );
  MUX2_X1 U10326 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8981), .S(n10204), .Z(
        P2_U3516) );
  MUX2_X1 U10327 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8982), .S(n10204), .Z(
        P2_U3515) );
  MUX2_X1 U10328 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8983), .S(n10204), .Z(
        P2_U3514) );
  MUX2_X1 U10329 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8984), .S(n10204), .Z(
        P2_U3513) );
  MUX2_X1 U10330 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8985), .S(n10204), .Z(
        P2_U3512) );
  MUX2_X1 U10331 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8986), .S(n10204), .Z(
        P2_U3511) );
  MUX2_X1 U10332 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8987), .S(n10204), .Z(
        P2_U3510) );
  MUX2_X1 U10333 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8988), .S(n10204), .Z(
        P2_U3509) );
  MUX2_X1 U10334 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8989), .S(n10204), .Z(
        P2_U3508) );
  MUX2_X1 U10335 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8990), .S(n10204), .Z(
        P2_U3507) );
  MUX2_X1 U10336 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8991), .S(n10204), .Z(
        P2_U3505) );
  MUX2_X1 U10337 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8992), .S(n10204), .Z(
        P2_U3502) );
  MUX2_X1 U10338 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8993), .S(n10204), .Z(
        P2_U3499) );
  MUX2_X1 U10339 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8994), .S(n10204), .Z(
        P2_U3496) );
  MUX2_X1 U10340 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8995), .S(n10204), .Z(
        P2_U3493) );
  MUX2_X1 U10341 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8996), .S(n10204), .Z(
        P2_U3490) );
  INV_X1 U10342 ( .A(n9148), .ZN(n9797) );
  NOR4_X1 U10343 ( .A1(n8998), .A2(P2_IR_REG_30__SCAN_IN), .A3(n7777), .A4(
        n8997), .ZN(n8999) );
  AOI21_X1 U10344 ( .B1(n9000), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8999), .ZN(
        n9001) );
  OAI21_X1 U10345 ( .B1(n9797), .B2(n9002), .A(n9001), .ZN(P2_U3327) );
  MUX2_X1 U10346 ( .A(n9003), .B(n10129), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3358) );
  XNOR2_X1 U10347 ( .A(n9005), .B(n9004), .ZN(n9006) );
  XNOR2_X1 U10348 ( .A(n9007), .B(n9006), .ZN(n9013) );
  OAI22_X1 U10349 ( .A1(n9137), .A2(n8404), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9008), .ZN(n9009) );
  AOI21_X1 U10350 ( .B1(n9139), .B2(n9542), .A(n9009), .ZN(n9010) );
  OAI21_X1 U10351 ( .B1(n9142), .B2(n9536), .A(n9010), .ZN(n9011) );
  AOI21_X1 U10352 ( .B1(n9692), .B2(n9144), .A(n9011), .ZN(n9012) );
  OAI21_X1 U10353 ( .B1(n9013), .B2(n9146), .A(n9012), .ZN(P1_U3212) );
  INV_X1 U10354 ( .A(n9015), .ZN(n9016) );
  NOR2_X1 U10355 ( .A1(n9014), .A2(n9016), .ZN(n9018) );
  XNOR2_X1 U10356 ( .A(n9018), .B(n9017), .ZN(n9023) );
  AOI22_X1 U10357 ( .A1(n9128), .A2(n9634), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9020) );
  NAND2_X1 U10358 ( .A1(n9139), .A2(n9567), .ZN(n9019) );
  OAI211_X1 U10359 ( .C1(n9142), .C2(n9604), .A(n9020), .B(n9019), .ZN(n9021)
         );
  AOI21_X1 U10360 ( .B1(n9714), .B2(n9144), .A(n9021), .ZN(n9022) );
  OAI21_X1 U10361 ( .B1(n9023), .B2(n9146), .A(n9022), .ZN(P1_U3214) );
  INV_X1 U10362 ( .A(n9024), .ZN(n9026) );
  NAND2_X1 U10363 ( .A1(n9026), .A2(n9025), .ZN(n9110) );
  NAND2_X1 U10364 ( .A1(n9110), .A2(n9108), .ZN(n9107) );
  NAND2_X1 U10365 ( .A1(n9024), .A2(n9027), .ZN(n9109) );
  NAND2_X1 U10366 ( .A1(n9107), .A2(n9109), .ZN(n9031) );
  XNOR2_X1 U10367 ( .A(n9029), .B(n9028), .ZN(n9030) );
  XNOR2_X1 U10368 ( .A(n9031), .B(n9030), .ZN(n9037) );
  NAND2_X1 U10369 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9502) );
  OAI21_X1 U10370 ( .B1(n9032), .B2(n9125), .A(n9502), .ZN(n9033) );
  AOI21_X1 U10371 ( .B1(n9128), .B2(n9665), .A(n9033), .ZN(n9034) );
  OAI21_X1 U10372 ( .B1(n9142), .B2(n9657), .A(n9034), .ZN(n9035) );
  AOI21_X1 U10373 ( .B1(n9732), .B2(n9144), .A(n9035), .ZN(n9036) );
  OAI21_X1 U10374 ( .B1(n9037), .B2(n9146), .A(n9036), .ZN(P1_U3217) );
  XOR2_X1 U10375 ( .A(n4430), .B(n9038), .Z(n9044) );
  OAI22_X1 U10376 ( .A1(n9125), .A2(n9600), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9039), .ZN(n9040) );
  AOI21_X1 U10377 ( .B1(n9128), .B2(n9666), .A(n9040), .ZN(n9041) );
  OAI21_X1 U10378 ( .B1(n9142), .B2(n9627), .A(n9041), .ZN(n9042) );
  AOI21_X1 U10379 ( .B1(n9723), .B2(n9144), .A(n9042), .ZN(n9043) );
  OAI21_X1 U10380 ( .B1(n9044), .B2(n9146), .A(n9043), .ZN(P1_U3221) );
  XOR2_X1 U10381 ( .A(n9046), .B(n9045), .Z(n9051) );
  AOI22_X1 U10382 ( .A1(n9139), .A2(n9568), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9048) );
  NAND2_X1 U10383 ( .A1(n9128), .A2(n9567), .ZN(n9047) );
  OAI211_X1 U10384 ( .C1(n9142), .C2(n9561), .A(n9048), .B(n9047), .ZN(n9049)
         );
  AOI21_X1 U10385 ( .B1(n9703), .B2(n9144), .A(n9049), .ZN(n9050) );
  OAI21_X1 U10386 ( .B1(n9051), .B2(n9146), .A(n9050), .ZN(P1_U3223) );
  INV_X1 U10387 ( .A(n9052), .ZN(n9057) );
  AOI21_X1 U10388 ( .B1(n9055), .B2(n9053), .A(n9054), .ZN(n9056) );
  OAI21_X1 U10389 ( .B1(n9057), .B2(n9056), .A(n9119), .ZN(n9064) );
  INV_X1 U10390 ( .A(n9142), .ZN(n9092) );
  NOR2_X1 U10391 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9058), .ZN(n9995) );
  AOI21_X1 U10392 ( .B1(n9139), .B2(n9448), .A(n9995), .ZN(n9059) );
  OAI21_X1 U10393 ( .B1(n9060), .B2(n9137), .A(n9059), .ZN(n9061) );
  AOI21_X1 U10394 ( .B1(n9062), .B2(n9092), .A(n9061), .ZN(n9063) );
  OAI211_X1 U10395 ( .C1(n9065), .C2(n9131), .A(n9064), .B(n9063), .ZN(
        P1_U3224) );
  OAI21_X1 U10396 ( .B1(n9068), .B2(n9067), .A(n9066), .ZN(n9069) );
  NAND2_X1 U10397 ( .A1(n9069), .A2(n9119), .ZN(n9075) );
  NOR2_X1 U10398 ( .A1(n9142), .A2(n9070), .ZN(n9073) );
  NAND2_X1 U10399 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10009)
         );
  OAI21_X1 U10400 ( .B1(n9125), .B2(n9071), .A(n10009), .ZN(n9072) );
  AOI211_X1 U10401 ( .C1(n9128), .C2(n9449), .A(n9073), .B(n9072), .ZN(n9074)
         );
  OAI211_X1 U10402 ( .C1(n9076), .C2(n9131), .A(n9075), .B(n9074), .ZN(
        P1_U3226) );
  OAI21_X1 U10403 ( .B1(n9078), .B2(n4467), .A(n9077), .ZN(n9079) );
  NAND2_X1 U10404 ( .A1(n9079), .A2(n9119), .ZN(n9084) );
  NOR2_X1 U10405 ( .A1(n9142), .A2(n9586), .ZN(n9082) );
  INV_X1 U10406 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9080) );
  OAI22_X1 U10407 ( .A1(n9125), .A2(n9582), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9080), .ZN(n9081) );
  AOI211_X1 U10408 ( .C1(n9128), .C2(n8399), .A(n9082), .B(n9081), .ZN(n9083)
         );
  OAI211_X1 U10409 ( .C1(n9590), .C2(n9131), .A(n9084), .B(n9083), .ZN(
        P1_U3227) );
  OAI21_X1 U10410 ( .B1(n9086), .B2(n9088), .A(n9085), .ZN(n9087) );
  OAI21_X1 U10411 ( .B1(n4817), .B2(n9088), .A(n9087), .ZN(n9089) );
  NAND2_X1 U10412 ( .A1(n9089), .A2(n9119), .ZN(n9094) );
  AOI22_X1 U10413 ( .A1(n9649), .A2(n9139), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9090) );
  OAI21_X1 U10414 ( .B1(n9114), .B2(n9137), .A(n9090), .ZN(n9091) );
  AOI21_X1 U10415 ( .B1(n9642), .B2(n9092), .A(n9091), .ZN(n9093) );
  OAI211_X1 U10416 ( .C1(n9644), .C2(n9131), .A(n9094), .B(n9093), .ZN(
        P1_U3231) );
  INV_X1 U10417 ( .A(n9096), .ZN(n9097) );
  NOR2_X1 U10418 ( .A1(n9095), .A2(n9097), .ZN(n9099) );
  XNOR2_X1 U10419 ( .A(n9099), .B(n9098), .ZN(n9104) );
  AOI22_X1 U10420 ( .A1(n9649), .A2(n9128), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9101) );
  NAND2_X1 U10421 ( .A1(n9139), .A2(n8399), .ZN(n9100) );
  OAI211_X1 U10422 ( .C1(n9142), .C2(n9614), .A(n9101), .B(n9100), .ZN(n9102)
         );
  AOI21_X1 U10423 ( .B1(n9717), .B2(n9144), .A(n9102), .ZN(n9103) );
  OAI21_X1 U10424 ( .B1(n9104), .B2(n9146), .A(n9103), .ZN(P1_U3233) );
  INV_X1 U10425 ( .A(n9105), .ZN(n9738) );
  INV_X1 U10426 ( .A(n9109), .ZN(n9106) );
  NOR2_X1 U10427 ( .A1(n9107), .A2(n9106), .ZN(n9112) );
  AOI21_X1 U10428 ( .B1(n9110), .B2(n9109), .A(n9108), .ZN(n9111) );
  OAI21_X1 U10429 ( .B1(n9112), .B2(n9111), .A(n9119), .ZN(n9118) );
  NOR2_X1 U10430 ( .A1(n9142), .A2(n9113), .ZN(n9116) );
  NAND2_X1 U10431 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10019)
         );
  OAI21_X1 U10432 ( .B1(n9125), .B2(n9114), .A(n10019), .ZN(n9115) );
  AOI211_X1 U10433 ( .C1(n9128), .C2(n9448), .A(n9116), .B(n9115), .ZN(n9117)
         );
  OAI211_X1 U10434 ( .C1(n9738), .C2(n9131), .A(n9118), .B(n9117), .ZN(
        P1_U3236) );
  OAI211_X1 U10435 ( .C1(n9122), .C2(n9121), .A(n9120), .B(n9119), .ZN(n9130)
         );
  NOR2_X1 U10436 ( .A1(n9142), .A2(n9549), .ZN(n9127) );
  OAI22_X1 U10437 ( .A1(n9125), .A2(n9124), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9123), .ZN(n9126) );
  AOI211_X1 U10438 ( .C1(n9128), .C2(n8403), .A(n9127), .B(n9126), .ZN(n9129)
         );
  OAI211_X1 U10439 ( .C1(n8405), .C2(n9131), .A(n9130), .B(n9129), .ZN(
        P1_U3238) );
  NAND2_X1 U10440 ( .A1(n9132), .A2(n9053), .ZN(n9133) );
  XOR2_X1 U10441 ( .A(n9134), .B(n9133), .Z(n9147) );
  NOR2_X1 U10442 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9135), .ZN(n9985) );
  NOR2_X1 U10443 ( .A1(n9137), .A2(n9136), .ZN(n9138) );
  AOI211_X1 U10444 ( .C1(n9139), .C2(n9449), .A(n9985), .B(n9138), .ZN(n9140)
         );
  OAI21_X1 U10445 ( .B1(n9142), .B2(n9141), .A(n9140), .ZN(n9143) );
  AOI21_X1 U10446 ( .B1(n9754), .B2(n9144), .A(n9143), .ZN(n9145) );
  OAI21_X1 U10447 ( .B1(n9147), .B2(n9146), .A(n9145), .ZN(P1_U3239) );
  INV_X1 U10448 ( .A(n9507), .ZN(n9158) );
  NAND2_X1 U10449 ( .A1(n9148), .A2(n9151), .ZN(n9150) );
  OR2_X1 U10450 ( .A1(n9154), .A2(n6613), .ZN(n9149) );
  NAND2_X1 U10451 ( .A1(n9152), .A2(n9151), .ZN(n9156) );
  OR2_X1 U10452 ( .A1(n9154), .A2(n9153), .ZN(n9155) );
  NAND2_X1 U10453 ( .A1(n9513), .A2(n8431), .ZN(n9157) );
  NAND2_X1 U10454 ( .A1(n9394), .A2(n9157), .ZN(n9431) );
  NAND2_X1 U10455 ( .A1(n9192), .A2(n9158), .ZN(n9429) );
  INV_X1 U10456 ( .A(n9547), .ZN(n9552) );
  INV_X1 U10457 ( .A(n9340), .ZN(n9160) );
  NAND2_X1 U10458 ( .A1(n9298), .A2(n9162), .ZN(n9303) );
  INV_X1 U10459 ( .A(n9303), .ZN(n9215) );
  INV_X1 U10460 ( .A(n9166), .ZN(n9168) );
  NOR3_X1 U10461 ( .A1(n9169), .A2(n9168), .A3(n9167), .ZN(n9172) );
  NAND4_X1 U10462 ( .A1(n9172), .A2(n4580), .A3(n9171), .A4(n9170), .ZN(n9174)
         );
  NOR2_X1 U10463 ( .A1(n9174), .A2(n9173), .ZN(n9175) );
  AND4_X1 U10464 ( .A1(n9214), .A2(n9215), .A3(n9176), .A4(n9175), .ZN(n9177)
         );
  NAND4_X1 U10465 ( .A1(n7752), .A2(n4470), .A3(n9178), .A4(n9177), .ZN(n9179)
         );
  NOR2_X1 U10466 ( .A1(n9317), .A2(n9179), .ZN(n9180) );
  AND4_X1 U10467 ( .A1(n9664), .A2(n9325), .A3(n9181), .A4(n9180), .ZN(n9182)
         );
  NAND4_X1 U10468 ( .A1(n9618), .A2(n9633), .A3(n9647), .A4(n9182), .ZN(n9183)
         );
  OR2_X1 U10469 ( .A1(n9595), .A2(n9183), .ZN(n9184) );
  NOR2_X1 U10470 ( .A1(n9184), .A2(n9579), .ZN(n9185) );
  AND4_X1 U10471 ( .A1(n9423), .A2(n9552), .A3(n4923), .A4(n9185), .ZN(n9186)
         );
  AND2_X1 U10472 ( .A1(n9527), .A2(n9186), .ZN(n9188) );
  OR2_X1 U10473 ( .A1(n9513), .A2(n8431), .ZN(n9428) );
  NAND4_X1 U10474 ( .A1(n9429), .A2(n9188), .A3(n9428), .A4(n9187), .ZN(n9189)
         );
  NAND2_X1 U10475 ( .A1(n9191), .A2(n9190), .ZN(n9389) );
  NAND2_X1 U10476 ( .A1(n9428), .A2(n9507), .ZN(n9193) );
  NAND2_X1 U10477 ( .A1(n9193), .A2(n9192), .ZN(n9385) );
  NAND2_X1 U10478 ( .A1(n9447), .A2(n9507), .ZN(n9194) );
  NAND2_X1 U10479 ( .A1(n9513), .A2(n9194), .ZN(n9383) );
  INV_X1 U10480 ( .A(n9529), .ZN(n9380) );
  OR2_X1 U10481 ( .A1(n9682), .A2(n9380), .ZN(n9195) );
  NAND2_X1 U10482 ( .A1(n9195), .A2(n9365), .ZN(n9426) );
  NAND2_X1 U10483 ( .A1(n9361), .A2(n9351), .ZN(n9196) );
  NAND2_X1 U10484 ( .A1(n9196), .A2(n9362), .ZN(n9197) );
  AND2_X1 U10485 ( .A1(n9364), .A2(n9197), .ZN(n9198) );
  OR2_X1 U10486 ( .A1(n9426), .A2(n9198), .ZN(n9200) );
  NAND2_X1 U10487 ( .A1(n9682), .A2(n9380), .ZN(n9199) );
  AND2_X1 U10488 ( .A1(n9200), .A2(n9199), .ZN(n9424) );
  INV_X1 U10489 ( .A(n9426), .ZN(n9259) );
  INV_X1 U10490 ( .A(n9264), .ZN(n9574) );
  INV_X1 U10491 ( .A(n9201), .ZN(n9269) );
  AND2_X1 U10492 ( .A1(n9331), .A2(n9202), .ZN(n9334) );
  INV_X1 U10493 ( .A(n9334), .ZN(n9204) );
  NAND2_X1 U10494 ( .A1(n9210), .A2(n9206), .ZN(n9346) );
  INV_X1 U10495 ( .A(n9346), .ZN(n9203) );
  AND2_X1 U10496 ( .A1(n9344), .A2(n9329), .ZN(n9336) );
  OAI211_X1 U10497 ( .C1(n9269), .C2(n9204), .A(n9203), .B(n9336), .ZN(n9211)
         );
  INV_X1 U10498 ( .A(n9332), .ZN(n9205) );
  NAND2_X1 U10499 ( .A1(n9206), .A2(n9205), .ZN(n9207) );
  NAND2_X1 U10500 ( .A1(n9207), .A2(n9343), .ZN(n9208) );
  OR2_X1 U10501 ( .A1(n9209), .A2(n9208), .ZN(n9247) );
  NAND2_X1 U10502 ( .A1(n9247), .A2(n9210), .ZN(n9341) );
  NAND2_X1 U10503 ( .A1(n9211), .A2(n9341), .ZN(n9212) );
  NAND2_X1 U10504 ( .A1(n9574), .A2(n9212), .ZN(n9249) );
  NAND2_X1 U10505 ( .A1(n9312), .A2(n9216), .ZN(n9311) );
  INV_X1 U10506 ( .A(n9298), .ZN(n9213) );
  NOR2_X1 U10507 ( .A1(n9214), .A2(n9213), .ZN(n9305) );
  INV_X1 U10508 ( .A(n9305), .ZN(n9223) );
  NAND2_X1 U10509 ( .A1(n9297), .A2(n9292), .ZN(n9289) );
  INV_X1 U10510 ( .A(n9289), .ZN(n9217) );
  OAI211_X1 U10511 ( .C1(n4719), .C2(n9217), .A(n9216), .B(n9215), .ZN(n9240)
         );
  AND2_X1 U10512 ( .A1(n9294), .A2(n9218), .ZN(n9295) );
  AND2_X1 U10513 ( .A1(n9288), .A2(n9295), .ZN(n9219) );
  NOR2_X1 U10514 ( .A1(n9240), .A2(n9219), .ZN(n9221) );
  NAND2_X1 U10515 ( .A1(n9310), .A2(n9220), .ZN(n9313) );
  OAI21_X1 U10516 ( .B1(n9221), .B2(n9313), .A(n9312), .ZN(n9222) );
  OAI211_X1 U10517 ( .C1(n9311), .C2(n9223), .A(n9222), .B(n9318), .ZN(n9224)
         );
  NAND2_X1 U10518 ( .A1(n9224), .A2(n9319), .ZN(n9225) );
  NAND2_X1 U10519 ( .A1(n9225), .A2(n9323), .ZN(n9226) );
  AND2_X1 U10520 ( .A1(n9226), .A2(n9322), .ZN(n9227) );
  NAND2_X1 U10521 ( .A1(n9270), .A2(n9227), .ZN(n9243) );
  NAND2_X1 U10522 ( .A1(n9243), .A2(n9281), .ZN(n9228) );
  OR2_X1 U10523 ( .A1(n9249), .A2(n9228), .ZN(n9416) );
  INV_X1 U10524 ( .A(n9275), .ZN(n9238) );
  INV_X1 U10525 ( .A(n9229), .ZN(n9231) );
  NAND2_X1 U10526 ( .A1(n9231), .A2(n9230), .ZN(n9271) );
  OR2_X1 U10527 ( .A1(n9232), .A2(n4714), .ZN(n9233) );
  NAND2_X1 U10528 ( .A1(n9271), .A2(n9233), .ZN(n9272) );
  AND2_X1 U10529 ( .A1(n9235), .A2(n9234), .ZN(n9410) );
  NAND2_X1 U10530 ( .A1(n9236), .A2(n9410), .ZN(n9237) );
  OAI211_X1 U10531 ( .C1(n9238), .C2(n9272), .A(n9237), .B(n9279), .ZN(n9239)
         );
  INV_X1 U10532 ( .A(n9239), .ZN(n9250) );
  INV_X1 U10533 ( .A(n9240), .ZN(n9241) );
  AND4_X1 U10534 ( .A1(n9241), .A2(n9312), .A3(n9291), .A4(n9280), .ZN(n9242)
         );
  NAND4_X1 U10535 ( .A1(n9270), .A2(n9242), .A3(n9319), .A4(n9322), .ZN(n9244)
         );
  NAND2_X1 U10536 ( .A1(n9244), .A2(n9243), .ZN(n9245) );
  NAND2_X1 U10537 ( .A1(n9245), .A2(n9331), .ZN(n9246) );
  NOR2_X1 U10538 ( .A1(n9247), .A2(n9246), .ZN(n9248) );
  OR2_X1 U10539 ( .A1(n9249), .A2(n9248), .ZN(n9413) );
  OAI21_X1 U10540 ( .B1(n9416), .B2(n9250), .A(n9413), .ZN(n9255) );
  NAND2_X1 U10541 ( .A1(n9254), .A2(n9251), .ZN(n9266) );
  INV_X1 U10542 ( .A(n9266), .ZN(n9417) );
  NAND2_X1 U10543 ( .A1(n9565), .A2(n9340), .ZN(n9412) );
  NAND2_X1 U10544 ( .A1(n9412), .A2(n9251), .ZN(n9252) );
  AND2_X1 U10545 ( .A1(n9419), .A2(n9252), .ZN(n9268) );
  INV_X1 U10546 ( .A(n9268), .ZN(n9253) );
  AOI22_X1 U10547 ( .A1(n9255), .A2(n9417), .B1(n9254), .B2(n9253), .ZN(n9257)
         );
  INV_X1 U10548 ( .A(n9422), .ZN(n9256) );
  NOR2_X1 U10549 ( .A1(n9257), .A2(n9256), .ZN(n9258) );
  NAND3_X1 U10550 ( .A1(n9259), .A2(n9258), .A3(n9362), .ZN(n9260) );
  NAND3_X1 U10551 ( .A1(n9383), .A2(n9424), .A3(n9260), .ZN(n9261) );
  NAND2_X1 U10552 ( .A1(n9385), .A2(n9261), .ZN(n9262) );
  NAND3_X1 U10553 ( .A1(n9262), .A2(n5948), .A3(n9394), .ZN(n9263) );
  AND2_X1 U10554 ( .A1(n9389), .A2(n9263), .ZN(n9392) );
  AND2_X1 U10555 ( .A1(n9565), .A2(n9264), .ZN(n9265) );
  NOR2_X1 U10556 ( .A1(n9266), .A2(n9265), .ZN(n9267) );
  MUX2_X1 U10557 ( .A(n9268), .B(n9267), .S(n9373), .Z(n9349) );
  MUX2_X1 U10558 ( .A(n9270), .B(n9269), .S(n9373), .Z(n9328) );
  INV_X1 U10559 ( .A(n9271), .ZN(n9273) );
  OAI211_X1 U10560 ( .C1(n9274), .C2(n9273), .A(n4580), .B(n9272), .ZN(n9278)
         );
  AND2_X1 U10561 ( .A1(n9281), .A2(n9275), .ZN(n9277) );
  INV_X1 U10562 ( .A(n9280), .ZN(n9276) );
  AOI21_X1 U10563 ( .B1(n9278), .B2(n9277), .A(n9276), .ZN(n9286) );
  AND2_X1 U10564 ( .A1(n9280), .A2(n9279), .ZN(n9283) );
  INV_X1 U10565 ( .A(n9281), .ZN(n9282) );
  AOI21_X1 U10566 ( .B1(n9284), .B2(n9283), .A(n9282), .ZN(n9285) );
  MUX2_X1 U10567 ( .A(n9286), .B(n9285), .S(n9373), .Z(n9296) );
  INV_X1 U10568 ( .A(n9295), .ZN(n9287) );
  AOI21_X1 U10569 ( .B1(n9296), .B2(n9291), .A(n9287), .ZN(n9290) );
  OAI211_X1 U10570 ( .C1(n9290), .C2(n9289), .A(n9288), .B(n9302), .ZN(n9301)
         );
  NAND2_X1 U10571 ( .A1(n9292), .A2(n9291), .ZN(n9293) );
  AOI22_X1 U10572 ( .A1(n9296), .A2(n9295), .B1(n9294), .B2(n9293), .ZN(n9299)
         );
  OAI211_X1 U10573 ( .C1(n9299), .C2(n4719), .A(n9298), .B(n9297), .ZN(n9300)
         );
  AND2_X1 U10574 ( .A1(n9303), .A2(n9302), .ZN(n9304) );
  NOR2_X1 U10575 ( .A1(n9311), .A2(n9304), .ZN(n9307) );
  NOR2_X1 U10576 ( .A1(n9313), .A2(n9305), .ZN(n9306) );
  MUX2_X1 U10577 ( .A(n9307), .B(n9306), .S(n9373), .Z(n9308) );
  NAND2_X1 U10578 ( .A1(n9311), .A2(n9310), .ZN(n9315) );
  NAND2_X1 U10579 ( .A1(n9313), .A2(n9312), .ZN(n9314) );
  INV_X1 U10580 ( .A(n9373), .ZN(n9379) );
  MUX2_X1 U10581 ( .A(n9315), .B(n9314), .S(n9379), .Z(n9316) );
  INV_X1 U10582 ( .A(n9317), .ZN(n9321) );
  MUX2_X1 U10583 ( .A(n9319), .B(n9318), .S(n9373), .Z(n9320) );
  MUX2_X1 U10584 ( .A(n9323), .B(n9322), .S(n9373), .Z(n9324) );
  NAND3_X1 U10585 ( .A1(n9326), .A2(n9325), .A3(n9324), .ZN(n9327) );
  NAND2_X1 U10586 ( .A1(n9328), .A2(n9327), .ZN(n9335) );
  NAND3_X1 U10587 ( .A1(n9335), .A2(n9330), .A3(n9329), .ZN(n9333) );
  NAND3_X1 U10588 ( .A1(n9333), .A2(n9332), .A3(n9331), .ZN(n9339) );
  NAND2_X1 U10589 ( .A1(n9335), .A2(n9334), .ZN(n9337) );
  NAND2_X1 U10590 ( .A1(n9337), .A2(n9336), .ZN(n9338) );
  MUX2_X1 U10591 ( .A(n9339), .B(n9338), .S(n9373), .Z(n9345) );
  OAI211_X1 U10592 ( .C1(n9346), .C2(n9345), .A(n9341), .B(n9340), .ZN(n9342)
         );
  AOI21_X1 U10593 ( .B1(n9345), .B2(n9344), .A(n4712), .ZN(n9347) );
  OAI22_X1 U10594 ( .A1(n9359), .A2(n9698), .B1(n9379), .B2(n9419), .ZN(n9350)
         );
  OAI21_X1 U10595 ( .B1(n9354), .B2(n9568), .A(n9351), .ZN(n9352) );
  MUX2_X1 U10596 ( .A(n9352), .B(n8405), .S(n9373), .Z(n9353) );
  OAI21_X1 U10597 ( .B1(n8405), .B2(n9354), .A(n9361), .ZN(n9357) );
  NAND2_X1 U10598 ( .A1(n9419), .A2(n9568), .ZN(n9355) );
  NAND2_X1 U10599 ( .A1(n9362), .A2(n9355), .ZN(n9356) );
  MUX2_X1 U10600 ( .A(n9357), .B(n9356), .S(n9373), .Z(n9358) );
  OAI21_X1 U10601 ( .B1(n9359), .B2(n9540), .A(n9358), .ZN(n9360) );
  MUX2_X1 U10602 ( .A(n9362), .B(n9361), .S(n9373), .Z(n9363) );
  AND2_X1 U10603 ( .A1(n9527), .A2(n9363), .ZN(n9369) );
  INV_X1 U10604 ( .A(n9364), .ZN(n9367) );
  INV_X1 U10605 ( .A(n9365), .ZN(n9366) );
  NAND3_X1 U10606 ( .A1(n9383), .A2(n9372), .A3(n9529), .ZN(n9370) );
  NAND2_X1 U10607 ( .A1(n9385), .A2(n9370), .ZN(n9371) );
  NAND2_X1 U10608 ( .A1(n9371), .A2(n9379), .ZN(n9388) );
  INV_X1 U10609 ( .A(n9372), .ZN(n9382) );
  AND2_X1 U10610 ( .A1(n9529), .A2(n9373), .ZN(n9375) );
  NAND2_X1 U10611 ( .A1(n9382), .A2(n9375), .ZN(n9377) );
  NAND2_X1 U10612 ( .A1(n9682), .A2(n9373), .ZN(n9374) );
  OAI21_X1 U10613 ( .B1(n9682), .B2(n9375), .A(n9374), .ZN(n9376) );
  NAND3_X1 U10614 ( .A1(n9377), .A2(n9383), .A3(n9376), .ZN(n9378) );
  OAI21_X1 U10615 ( .B1(n9379), .B2(n9383), .A(n9378), .ZN(n9386) );
  NAND4_X1 U10616 ( .A1(n9383), .A2(n9382), .A3(n9381), .A4(n9380), .ZN(n9384)
         );
  NAND3_X1 U10617 ( .A1(n9386), .A2(n9385), .A3(n9384), .ZN(n9387) );
  NAND3_X1 U10618 ( .A1(n9388), .A2(n9394), .A3(n9387), .ZN(n9395) );
  OAI21_X1 U10619 ( .B1(n9395), .B2(n9390), .A(n9389), .ZN(n9391) );
  MUX2_X1 U10620 ( .A(n9392), .B(n9391), .S(n10039), .Z(n9436) );
  AND4_X1 U10621 ( .A1(n9395), .A2(n5948), .A3(n9394), .A4(n9393), .ZN(n9397)
         );
  OR2_X2 U10622 ( .A1(n9397), .A2(n7142), .ZN(n9435) );
  INV_X1 U10623 ( .A(n9398), .ZN(n9400) );
  NAND2_X1 U10624 ( .A1(n4400), .A2(n10045), .ZN(n9399) );
  NAND3_X1 U10625 ( .A1(n9400), .A2(n5948), .A3(n9399), .ZN(n9401) );
  NAND2_X1 U10626 ( .A1(n9402), .A2(n9401), .ZN(n9404) );
  OAI21_X1 U10627 ( .B1(n9405), .B2(n9404), .A(n9403), .ZN(n9407) );
  NAND2_X1 U10628 ( .A1(n9407), .A2(n9406), .ZN(n9411) );
  INV_X1 U10629 ( .A(n9408), .ZN(n9409) );
  AOI21_X1 U10630 ( .B1(n9411), .B2(n9410), .A(n9409), .ZN(n9415) );
  INV_X1 U10631 ( .A(n9412), .ZN(n9414) );
  OAI211_X1 U10632 ( .C1(n9416), .C2(n9415), .A(n9414), .B(n9413), .ZN(n9418)
         );
  NAND2_X1 U10633 ( .A1(n9418), .A2(n9417), .ZN(n9420) );
  NAND2_X1 U10634 ( .A1(n9420), .A2(n9419), .ZN(n9421) );
  NAND3_X1 U10635 ( .A1(n9423), .A2(n9422), .A3(n9421), .ZN(n9425) );
  OAI21_X1 U10636 ( .B1(n9426), .B2(n9425), .A(n9424), .ZN(n9427) );
  AND2_X1 U10637 ( .A1(n9428), .A2(n9427), .ZN(n9430) );
  OAI21_X1 U10638 ( .B1(n9431), .B2(n9430), .A(n9429), .ZN(n9432) );
  XNOR2_X1 U10639 ( .A(n9432), .B(n9499), .ZN(n9433) );
  NAND3_X1 U10640 ( .A1(n9439), .A2(n9438), .A3(n9437), .ZN(n9440) );
  NOR2_X1 U10641 ( .A1(n9441), .A2(n9440), .ZN(n9444) );
  OAI21_X1 U10642 ( .B1(n9442), .B2(n9445), .A(P1_B_REG_SCAN_IN), .ZN(n9443)
         );
  OAI22_X1 U10643 ( .A1(n9446), .A2(n9445), .B1(n9444), .B2(n9443), .ZN(
        P1_U3240) );
  MUX2_X1 U10644 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9447), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10645 ( .A(n9529), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9462), .Z(
        P1_U3584) );
  MUX2_X1 U10646 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9542), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10647 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9554), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10648 ( .A(n9568), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9462), .Z(
        P1_U3581) );
  MUX2_X1 U10649 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n8403), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10650 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9567), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10651 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n8399), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10652 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9634), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10653 ( .A(n9649), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9462), .Z(
        P1_U3576) );
  MUX2_X1 U10654 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9666), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10655 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9648), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10656 ( .A(n9665), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9462), .Z(
        P1_U3573) );
  MUX2_X1 U10657 ( .A(n9448), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9462), .Z(
        P1_U3572) );
  MUX2_X1 U10658 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9449), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10659 ( .A(n9450), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9462), .Z(
        P1_U3570) );
  MUX2_X1 U10660 ( .A(n9451), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9462), .Z(
        P1_U3569) );
  MUX2_X1 U10661 ( .A(n9868), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9462), .Z(
        P1_U3568) );
  MUX2_X1 U10662 ( .A(n9452), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9462), .Z(
        P1_U3567) );
  MUX2_X1 U10663 ( .A(n9866), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9462), .Z(
        P1_U3566) );
  MUX2_X1 U10664 ( .A(n9453), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9462), .Z(
        P1_U3565) );
  MUX2_X1 U10665 ( .A(n9454), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9462), .Z(
        P1_U3564) );
  MUX2_X1 U10666 ( .A(n9455), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9462), .Z(
        P1_U3563) );
  MUX2_X1 U10667 ( .A(n9456), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9462), .Z(
        P1_U3562) );
  MUX2_X1 U10668 ( .A(n9457), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9462), .Z(
        P1_U3561) );
  MUX2_X1 U10669 ( .A(n9458), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9462), .Z(
        P1_U3560) );
  MUX2_X1 U10670 ( .A(n9459), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9462), .Z(
        P1_U3559) );
  MUX2_X1 U10671 ( .A(n9460), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9462), .Z(
        P1_U3558) );
  MUX2_X1 U10672 ( .A(n9461), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9462), .Z(
        P1_U3557) );
  MUX2_X1 U10673 ( .A(n4400), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9462), .Z(
        P1_U3556) );
  XNOR2_X1 U10674 ( .A(n9956), .B(n9463), .ZN(n9960) );
  NAND2_X1 U10675 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9947), .ZN(n9465) );
  OAI21_X1 U10676 ( .B1(n9947), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9465), .ZN(
        n9943) );
  OAI21_X1 U10677 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9476), .A(n9464), .ZN(
        n9944) );
  NOR2_X1 U10678 ( .A1(n9943), .A2(n9944), .ZN(n9942) );
  NOR2_X1 U10679 ( .A1(n9466), .A2(n9483), .ZN(n9467) );
  XNOR2_X1 U10680 ( .A(n9466), .B(n9483), .ZN(n9971) );
  NOR2_X1 U10681 ( .A1(n7590), .A2(n9971), .ZN(n9970) );
  NOR2_X1 U10682 ( .A1(n9467), .A2(n9970), .ZN(n9468) );
  NOR2_X1 U10683 ( .A1(n9468), .A2(n9485), .ZN(n9469) );
  NAND2_X1 U10684 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9996), .ZN(n9470) );
  OAI21_X1 U10685 ( .B1(n9996), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9470), .ZN(
        n9993) );
  AOI21_X1 U10686 ( .B1(n9996), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9992), .ZN(
        n10004) );
  OR2_X1 U10687 ( .A1(n10008), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9472) );
  NAND2_X1 U10688 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n10008), .ZN(n9471) );
  NAND2_X1 U10689 ( .A1(n9472), .A2(n9471), .ZN(n10005) );
  NOR2_X1 U10690 ( .A1(n10004), .A2(n10005), .ZN(n10003) );
  NOR2_X1 U10691 ( .A1(n10027), .A2(n9473), .ZN(n9474) );
  AOI21_X1 U10692 ( .B1(n10027), .B2(n9473), .A(n9474), .ZN(n10023) );
  NAND2_X1 U10693 ( .A1(n9498), .A2(n9475), .ZN(n9496) );
  XNOR2_X1 U10694 ( .A(n10027), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n10030) );
  INV_X1 U10695 ( .A(n10008), .ZN(n9490) );
  INV_X1 U10696 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9489) );
  XNOR2_X1 U10697 ( .A(n9490), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n10015) );
  INV_X1 U10698 ( .A(n9996), .ZN(n9488) );
  XOR2_X1 U10699 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9996), .Z(n9998) );
  INV_X1 U10700 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9482) );
  INV_X1 U10701 ( .A(n9956), .ZN(n9481) );
  MUX2_X1 U10702 ( .A(n9482), .B(P1_REG1_REG_13__SCAN_IN), .S(n9956), .Z(n9964) );
  INV_X1 U10703 ( .A(n9947), .ZN(n9480) );
  NOR2_X1 U10704 ( .A1(n9476), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9477) );
  NOR2_X1 U10705 ( .A1(n9478), .A2(n9477), .ZN(n9950) );
  MUX2_X1 U10706 ( .A(n9479), .B(P1_REG1_REG_12__SCAN_IN), .S(n9947), .Z(n9949) );
  NOR2_X1 U10707 ( .A1(n9950), .A2(n9949), .ZN(n9948) );
  AOI21_X1 U10708 ( .B1(n9480), .B2(n9479), .A(n9948), .ZN(n9965) );
  NOR2_X1 U10709 ( .A1(n9964), .A2(n9965), .ZN(n9963) );
  AOI21_X1 U10710 ( .B1(n9482), .B2(n9481), .A(n9963), .ZN(n9977) );
  MUX2_X1 U10711 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9893), .S(n9483), .Z(n9976) );
  NOR2_X1 U10712 ( .A1(n9977), .A2(n9976), .ZN(n9975) );
  AOI21_X1 U10713 ( .B1(n9483), .B2(n9893), .A(n9975), .ZN(n9484) );
  NAND2_X1 U10714 ( .A1(n9986), .A2(n9484), .ZN(n9486) );
  XNOR2_X1 U10715 ( .A(n9485), .B(n9484), .ZN(n9988) );
  NAND2_X1 U10716 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9988), .ZN(n9987) );
  NAND2_X1 U10717 ( .A1(n9486), .A2(n9987), .ZN(n9999) );
  NAND2_X1 U10718 ( .A1(n9998), .A2(n9999), .ZN(n9997) );
  OAI21_X1 U10719 ( .B1(n9488), .B2(n9487), .A(n9997), .ZN(n10014) );
  NAND2_X1 U10720 ( .A1(n10015), .A2(n10014), .ZN(n10013) );
  OAI21_X1 U10721 ( .B1(n9490), .B2(n9489), .A(n10013), .ZN(n10029) );
  NOR2_X1 U10722 ( .A1(n10030), .A2(n10029), .ZN(n10028) );
  AOI21_X1 U10723 ( .B1(n9492), .B2(n9491), .A(n10028), .ZN(n9494) );
  XOR2_X1 U10724 ( .A(n9494), .B(n9493), .Z(n9497) );
  AOI21_X1 U10725 ( .B1(n9497), .B2(n10012), .A(n10026), .ZN(n9495) );
  NAND2_X1 U10726 ( .A1(n9496), .A2(n9495), .ZN(n9501) );
  OAI22_X1 U10727 ( .A1(n9498), .A2(n10020), .B1(n9497), .B2(n10032), .ZN(
        n9500) );
  MUX2_X1 U10728 ( .A(n9501), .B(n9500), .S(n9499), .Z(n9504) );
  OAI21_X1 U10729 ( .B1(n10035), .B2(n4506), .A(n9502), .ZN(n9503) );
  NAND2_X1 U10730 ( .A1(n9679), .A2(n9511), .ZN(n9676) );
  XNOR2_X1 U10731 ( .A(n9676), .B(n9192), .ZN(n9674) );
  NOR2_X1 U10732 ( .A1(n9610), .A2(n9505), .ZN(n9508) );
  NAND2_X1 U10733 ( .A1(n9507), .A2(n9506), .ZN(n9677) );
  NOR2_X1 U10734 ( .A1(n4399), .A2(n9677), .ZN(n9514) );
  AOI211_X1 U10735 ( .C1(n9192), .C2(n9874), .A(n9508), .B(n9514), .ZN(n9509)
         );
  OAI21_X1 U10736 ( .B1(n9674), .B2(n9510), .A(n9509), .ZN(P1_U3261) );
  INV_X1 U10737 ( .A(n9511), .ZN(n9512) );
  NAND2_X1 U10738 ( .A1(n9513), .A2(n9512), .ZN(n9675) );
  NAND3_X1 U10739 ( .A1(n9676), .A2(n9670), .A3(n9675), .ZN(n9516) );
  AOI21_X1 U10740 ( .B1(n4399), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9514), .ZN(
        n9515) );
  OAI211_X1 U10741 ( .C1(n9679), .C2(n9660), .A(n9516), .B(n9515), .ZN(
        P1_U3262) );
  AOI21_X1 U10742 ( .B1(n9527), .B2(n9518), .A(n9517), .ZN(n9519) );
  INV_X1 U10743 ( .A(n9519), .ZN(n9691) );
  INV_X1 U10744 ( .A(n9534), .ZN(n9522) );
  INV_X1 U10745 ( .A(n9520), .ZN(n9521) );
  AOI211_X1 U10746 ( .C1(n9688), .C2(n9522), .A(n10101), .B(n9521), .ZN(n9687)
         );
  INV_X1 U10747 ( .A(n9523), .ZN(n9524) );
  AOI22_X1 U10748 ( .A1(n4399), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9524), .B2(
        n9872), .ZN(n9525) );
  OAI21_X1 U10749 ( .B1(n9526), .B2(n9660), .A(n9525), .ZN(n9531) );
  OAI21_X1 U10750 ( .B1(n9691), .B2(n9672), .A(n9532), .ZN(P1_U3263) );
  XNOR2_X1 U10751 ( .A(n9533), .B(n9540), .ZN(n9696) );
  INV_X1 U10752 ( .A(n9548), .ZN(n9535) );
  AOI21_X1 U10753 ( .B1(n9692), .B2(n9535), .A(n9534), .ZN(n9693) );
  INV_X1 U10754 ( .A(n9536), .ZN(n9537) );
  AOI22_X1 U10755 ( .A1(n4399), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9537), .B2(
        n9872), .ZN(n9538) );
  OAI21_X1 U10756 ( .B1(n9539), .B2(n9660), .A(n9538), .ZN(n9545) );
  XNOR2_X1 U10757 ( .A(n9541), .B(n9540), .ZN(n9543) );
  AOI222_X1 U10758 ( .A1(n9870), .A2(n9543), .B1(n9542), .B2(n9867), .C1(n9568), .C2(n9865), .ZN(n9695) );
  NOR2_X1 U10759 ( .A1(n9695), .A2(n4399), .ZN(n9544) );
  AOI211_X1 U10760 ( .C1(n9670), .C2(n9693), .A(n9545), .B(n9544), .ZN(n9546)
         );
  OAI21_X1 U10761 ( .B1(n9696), .B2(n9672), .A(n9546), .ZN(P1_U3264) );
  XNOR2_X1 U10762 ( .A(n4461), .B(n9547), .ZN(n9701) );
  AOI211_X1 U10763 ( .C1(n9698), .C2(n9560), .A(n10101), .B(n9548), .ZN(n9697)
         );
  INV_X1 U10764 ( .A(n9549), .ZN(n9550) );
  AOI22_X1 U10765 ( .A1(n4399), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9550), .B2(
        n9872), .ZN(n9551) );
  OAI21_X1 U10766 ( .B1(n8405), .B2(n9660), .A(n9551), .ZN(n9557) );
  XNOR2_X1 U10767 ( .A(n9553), .B(n9552), .ZN(n9555) );
  AOI222_X1 U10768 ( .A1(n9870), .A2(n9555), .B1(n9554), .B2(n9867), .C1(n8403), .C2(n9865), .ZN(n9700) );
  NOR2_X1 U10769 ( .A1(n9700), .A2(n4399), .ZN(n9556) );
  AOI211_X1 U10770 ( .C1(n9697), .C2(n9884), .A(n9557), .B(n9556), .ZN(n9558)
         );
  OAI21_X1 U10771 ( .B1(n9701), .B2(n9672), .A(n9558), .ZN(P1_U3265) );
  XNOR2_X1 U10772 ( .A(n9559), .B(n4923), .ZN(n9706) );
  AOI211_X1 U10773 ( .C1(n9703), .C2(n9583), .A(n10101), .B(n4766), .ZN(n9702)
         );
  INV_X1 U10774 ( .A(n9561), .ZN(n9562) );
  AOI22_X1 U10775 ( .A1(n4399), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9562), .B2(
        n9872), .ZN(n9563) );
  OAI21_X1 U10776 ( .B1(n9564), .B2(n9660), .A(n9563), .ZN(n9571) );
  NAND2_X1 U10777 ( .A1(n9576), .A2(n9565), .ZN(n9566) );
  XNOR2_X1 U10778 ( .A(n9566), .B(n4923), .ZN(n9569) );
  AOI222_X1 U10779 ( .A1(n9870), .A2(n9569), .B1(n9568), .B2(n9867), .C1(n9567), .C2(n9865), .ZN(n9705) );
  NOR2_X1 U10780 ( .A1(n9705), .A2(n4399), .ZN(n9570) );
  AOI211_X1 U10781 ( .C1(n9702), .C2(n9884), .A(n9571), .B(n9570), .ZN(n9572)
         );
  OAI21_X1 U10782 ( .B1(n9706), .B2(n9672), .A(n9572), .ZN(P1_U3266) );
  XOR2_X1 U10783 ( .A(n9573), .B(n9579), .Z(n9711) );
  NAND2_X1 U10784 ( .A1(n9575), .A2(n9574), .ZN(n9578) );
  INV_X1 U10785 ( .A(n9576), .ZN(n9577) );
  AOI21_X1 U10786 ( .B1(n9579), .B2(n9578), .A(n9577), .ZN(n9580) );
  OAI222_X1 U10787 ( .A1(n9599), .A2(n9582), .B1(n9601), .B2(n9581), .C1(n9596), .C2(n9580), .ZN(n9707) );
  INV_X1 U10788 ( .A(n9602), .ZN(n9585) );
  INV_X1 U10789 ( .A(n9583), .ZN(n9584) );
  AOI211_X1 U10790 ( .C1(n9709), .C2(n9585), .A(n10101), .B(n9584), .ZN(n9708)
         );
  NAND2_X1 U10791 ( .A1(n9708), .A2(n9884), .ZN(n9589) );
  INV_X1 U10792 ( .A(n9586), .ZN(n9587) );
  AOI22_X1 U10793 ( .A1(n4399), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9587), .B2(
        n9872), .ZN(n9588) );
  OAI211_X1 U10794 ( .C1(n9590), .C2(n9660), .A(n9589), .B(n9588), .ZN(n9591)
         );
  AOI21_X1 U10795 ( .B1(n9707), .B2(n9610), .A(n9591), .ZN(n9592) );
  OAI21_X1 U10796 ( .B1(n9711), .B2(n9672), .A(n9592), .ZN(P1_U3267) );
  XOR2_X1 U10797 ( .A(n9593), .B(n9595), .Z(n9716) );
  XOR2_X1 U10798 ( .A(n9595), .B(n9594), .Z(n9597) );
  OAI222_X1 U10799 ( .A1(n9601), .A2(n9600), .B1(n9599), .B2(n9598), .C1(n9597), .C2(n9596), .ZN(n9712) );
  INV_X1 U10800 ( .A(n9613), .ZN(n9603) );
  AOI211_X1 U10801 ( .C1(n9714), .C2(n9603), .A(n10101), .B(n9602), .ZN(n9713)
         );
  NAND2_X1 U10802 ( .A1(n9713), .A2(n9884), .ZN(n9607) );
  INV_X1 U10803 ( .A(n9604), .ZN(n9605) );
  AOI22_X1 U10804 ( .A1(n4399), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9605), .B2(
        n9872), .ZN(n9606) );
  OAI211_X1 U10805 ( .C1(n9608), .C2(n9660), .A(n9607), .B(n9606), .ZN(n9609)
         );
  AOI21_X1 U10806 ( .B1(n9712), .B2(n9610), .A(n9609), .ZN(n9611) );
  OAI21_X1 U10807 ( .B1(n9716), .B2(n9672), .A(n9611), .ZN(P1_U3268) );
  XNOR2_X1 U10808 ( .A(n9612), .B(n9618), .ZN(n9721) );
  AOI21_X1 U10809 ( .B1(n9717), .B2(n9626), .A(n9613), .ZN(n9718) );
  INV_X1 U10810 ( .A(n9614), .ZN(n9615) );
  AOI22_X1 U10811 ( .A1(n4399), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9615), .B2(
        n9872), .ZN(n9616) );
  OAI21_X1 U10812 ( .B1(n9617), .B2(n9660), .A(n9616), .ZN(n9622) );
  XNOR2_X1 U10813 ( .A(n9619), .B(n9618), .ZN(n9620) );
  AOI222_X1 U10814 ( .A1(n9870), .A2(n9620), .B1(n8399), .B2(n9867), .C1(n9649), .C2(n9865), .ZN(n9720) );
  NOR2_X1 U10815 ( .A1(n9720), .A2(n4399), .ZN(n9621) );
  AOI211_X1 U10816 ( .C1(n9718), .C2(n9670), .A(n9622), .B(n9621), .ZN(n9623)
         );
  OAI21_X1 U10817 ( .B1(n9721), .B2(n9672), .A(n9623), .ZN(P1_U3269) );
  XNOR2_X1 U10818 ( .A(n9625), .B(n9624), .ZN(n9726) );
  AOI211_X1 U10819 ( .C1(n9723), .C2(n9640), .A(n10101), .B(n4767), .ZN(n9722)
         );
  INV_X1 U10820 ( .A(n9723), .ZN(n9630) );
  INV_X1 U10821 ( .A(n9627), .ZN(n9628) );
  AOI22_X1 U10822 ( .A1(n9628), .A2(n9872), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n4399), .ZN(n9629) );
  OAI21_X1 U10823 ( .B1(n9630), .B2(n9660), .A(n9629), .ZN(n9637) );
  OAI21_X1 U10824 ( .B1(n9633), .B2(n9632), .A(n9631), .ZN(n9635) );
  AOI222_X1 U10825 ( .A1(n9870), .A2(n9635), .B1(n9634), .B2(n9867), .C1(n9666), .C2(n9865), .ZN(n9725) );
  NOR2_X1 U10826 ( .A1(n9725), .A2(n4399), .ZN(n9636) );
  AOI211_X1 U10827 ( .C1(n9722), .C2(n9884), .A(n9637), .B(n9636), .ZN(n9638)
         );
  OAI21_X1 U10828 ( .B1(n9726), .B2(n9672), .A(n9638), .ZN(P1_U3270) );
  XOR2_X1 U10829 ( .A(n9647), .B(n9639), .Z(n9731) );
  INV_X1 U10830 ( .A(n9655), .ZN(n9641) );
  AOI211_X1 U10831 ( .C1(n9728), .C2(n9641), .A(n10101), .B(n4768), .ZN(n9727)
         );
  AOI22_X1 U10832 ( .A1(n9642), .A2(n9872), .B1(n4399), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9643) );
  OAI21_X1 U10833 ( .B1(n9644), .B2(n9660), .A(n9643), .ZN(n9652) );
  OAI21_X1 U10834 ( .B1(n9647), .B2(n9646), .A(n9645), .ZN(n9650) );
  AOI222_X1 U10835 ( .A1(n9870), .A2(n9650), .B1(n9649), .B2(n9867), .C1(n9648), .C2(n9865), .ZN(n9730) );
  NOR2_X1 U10836 ( .A1(n9730), .A2(n4399), .ZN(n9651) );
  AOI211_X1 U10837 ( .C1(n9727), .C2(n9884), .A(n9652), .B(n9651), .ZN(n9653)
         );
  OAI21_X1 U10838 ( .B1(n9731), .B2(n9672), .A(n9653), .ZN(P1_U3271) );
  XNOR2_X1 U10839 ( .A(n4474), .B(n9664), .ZN(n9736) );
  INV_X1 U10840 ( .A(n9654), .ZN(n9656) );
  AOI21_X1 U10841 ( .B1(n9732), .B2(n9656), .A(n9655), .ZN(n9733) );
  INV_X1 U10842 ( .A(n9657), .ZN(n9658) );
  AOI22_X1 U10843 ( .A1(n4399), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9658), .B2(
        n9872), .ZN(n9659) );
  OAI21_X1 U10844 ( .B1(n9661), .B2(n9660), .A(n9659), .ZN(n9669) );
  OAI21_X1 U10845 ( .B1(n9664), .B2(n9663), .A(n9662), .ZN(n9667) );
  AOI222_X1 U10846 ( .A1(n9870), .A2(n9667), .B1(n9666), .B2(n9867), .C1(n9665), .C2(n9865), .ZN(n9735) );
  NOR2_X1 U10847 ( .A1(n9735), .A2(n4399), .ZN(n9668) );
  AOI211_X1 U10848 ( .C1(n9733), .C2(n9670), .A(n9669), .B(n9668), .ZN(n9671)
         );
  OAI21_X1 U10849 ( .B1(n9736), .B2(n9672), .A(n9671), .ZN(P1_U3272) );
  NAND2_X1 U10850 ( .A1(n9192), .A2(n9766), .ZN(n9673) );
  OAI211_X1 U10851 ( .C1(n9674), .C2(n10101), .A(n9673), .B(n9677), .ZN(n9771)
         );
  MUX2_X1 U10852 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9771), .S(n10117), .Z(
        P1_U3554) );
  NAND3_X1 U10853 ( .A1(n9676), .A2(n9881), .A3(n9675), .ZN(n9678) );
  OAI211_X1 U10854 ( .C1(n9679), .C2(n10093), .A(n9678), .B(n9677), .ZN(n9772)
         );
  MUX2_X1 U10855 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9772), .S(n10117), .Z(
        P1_U3553) );
  AOI21_X1 U10856 ( .B1(n9766), .B2(n9682), .A(n9681), .ZN(n9683) );
  AND2_X1 U10857 ( .A1(n9684), .A2(n9683), .ZN(n9685) );
  AOI21_X1 U10858 ( .B1(n9766), .B2(n9688), .A(n9687), .ZN(n9689) );
  OAI211_X1 U10859 ( .C1(n9691), .C2(n9822), .A(n9690), .B(n9689), .ZN(n9774)
         );
  MUX2_X1 U10860 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9774), .S(n10117), .Z(
        P1_U3551) );
  AOI22_X1 U10861 ( .A1(n9693), .A2(n9881), .B1(n9766), .B2(n9692), .ZN(n9694)
         );
  OAI211_X1 U10862 ( .C1(n9696), .C2(n9822), .A(n9695), .B(n9694), .ZN(n9775)
         );
  MUX2_X1 U10863 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9775), .S(n10117), .Z(
        P1_U3550) );
  AOI21_X1 U10864 ( .B1(n9766), .B2(n9698), .A(n9697), .ZN(n9699) );
  OAI211_X1 U10865 ( .C1(n9701), .C2(n9822), .A(n9700), .B(n9699), .ZN(n9776)
         );
  MUX2_X1 U10866 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9776), .S(n10117), .Z(
        P1_U3549) );
  AOI21_X1 U10867 ( .B1(n9766), .B2(n9703), .A(n9702), .ZN(n9704) );
  OAI211_X1 U10868 ( .C1(n9706), .C2(n9822), .A(n9705), .B(n9704), .ZN(n9777)
         );
  MUX2_X1 U10869 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9777), .S(n10117), .Z(
        P1_U3548) );
  AOI211_X1 U10870 ( .C1(n9766), .C2(n9709), .A(n9708), .B(n9707), .ZN(n9710)
         );
  OAI21_X1 U10871 ( .B1(n9711), .B2(n9822), .A(n9710), .ZN(n9778) );
  MUX2_X1 U10872 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9778), .S(n10117), .Z(
        P1_U3547) );
  AOI211_X1 U10873 ( .C1(n9766), .C2(n9714), .A(n9713), .B(n9712), .ZN(n9715)
         );
  OAI21_X1 U10874 ( .B1(n9716), .B2(n9822), .A(n9715), .ZN(n9779) );
  MUX2_X1 U10875 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9779), .S(n10117), .Z(
        P1_U3546) );
  AOI22_X1 U10876 ( .A1(n9718), .A2(n9881), .B1(n9766), .B2(n9717), .ZN(n9719)
         );
  OAI211_X1 U10877 ( .C1(n9721), .C2(n9822), .A(n9720), .B(n9719), .ZN(n9780)
         );
  MUX2_X1 U10878 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9780), .S(n10117), .Z(
        P1_U3545) );
  AOI21_X1 U10879 ( .B1(n9766), .B2(n9723), .A(n9722), .ZN(n9724) );
  OAI211_X1 U10880 ( .C1(n9726), .C2(n9822), .A(n9725), .B(n9724), .ZN(n9781)
         );
  MUX2_X1 U10881 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9781), .S(n10117), .Z(
        P1_U3544) );
  AOI21_X1 U10882 ( .B1(n9766), .B2(n9728), .A(n9727), .ZN(n9729) );
  OAI211_X1 U10883 ( .C1(n9731), .C2(n9822), .A(n9730), .B(n9729), .ZN(n9782)
         );
  MUX2_X1 U10884 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9782), .S(n10117), .Z(
        P1_U3543) );
  AOI22_X1 U10885 ( .A1(n9733), .A2(n9881), .B1(n9766), .B2(n9732), .ZN(n9734)
         );
  OAI211_X1 U10886 ( .C1(n9736), .C2(n9822), .A(n9735), .B(n9734), .ZN(n9783)
         );
  MUX2_X1 U10887 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9783), .S(n10117), .Z(
        P1_U3542) );
  OAI21_X1 U10888 ( .B1(n9738), .B2(n10093), .A(n9737), .ZN(n9739) );
  NOR2_X1 U10889 ( .A1(n9740), .A2(n9739), .ZN(n9741) );
  OAI21_X1 U10890 ( .B1(n9742), .B2(n9822), .A(n9741), .ZN(n9784) );
  MUX2_X1 U10891 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9784), .S(n10117), .Z(
        P1_U3541) );
  AOI211_X1 U10892 ( .C1(n9766), .C2(n9745), .A(n9744), .B(n9743), .ZN(n9746)
         );
  OAI21_X1 U10893 ( .B1(n9747), .B2(n9822), .A(n9746), .ZN(n9785) );
  MUX2_X1 U10894 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9785), .S(n10117), .Z(
        P1_U3540) );
  AOI211_X1 U10895 ( .C1(n9766), .C2(n9750), .A(n9749), .B(n9748), .ZN(n9751)
         );
  OAI21_X1 U10896 ( .B1(n9752), .B2(n9822), .A(n9751), .ZN(n9786) );
  MUX2_X1 U10897 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9786), .S(n10117), .Z(
        P1_U3539) );
  INV_X1 U10898 ( .A(n9753), .ZN(n9758) );
  AOI22_X1 U10899 ( .A1(n9755), .A2(n9881), .B1(n9766), .B2(n9754), .ZN(n9756)
         );
  OAI211_X1 U10900 ( .C1(n9758), .C2(n10065), .A(n9757), .B(n9756), .ZN(n9787)
         );
  MUX2_X1 U10901 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9787), .S(n10117), .Z(
        P1_U3538) );
  AOI22_X1 U10902 ( .A1(n9760), .A2(n9881), .B1(n9766), .B2(n9759), .ZN(n9761)
         );
  OAI211_X1 U10903 ( .C1(n9763), .C2(n9822), .A(n9762), .B(n9761), .ZN(n9788)
         );
  MUX2_X1 U10904 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9788), .S(n10117), .Z(
        P1_U3536) );
  INV_X1 U10905 ( .A(n9764), .ZN(n9770) );
  AOI22_X1 U10906 ( .A1(n9767), .A2(n9881), .B1(n9766), .B2(n9765), .ZN(n9768)
         );
  OAI211_X1 U10907 ( .C1(n9770), .C2(n10065), .A(n9769), .B(n9768), .ZN(n9789)
         );
  MUX2_X1 U10908 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9789), .S(n10117), .Z(
        P1_U3534) );
  MUX2_X1 U10909 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9771), .S(n10107), .Z(
        P1_U3522) );
  MUX2_X1 U10910 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9772), .S(n10107), .Z(
        P1_U3521) );
  MUX2_X1 U10911 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9774), .S(n10107), .Z(
        P1_U3519) );
  MUX2_X1 U10912 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9775), .S(n10107), .Z(
        P1_U3518) );
  MUX2_X1 U10913 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9776), .S(n10107), .Z(
        P1_U3517) );
  MUX2_X1 U10914 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9777), .S(n10107), .Z(
        P1_U3516) );
  MUX2_X1 U10915 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9778), .S(n10107), .Z(
        P1_U3515) );
  MUX2_X1 U10916 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9779), .S(n10107), .Z(
        P1_U3514) );
  MUX2_X1 U10917 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9780), .S(n10107), .Z(
        P1_U3513) );
  MUX2_X1 U10918 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9781), .S(n10107), .Z(
        P1_U3512) );
  MUX2_X1 U10919 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9782), .S(n10107), .Z(
        P1_U3511) );
  MUX2_X1 U10920 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9783), .S(n10107), .Z(
        P1_U3510) );
  MUX2_X1 U10921 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9784), .S(n10107), .Z(
        P1_U3508) );
  MUX2_X1 U10922 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9785), .S(n10107), .Z(
        P1_U3505) );
  MUX2_X1 U10923 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9786), .S(n10107), .Z(
        P1_U3502) );
  MUX2_X1 U10924 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9787), .S(n10107), .Z(
        P1_U3499) );
  MUX2_X1 U10925 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9788), .S(n10107), .Z(
        P1_U3493) );
  MUX2_X1 U10926 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n9789), .S(n10107), .Z(
        P1_U3487) );
  NAND3_X1 U10927 ( .A1(n9790), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9792) );
  OAI22_X1 U10928 ( .A1(n9793), .A2(n9792), .B1(n6613), .B2(n9791), .ZN(n9794)
         );
  INV_X1 U10929 ( .A(n9794), .ZN(n9795) );
  OAI21_X1 U10930 ( .B1(n9797), .B2(n9796), .A(n9795), .ZN(P1_U3322) );
  MUX2_X1 U10931 ( .A(n9798), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10932 ( .A1(n10124), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n7777), .ZN(n9809) );
  NAND2_X1 U10933 ( .A1(n10129), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9801) );
  AOI211_X1 U10934 ( .C1(n9801), .C2(n9800), .A(n9799), .B(n10122), .ZN(n9802)
         );
  AOI21_X1 U10935 ( .B1(n9815), .B2(n9803), .A(n9802), .ZN(n9808) );
  NOR2_X1 U10936 ( .A1(n10127), .A2(n10205), .ZN(n9806) );
  OAI211_X1 U10937 ( .C1(n9806), .C2(n9805), .A(n10119), .B(n9804), .ZN(n9807)
         );
  NAND3_X1 U10938 ( .A1(n9809), .A2(n9808), .A3(n9807), .ZN(P2_U3246) );
  AOI22_X1 U10939 ( .A1(n10124), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9821) );
  AOI211_X1 U10940 ( .C1(n9812), .C2(n9811), .A(n9810), .B(n10122), .ZN(n9813)
         );
  AOI21_X1 U10941 ( .B1(n9815), .B2(n9814), .A(n9813), .ZN(n9820) );
  OAI211_X1 U10942 ( .C1(n9818), .C2(n9817), .A(n10119), .B(n9816), .ZN(n9819)
         );
  NAND3_X1 U10943 ( .A1(n9821), .A2(n9820), .A3(n9819), .ZN(P2_U3247) );
  INV_X1 U10944 ( .A(n9822), .ZN(n10103) );
  OAI21_X1 U10945 ( .B1(n9824), .B2(n10093), .A(n9823), .ZN(n9825) );
  AOI211_X1 U10946 ( .C1(n9827), .C2(n10103), .A(n9826), .B(n9825), .ZN(n9830)
         );
  INV_X1 U10947 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9828) );
  AOI22_X1 U10948 ( .A1(n10107), .A2(n9830), .B1(n9828), .B2(n10105), .ZN(
        P1_U3484) );
  AOI22_X1 U10949 ( .A1(n10117), .A2(n9830), .B1(n9829), .B2(n4906), .ZN(
        P1_U3533) );
  INV_X1 U10950 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10257) );
  NOR2_X1 U10951 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9831) );
  AOI21_X1 U10952 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9831), .ZN(n10225) );
  NOR2_X1 U10953 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9832) );
  AOI21_X1 U10954 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9832), .ZN(n10228) );
  NOR2_X1 U10955 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9833) );
  AOI21_X1 U10956 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9833), .ZN(n10231) );
  NOR2_X1 U10957 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9834) );
  AOI21_X1 U10958 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9834), .ZN(n10234) );
  NOR2_X1 U10959 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9835) );
  AOI21_X1 U10960 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9835), .ZN(n10237) );
  NOR2_X1 U10961 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9842) );
  XNOR2_X1 U10962 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10265) );
  NAND2_X1 U10963 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9840) );
  XOR2_X1 U10964 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10263) );
  NAND2_X1 U10965 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9838) );
  XOR2_X1 U10966 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10260) );
  AOI21_X1 U10967 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10218) );
  INV_X1 U10968 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9836) );
  NAND3_X1 U10969 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10220) );
  OAI21_X1 U10970 ( .B1(n10218), .B2(n9836), .A(n10220), .ZN(n10259) );
  NAND2_X1 U10971 ( .A1(n10260), .A2(n10259), .ZN(n9837) );
  NAND2_X1 U10972 ( .A1(n9838), .A2(n9837), .ZN(n10262) );
  NAND2_X1 U10973 ( .A1(n10263), .A2(n10262), .ZN(n9839) );
  NAND2_X1 U10974 ( .A1(n9840), .A2(n9839), .ZN(n10264) );
  NOR2_X1 U10975 ( .A1(n10265), .A2(n10264), .ZN(n9841) );
  NOR2_X1 U10976 ( .A1(n9842), .A2(n9841), .ZN(n9843) );
  NOR2_X1 U10977 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9843), .ZN(n10253) );
  AND2_X1 U10978 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9843), .ZN(n10252) );
  NOR2_X1 U10979 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10252), .ZN(n9844) );
  NOR2_X1 U10980 ( .A1(n10253), .A2(n9844), .ZN(n9845) );
  NAND2_X1 U10981 ( .A1(n9845), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9847) );
  XOR2_X1 U10982 ( .A(n9845), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10251) );
  NAND2_X1 U10983 ( .A1(n10251), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9846) );
  NAND2_X1 U10984 ( .A1(n9847), .A2(n9846), .ZN(n9848) );
  NAND2_X1 U10985 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9848), .ZN(n9850) );
  XOR2_X1 U10986 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9848), .Z(n10247) );
  NAND2_X1 U10987 ( .A1(n10247), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n9849) );
  NAND2_X1 U10988 ( .A1(n9850), .A2(n9849), .ZN(n9851) );
  NAND2_X1 U10989 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9851), .ZN(n9853) );
  XOR2_X1 U10990 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9851), .Z(n10261) );
  NAND2_X1 U10991 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10261), .ZN(n9852) );
  NAND2_X1 U10992 ( .A1(n9853), .A2(n9852), .ZN(n9854) );
  AND2_X1 U10993 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9854), .ZN(n9855) );
  XNOR2_X1 U10994 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9854), .ZN(n10250) );
  INV_X1 U10995 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10249) );
  NOR2_X1 U10996 ( .A1(n10250), .A2(n10249), .ZN(n10248) );
  NOR2_X1 U10997 ( .A1(n9855), .A2(n10248), .ZN(n10246) );
  NAND2_X1 U10998 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9856) );
  OAI21_X1 U10999 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9856), .ZN(n10245) );
  NOR2_X1 U11000 ( .A1(n10246), .A2(n10245), .ZN(n10244) );
  AOI21_X1 U11001 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10244), .ZN(n10243) );
  NAND2_X1 U11002 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9857) );
  OAI21_X1 U11003 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9857), .ZN(n10242) );
  NOR2_X1 U11004 ( .A1(n10243), .A2(n10242), .ZN(n10241) );
  AOI21_X1 U11005 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10241), .ZN(n10240) );
  NOR2_X1 U11006 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9858) );
  AOI21_X1 U11007 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9858), .ZN(n10239) );
  NAND2_X1 U11008 ( .A1(n10240), .A2(n10239), .ZN(n10238) );
  OAI21_X1 U11009 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10238), .ZN(n10236) );
  NAND2_X1 U11010 ( .A1(n10237), .A2(n10236), .ZN(n10235) );
  OAI21_X1 U11011 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10235), .ZN(n10233) );
  NAND2_X1 U11012 ( .A1(n10234), .A2(n10233), .ZN(n10232) );
  OAI21_X1 U11013 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10232), .ZN(n10230) );
  NAND2_X1 U11014 ( .A1(n10231), .A2(n10230), .ZN(n10229) );
  OAI21_X1 U11015 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10229), .ZN(n10227) );
  NAND2_X1 U11016 ( .A1(n10228), .A2(n10227), .ZN(n10226) );
  OAI21_X1 U11017 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10226), .ZN(n10224) );
  NAND2_X1 U11018 ( .A1(n10225), .A2(n10224), .ZN(n10223) );
  OAI21_X1 U11019 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10223), .ZN(n10256) );
  NOR2_X1 U11020 ( .A1(n10257), .A2(n10256), .ZN(n9859) );
  NAND2_X1 U11021 ( .A1(n10257), .A2(n10256), .ZN(n10255) );
  OAI21_X1 U11022 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9859), .A(n10255), .ZN(
        n9861) );
  XOR2_X1 U11023 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n9860) );
  XNOR2_X1 U11024 ( .A(n9861), .B(n9860), .ZN(ADD_1071_U4) );
  NAND2_X1 U11025 ( .A1(n9863), .A2(n9862), .ZN(n9864) );
  XOR2_X1 U11026 ( .A(n9879), .B(n9864), .Z(n9869) );
  AOI222_X1 U11027 ( .A1(n9870), .A2(n9869), .B1(n9868), .B2(n9867), .C1(n9866), .C2(n9865), .ZN(n9895) );
  INV_X1 U11028 ( .A(n9871), .ZN(n9873) );
  AOI222_X1 U11029 ( .A1(n9875), .A2(n9874), .B1(n9873), .B2(n9872), .C1(
        P1_REG2_REG_12__SCAN_IN), .C2(n4399), .ZN(n9887) );
  INV_X1 U11030 ( .A(n9876), .ZN(n9877) );
  AOI21_X1 U11031 ( .B1(n9879), .B2(n9878), .A(n9877), .ZN(n9898) );
  OAI211_X1 U11032 ( .C1(n9882), .C2(n9896), .A(n9881), .B(n9880), .ZN(n9894)
         );
  INV_X1 U11033 ( .A(n9894), .ZN(n9883) );
  AOI22_X1 U11034 ( .A1(n9898), .A2(n9885), .B1(n9884), .B2(n9883), .ZN(n9886)
         );
  OAI211_X1 U11035 ( .C1(n4399), .C2(n9895), .A(n9887), .B(n9886), .ZN(
        P1_U3279) );
  OAI21_X1 U11036 ( .B1(n9889), .B2(n10093), .A(n9888), .ZN(n9890) );
  AOI211_X1 U11037 ( .C1(n9892), .C2(n10103), .A(n9891), .B(n9890), .ZN(n9899)
         );
  AOI22_X1 U11038 ( .A1(n10117), .A2(n9899), .B1(n9893), .B2(n4906), .ZN(
        P1_U3537) );
  OAI211_X1 U11039 ( .C1(n9896), .C2(n10093), .A(n9895), .B(n9894), .ZN(n9897)
         );
  AOI21_X1 U11040 ( .B1(n9898), .B2(n10103), .A(n9897), .ZN(n9901) );
  AOI22_X1 U11041 ( .A1(n10117), .A2(n9901), .B1(n9479), .B2(n4906), .ZN(
        P1_U3535) );
  AOI22_X1 U11042 ( .A1(n10107), .A2(n9899), .B1(n7572), .B2(n10105), .ZN(
        P1_U3496) );
  INV_X1 U11043 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9900) );
  AOI22_X1 U11044 ( .A1(n10107), .A2(n9901), .B1(n9900), .B2(n10105), .ZN(
        P1_U3490) );
  XNOR2_X1 U11045 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11046 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U11047 ( .B1(n9904), .B2(n9903), .A(n9902), .ZN(n9905) );
  AOI22_X1 U11048 ( .A1(n9905), .A2(n10007), .B1(n9907), .B2(n10026), .ZN(
        n9917) );
  INV_X1 U11049 ( .A(n9906), .ZN(n9910) );
  MUX2_X1 U11050 ( .A(n9908), .B(P1_REG1_REG_4__SCAN_IN), .S(n9907), .Z(n9909)
         );
  NAND2_X1 U11051 ( .A1(n9910), .A2(n9909), .ZN(n9911) );
  AOI21_X1 U11052 ( .B1(n9912), .B2(n9911), .A(n10032), .ZN(n9913) );
  AOI211_X1 U11053 ( .C1(P1_ADDR_REG_4__SCAN_IN), .C2(n9930), .A(n9914), .B(
        n9913), .ZN(n9916) );
  NAND3_X1 U11054 ( .A1(n9917), .A2(n9916), .A3(n9915), .ZN(P1_U3245) );
  AOI22_X1 U11055 ( .A1(n9930), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n9918), .B2(
        n10026), .ZN(n9928) );
  XNOR2_X1 U11056 ( .A(n9920), .B(n9919), .ZN(n9921) );
  NAND2_X1 U11057 ( .A1(n10007), .A2(n9921), .ZN(n9926) );
  OAI211_X1 U11058 ( .C1(n9924), .C2(n9923), .A(n10012), .B(n9922), .ZN(n9925)
         );
  NAND4_X1 U11059 ( .A1(n9928), .A2(n9927), .A3(n9926), .A4(n9925), .ZN(
        P1_U3246) );
  AOI22_X1 U11060 ( .A1(n9930), .A2(P1_ADDR_REG_8__SCAN_IN), .B1(n9929), .B2(
        n10026), .ZN(n9941) );
  OAI21_X1 U11061 ( .B1(n9933), .B2(n9932), .A(n9931), .ZN(n9934) );
  NAND2_X1 U11062 ( .A1(n9934), .A2(n10007), .ZN(n9939) );
  OAI211_X1 U11063 ( .C1(n9937), .C2(n9936), .A(n10012), .B(n9935), .ZN(n9938)
         );
  NAND4_X1 U11064 ( .A1(n9941), .A2(n9940), .A3(n9939), .A4(n9938), .ZN(
        P1_U3249) );
  INV_X1 U11065 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9954) );
  AOI211_X1 U11066 ( .C1(n9944), .C2(n9943), .A(n9942), .B(n10020), .ZN(n9945)
         );
  AOI211_X1 U11067 ( .C1(n10026), .C2(n9947), .A(n9946), .B(n9945), .ZN(n9953)
         );
  AOI21_X1 U11068 ( .B1(n9950), .B2(n9949), .A(n9948), .ZN(n9951) );
  OR2_X1 U11069 ( .A1(n9951), .A2(n10032), .ZN(n9952) );
  OAI211_X1 U11070 ( .C1(n9954), .C2(n10035), .A(n9953), .B(n9952), .ZN(
        P1_U3253) );
  INV_X1 U11071 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9969) );
  AOI21_X1 U11072 ( .B1(n10026), .B2(n9956), .A(n9955), .ZN(n9962) );
  INV_X1 U11073 ( .A(n9957), .ZN(n9958) );
  OAI211_X1 U11074 ( .C1(n9960), .C2(n9959), .A(n10007), .B(n9958), .ZN(n9961)
         );
  AND2_X1 U11075 ( .A1(n9962), .A2(n9961), .ZN(n9968) );
  AOI21_X1 U11076 ( .B1(n9965), .B2(n9964), .A(n9963), .ZN(n9966) );
  OR2_X1 U11077 ( .A1(n10032), .A2(n9966), .ZN(n9967) );
  OAI211_X1 U11078 ( .C1(n9969), .C2(n10035), .A(n9968), .B(n9967), .ZN(
        P1_U3254) );
  AOI211_X1 U11079 ( .C1(n9971), .C2(n7590), .A(n9970), .B(n10020), .ZN(n9972)
         );
  AOI211_X1 U11080 ( .C1(n10026), .C2(n9974), .A(n9973), .B(n9972), .ZN(n9980)
         );
  AOI21_X1 U11081 ( .B1(n9977), .B2(n9976), .A(n9975), .ZN(n9978) );
  OR2_X1 U11082 ( .A1(n9978), .A2(n10032), .ZN(n9979) );
  OAI211_X1 U11083 ( .C1(n9981), .C2(n10035), .A(n9980), .B(n9979), .ZN(
        P1_U3255) );
  INV_X1 U11084 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9991) );
  AOI211_X1 U11085 ( .C1(n9983), .C2(n7767), .A(n9982), .B(n10020), .ZN(n9984)
         );
  AOI211_X1 U11086 ( .C1(n10026), .C2(n9986), .A(n9985), .B(n9984), .ZN(n9990)
         );
  OAI211_X1 U11087 ( .C1(n9988), .C2(P1_REG1_REG_15__SCAN_IN), .A(n10012), .B(
        n9987), .ZN(n9989) );
  OAI211_X1 U11088 ( .C1(n9991), .C2(n10035), .A(n9990), .B(n9989), .ZN(
        P1_U3256) );
  INV_X1 U11089 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10002) );
  AOI211_X1 U11090 ( .C1(n4442), .C2(n9993), .A(n9992), .B(n10020), .ZN(n9994)
         );
  AOI211_X1 U11091 ( .C1(n10026), .C2(n9996), .A(n9995), .B(n9994), .ZN(n10001) );
  OAI211_X1 U11092 ( .C1(n9999), .C2(n9998), .A(n10012), .B(n9997), .ZN(n10000) );
  OAI211_X1 U11093 ( .C1(n10002), .C2(n10035), .A(n10001), .B(n10000), .ZN(
        P1_U3257) );
  AOI21_X1 U11094 ( .B1(n10005), .B2(n10004), .A(n10003), .ZN(n10006) );
  NAND2_X1 U11095 ( .A1(n10007), .A2(n10006), .ZN(n10011) );
  NAND2_X1 U11096 ( .A1(n10026), .A2(n10008), .ZN(n10010) );
  AND3_X1 U11097 ( .A1(n10011), .A2(n10010), .A3(n10009), .ZN(n10017) );
  OAI211_X1 U11098 ( .C1(n10015), .C2(n10014), .A(n10013), .B(n10012), .ZN(
        n10016) );
  OAI211_X1 U11099 ( .C1(n10018), .C2(n10035), .A(n10017), .B(n10016), .ZN(
        P1_U3258) );
  INV_X1 U11100 ( .A(n10019), .ZN(n10025) );
  AOI211_X1 U11101 ( .C1(n10023), .C2(n10022), .A(n10021), .B(n10020), .ZN(
        n10024) );
  AOI211_X1 U11102 ( .C1(n10027), .C2(n10026), .A(n10025), .B(n10024), .ZN(
        n10034) );
  AOI21_X1 U11103 ( .B1(n10030), .B2(n10029), .A(n10028), .ZN(n10031) );
  OR2_X1 U11104 ( .A1(n10032), .A2(n10031), .ZN(n10033) );
  OAI211_X1 U11105 ( .C1(n10036), .C2(n10035), .A(n10034), .B(n10033), .ZN(
        P1_U3259) );
  INV_X1 U11106 ( .A(n10037), .ZN(n10041) );
  NOR2_X1 U11107 ( .A1(n10038), .A2(n6100), .ZN(n10040) );
  MUX2_X1 U11108 ( .A(n10041), .B(n10040), .S(n10039), .Z(n10048) );
  OAI22_X1 U11109 ( .A1(n10045), .A2(n10044), .B1(n10043), .B2(n10042), .ZN(
        n10046) );
  NOR3_X1 U11110 ( .A1(n10048), .A2(n10047), .A3(n10046), .ZN(n10049) );
  AOI22_X1 U11111 ( .A1(n4399), .A2(n5939), .B1(n10049), .B2(n9610), .ZN(
        P1_U3290) );
  AND2_X1 U11112 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10058), .ZN(P1_U3292) );
  AND2_X1 U11113 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10058), .ZN(P1_U3293) );
  AND2_X1 U11114 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10058), .ZN(P1_U3294) );
  AND2_X1 U11115 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10058), .ZN(P1_U3295) );
  AND2_X1 U11116 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10058), .ZN(P1_U3296) );
  AND2_X1 U11117 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10058), .ZN(P1_U3297) );
  AND2_X1 U11118 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10058), .ZN(P1_U3298) );
  NOR2_X1 U11119 ( .A1(n10057), .A2(n10050), .ZN(P1_U3299) );
  AND2_X1 U11120 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10058), .ZN(P1_U3300) );
  NOR2_X1 U11121 ( .A1(n10057), .A2(n10051), .ZN(P1_U3301) );
  AND2_X1 U11122 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10058), .ZN(P1_U3302) );
  AND2_X1 U11123 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10058), .ZN(P1_U3303) );
  NOR2_X1 U11124 ( .A1(n10057), .A2(n10052), .ZN(P1_U3304) );
  AND2_X1 U11125 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10058), .ZN(P1_U3305) );
  AND2_X1 U11126 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10058), .ZN(P1_U3306) );
  AND2_X1 U11127 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10058), .ZN(P1_U3307) );
  AND2_X1 U11128 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10058), .ZN(P1_U3308) );
  AND2_X1 U11129 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10058), .ZN(P1_U3309) );
  AND2_X1 U11130 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10058), .ZN(P1_U3310) );
  NOR2_X1 U11131 ( .A1(n10057), .A2(n10053), .ZN(P1_U3311) );
  AND2_X1 U11132 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10058), .ZN(P1_U3312) );
  AND2_X1 U11133 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10058), .ZN(P1_U3313) );
  NOR2_X1 U11134 ( .A1(n10057), .A2(n10054), .ZN(P1_U3314) );
  AND2_X1 U11135 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10058), .ZN(P1_U3315) );
  NOR2_X1 U11136 ( .A1(n10057), .A2(n10055), .ZN(P1_U3316) );
  AND2_X1 U11137 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10058), .ZN(P1_U3317) );
  AND2_X1 U11138 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10058), .ZN(P1_U3318) );
  NOR2_X1 U11139 ( .A1(n10057), .A2(n10056), .ZN(P1_U3319) );
  AND2_X1 U11140 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10058), .ZN(P1_U3320) );
  AND2_X1 U11141 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10058), .ZN(P1_U3321) );
  AOI22_X1 U11142 ( .A1(n10107), .A2(n10059), .B1(n5937), .B2(n10105), .ZN(
        P1_U3457) );
  OAI21_X1 U11143 ( .B1(n10061), .B2(n10101), .A(n10060), .ZN(n10063) );
  AOI211_X1 U11144 ( .C1(n10103), .C2(n10064), .A(n10063), .B(n10062), .ZN(
        n10108) );
  AOI22_X1 U11145 ( .A1(n10107), .A2(n10108), .B1(n5979), .B2(n10105), .ZN(
        P1_U3460) );
  INV_X1 U11146 ( .A(n10065), .ZN(n10077) );
  OAI22_X1 U11147 ( .A1(n10067), .A2(n10101), .B1(n10066), .B2(n10093), .ZN(
        n10069) );
  AOI211_X1 U11148 ( .C1(n10077), .C2(n10070), .A(n10069), .B(n10068), .ZN(
        n10109) );
  AOI22_X1 U11149 ( .A1(n10107), .A2(n10109), .B1(n5997), .B2(n10105), .ZN(
        P1_U3463) );
  INV_X1 U11150 ( .A(n10071), .ZN(n10076) );
  OAI22_X1 U11151 ( .A1(n10073), .A2(n10101), .B1(n10072), .B2(n10093), .ZN(
        n10075) );
  AOI211_X1 U11152 ( .C1(n10077), .C2(n10076), .A(n10075), .B(n10074), .ZN(
        n10110) );
  AOI22_X1 U11153 ( .A1(n10107), .A2(n10110), .B1(n6015), .B2(n10105), .ZN(
        P1_U3466) );
  NAND2_X1 U11154 ( .A1(n10079), .A2(n10078), .ZN(n10080) );
  AOI21_X1 U11155 ( .B1(n10081), .B2(n10103), .A(n10080), .ZN(n10083) );
  AND2_X1 U11156 ( .A1(n10083), .A2(n10082), .ZN(n10112) );
  AOI22_X1 U11157 ( .A1(n10107), .A2(n10112), .B1(n6032), .B2(n10105), .ZN(
        P1_U3469) );
  INV_X1 U11158 ( .A(n10084), .ZN(n10085) );
  OAI211_X1 U11159 ( .C1(n10101), .C2(n10087), .A(n10086), .B(n10085), .ZN(
        n10088) );
  AOI21_X1 U11160 ( .B1(n10103), .B2(n10089), .A(n10088), .ZN(n10113) );
  INV_X1 U11161 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10090) );
  AOI22_X1 U11162 ( .A1(n10107), .A2(n10113), .B1(n10090), .B2(n10105), .ZN(
        P1_U3472) );
  OAI211_X1 U11163 ( .C1(n10094), .C2(n10093), .A(n10092), .B(n10091), .ZN(
        n10095) );
  AOI21_X1 U11164 ( .B1(n10096), .B2(n10103), .A(n10095), .ZN(n10115) );
  AOI22_X1 U11165 ( .A1(n10107), .A2(n10115), .B1(n10097), .B2(n10105), .ZN(
        P1_U3475) );
  OAI211_X1 U11166 ( .C1(n10101), .C2(n10100), .A(n10099), .B(n10098), .ZN(
        n10102) );
  AOI21_X1 U11167 ( .B1(n10104), .B2(n10103), .A(n10102), .ZN(n10116) );
  INV_X1 U11168 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10106) );
  AOI22_X1 U11169 ( .A1(n10107), .A2(n10116), .B1(n10106), .B2(n10105), .ZN(
        P1_U3478) );
  AOI22_X1 U11170 ( .A1(n10117), .A2(n10108), .B1(n6260), .B2(n4906), .ZN(
        P1_U3525) );
  AOI22_X1 U11171 ( .A1(n10117), .A2(n10109), .B1(n6261), .B2(n4906), .ZN(
        P1_U3526) );
  AOI22_X1 U11172 ( .A1(n10117), .A2(n10110), .B1(n9908), .B2(n4906), .ZN(
        P1_U3527) );
  AOI22_X1 U11173 ( .A1(n10117), .A2(n10112), .B1(n10111), .B2(n4906), .ZN(
        P1_U3528) );
  AOI22_X1 U11174 ( .A1(n10117), .A2(n10113), .B1(n6053), .B2(n4906), .ZN(
        P1_U3529) );
  AOI22_X1 U11175 ( .A1(n10117), .A2(n10115), .B1(n10114), .B2(n4906), .ZN(
        P1_U3530) );
  AOI22_X1 U11176 ( .A1(n10117), .A2(n10116), .B1(n6662), .B2(n4906), .ZN(
        P1_U3531) );
  AOI22_X1 U11177 ( .A1(n10118), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10119), .ZN(n10128) );
  NAND2_X1 U11178 ( .A1(n10119), .A2(n10205), .ZN(n10120) );
  OAI211_X1 U11179 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n10122), .A(n10121), .B(
        n10120), .ZN(n10123) );
  INV_X1 U11180 ( .A(n10123), .ZN(n10126) );
  AOI22_X1 U11181 ( .A1(n10124), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10125) );
  OAI221_X1 U11182 ( .B1(n10129), .B2(n10128), .C1(n10127), .C2(n10126), .A(
        n10125), .ZN(P2_U3245) );
  NOR2_X1 U11183 ( .A1(n10131), .A2(n10130), .ZN(n10138) );
  AND2_X1 U11184 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10141), .ZN(P2_U3297) );
  AND2_X1 U11185 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10141), .ZN(P2_U3298) );
  NOR2_X1 U11186 ( .A1(n10138), .A2(n10132), .ZN(P2_U3299) );
  AND2_X1 U11187 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10141), .ZN(P2_U3300) );
  NOR2_X1 U11188 ( .A1(n10138), .A2(n10133), .ZN(P2_U3301) );
  AND2_X1 U11189 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10141), .ZN(P2_U3302) );
  AND2_X1 U11190 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10141), .ZN(P2_U3303) );
  AND2_X1 U11191 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10141), .ZN(P2_U3304) );
  AND2_X1 U11192 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10141), .ZN(P2_U3305) );
  AND2_X1 U11193 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10141), .ZN(P2_U3306) );
  AND2_X1 U11194 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10141), .ZN(P2_U3307) );
  NOR2_X1 U11195 ( .A1(n10138), .A2(n10134), .ZN(P2_U3308) );
  NOR2_X1 U11196 ( .A1(n10138), .A2(n10135), .ZN(P2_U3309) );
  AND2_X1 U11197 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10141), .ZN(P2_U3310) );
  AND2_X1 U11198 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10141), .ZN(P2_U3311) );
  AND2_X1 U11199 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10141), .ZN(P2_U3312) );
  NOR2_X1 U11200 ( .A1(n10138), .A2(n10136), .ZN(P2_U3313) );
  AND2_X1 U11201 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10141), .ZN(P2_U3314) );
  AND2_X1 U11202 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10141), .ZN(P2_U3315) );
  NOR2_X1 U11203 ( .A1(n10138), .A2(n10137), .ZN(P2_U3316) );
  AND2_X1 U11204 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10141), .ZN(P2_U3317) );
  AND2_X1 U11205 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10141), .ZN(P2_U3318) );
  AND2_X1 U11206 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10141), .ZN(P2_U3319) );
  AND2_X1 U11207 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10141), .ZN(P2_U3320) );
  AND2_X1 U11208 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10141), .ZN(P2_U3321) );
  AND2_X1 U11209 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10141), .ZN(P2_U3322) );
  AND2_X1 U11210 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10141), .ZN(P2_U3323) );
  AND2_X1 U11211 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10141), .ZN(P2_U3324) );
  AND2_X1 U11212 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10141), .ZN(P2_U3325) );
  AND2_X1 U11213 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10141), .ZN(P2_U3326) );
  AOI22_X1 U11214 ( .A1(n10140), .A2(n10141), .B1(n10144), .B2(n10139), .ZN(
        P2_U3437) );
  AOI22_X1 U11215 ( .A1(n10144), .A2(n10143), .B1(n10142), .B2(n10141), .ZN(
        P2_U3438) );
  AOI22_X1 U11216 ( .A1(n10147), .A2(n10177), .B1(n10146), .B2(n10145), .ZN(
        n10148) );
  AND2_X1 U11217 ( .A1(n10149), .A2(n10148), .ZN(n10206) );
  AOI22_X1 U11218 ( .A1(n10204), .A2(n10206), .B1(n5198), .B2(n10202), .ZN(
        P2_U3451) );
  OAI22_X1 U11219 ( .A1(n10151), .A2(n10187), .B1(n10150), .B2(n10186), .ZN(
        n10153) );
  AOI211_X1 U11220 ( .C1(n10177), .C2(n10154), .A(n10153), .B(n10152), .ZN(
        n10207) );
  INV_X1 U11221 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U11222 ( .A1(n10204), .A2(n10207), .B1(n10155), .B2(n10202), .ZN(
        P2_U3454) );
  OAI22_X1 U11223 ( .A1(n10157), .A2(n10187), .B1(n10156), .B2(n10186), .ZN(
        n10159) );
  AOI211_X1 U11224 ( .C1(n10177), .C2(n10160), .A(n10159), .B(n10158), .ZN(
        n10208) );
  AOI22_X1 U11225 ( .A1(n10204), .A2(n10208), .B1(n10161), .B2(n10202), .ZN(
        P2_U3457) );
  OAI22_X1 U11226 ( .A1(n10163), .A2(n10187), .B1(n10162), .B2(n10186), .ZN(
        n10165) );
  AOI211_X1 U11227 ( .C1(n10177), .C2(n10166), .A(n10165), .B(n10164), .ZN(
        n10209) );
  AOI22_X1 U11228 ( .A1(n10204), .A2(n10209), .B1(n5152), .B2(n10202), .ZN(
        P2_U3463) );
  OAI211_X1 U11229 ( .C1(n10169), .C2(n10186), .A(n10168), .B(n10167), .ZN(
        n10170) );
  AOI21_X1 U11230 ( .B1(n10177), .B2(n10171), .A(n10170), .ZN(n10210) );
  AOI22_X1 U11231 ( .A1(n10204), .A2(n10210), .B1(n5142), .B2(n10202), .ZN(
        P2_U3466) );
  OAI22_X1 U11232 ( .A1(n10173), .A2(n10187), .B1(n10172), .B2(n10186), .ZN(
        n10175) );
  AOI211_X1 U11233 ( .C1(n10177), .C2(n10176), .A(n10175), .B(n10174), .ZN(
        n10211) );
  AOI22_X1 U11234 ( .A1(n10204), .A2(n10211), .B1(n5185), .B2(n10202), .ZN(
        P2_U3469) );
  INV_X1 U11235 ( .A(n10178), .ZN(n10183) );
  OAI22_X1 U11236 ( .A1(n10180), .A2(n10187), .B1(n10179), .B2(n10186), .ZN(
        n10182) );
  AOI211_X1 U11237 ( .C1(n10192), .C2(n10183), .A(n10182), .B(n10181), .ZN(
        n10212) );
  AOI22_X1 U11238 ( .A1(n10204), .A2(n10212), .B1(n5266), .B2(n10202), .ZN(
        P2_U3475) );
  INV_X1 U11239 ( .A(n10184), .ZN(n10191) );
  OAI22_X1 U11240 ( .A1(n10188), .A2(n10187), .B1(n4655), .B2(n10186), .ZN(
        n10190) );
  AOI211_X1 U11241 ( .C1(n10192), .C2(n10191), .A(n10190), .B(n10189), .ZN(
        n10214) );
  AOI22_X1 U11242 ( .A1(n10204), .A2(n10214), .B1(n5307), .B2(n10202), .ZN(
        P2_U3481) );
  AOI22_X1 U11243 ( .A1(n10196), .A2(n10195), .B1(n10194), .B2(n10193), .ZN(
        n10197) );
  OAI211_X1 U11244 ( .C1(n10200), .C2(n10199), .A(n10198), .B(n10197), .ZN(
        n10201) );
  INV_X1 U11245 ( .A(n10201), .ZN(n10216) );
  INV_X1 U11246 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U11247 ( .A1(n10204), .A2(n10216), .B1(n10203), .B2(n10202), .ZN(
        P2_U3487) );
  AOI22_X1 U11248 ( .A1(n10217), .A2(n10206), .B1(n10205), .B2(n10215), .ZN(
        P2_U3520) );
  AOI22_X1 U11249 ( .A1(n10217), .A2(n10207), .B1(n6718), .B2(n10215), .ZN(
        P2_U3521) );
  AOI22_X1 U11250 ( .A1(n10217), .A2(n10208), .B1(n6717), .B2(n10215), .ZN(
        P2_U3522) );
  AOI22_X1 U11251 ( .A1(n10217), .A2(n10209), .B1(n6715), .B2(n10215), .ZN(
        P2_U3524) );
  AOI22_X1 U11252 ( .A1(n10217), .A2(n10210), .B1(n6714), .B2(n10215), .ZN(
        P2_U3525) );
  AOI22_X1 U11253 ( .A1(n10217), .A2(n10211), .B1(n6713), .B2(n10215), .ZN(
        P2_U3526) );
  AOI22_X1 U11254 ( .A1(n10217), .A2(n10212), .B1(n6711), .B2(n10215), .ZN(
        P2_U3528) );
  AOI22_X1 U11255 ( .A1(n10217), .A2(n10214), .B1(n10213), .B2(n10215), .ZN(
        P2_U3530) );
  AOI22_X1 U11256 ( .A1(n10217), .A2(n10216), .B1(n6924), .B2(n10215), .ZN(
        P2_U3532) );
  INV_X1 U11257 ( .A(n10218), .ZN(n10219) );
  NAND2_X1 U11258 ( .A1(n10220), .A2(n10219), .ZN(n10221) );
  XNOR2_X1 U11259 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10221), .ZN(ADD_1071_U5)
         );
  AOI22_X1 U11260 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n10222), .B2(n6218), .ZN(ADD_1071_U46) );
  OAI21_X1 U11261 ( .B1(n10225), .B2(n10224), .A(n10223), .ZN(ADD_1071_U56) );
  OAI21_X1 U11262 ( .B1(n10228), .B2(n10227), .A(n10226), .ZN(ADD_1071_U57) );
  OAI21_X1 U11263 ( .B1(n10231), .B2(n10230), .A(n10229), .ZN(ADD_1071_U58) );
  OAI21_X1 U11264 ( .B1(n10234), .B2(n10233), .A(n10232), .ZN(ADD_1071_U59) );
  OAI21_X1 U11265 ( .B1(n10237), .B2(n10236), .A(n10235), .ZN(ADD_1071_U60) );
  OAI21_X1 U11266 ( .B1(n10240), .B2(n10239), .A(n10238), .ZN(ADD_1071_U61) );
  AOI21_X1 U11267 ( .B1(n10243), .B2(n10242), .A(n10241), .ZN(ADD_1071_U62) );
  AOI21_X1 U11268 ( .B1(n10246), .B2(n10245), .A(n10244), .ZN(ADD_1071_U63) );
  XOR2_X1 U11269 ( .A(n10247), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  AOI21_X1 U11270 ( .B1(n10250), .B2(n10249), .A(n10248), .ZN(ADD_1071_U47) );
  XOR2_X1 U11271 ( .A(n10251), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11272 ( .A1(n10253), .A2(n10252), .ZN(n10254) );
  XOR2_X1 U11273 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10254), .Z(ADD_1071_U51) );
  OAI21_X1 U11274 ( .B1(n10257), .B2(n10256), .A(n10255), .ZN(n10258) );
  XNOR2_X1 U11275 ( .A(n10258), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11276 ( .A(n10260), .B(n10259), .Z(ADD_1071_U54) );
  XOR2_X1 U11277 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10261), .Z(ADD_1071_U48) );
  XOR2_X1 U11278 ( .A(n10263), .B(n10262), .Z(ADD_1071_U53) );
  XNOR2_X1 U11279 ( .A(n10265), .B(n10264), .ZN(ADD_1071_U52) );
  CLKBUF_X3 U4900 ( .A(n5886), .Z(n8376) );
  INV_X1 U4902 ( .A(n5938), .ZN(n5941) );
  INV_X2 U4910 ( .A(P2_STATE_REG_SCAN_IN), .ZN(n7777) );
endmodule

