

module b14_C_SARLock_k_128_6 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870;

  CLKBUF_X2 U2397 ( .A(n2411), .Z(n3783) );
  INV_X1 U2398 ( .A(n2819), .ZN(n2832) );
  INV_X2 U2399 ( .A(n3879), .ZN(n2804) );
  OAI21_X1 U2400 ( .B1(n4328), .B2(n3015), .A(n3017), .ZN(n3053) );
  OR2_X1 U2401 ( .A1(n3950), .A2(n3937), .ZN(n3781) );
  NAND2_X1 U2402 ( .A1(n3725), .A2(n2934), .ZN(n2932) );
  INV_X2 U2403 ( .A(n2742), .ZN(n3879) );
  INV_X1 U2405 ( .A(n4506), .ZN(n4512) );
  AND2_X1 U2406 ( .A1(n3132), .A2(n2884), .ZN(n4506) );
  XNOR2_X1 U2407 ( .A(n2384), .B(IR_REG_22__SCAN_IN), .ZN(n3880) );
  NAND2_X1 U2408 ( .A1(n3364), .A2(n3346), .ZN(n3378) );
  XNOR2_X2 U2409 ( .A(n2347), .B(IR_REG_30__SCAN_IN), .ZN(n4252) );
  NOR2_X2 U2410 ( .A1(n2691), .A2(n3689), .ZN(n2709) );
  AND2_X4 U2411 ( .A1(n2816), .A2(n4512), .ZN(n2651) );
  XNOR2_X1 U2412 ( .A(n2400), .B(IR_REG_1__SCAN_IN), .ZN(n3064) );
  XNOR2_X2 U2413 ( .A(n2417), .B(IR_REG_2__SCAN_IN), .ZN(n3028) );
  NAND2_X1 U2414 ( .A1(n3203), .A2(n3204), .ZN(n2480) );
  NAND3_X1 U2415 ( .A1(n2358), .A2(n2357), .A3(n2330), .ZN(n3895) );
  NAND4_X2 U2416 ( .A1(n2435), .A2(n2434), .A3(n2433), .A4(n2432), .ZN(n3894)
         );
  INV_X1 U2417 ( .A(n3222), .ZN(n3173) );
  NAND4_X2 U2418 ( .A1(n2399), .A2(n2398), .A3(n2397), .A4(n2396), .ZN(n3155)
         );
  AND4_X1 U2419 ( .A1(n2415), .A2(n2414), .A3(n2413), .A4(n2412), .ZN(n3222)
         );
  BUF_X2 U2420 ( .A(n2429), .Z(n2773) );
  INV_X2 U2421 ( .A(n3900), .ZN(U4043) );
  INV_X2 U2422 ( .A(n2395), .ZN(n2877) );
  AND2_X1 U2423 ( .A1(n3053), .A2(n3018), .ZN(n3054) );
  CLKBUF_X1 U2424 ( .A(n2792), .Z(n2876) );
  AND2_X1 U2425 ( .A1(n4255), .A2(n2992), .ZN(n2365) );
  NAND2_X2 U2427 ( .A1(n3877), .A2(n3216), .ZN(n2819) );
  NAND2_X1 U2428 ( .A1(n2348), .A2(n2351), .ZN(n2354) );
  NAND2_X1 U2429 ( .A1(n2348), .A2(IR_REG_31__SCAN_IN), .ZN(n2347) );
  AND2_X1 U2430 ( .A1(n2866), .A2(n2867), .ZN(n3132) );
  NAND2_X1 U2431 ( .A1(n2884), .A2(n4256), .ZN(n3216) );
  XNOR2_X1 U2432 ( .A(n2359), .B(IR_REG_26__SCAN_IN), .ZN(n4254) );
  OR2_X1 U2433 ( .A1(n2374), .A2(n2373), .ZN(n2199) );
  XNOR2_X1 U2434 ( .A(n2370), .B(IR_REG_21__SCAN_IN), .ZN(n4256) );
  OAI21_X1 U2435 ( .B1(n2363), .B2(IR_REG_25__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2359) );
  NAND2_X1 U2436 ( .A1(n2175), .A2(IR_REG_31__SCAN_IN), .ZN(n2384) );
  NOR2_X1 U2437 ( .A1(IR_REG_18__SCAN_IN), .A2(n2177), .ZN(n2328) );
  INV_X1 U2438 ( .A(IR_REG_2__SCAN_IN), .ZN(n4663) );
  NOR2_X1 U2439 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2335)
         );
  NOR2_X1 U2440 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2336)
         );
  NOR2_X1 U2441 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2337)
         );
  INV_X1 U2442 ( .A(IR_REG_3__SCAN_IN), .ZN(n2467) );
  NOR2_X1 U2443 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2539)
         );
  NOR2_X1 U2444 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2340)
         );
  AND2_X1 U2445 ( .A1(n2158), .A2(n2188), .ZN(n2345) );
  AND2_X1 U2446 ( .A1(n2342), .A2(n2681), .ZN(n2188) );
  INV_X1 U2447 ( .A(n2910), .ZN(n2316) );
  NAND2_X1 U2448 ( .A1(n3014), .A2(n3013), .ZN(n3016) );
  OAI21_X1 U2449 ( .B1(n3358), .B2(n2908), .A(n2907), .ZN(n3388) );
  NAND2_X1 U2450 ( .A1(n2327), .A2(n2326), .ZN(n2325) );
  INV_X1 U2451 ( .A(IR_REG_26__SCAN_IN), .ZN(n2327) );
  INV_X1 U2452 ( .A(IR_REG_25__SCAN_IN), .ZN(n2326) );
  NOR2_X1 U2453 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_21__SCAN_IN), .ZN(n2249)
         );
  NOR2_X1 U2454 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2338)
         );
  NOR2_X1 U2455 ( .A1(n2660), .A2(n2659), .ZN(n3707) );
  AND2_X1 U2456 ( .A1(n4252), .A2(n2354), .ZN(n2431) );
  XNOR2_X1 U2457 ( .A(n3029), .B(n4262), .ZN(n3044) );
  XNOR2_X1 U2458 ( .A(n3016), .B(n4336), .ZN(n4328) );
  NAND2_X1 U2459 ( .A1(n2276), .A2(n2277), .ZN(n2275) );
  OAI22_X1 U2460 ( .A1(n4384), .A2(n4381), .B1(REG2_REG_13__SCAN_IN), .B2(
        n4292), .ZN(n4273) );
  AOI22_X1 U2461 ( .A1(n4002), .A2(n2926), .B1(n4014), .B2(n4028), .ZN(n3982)
         );
  NOR2_X1 U2462 ( .A1(n2874), .A2(IR_REG_28__SCAN_IN), .ZN(n2349) );
  NOR2_X1 U2463 ( .A1(n3260), .A2(n2242), .ZN(n2241) );
  INV_X1 U2464 ( .A(n2479), .ZN(n2242) );
  INV_X1 U2465 ( .A(n3457), .ZN(n2257) );
  INV_X1 U2466 ( .A(n2241), .ZN(n2236) );
  OR2_X1 U2467 ( .A1(n2199), .A2(n2375), .ZN(n2377) );
  NOR2_X1 U2468 ( .A1(n3911), .A2(n2218), .ZN(n3029) );
  NOR2_X1 U2469 ( .A1(n4406), .A2(n2219), .ZN(n4275) );
  AND2_X1 U2470 ( .A1(n4296), .A2(REG2_REG_15__SCAN_IN), .ZN(n2219) );
  AOI21_X1 U2471 ( .B1(n3807), .B2(n2906), .A(n2159), .ZN(n2288) );
  NAND2_X1 U2472 ( .A1(n3296), .A2(n3252), .ZN(n3735) );
  AND2_X1 U2473 ( .A1(n3880), .A2(n4256), .ZN(n3021) );
  AND2_X1 U2474 ( .A1(n3787), .A2(DATAI_21_), .ZN(n2974) );
  OR2_X1 U2475 ( .A1(n4141), .A2(n2951), .ZN(n2205) );
  AND2_X1 U2476 ( .A1(n3407), .A2(n3431), .ZN(n2207) );
  INV_X1 U2477 ( .A(IR_REG_6__SCAN_IN), .ZN(n2538) );
  NOR2_X1 U2478 ( .A1(n3330), .A2(n2239), .ZN(n2238) );
  OR2_X1 U2479 ( .A1(n3456), .A2(n2257), .ZN(n2256) );
  NAND2_X1 U2480 ( .A1(n3351), .A2(n3352), .ZN(n2243) );
  NAND2_X1 U2481 ( .A1(n2799), .A2(n2246), .ZN(n2245) );
  NOR2_X1 U2482 ( .A1(n3696), .A2(n2247), .ZN(n2246) );
  INV_X1 U2483 ( .A(n3628), .ZN(n2247) );
  AOI21_X1 U2484 ( .B1(n3895), .B2(n2742), .A(n2381), .ZN(n2392) );
  NAND2_X1 U2485 ( .A1(n2226), .A2(n2746), .ZN(n2225) );
  AOI21_X1 U2486 ( .B1(n2160), .B2(n2226), .A(n2183), .ZN(n2224) );
  XNOR2_X1 U2487 ( .A(n2420), .B(n2832), .ZN(n2421) );
  INV_X1 U2488 ( .A(n2431), .ZN(n2881) );
  NAND2_X1 U2489 ( .A1(n2410), .A2(REG0_REG_1__SCAN_IN), .ZN(n2399) );
  INV_X1 U2490 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2259) );
  NAND2_X1 U2491 ( .A1(n3077), .A2(n2214), .ZN(n2211) );
  NOR2_X1 U2492 ( .A1(n3078), .A2(n2215), .ZN(n2214) );
  OR2_X1 U2493 ( .A1(n2217), .A2(n3078), .ZN(n2213) );
  NOR2_X1 U2494 ( .A1(n4339), .A2(n2181), .ZN(n4284) );
  XNOR2_X1 U2495 ( .A(n4273), .B(n2223), .ZN(n4389) );
  NOR2_X1 U2496 ( .A1(n4389), .A2(n4390), .ZN(n4388) );
  XNOR2_X1 U2497 ( .A(n4297), .B(n2655), .ZN(n4418) );
  NOR2_X1 U2498 ( .A1(n4401), .A2(n2261), .ZN(n4297) );
  AND2_X1 U2499 ( .A1(n4296), .A2(REG1_REG_15__SCAN_IN), .ZN(n2261) );
  NAND2_X1 U2500 ( .A1(n4418), .A2(n4792), .ZN(n4417) );
  NAND2_X1 U2501 ( .A1(n4427), .A2(n2285), .ZN(n2284) );
  OR2_X1 U2502 ( .A1(n4299), .A2(REG1_REG_17__SCAN_IN), .ZN(n2285) );
  NAND2_X1 U2503 ( .A1(n4424), .A2(n2222), .ZN(n4443) );
  OR2_X1 U2504 ( .A1(n4299), .A2(REG2_REG_17__SCAN_IN), .ZN(n2222) );
  NOR2_X1 U2505 ( .A1(n4443), .A2(n4444), .ZN(n4442) );
  AND2_X1 U2506 ( .A1(n3973), .A2(n2186), .ZN(n4157) );
  NOR2_X1 U2507 ( .A1(n2811), .A2(n4847), .ZN(n2822) );
  NAND2_X1 U2508 ( .A1(n3635), .A2(n3956), .ZN(n2307) );
  NAND2_X1 U2509 ( .A1(n2919), .A2(n2320), .ZN(n4103) );
  NOR2_X1 U2510 ( .A1(n4107), .A2(n2321), .ZN(n2320) );
  INV_X1 U2511 ( .A(n2918), .ZN(n2321) );
  AND2_X1 U2512 ( .A1(n2313), .A2(n2912), .ZN(n2312) );
  OAI21_X1 U2513 ( .B1(n2155), .B2(n2311), .A(n2174), .ZN(n2310) );
  NAND2_X1 U2514 ( .A1(n2309), .A2(n2155), .ZN(n3478) );
  NAND2_X1 U2515 ( .A1(n3422), .A2(n2313), .ZN(n2309) );
  NOR2_X1 U2516 ( .A1(n3364), .A2(n3365), .ZN(n3396) );
  AND2_X1 U2517 ( .A1(n3895), .A2(n3115), .ZN(n3141) );
  NOR2_X1 U2518 ( .A1(n3512), .A2(n3511), .ZN(n3510) );
  INV_X1 U2519 ( .A(n2852), .ZN(n2997) );
  NAND2_X1 U2520 ( .A1(n2984), .A2(n4461), .ZN(n3024) );
  MUX2_X1 U2521 ( .A(IR_REG_31__SCAN_IN), .B(n2350), .S(IR_REG_29__SCAN_IN), 
        .Z(n2351) );
  OR2_X1 U2522 ( .A1(n2349), .A2(n2373), .ZN(n2350) );
  NOR2_X1 U2523 ( .A1(n2323), .A2(IR_REG_27__SCAN_IN), .ZN(n2322) );
  NAND2_X1 U2524 ( .A1(n2324), .A2(n2329), .ZN(n2323) );
  INV_X1 U2525 ( .A(n2325), .ZN(n2324) );
  AND3_X1 U2526 ( .A1(n2342), .A2(n2681), .A3(n2329), .ZN(n2187) );
  INV_X1 U2527 ( .A(IR_REG_23__SCAN_IN), .ZN(n2853) );
  XNOR2_X1 U2528 ( .A(n2368), .B(n2367), .ZN(n2884) );
  NAND2_X1 U2529 ( .A1(n2665), .A2(n2664), .ZN(n2666) );
  OAI211_X1 U2530 ( .C1(n3707), .C2(n3710), .A(n3640), .B(n3708), .ZN(n2250)
         );
  INV_X1 U2531 ( .A(n4028), .ZN(n3993) );
  AOI22_X1 U2532 ( .A1(n4327), .A2(REG2_REG_4__SCAN_IN), .B1(n4336), .B2(n3032), .ZN(n3052) );
  NAND2_X1 U2533 ( .A1(n3020), .A2(n3038), .ZN(n2276) );
  NAND2_X1 U2534 ( .A1(n2279), .A2(n4260), .ZN(n2277) );
  NAND2_X1 U2535 ( .A1(n4373), .A2(n4272), .ZN(n4384) );
  NOR2_X1 U2536 ( .A1(n2284), .A2(n4438), .ZN(n4437) );
  INV_X1 U2537 ( .A(n2283), .ZN(n2282) );
  AOI21_X1 U2538 ( .B1(n2284), .B2(n4438), .A(n4436), .ZN(n2283) );
  OR2_X1 U2539 ( .A1(n4325), .A2(n3904), .ZN(n4441) );
  INV_X1 U2540 ( .A(n4436), .ZN(n4431) );
  OR2_X1 U2541 ( .A1(n4442), .A2(n2221), .ZN(n2220) );
  NOR2_X1 U2542 ( .A1(n4462), .A2(n4823), .ZN(n2221) );
  NAND2_X1 U2543 ( .A1(n2295), .A2(n2293), .ZN(n3587) );
  AOI21_X1 U2544 ( .B1(n2294), .B2(n2297), .A(n2173), .ZN(n2293) );
  OAI21_X1 U2545 ( .B1(n3599), .B2(n4139), .A(n2182), .ZN(n4165) );
  OAI21_X1 U2546 ( .B1(n3963), .B2(n2300), .A(n2297), .ZN(n3586) );
  INV_X2 U2547 ( .A(n4530), .ZN(n4533) );
  INV_X1 U2548 ( .A(n4255), .ZN(n2998) );
  NAND2_X1 U2549 ( .A1(n2391), .A2(n2390), .ZN(n4305) );
  NAND2_X1 U2550 ( .A1(n3054), .A2(n2269), .ZN(n2267) );
  OAI21_X1 U2551 ( .B1(n2167), .B2(n2270), .A(n3038), .ZN(n2269) );
  NAND2_X1 U2552 ( .A1(n2275), .A2(REG1_REG_6__SCAN_IN), .ZN(n2272) );
  NOR2_X1 U2553 ( .A1(n2232), .A2(n3667), .ZN(n2231) );
  INV_X1 U2554 ( .A(n3614), .ZN(n2232) );
  AOI21_X1 U2555 ( .B1(n4287), .B2(REG1_REG_11__SCAN_IN), .A(n4358), .ZN(n4289) );
  INV_X1 U2556 ( .A(n2928), .ZN(n2299) );
  NAND2_X1 U2557 ( .A1(n3965), .A2(n3856), .ZN(n3946) );
  NAND2_X1 U2558 ( .A1(n3985), .A2(n3859), .ZN(n3965) );
  OAI21_X1 U2559 ( .B1(n4040), .B2(n3855), .A(n3853), .ZN(n3985) );
  INV_X1 U2560 ( .A(n2912), .ZN(n2311) );
  INV_X1 U2561 ( .A(n2315), .ZN(n2314) );
  OAI21_X1 U2562 ( .B1(n2317), .B2(n2316), .A(n2911), .ZN(n2315) );
  NOR2_X1 U2563 ( .A1(n2316), .A2(n2166), .ZN(n2313) );
  INV_X1 U2564 ( .A(n3816), .ZN(n2317) );
  OAI211_X1 U2565 ( .C1(n2292), .C2(n2291), .A(n2290), .B(n2896), .ZN(n3242)
         );
  NAND2_X1 U2566 ( .A1(n2932), .A2(n2172), .ZN(n2290) );
  CLKBUF_X1 U2567 ( .A(n2934), .Z(n3728) );
  AND2_X1 U2568 ( .A1(n2935), .A2(n3181), .ZN(n2292) );
  NOR2_X1 U2569 ( .A1(n2975), .A2(n2210), .ZN(n2208) );
  AND2_X1 U2570 ( .A1(n2838), .A2(n4254), .ZN(n2852) );
  INV_X1 U2571 ( .A(IR_REG_20__SCAN_IN), .ZN(n2367) );
  NAND2_X1 U2572 ( .A1(n2480), .A2(n2241), .ZN(n2240) );
  NAND2_X1 U2573 ( .A1(n2401), .A2(DATAI_27_), .ZN(n3937) );
  INV_X1 U2574 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2616) );
  NAND2_X1 U2575 ( .A1(n2401), .A2(DATAI_23_), .ZN(n3803) );
  AND2_X1 U2576 ( .A1(n2228), .A2(n2227), .ZN(n2226) );
  INV_X1 U2577 ( .A(n2662), .ZN(n2665) );
  NAND2_X1 U2578 ( .A1(n2771), .A2(REG3_REG_24__SCAN_IN), .ZN(n2790) );
  AND2_X1 U2579 ( .A1(n2756), .A2(REG3_REG_23__SCAN_IN), .ZN(n2771) );
  OAI21_X1 U2580 ( .B1(n2480), .B2(n2237), .A(n2235), .ZN(n4538) );
  INV_X1 U2581 ( .A(n2238), .ZN(n2237) );
  AOI21_X1 U2582 ( .B1(n2238), .B2(n2236), .A(n2178), .ZN(n2235) );
  NAND2_X1 U2583 ( .A1(n2229), .A2(n2332), .ZN(n2228) );
  INV_X1 U2584 ( .A(n3667), .ZN(n2229) );
  NAND2_X1 U2585 ( .A1(n3613), .A2(n2231), .ZN(n2230) );
  OR2_X1 U2586 ( .A1(n2599), .A2(n3460), .ZN(n2617) );
  OR2_X1 U2587 ( .A1(n2670), .A2(n2669), .ZN(n2691) );
  NOR2_X1 U2588 ( .A1(n2481), .A2(n3036), .ZN(n2497) );
  INV_X1 U2589 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3036) );
  AND3_X1 U2590 ( .A1(n2795), .A2(n2794), .A3(n2793), .ZN(n3699) );
  OR2_X1 U2591 ( .A1(n3632), .A2(n2876), .ZN(n2794) );
  NAND2_X1 U2592 ( .A1(n3026), .A2(n2171), .ZN(n3907) );
  AOI21_X1 U2593 ( .B1(n3907), .B2(n3908), .A(n3909), .ZN(n3911) );
  INV_X1 U2594 ( .A(REG3_REG_8__SCAN_IN), .ZN(n3085) );
  AND3_X1 U2595 ( .A1(n2211), .A2(n2184), .A3(n2213), .ZN(n4265) );
  INV_X1 U2596 ( .A(n4259), .ZN(n2216) );
  XNOR2_X1 U2597 ( .A(n4284), .B(n2262), .ZN(n4350) );
  XNOR2_X1 U2598 ( .A(n4289), .B(n4469), .ZN(n4369) );
  OAI21_X1 U2599 ( .B1(n4369), .B2(n2265), .A(n2264), .ZN(n4377) );
  NAND2_X1 U2600 ( .A1(n2266), .A2(REG1_REG_12__SCAN_IN), .ZN(n2265) );
  NAND2_X1 U2601 ( .A1(n4290), .A2(n2266), .ZN(n2264) );
  INV_X1 U2602 ( .A(n4378), .ZN(n2266) );
  NOR2_X1 U2603 ( .A1(n4369), .A2(n4743), .ZN(n4368) );
  INV_X1 U2604 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3460) );
  NAND2_X1 U2605 ( .A1(n4363), .A2(n4270), .ZN(n4271) );
  NOR2_X1 U2606 ( .A1(n2623), .A2(IR_REG_13__SCAN_IN), .ZN(n2639) );
  AOI21_X1 U2607 ( .B1(n4292), .B2(REG1_REG_13__SCAN_IN), .A(n4377), .ZN(n4293) );
  XNOR2_X1 U2608 ( .A(n4275), .B(n2655), .ZN(n4416) );
  NAND2_X1 U2609 ( .A1(n4416), .A2(n4415), .ZN(n4414) );
  AND2_X1 U2610 ( .A1(n3787), .A2(n3022), .ZN(n3034) );
  AND2_X1 U2611 ( .A1(n2297), .A2(n3584), .ZN(n2296) );
  NOR2_X1 U2612 ( .A1(n2302), .A2(n3830), .ZN(n2294) );
  AND2_X1 U2613 ( .A1(n2301), .A2(n2298), .ZN(n2297) );
  OR2_X1 U2614 ( .A1(n2306), .A2(n2157), .ZN(n2301) );
  NAND2_X1 U2615 ( .A1(n2302), .A2(n2299), .ZN(n2298) );
  AND2_X1 U2616 ( .A1(n2930), .A2(n2307), .ZN(n2306) );
  AND2_X1 U2617 ( .A1(n3787), .A2(DATAI_28_), .ZN(n2975) );
  AND2_X1 U2618 ( .A1(n2830), .A2(n2829), .ZN(n3930) );
  OR2_X1 U2619 ( .A1(n3920), .A2(n2876), .ZN(n2830) );
  OR2_X1 U2620 ( .A1(n2790), .A2(n3633), .ZN(n2800) );
  AND2_X1 U2621 ( .A1(n3800), .A2(n3945), .ZN(n3966) );
  AND2_X1 U2622 ( .A1(n3787), .A2(DATAI_25_), .ZN(n3968) );
  INV_X1 U2623 ( .A(n3995), .ZN(n3989) );
  NAND2_X1 U2624 ( .A1(n4039), .A2(n2922), .ZN(n2319) );
  OR2_X1 U2625 ( .A1(n2733), .A2(n3623), .ZN(n2747) );
  NAND2_X1 U2626 ( .A1(n4103), .A2(n2920), .ZN(n4081) );
  INV_X1 U2627 ( .A(n3887), .ZN(n4113) );
  AOI21_X1 U2628 ( .B1(n3550), .B2(n3547), .A(n3768), .ZN(n4130) );
  OAI21_X1 U2629 ( .B1(n3466), .B2(n3809), .A(n3747), .ZN(n3550) );
  AOI21_X1 U2630 ( .B1(n3465), .B2(n2914), .A(n2331), .ZN(n3549) );
  NAND2_X1 U2631 ( .A1(n3503), .A2(n3766), .ZN(n3466) );
  NAND2_X1 U2632 ( .A1(n2566), .A2(REG3_REG_11__SCAN_IN), .ZN(n2580) );
  INV_X1 U2633 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2579) );
  INV_X1 U2634 ( .A(n3425), .ZN(n3431) );
  OAI22_X1 U2635 ( .A1(n3388), .A2(n2909), .B1(n3427), .B2(n3407), .ZN(n3422)
         );
  NAND2_X1 U2636 ( .A1(n2318), .A2(n2317), .ZN(n3424) );
  INV_X1 U2637 ( .A(n3422), .ZN(n2318) );
  AND2_X1 U2638 ( .A1(n3437), .A2(n3440), .ZN(n3816) );
  NAND2_X1 U2639 ( .A1(n2287), .A2(n2286), .ZN(n3358) );
  AOI21_X1 U2640 ( .B1(n2288), .B2(n2289), .A(n2169), .ZN(n2286) );
  INV_X1 U2641 ( .A(n3890), .ZN(n3427) );
  AOI21_X1 U2642 ( .B1(n2196), .B2(n2195), .A(n2194), .ZN(n2193) );
  INV_X1 U2643 ( .A(n3753), .ZN(n2194) );
  INV_X1 U2644 ( .A(n3331), .ZN(n3310) );
  OAI21_X1 U2645 ( .B1(n3240), .B2(n2937), .A(n3738), .ZN(n3294) );
  NAND2_X1 U2646 ( .A1(n3227), .A2(n2201), .ZN(n3300) );
  AND2_X1 U2647 ( .A1(n3226), .A2(n3165), .ZN(n2201) );
  AND2_X1 U2648 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2460) );
  NAND2_X1 U2649 ( .A1(n3218), .A2(n3734), .ZN(n3240) );
  INV_X1 U2650 ( .A(n4112), .ZN(n4137) );
  NAND2_X1 U2651 ( .A1(n3227), .A2(n3226), .ZN(n3251) );
  NAND2_X1 U2652 ( .A1(n3219), .A2(n3810), .ZN(n3218) );
  NAND2_X1 U2653 ( .A1(n2932), .A2(n3141), .ZN(n3182) );
  INV_X1 U2654 ( .A(n4162), .ZN(n4132) );
  INV_X1 U2655 ( .A(n3122), .ZN(n3146) );
  INV_X1 U2656 ( .A(n4305), .ZN(n2961) );
  INV_X1 U2657 ( .A(n4139), .ZN(n4115) );
  AND2_X1 U2658 ( .A1(n3787), .A2(DATAI_30_), .ZN(n4163) );
  AND2_X1 U2659 ( .A1(n3132), .A2(n4257), .ZN(n4162) );
  INV_X1 U2660 ( .A(n2975), .ZN(n3585) );
  NAND2_X1 U2661 ( .A1(n3973), .A2(n2209), .ZN(n3936) );
  NAND2_X1 U2662 ( .A1(n2401), .A2(DATAI_26_), .ZN(n3956) );
  INV_X1 U2663 ( .A(n3968), .ZN(n3975) );
  NOR2_X1 U2664 ( .A1(n3994), .A2(n3968), .ZN(n3973) );
  NAND2_X1 U2665 ( .A1(n2401), .A2(DATAI_24_), .ZN(n3995) );
  OR2_X1 U2666 ( .A1(n4016), .A2(n3989), .ZN(n3994) );
  OR2_X1 U2667 ( .A1(n4188), .A2(n4014), .ZN(n4016) );
  INV_X1 U2668 ( .A(n3803), .ZN(n4014) );
  NAND2_X1 U2669 ( .A1(n4047), .A2(n4034), .ZN(n4188) );
  NAND2_X1 U2670 ( .A1(n2204), .A2(n2203), .ZN(n2202) );
  NOR2_X1 U2671 ( .A1(n4108), .A2(n4075), .ZN(n2203) );
  INV_X1 U2672 ( .A(n2205), .ZN(n2204) );
  NOR2_X1 U2673 ( .A1(n4197), .A2(n2974), .ZN(n4047) );
  NOR3_X1 U2674 ( .A1(n4213), .A2(n4108), .A3(n4141), .ZN(n4118) );
  NOR2_X1 U2675 ( .A1(n4213), .A2(n4141), .ZN(n4142) );
  OR2_X1 U2676 ( .A1(n3557), .A2(n3556), .ZN(n4213) );
  INV_X1 U2677 ( .A(n3713), .ZN(n3470) );
  NAND2_X1 U2678 ( .A1(n3396), .A2(n2180), .ZN(n3512) );
  NAND2_X1 U2679 ( .A1(n3396), .A2(n2163), .ZN(n3492) );
  NAND2_X1 U2680 ( .A1(n3396), .A2(n2207), .ZN(n3450) );
  AND2_X1 U2681 ( .A1(n3396), .A2(n3407), .ZN(n4507) );
  INV_X1 U2682 ( .A(n3340), .ZN(n4541) );
  OR2_X1 U2683 ( .A1(n3345), .A2(n4541), .ZN(n3364) );
  INV_X1 U2684 ( .A(n3276), .ZN(n3284) );
  NOR2_X1 U2685 ( .A1(n2200), .A2(n3300), .ZN(n3311) );
  NAND2_X1 U2686 ( .A1(n2938), .A2(n3284), .ZN(n2200) );
  NOR2_X1 U2687 ( .A1(n3300), .A2(n3301), .ZN(n3299) );
  NAND2_X1 U2688 ( .A1(n3508), .A2(n4480), .ZN(n4496) );
  NOR2_X1 U2689 ( .A1(n3194), .A2(n3193), .ZN(n3227) );
  OR2_X1 U2690 ( .A1(n3213), .A2(n2972), .ZN(n2980) );
  AND2_X1 U2691 ( .A1(n4449), .A2(n2866), .ZN(n4517) );
  NOR2_X1 U2692 ( .A1(n2363), .A2(n2325), .ZN(n2374) );
  INV_X1 U2693 ( .A(IR_REG_19__SCAN_IN), .ZN(n2388) );
  AND2_X1 U2694 ( .A1(n2342), .A2(n2681), .ZN(n2698) );
  AND2_X1 U2695 ( .A1(n2652), .A2(n2643), .ZN(n4296) );
  AND2_X1 U2696 ( .A1(n2542), .A2(n2608), .ZN(n4283) );
  OR2_X1 U2697 ( .A1(n2503), .A2(n2373), .ZN(n2517) );
  INV_X1 U2698 ( .A(n2254), .ZN(n2253) );
  AOI21_X1 U2699 ( .B1(n2254), .B2(n2252), .A(n2165), .ZN(n2251) );
  AND2_X1 U2700 ( .A1(n2256), .A2(n2255), .ZN(n2254) );
  AND2_X1 U2701 ( .A1(n3606), .A2(n3607), .ZN(n2770) );
  NAND2_X1 U2702 ( .A1(n2243), .A2(n2549), .ZN(n3405) );
  INV_X1 U2703 ( .A(n3103), .ZN(n4544) );
  INV_X1 U2704 ( .A(n3390), .ZN(n3407) );
  INV_X1 U2705 ( .A(n3442), .ZN(n3417) );
  INV_X1 U2706 ( .A(n3220), .ZN(n3226) );
  NOR2_X1 U2707 ( .A1(n2248), .A2(n3695), .ZN(n2244) );
  INV_X1 U2708 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3623) );
  AOI21_X1 U2709 ( .B1(n3613), .B2(n3614), .A(n2332), .ZN(n3669) );
  NAND2_X1 U2710 ( .A1(n2230), .A2(n2228), .ZN(n3670) );
  INV_X1 U2711 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4850) );
  NAND2_X1 U2712 ( .A1(n2882), .A2(n3897), .ZN(n3715) );
  OAI22_X1 U2713 ( .A1(n3649), .A2(n2690), .B1(n3651), .B2(n3650), .ZN(n3688)
         );
  NAND2_X1 U2714 ( .A1(n2799), .A2(n3628), .ZN(n3698) );
  INV_X1 U2715 ( .A(n3700), .ZN(n4542) );
  INV_X1 U2716 ( .A(n4543), .ZN(n3712) );
  OAI211_X1 U2717 ( .C1(n3939), .C2(n2876), .A(n2814), .B(n2813), .ZN(n3950)
         );
  OAI211_X1 U2718 ( .C1(n3958), .C2(n2876), .A(n2803), .B(n2802), .ZN(n3969)
         );
  INV_X1 U2719 ( .A(n3699), .ZN(n3990) );
  NAND4_X1 U2720 ( .A1(n2761), .A2(n2760), .A3(n2759), .A4(n2758), .ZN(n4028)
         );
  NAND4_X1 U2721 ( .A1(n2714), .A2(n2713), .A3(n2712), .A4(n2711), .ZN(n4110)
         );
  NAND4_X2 U2722 ( .A1(n2446), .A2(n2445), .A3(n2444), .A4(n2443), .ZN(n3893)
         );
  NAND2_X1 U2723 ( .A1(n2411), .A2(REG1_REG_1__SCAN_IN), .ZN(n2396) );
  NAND2_X1 U2724 ( .A1(n2429), .A2(REG3_REG_1__SCAN_IN), .ZN(n2398) );
  OR2_X1 U2725 ( .A1(n2395), .A2(n2353), .ZN(n2357) );
  OR2_X1 U2726 ( .A1(n2984), .A2(n3878), .ZN(n3900) );
  NAND2_X1 U2727 ( .A1(n3054), .A2(n3038), .ZN(n2274) );
  AND2_X1 U2728 ( .A1(n2212), .A2(n2217), .ZN(n3079) );
  NAND2_X1 U2729 ( .A1(n2211), .A2(n2213), .ZN(n3084) );
  NAND2_X1 U2730 ( .A1(n3077), .A2(REG2_REG_6__SCAN_IN), .ZN(n2212) );
  AND2_X1 U2731 ( .A1(n2273), .A2(n2278), .ZN(n3087) );
  OAI211_X1 U2732 ( .C1(n3054), .C2(n2275), .A(REG1_REG_6__SCAN_IN), .B(n2268), 
        .ZN(n2273) );
  NAND2_X1 U2733 ( .A1(n3054), .A2(n2167), .ZN(n2268) );
  OR2_X1 U2734 ( .A1(n3090), .A2(n3374), .ZN(n4279) );
  AND2_X1 U2735 ( .A1(n4282), .A2(n2263), .ZN(n4339) );
  INV_X1 U2736 ( .A(n4340), .ZN(n2263) );
  INV_X1 U2737 ( .A(n4282), .ZN(n4341) );
  NAND2_X1 U2738 ( .A1(n4354), .A2(n4269), .ZN(n4364) );
  NAND2_X1 U2739 ( .A1(n4364), .A2(n4365), .ZN(n4363) );
  XNOR2_X1 U2740 ( .A(n4271), .B(n4469), .ZN(n4374) );
  NOR2_X1 U2741 ( .A1(n4274), .A2(n4388), .ZN(n4407) );
  NOR2_X1 U2742 ( .A1(n4407), .A2(n4408), .ZN(n4406) );
  NAND2_X1 U2743 ( .A1(n4417), .A2(n4298), .ZN(n4428) );
  AND2_X1 U2744 ( .A1(n2308), .A2(n2307), .ZN(n3934) );
  NAND2_X1 U2745 ( .A1(n2305), .A2(n2303), .ZN(n2308) );
  NAND2_X1 U2746 ( .A1(n2919), .A2(n2918), .ZN(n4105) );
  NAND2_X1 U2747 ( .A1(n3316), .A2(n2906), .ZN(n3344) );
  AND2_X1 U2748 ( .A1(n4125), .A2(n4305), .ZN(n4120) );
  AND2_X1 U2749 ( .A1(n4120), .A2(n4506), .ZN(n4316) );
  OR2_X1 U2750 ( .A1(n3214), .A2(n3213), .ZN(n3215) );
  OR2_X1 U2751 ( .A1(n2980), .A2(n3211), .ZN(n4530) );
  OAI21_X1 U2752 ( .B1(n4167), .B2(n4501), .A(n2192), .ZN(n2191) );
  NAND2_X1 U2753 ( .A1(n4166), .A2(n4506), .ZN(n2192) );
  INV_X2 U2754 ( .A(n4518), .ZN(n4520) );
  NAND2_X1 U2755 ( .A1(n2997), .A2(n2996), .ZN(n4459) );
  INV_X1 U2756 ( .A(IR_REG_29__SCAN_IN), .ZN(n2346) );
  INV_X1 U2757 ( .A(n2354), .ZN(n4253) );
  XNOR2_X1 U2758 ( .A(n2875), .B(n2375), .ZN(n4311) );
  XNOR2_X1 U2759 ( .A(n2364), .B(IR_REG_25__SCAN_IN), .ZN(n2992) );
  XNOR2_X1 U2760 ( .A(n2362), .B(IR_REG_24__SCAN_IN), .ZN(n4255) );
  AND2_X1 U2761 ( .A1(n3023), .A2(STATE_REG_SCAN_IN), .ZN(n4461) );
  INV_X1 U2762 ( .A(n4283), .ZN(n4475) );
  XNOR2_X1 U2763 ( .A(n2448), .B(IR_REG_4__SCAN_IN), .ZN(n4336) );
  AND2_X1 U2764 ( .A1(n2447), .A2(n2438), .ZN(n4262) );
  OAI211_X1 U2765 ( .C1(n3054), .C2(n2277), .A(n2276), .B(n2274), .ZN(n3072)
         );
  INV_X1 U2766 ( .A(n2280), .ZN(n4447) );
  OAI21_X1 U2767 ( .B1(n4437), .B2(n2282), .A(n2281), .ZN(n2280) );
  XNOR2_X1 U2768 ( .A(n2220), .B(n4277), .ZN(n4309) );
  NAND2_X1 U2769 ( .A1(n2190), .A2(n2189), .ZN(U3547) );
  OR2_X1 U2770 ( .A1(n4533), .A2(n4634), .ZN(n2189) );
  NAND2_X1 U2771 ( .A1(n4221), .A2(n4533), .ZN(n2190) );
  OR2_X1 U2772 ( .A1(n3918), .A2(n4211), .ZN(n2977) );
  MUX2_X1 U2773 ( .A(n2973), .B(n2981), .S(n4533), .Z(n2978) );
  MUX2_X1 U2774 ( .A(n4630), .B(n2981), .S(n4520), .Z(n2983) );
  INV_X1 U2775 ( .A(n2906), .ZN(n2289) );
  OR2_X1 U2776 ( .A1(n2314), .A2(n2166), .ZN(n2155) );
  AND2_X1 U2777 ( .A1(n4259), .A2(REG1_REG_7__SCAN_IN), .ZN(n2156) );
  AND2_X1 U2778 ( .A1(n3950), .A2(n3928), .ZN(n2157) );
  AND2_X1 U2779 ( .A1(n2328), .A2(n2249), .ZN(n2158) );
  AND2_X1 U2780 ( .A1(n3353), .A2(n3340), .ZN(n2159) );
  NOR2_X1 U2781 ( .A1(n2231), .A2(n2234), .ZN(n2160) );
  AND2_X1 U2782 ( .A1(n2924), .A2(n2923), .ZN(n2161) );
  AND2_X1 U2783 ( .A1(n2560), .A2(n2549), .ZN(n2162) );
  AND2_X1 U2784 ( .A1(n2207), .A2(n3445), .ZN(n2163) );
  OR3_X1 U2785 ( .A1(n4213), .A2(n2205), .A3(n4108), .ZN(n2164) );
  AND2_X1 U2786 ( .A1(n3456), .A2(n2257), .ZN(n2165) );
  NAND2_X1 U2787 ( .A1(n2905), .A2(n2904), .ZN(n3316) );
  NAND2_X1 U2788 ( .A1(n2240), .A2(n3259), .ZN(n3329) );
  NOR2_X1 U2789 ( .A1(n3889), .A2(n3449), .ZN(n2166) );
  AND2_X1 U2790 ( .A1(n2276), .A2(n4260), .ZN(n2167) );
  AND2_X1 U2791 ( .A1(n2230), .A2(n2226), .ZN(n2168) );
  AND2_X1 U2792 ( .A1(n3891), .A2(n4541), .ZN(n2169) );
  NAND2_X1 U2793 ( .A1(n3990), .A2(n3968), .ZN(n2170) );
  NAND2_X1 U2794 ( .A1(n2187), .A2(n2158), .ZN(n2363) );
  NAND2_X1 U2795 ( .A1(n2319), .A2(n2923), .ZN(n4022) );
  INV_X1 U2796 ( .A(n2345), .ZN(n2360) );
  INV_X1 U2797 ( .A(n2302), .ZN(n2300) );
  NOR2_X1 U2798 ( .A1(n2157), .A2(n2304), .ZN(n2302) );
  AND2_X1 U2799 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2171)
         );
  AND2_X1 U2800 ( .A1(n3141), .A2(n2895), .ZN(n2172) );
  NOR2_X1 U2801 ( .A1(n3930), .A2(n3585), .ZN(n2173) );
  INV_X1 U2802 ( .A(n2938), .ZN(n3301) );
  NAND2_X1 U2803 ( .A1(n3477), .A2(n3485), .ZN(n2174) );
  AND2_X1 U2804 ( .A1(n2940), .A2(n3750), .ZN(n3807) );
  OR2_X1 U2805 ( .A1(n2369), .A2(IR_REG_21__SCAN_IN), .ZN(n2175) );
  INV_X1 U2806 ( .A(IR_REG_27__SCAN_IN), .ZN(n2378) );
  INV_X1 U2807 ( .A(n2304), .ZN(n2303) );
  NAND2_X1 U2808 ( .A1(n2170), .A2(n2929), .ZN(n2304) );
  OR2_X1 U2809 ( .A1(n2436), .A2(n2468), .ZN(n2176) );
  OR2_X1 U2810 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2177)
         );
  AND2_X1 U2811 ( .A1(n2510), .A2(n2509), .ZN(n2178) );
  INV_X1 U2812 ( .A(n2197), .ZN(n2196) );
  NAND2_X1 U2813 ( .A1(n2198), .A2(n3743), .ZN(n2197) );
  INV_X1 U2814 ( .A(n4023), .ZN(n2924) );
  INV_X1 U2815 ( .A(n4285), .ZN(n2262) );
  INV_X1 U2816 ( .A(n3750), .ZN(n2195) );
  NAND2_X1 U2817 ( .A1(n2250), .A2(n2666), .ZN(n3649) );
  NAND2_X1 U2818 ( .A1(n3424), .A2(n2910), .ZN(n3448) );
  NOR2_X1 U2819 ( .A1(n4213), .A2(n2202), .ZN(n2206) );
  NOR2_X1 U2820 ( .A1(n4368), .A2(n4290), .ZN(n2179) );
  AND2_X1 U2821 ( .A1(n3844), .A2(n3847), .ZN(n3547) );
  AND2_X1 U2822 ( .A1(n2163), .A2(n3493), .ZN(n2180) );
  AND2_X1 U2823 ( .A1(n4283), .A2(REG1_REG_9__SCAN_IN), .ZN(n2181) );
  INV_X1 U2824 ( .A(n2746), .ZN(n2234) );
  AND2_X1 U2825 ( .A1(n3597), .A2(n3598), .ZN(n2182) );
  AND2_X1 U2826 ( .A1(n2745), .A2(n3620), .ZN(n2183) );
  OR2_X1 U2827 ( .A1(n2216), .A2(n3313), .ZN(n2184) );
  INV_X1 U2828 ( .A(n4108), .ZN(n4117) );
  INV_X1 U2829 ( .A(n4396), .ZN(n2223) );
  OAI21_X1 U2830 ( .B1(n4538), .B2(n4535), .A(n4534), .ZN(n3351) );
  NAND2_X1 U2831 ( .A1(n2480), .A2(n2479), .ZN(n3258) );
  INV_X1 U2832 ( .A(n3414), .ZN(n2252) );
  INV_X1 U2833 ( .A(n3259), .ZN(n2239) );
  AND2_X1 U2834 ( .A1(n2240), .A2(n2238), .ZN(n2185) );
  INV_X1 U2835 ( .A(n3666), .ZN(n2227) );
  INV_X1 U2836 ( .A(n2956), .ZN(n4034) );
  AND2_X1 U2837 ( .A1(n3787), .A2(DATAI_22_), .ZN(n2956) );
  INV_X1 U2838 ( .A(n2951), .ZN(n4095) );
  XNOR2_X1 U2839 ( .A(n2654), .B(n2653), .ZN(n4465) );
  INV_X1 U2840 ( .A(n2210), .ZN(n2209) );
  NAND2_X1 U2841 ( .A1(n3956), .A2(n3937), .ZN(n2210) );
  INV_X1 U2842 ( .A(n3789), .ZN(n3596) );
  AND2_X1 U2843 ( .A1(n3789), .A2(n2208), .ZN(n2186) );
  INV_X1 U2844 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2215) );
  INV_X1 U2845 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2270) );
  OAI21_X1 U2846 ( .B1(n3054), .B2(n3020), .A(n4260), .ZN(n2278) );
  XNOR2_X1 U2847 ( .A(n3075), .B(n4260), .ZN(n3077) );
  AOI21_X1 U2848 ( .B1(n3020), .B2(n4260), .A(n2156), .ZN(n2271) );
  AOI21_X1 U2849 ( .B1(n4440), .B2(ADDR_REG_18__SCAN_IN), .A(n4439), .ZN(n2281) );
  AOI21_X4 U2850 ( .B1(n3114), .B2(n2871), .A(U3149), .ZN(n4547) );
  AOI21_X2 U2851 ( .B1(n4063), .B2(n3851), .A(n3850), .ZN(n4040) );
  NOR2_X4 U2852 ( .A1(n2436), .A2(n2341), .ZN(n2681) );
  NOR2_X2 U2853 ( .A1(n2677), .A2(n2339), .ZN(n2342) );
  OR2_X2 U2854 ( .A1(n4165), .A2(n2191), .ZN(n4221) );
  OAI21_X1 U2855 ( .B1(n3305), .B2(n2197), .A(n2193), .ZN(n3359) );
  OAI21_X1 U2856 ( .B1(n3305), .B2(n2941), .A(n3750), .ZN(n3339) );
  NAND2_X1 U2857 ( .A1(n2941), .A2(n3750), .ZN(n2198) );
  NAND2_X1 U2858 ( .A1(n2199), .A2(n2378), .ZN(n2376) );
  XNOR2_X1 U2859 ( .A(n2199), .B(IR_REG_27__SCAN_IN), .ZN(n4322) );
  INV_X1 U2860 ( .A(n2206), .ZN(n4197) );
  NAND2_X1 U2861 ( .A1(n3973), .A2(n2208), .ZN(n3588) );
  AND2_X1 U2862 ( .A1(n3973), .A2(n3956), .ZN(n3954) );
  NAND2_X1 U2863 ( .A1(n3076), .A2(n4260), .ZN(n2217) );
  AND2_X1 U2864 ( .A1(n3028), .A2(REG2_REG_2__SCAN_IN), .ZN(n2218) );
  MUX2_X1 U2865 ( .A(n3027), .B(REG2_REG_2__SCAN_IN), .S(n3028), .Z(n3909) );
  NAND2_X1 U2866 ( .A1(n2377), .A2(n2376), .ZN(n2380) );
  OAI21_X1 U2867 ( .B1(n3613), .B2(n2225), .A(n2224), .ZN(n2233) );
  INV_X1 U2868 ( .A(n2233), .ZN(n3676) );
  NAND2_X1 U2869 ( .A1(n2243), .A2(n2162), .ZN(n3403) );
  NAND2_X1 U2870 ( .A1(n2245), .A2(n3694), .ZN(n3577) );
  NAND2_X1 U2871 ( .A1(n2245), .A2(n2244), .ZN(n2893) );
  INV_X1 U2872 ( .A(n3576), .ZN(n2248) );
  NAND3_X1 U2873 ( .A1(n2342), .A2(n2681), .A3(n2328), .ZN(n2369) );
  OAI21_X1 U2874 ( .B1(n3413), .B2(n2253), .A(n2251), .ZN(n3528) );
  OAI21_X1 U2875 ( .B1(n3413), .B2(n3415), .A(n3414), .ZN(n3459) );
  NAND2_X1 U2876 ( .A1(n3415), .A2(n3414), .ZN(n2255) );
  XNOR2_X1 U2877 ( .A(n3905), .B(n2258), .ZN(n3914) );
  INV_X1 U2878 ( .A(n3009), .ZN(n2258) );
  XNOR2_X1 U2879 ( .A(n3028), .B(n2259), .ZN(n3009) );
  NAND2_X1 U2880 ( .A1(n2260), .A2(IR_REG_31__SCAN_IN), .ZN(n2417) );
  INV_X1 U2881 ( .A(n2416), .ZN(n2260) );
  OAI211_X1 U2882 ( .C1(n3054), .C2(n2272), .A(n2271), .B(n2267), .ZN(n3089)
         );
  INV_X1 U2883 ( .A(n3020), .ZN(n2279) );
  NAND2_X1 U2884 ( .A1(n2905), .A2(n2288), .ZN(n2287) );
  NAND2_X1 U2885 ( .A1(n3183), .A2(n2895), .ZN(n3210) );
  NAND2_X1 U2886 ( .A1(n2292), .A2(n3182), .ZN(n3183) );
  INV_X1 U2887 ( .A(n2895), .ZN(n2291) );
  NAND2_X1 U2888 ( .A1(n3963), .A2(n2296), .ZN(n2295) );
  NAND2_X1 U2889 ( .A1(n3963), .A2(n2928), .ZN(n2305) );
  AND2_X1 U2890 ( .A1(n2305), .A2(n2170), .ZN(n3944) );
  AOI21_X1 U2891 ( .B1(n3422), .B2(n2312), .A(n2310), .ZN(n3502) );
  NAND2_X1 U2892 ( .A1(n2319), .A2(n2161), .ZN(n4025) );
  NAND2_X1 U2893 ( .A1(n2345), .A2(n2322), .ZN(n2874) );
  NAND3_X1 U2894 ( .A1(n2342), .A2(n2681), .A3(n2343), .ZN(n2366) );
  INV_X2 U2895 ( .A(n2792), .ZN(n2429) );
  INV_X1 U2896 ( .A(n2935), .ZN(n3832) );
  NAND2_X1 U2897 ( .A1(n3222), .A2(n3193), .ZN(n3729) );
  XNOR2_X1 U2898 ( .A(n3587), .B(n3836), .ZN(n4167) );
  NAND2_X1 U2899 ( .A1(n2421), .A2(n2422), .ZN(n2428) );
  INV_X1 U2900 ( .A(n3155), .ZN(n3186) );
  NAND2_X1 U2901 ( .A1(n3186), .A2(n3122), .ZN(n2934) );
  OAI21_X2 U2902 ( .B1(n2788), .B2(n2787), .A(n2786), .ZN(n3659) );
  XNOR2_X1 U2903 ( .A(n2404), .B(n2819), .ZN(n2405) );
  OAI21_X2 U2904 ( .B1(n3688), .B2(n3685), .A(n3684), .ZN(n3613) );
  AND2_X1 U2905 ( .A1(n2853), .A2(n2344), .ZN(n2329) );
  INV_X1 U2906 ( .A(n4010), .ZN(n4042) );
  AND2_X1 U2907 ( .A1(n2356), .A2(n2355), .ZN(n2330) );
  AND2_X1 U2908 ( .A1(n3642), .A2(n3470), .ZN(n2331) );
  AND2_X1 U2909 ( .A1(n2720), .A2(n2719), .ZN(n2332) );
  XNOR2_X1 U2910 ( .A(n2451), .B(n2819), .ZN(n2456) );
  INV_X1 U2911 ( .A(IR_REG_31__SCAN_IN), .ZN(n2373) );
  NOR2_X2 U2912 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2605)
         );
  NOR2_X1 U2913 ( .A1(n3024), .A2(n2968), .ZN(n2333) );
  OR2_X1 U2914 ( .A1(n3024), .A2(n2872), .ZN(n2334) );
  NOR2_X1 U2915 ( .A1(n2883), .A2(n2856), .ZN(n3678) );
  NAND2_X2 U2916 ( .A1(n3215), .A2(n4096), .ZN(n4125) );
  INV_X1 U2917 ( .A(n4125), .ZN(n4458) );
  INV_X1 U2918 ( .A(n4125), .ZN(n4315) );
  INV_X1 U2919 ( .A(IR_REG_18__SCAN_IN), .ZN(n2343) );
  INV_X1 U2920 ( .A(IR_REG_24__SCAN_IN), .ZN(n2344) );
  INV_X1 U2921 ( .A(IR_REG_28__SCAN_IN), .ZN(n2375) );
  INV_X1 U2922 ( .A(IR_REG_4__SCAN_IN), .ZN(n2466) );
  INV_X1 U2923 ( .A(n2457), .ZN(n2458) );
  INV_X1 U2924 ( .A(n2372), .ZN(n2815) );
  INV_X1 U2925 ( .A(n2663), .ZN(n2664) );
  AND2_X1 U2926 ( .A1(n4062), .A2(n2955), .ZN(n3851) );
  INV_X1 U2927 ( .A(n3807), .ZN(n2904) );
  NAND2_X1 U2928 ( .A1(n2456), .A2(n2458), .ZN(n2459) );
  INV_X1 U2929 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2531) );
  INV_X1 U2930 ( .A(n3406), .ZN(n2560) );
  OR2_X1 U2931 ( .A1(n2511), .A2(n3085), .ZN(n2532) );
  NAND2_X1 U2932 ( .A1(n4010), .A2(n2956), .ZN(n2925) );
  AND2_X1 U2933 ( .A1(n2709), .A2(REG3_REG_19__SCAN_IN), .ZN(n2721) );
  AND2_X1 U2934 ( .A1(n2550), .A2(REG3_REG_10__SCAN_IN), .ZN(n2566) );
  INV_X1 U2935 ( .A(n3239), .ZN(n3815) );
  AND2_X1 U2936 ( .A1(n3787), .A2(DATAI_20_), .ZN(n4075) );
  AND2_X1 U2937 ( .A1(n4311), .A2(n3021), .ZN(n4109) );
  OR2_X1 U2938 ( .A1(n2608), .A2(n2607), .ZN(n2623) );
  NOR2_X1 U2939 ( .A1(n2617), .A2(n2616), .ZN(n2632) );
  NOR2_X1 U2940 ( .A1(n2861), .A2(n4551), .ZN(n2862) );
  OR2_X1 U2941 ( .A1(n2580), .A2(n2579), .ZN(n2599) );
  NOR2_X1 U2942 ( .A1(n2532), .A2(n2531), .ZN(n2550) );
  NAND2_X1 U2943 ( .A1(n2721), .A2(REG3_REG_20__SCAN_IN), .ZN(n2733) );
  NOR2_X1 U2944 ( .A1(n2747), .A2(n4850), .ZN(n2756) );
  NAND2_X1 U2945 ( .A1(n2632), .A2(REG3_REG_15__SCAN_IN), .ZN(n2670) );
  OR2_X1 U2946 ( .A1(n2800), .A2(n4844), .ZN(n2811) );
  INV_X1 U2947 ( .A(n2881), .ZN(n2672) );
  NOR2_X1 U2948 ( .A1(n4286), .A2(n4349), .ZN(n4360) );
  NOR2_X1 U2949 ( .A1(n4294), .A2(n4391), .ZN(n4403) );
  INV_X1 U2950 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3689) );
  AND2_X1 U2951 ( .A1(n2960), .A2(n3781), .ZN(n3933) );
  AND2_X1 U2952 ( .A1(n4005), .A2(n4003), .ZN(n4041) );
  INV_X1 U2953 ( .A(n3547), .ZN(n2915) );
  OR2_X1 U2954 ( .A1(n4311), .A2(n2964), .ZN(n4112) );
  INV_X1 U2955 ( .A(n4316), .ZN(n4146) );
  OR2_X1 U2956 ( .A1(n3024), .A2(n2970), .ZN(n4096) );
  AND2_X1 U2957 ( .A1(n2963), .A2(n2962), .ZN(n4139) );
  INV_X1 U2958 ( .A(n4109), .ZN(n4133) );
  INV_X1 U2959 ( .A(n3115), .ZN(n3145) );
  OR2_X1 U2960 ( .A1(n2541), .A2(IR_REG_9__SCAN_IN), .ZN(n2608) );
  NAND2_X1 U2961 ( .A1(n2882), .A2(n4311), .ZN(n4543) );
  XNOR2_X1 U2962 ( .A(n2405), .B(n2406), .ZN(n3120) );
  INV_X1 U2963 ( .A(n4131), .ZN(n4141) );
  INV_X1 U2964 ( .A(n3493), .ZN(n3485) );
  OR2_X1 U2965 ( .A1(n2812), .A2(n2822), .ZN(n3939) );
  INV_X1 U2966 ( .A(n4441), .ZN(n4433) );
  INV_X1 U2967 ( .A(n4311), .ZN(n3897) );
  AND2_X1 U2968 ( .A1(n4087), .A2(n4085), .ZN(n4107) );
  AND2_X1 U2969 ( .A1(n3734), .A2(n3731), .ZN(n3810) );
  INV_X1 U2970 ( .A(n4096), .ZN(n4453) );
  NAND2_X1 U2971 ( .A1(n2841), .A2(n2840), .ZN(n3211) );
  INV_X1 U2972 ( .A(n4517), .ZN(n4480) );
  INV_X1 U2973 ( .A(n4496), .ZN(n4501) );
  INV_X1 U2974 ( .A(n3211), .ZN(n2979) );
  INV_X1 U2975 ( .A(n4461), .ZN(n3878) );
  XNOR2_X1 U2976 ( .A(n2854), .B(n2853), .ZN(n3023) );
  NOR2_X2 U2977 ( .A1(n3035), .A2(n3034), .ZN(n4440) );
  NAND2_X1 U2978 ( .A1(n2893), .A2(n2863), .ZN(n2891) );
  INV_X1 U2979 ( .A(n3678), .ZN(n4551) );
  INV_X1 U2980 ( .A(n3930), .ZN(n3886) );
  OR2_X1 U2981 ( .A1(n4325), .A2(n4322), .ZN(n4436) );
  OR2_X1 U2982 ( .A1(n4325), .A2(n3897), .ZN(n4448) );
  NAND2_X1 U2983 ( .A1(n4125), .A2(n3283), .ZN(n4149) );
  NAND2_X1 U2984 ( .A1(n4533), .A2(n4506), .ZN(n4211) );
  OR2_X1 U2985 ( .A1(n3918), .A2(n4249), .ZN(n2982) );
  NAND2_X1 U2986 ( .A1(n4520), .A2(n4506), .ZN(n4249) );
  OR2_X1 U2987 ( .A1(n2980), .A2(n2979), .ZN(n4518) );
  INV_X1 U2988 ( .A(n4459), .ZN(n4460) );
  INV_X1 U2989 ( .A(n4292), .ZN(n4468) );
  XNOR2_X1 U2990 ( .A(n2517), .B(IR_REG_7__SCAN_IN), .ZN(n4259) );
  NAND4_X1 U2991 ( .A1(n2605), .A2(n2337), .A3(n2336), .A4(n2335), .ZN(n2677)
         );
  NAND2_X1 U2992 ( .A1(n2539), .A2(n2338), .ZN(n2339) );
  NAND2_X1 U2993 ( .A1(n2467), .A2(n2340), .ZN(n2341) );
  NOR2_X2 U2994 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2416)
         );
  NAND2_X1 U2995 ( .A1(n2416), .A2(n4663), .ZN(n2436) );
  NAND2_X1 U2996 ( .A1(n2349), .A2(n2346), .ZN(n2348) );
  INV_X1 U2997 ( .A(n4252), .ZN(n2352) );
  AND2_X2 U2998 ( .A1(n2352), .A2(n4253), .ZN(n2411) );
  NAND2_X1 U2999 ( .A1(n2411), .A2(REG1_REG_0__SCAN_IN), .ZN(n2358) );
  NAND2_X2 U3000 ( .A1(n2352), .A2(n2354), .ZN(n2395) );
  INV_X1 U3001 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2353) );
  NAND2_X1 U3002 ( .A1(n4253), .A2(n4252), .ZN(n2792) );
  NAND2_X1 U3003 ( .A1(n2429), .A2(REG3_REG_0__SCAN_IN), .ZN(n2356) );
  NAND2_X1 U3004 ( .A1(n2431), .A2(REG2_REG_0__SCAN_IN), .ZN(n2355) );
  NAND2_X1 U3005 ( .A1(n2360), .A2(IR_REG_31__SCAN_IN), .ZN(n2854) );
  NAND2_X1 U3006 ( .A1(n2854), .A2(n2853), .ZN(n2361) );
  NAND2_X1 U3007 ( .A1(n2361), .A2(IR_REG_31__SCAN_IN), .ZN(n2362) );
  NAND2_X1 U3008 ( .A1(n2363), .A2(IR_REG_31__SCAN_IN), .ZN(n2364) );
  NAND2_X2 U3009 ( .A1(n4254), .A2(n2365), .ZN(n2984) );
  NAND2_X1 U3010 ( .A1(n2366), .A2(IR_REG_31__SCAN_IN), .ZN(n2389) );
  NAND2_X1 U3011 ( .A1(n2389), .A2(n2388), .ZN(n2391) );
  NAND2_X1 U3012 ( .A1(n2391), .A2(IR_REG_31__SCAN_IN), .ZN(n2368) );
  NAND2_X1 U3013 ( .A1(n2369), .A2(IR_REG_31__SCAN_IN), .ZN(n2370) );
  INV_X1 U3014 ( .A(n3216), .ZN(n2371) );
  AND2_X2 U3015 ( .A1(n2984), .A2(n2371), .ZN(n2742) );
  INV_X1 U3016 ( .A(n2742), .ZN(n2372) );
  NAND2_X1 U3017 ( .A1(n2378), .A2(IR_REG_28__SCAN_IN), .ZN(n2379) );
  NAND2_X2 U3018 ( .A1(n2380), .A2(n2379), .ZN(n2401) );
  MUX2_X1 U3019 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2401), .Z(n3115) );
  AND2_X4 U3020 ( .A1(n2984), .A2(n3216), .ZN(n2816) );
  AND2_X1 U3021 ( .A1(n3115), .A2(n2816), .ZN(n2381) );
  INV_X1 U3022 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2382) );
  OR2_X1 U3023 ( .A1(n2984), .A2(n2382), .ZN(n2383) );
  NAND2_X1 U3024 ( .A1(n2392), .A2(n2383), .ZN(n3113) );
  INV_X1 U3025 ( .A(n3880), .ZN(n2866) );
  INV_X1 U3026 ( .A(n4256), .ZN(n2867) );
  NAND2_X1 U3027 ( .A1(n3895), .A2(n2651), .ZN(n2387) );
  INV_X1 U3028 ( .A(IR_REG_0__SCAN_IN), .ZN(n4830) );
  NOR2_X1 U3029 ( .A1(n2984), .A2(n4830), .ZN(n2385) );
  AOI21_X1 U3030 ( .B1(n3115), .B2(n2742), .A(n2385), .ZN(n2386) );
  NAND2_X1 U3031 ( .A1(n2387), .A2(n2386), .ZN(n3112) );
  NAND2_X1 U3032 ( .A1(n3113), .A2(n3112), .ZN(n2394) );
  OR2_X1 U3033 ( .A1(n2389), .A2(n2388), .ZN(n2390) );
  NAND2_X1 U3034 ( .A1(n3880), .A2(n4305), .ZN(n3877) );
  NAND2_X1 U3035 ( .A1(n2392), .A2(n2832), .ZN(n2393) );
  NAND2_X1 U3036 ( .A1(n2394), .A2(n2393), .ZN(n3121) );
  INV_X1 U3037 ( .A(n2395), .ZN(n2410) );
  NAND2_X1 U3038 ( .A1(n2431), .A2(REG2_REG_1__SCAN_IN), .ZN(n2397) );
  NAND2_X1 U3039 ( .A1(n3155), .A2(n2742), .ZN(n2403) );
  NAND2_X1 U3040 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2400)
         );
  MUX2_X1 U3041 ( .A(n2154), .B(DATAI_1_), .S(n2401), .Z(n3122) );
  NAND2_X1 U3042 ( .A1(n3122), .A2(n2816), .ZN(n2402) );
  NAND2_X1 U3043 ( .A1(n2403), .A2(n2402), .ZN(n2404) );
  AOI22_X1 U3044 ( .A1(n3155), .A2(n2651), .B1(n2742), .B2(n3122), .ZN(n2406)
         );
  NAND2_X1 U3045 ( .A1(n3121), .A2(n3120), .ZN(n2409) );
  INV_X1 U3046 ( .A(n2406), .ZN(n2407) );
  NAND2_X1 U3047 ( .A1(n2405), .A2(n2407), .ZN(n2408) );
  NAND2_X1 U3048 ( .A1(n2409), .A2(n2408), .ZN(n3150) );
  INV_X1 U3049 ( .A(n3150), .ZN(n2427) );
  NAND2_X1 U3050 ( .A1(n2410), .A2(REG0_REG_2__SCAN_IN), .ZN(n2415) );
  NAND2_X1 U3051 ( .A1(n2429), .A2(REG3_REG_2__SCAN_IN), .ZN(n2414) );
  NAND2_X1 U3052 ( .A1(n2411), .A2(REG1_REG_2__SCAN_IN), .ZN(n2413) );
  NAND2_X1 U3053 ( .A1(n2431), .A2(REG2_REG_2__SCAN_IN), .ZN(n2412) );
  NAND2_X1 U3054 ( .A1(n3173), .A2(n2815), .ZN(n2419) );
  MUX2_X1 U3055 ( .A(n3028), .B(DATAI_2_), .S(n2401), .Z(n3193) );
  NAND2_X1 U3056 ( .A1(n3193), .A2(n2816), .ZN(n2418) );
  NAND2_X1 U3057 ( .A1(n2419), .A2(n2418), .ZN(n2420) );
  AOI22_X1 U3058 ( .A1(n3173), .A2(n2651), .B1(n2742), .B2(n3193), .ZN(n2422)
         );
  INV_X1 U3059 ( .A(n2421), .ZN(n2424) );
  INV_X1 U3060 ( .A(n2422), .ZN(n2423) );
  NAND2_X1 U3061 ( .A1(n2424), .A2(n2423), .ZN(n2425) );
  NAND2_X1 U3062 ( .A1(n2428), .A2(n2425), .ZN(n3153) );
  INV_X1 U3063 ( .A(n3153), .ZN(n2426) );
  NAND2_X1 U3064 ( .A1(n2427), .A2(n2426), .ZN(n3151) );
  NAND2_X1 U3065 ( .A1(n3151), .A2(n2428), .ZN(n3171) );
  INV_X1 U3066 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2430) );
  NAND2_X1 U3067 ( .A1(n2773), .A2(n2430), .ZN(n2435) );
  NAND2_X1 U3068 ( .A1(n2877), .A2(REG0_REG_3__SCAN_IN), .ZN(n2434) );
  NAND2_X1 U3069 ( .A1(n2672), .A2(REG2_REG_3__SCAN_IN), .ZN(n2433) );
  NAND2_X1 U3070 ( .A1(n2411), .A2(REG1_REG_3__SCAN_IN), .ZN(n2432) );
  NAND2_X1 U3071 ( .A1(n3894), .A2(n2804), .ZN(n2440) );
  NAND2_X1 U3072 ( .A1(n2436), .A2(IR_REG_31__SCAN_IN), .ZN(n2437) );
  NAND2_X1 U3073 ( .A1(n2437), .A2(n2467), .ZN(n2447) );
  OR2_X1 U3074 ( .A1(n2437), .A2(n2467), .ZN(n2438) );
  MUX2_X1 U3075 ( .A(n4262), .B(DATAI_3_), .S(n2401), .Z(n3220) );
  NAND2_X1 U3076 ( .A1(n3220), .A2(n2816), .ZN(n2439) );
  NAND2_X1 U3077 ( .A1(n2440), .A2(n2439), .ZN(n2441) );
  XNOR2_X1 U3078 ( .A(n2441), .B(n2819), .ZN(n2452) );
  AOI22_X1 U3079 ( .A1(n3894), .A2(n2651), .B1(n2742), .B2(n3220), .ZN(n2453)
         );
  XNOR2_X1 U3080 ( .A(n2452), .B(n2453), .ZN(n3172) );
  NAND2_X1 U3081 ( .A1(n3171), .A2(n3172), .ZN(n3160) );
  NOR2_X1 U3082 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2442) );
  NOR2_X1 U3083 ( .A1(n2460), .A2(n2442), .ZN(n3253) );
  NAND2_X1 U3084 ( .A1(n2773), .A2(n3253), .ZN(n2446) );
  NAND2_X1 U3085 ( .A1(n2877), .A2(REG0_REG_4__SCAN_IN), .ZN(n2445) );
  NAND2_X1 U3086 ( .A1(n2411), .A2(REG1_REG_4__SCAN_IN), .ZN(n2444) );
  NAND2_X1 U3087 ( .A1(n2672), .A2(REG2_REG_4__SCAN_IN), .ZN(n2443) );
  NAND2_X1 U3088 ( .A1(n3893), .A2(n2804), .ZN(n2450) );
  NAND2_X1 U3089 ( .A1(n2447), .A2(IR_REG_31__SCAN_IN), .ZN(n2448) );
  MUX2_X1 U3090 ( .A(n4336), .B(DATAI_4_), .S(n2401), .Z(n3252) );
  NAND2_X1 U3091 ( .A1(n3252), .A2(n2816), .ZN(n2449) );
  NAND2_X1 U3092 ( .A1(n2450), .A2(n2449), .ZN(n2451) );
  AOI22_X1 U3093 ( .A1(n3893), .A2(n2651), .B1(n2742), .B2(n3252), .ZN(n2457)
         );
  XNOR2_X1 U3094 ( .A(n2456), .B(n2457), .ZN(n3161) );
  INV_X1 U3095 ( .A(n2452), .ZN(n2454) );
  NAND2_X1 U3096 ( .A1(n2454), .A2(n2453), .ZN(n3162) );
  AND2_X1 U3097 ( .A1(n3161), .A2(n3162), .ZN(n2455) );
  NAND2_X1 U3098 ( .A1(n3160), .A2(n2455), .ZN(n3159) );
  NAND2_X1 U3099 ( .A1(n3159), .A2(n2459), .ZN(n3203) );
  NAND2_X1 U3100 ( .A1(n2460), .A2(REG3_REG_5__SCAN_IN), .ZN(n2481) );
  OAI21_X1 U3101 ( .B1(n2460), .B2(REG3_REG_5__SCAN_IN), .A(n2481), .ZN(n2461)
         );
  INV_X1 U3102 ( .A(n2461), .ZN(n3302) );
  NAND2_X1 U3103 ( .A1(n2773), .A2(n3302), .ZN(n2465) );
  NAND2_X1 U3104 ( .A1(n2877), .A2(REG0_REG_5__SCAN_IN), .ZN(n2464) );
  NAND2_X1 U3105 ( .A1(n3783), .A2(REG1_REG_5__SCAN_IN), .ZN(n2463) );
  INV_X2 U3106 ( .A(n2881), .ZN(n2693) );
  NAND2_X1 U3107 ( .A1(n2693), .A2(REG2_REG_5__SCAN_IN), .ZN(n2462) );
  NAND4_X1 U3108 ( .A1(n2465), .A2(n2464), .A3(n2463), .A4(n2462), .ZN(n3277)
         );
  NAND2_X1 U3109 ( .A1(n3277), .A2(n2804), .ZN(n2473) );
  NAND2_X1 U3110 ( .A1(n2467), .A2(n2466), .ZN(n2468) );
  NAND2_X1 U3111 ( .A1(n2176), .A2(IR_REG_31__SCAN_IN), .ZN(n2470) );
  INV_X1 U3112 ( .A(IR_REG_5__SCAN_IN), .ZN(n2469) );
  XNOR2_X1 U3113 ( .A(n2470), .B(n2469), .ZN(n3061) );
  INV_X1 U3114 ( .A(DATAI_5_), .ZN(n2471) );
  MUX2_X1 U3115 ( .A(n3061), .B(n2471), .S(n3787), .Z(n2938) );
  NAND2_X1 U3116 ( .A1(n3301), .A2(n2816), .ZN(n2472) );
  NAND2_X1 U3117 ( .A1(n2473), .A2(n2472), .ZN(n2474) );
  XNOR2_X1 U3118 ( .A(n2474), .B(n2819), .ZN(n2478) );
  NOR2_X1 U3119 ( .A1(n2938), .A2(n3879), .ZN(n2475) );
  AOI21_X1 U3120 ( .B1(n3277), .B2(n2651), .A(n2475), .ZN(n2476) );
  XNOR2_X1 U3121 ( .A(n2478), .B(n2476), .ZN(n3204) );
  INV_X1 U3122 ( .A(n2476), .ZN(n2477) );
  NAND2_X1 U3123 ( .A1(n2478), .A2(n2477), .ZN(n2479) );
  AND2_X1 U3124 ( .A1(n2481), .A2(n3036), .ZN(n2482) );
  NOR2_X1 U3125 ( .A1(n2497), .A2(n2482), .ZN(n3286) );
  NAND2_X1 U3126 ( .A1(n2773), .A2(n3286), .ZN(n2486) );
  NAND2_X1 U3127 ( .A1(n2877), .A2(REG0_REG_6__SCAN_IN), .ZN(n2485) );
  NAND2_X1 U3128 ( .A1(n3783), .A2(REG1_REG_6__SCAN_IN), .ZN(n2484) );
  NAND2_X1 U3129 ( .A1(n2693), .A2(REG2_REG_6__SCAN_IN), .ZN(n2483) );
  NAND4_X1 U3130 ( .A1(n2486), .A2(n2485), .A3(n2484), .A4(n2483), .ZN(n3892)
         );
  NAND2_X1 U3131 ( .A1(n3892), .A2(n2815), .ZN(n2489) );
  OR2_X1 U3132 ( .A1(n2681), .A2(n2373), .ZN(n2487) );
  XNOR2_X1 U3133 ( .A(n2487), .B(IR_REG_6__SCAN_IN), .ZN(n4260) );
  MUX2_X1 U3134 ( .A(n4260), .B(DATAI_6_), .S(n3787), .Z(n3276) );
  NAND2_X1 U3135 ( .A1(n3276), .A2(n2816), .ZN(n2488) );
  NAND2_X1 U3136 ( .A1(n2489), .A2(n2488), .ZN(n2490) );
  XNOR2_X1 U3137 ( .A(n2490), .B(n2819), .ZN(n2493) );
  NAND2_X1 U3138 ( .A1(n3892), .A2(n2651), .ZN(n2492) );
  NAND2_X1 U3139 ( .A1(n3276), .A2(n2742), .ZN(n2491) );
  NAND2_X1 U3140 ( .A1(n2492), .A2(n2491), .ZN(n2494) );
  AND2_X1 U3141 ( .A1(n2493), .A2(n2494), .ZN(n3260) );
  INV_X1 U3142 ( .A(n2493), .ZN(n2496) );
  INV_X1 U3143 ( .A(n2494), .ZN(n2495) );
  NAND2_X1 U3144 ( .A1(n2496), .A2(n2495), .ZN(n3259) );
  NAND2_X1 U3145 ( .A1(n2497), .A2(REG3_REG_7__SCAN_IN), .ZN(n2511) );
  OR2_X1 U3146 ( .A1(n2497), .A2(REG3_REG_7__SCAN_IN), .ZN(n2498) );
  AND2_X1 U3147 ( .A1(n2511), .A2(n2498), .ZN(n3312) );
  NAND2_X1 U31480 ( .A1(n2773), .A2(n3312), .ZN(n2502) );
  NAND2_X1 U31490 ( .A1(n2877), .A2(REG0_REG_7__SCAN_IN), .ZN(n2501) );
  NAND2_X1 U3150 ( .A1(n3783), .A2(REG1_REG_7__SCAN_IN), .ZN(n2500) );
  NAND2_X1 U3151 ( .A1(n2693), .A2(REG2_REG_7__SCAN_IN), .ZN(n2499) );
  NAND4_X1 U3152 ( .A1(n2502), .A2(n2501), .A3(n2500), .A4(n2499), .ZN(n4539)
         );
  NAND2_X1 U3153 ( .A1(n4539), .A2(n2742), .ZN(n2505) );
  AND2_X1 U3154 ( .A1(n2681), .A2(n2538), .ZN(n2503) );
  MUX2_X1 U3155 ( .A(n4259), .B(DATAI_7_), .S(n3787), .Z(n3331) );
  NAND2_X1 U3156 ( .A1(n3331), .A2(n2816), .ZN(n2504) );
  NAND2_X1 U3157 ( .A1(n2505), .A2(n2504), .ZN(n2506) );
  XNOR2_X1 U3158 ( .A(n2506), .B(n2832), .ZN(n2507) );
  AOI22_X1 U3159 ( .A1(n4539), .A2(n2651), .B1(n2742), .B2(n3331), .ZN(n2508)
         );
  XNOR2_X1 U3160 ( .A(n2507), .B(n2508), .ZN(n3330) );
  INV_X1 U3161 ( .A(n2507), .ZN(n2510) );
  INV_X1 U3162 ( .A(n2508), .ZN(n2509) );
  NAND2_X1 U3163 ( .A1(n2511), .A2(n3085), .ZN(n2512) );
  AND2_X1 U3164 ( .A1(n2532), .A2(n2512), .ZN(n4548) );
  NAND2_X1 U3165 ( .A1(n2773), .A2(n4548), .ZN(n2516) );
  NAND2_X1 U3166 ( .A1(n2877), .A2(REG0_REG_8__SCAN_IN), .ZN(n2515) );
  NAND2_X1 U3167 ( .A1(n3783), .A2(REG1_REG_8__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U3168 ( .A1(n2693), .A2(REG2_REG_8__SCAN_IN), .ZN(n2513) );
  NAND4_X1 U3169 ( .A1(n2516), .A2(n2515), .A3(n2514), .A4(n2513), .ZN(n3891)
         );
  NAND2_X1 U3170 ( .A1(n3891), .A2(n2815), .ZN(n2523) );
  INV_X1 U3171 ( .A(IR_REG_7__SCAN_IN), .ZN(n4713) );
  NAND2_X1 U3172 ( .A1(n2517), .A2(n4713), .ZN(n2518) );
  NAND2_X1 U3173 ( .A1(n2518), .A2(IR_REG_31__SCAN_IN), .ZN(n2520) );
  INV_X1 U3174 ( .A(IR_REG_8__SCAN_IN), .ZN(n2519) );
  XNOR2_X1 U3175 ( .A(n2520), .B(n2519), .ZN(n4280) );
  INV_X1 U3176 ( .A(DATAI_8_), .ZN(n2521) );
  MUX2_X1 U3177 ( .A(n4280), .B(n2521), .S(n3787), .Z(n3340) );
  NAND2_X1 U3178 ( .A1(n4541), .A2(n2816), .ZN(n2522) );
  NAND2_X1 U3179 ( .A1(n2523), .A2(n2522), .ZN(n2524) );
  XNOR2_X1 U3180 ( .A(n2524), .B(n2819), .ZN(n2527) );
  NAND2_X1 U3181 ( .A1(n3891), .A2(n2651), .ZN(n2526) );
  NAND2_X1 U3182 ( .A1(n4541), .A2(n2815), .ZN(n2525) );
  NAND2_X1 U3183 ( .A1(n2526), .A2(n2525), .ZN(n2528) );
  AND2_X1 U3184 ( .A1(n2527), .A2(n2528), .ZN(n4535) );
  INV_X1 U3185 ( .A(n2527), .ZN(n2530) );
  INV_X1 U3186 ( .A(n2528), .ZN(n2529) );
  NAND2_X1 U3187 ( .A1(n2530), .A2(n2529), .ZN(n4534) );
  AND2_X1 U3188 ( .A1(n2532), .A2(n2531), .ZN(n2533) );
  NOR2_X1 U3189 ( .A1(n2550), .A2(n2533), .ZN(n3366) );
  NAND2_X1 U3190 ( .A1(n2773), .A2(n3366), .ZN(n2537) );
  NAND2_X1 U3191 ( .A1(n2877), .A2(REG0_REG_9__SCAN_IN), .ZN(n2536) );
  NAND2_X1 U3192 ( .A1(n3783), .A2(REG1_REG_9__SCAN_IN), .ZN(n2535) );
  NAND2_X1 U3193 ( .A1(n2693), .A2(REG2_REG_9__SCAN_IN), .ZN(n2534) );
  NAND4_X1 U3194 ( .A1(n2537), .A2(n2536), .A3(n2535), .A4(n2534), .ZN(n3103)
         );
  NAND2_X1 U3195 ( .A1(n3103), .A2(n2815), .ZN(n2544) );
  AND2_X1 U3196 ( .A1(n2539), .A2(n2538), .ZN(n2678) );
  NAND2_X1 U3197 ( .A1(n2681), .A2(n2678), .ZN(n2541) );
  NAND2_X1 U3198 ( .A1(n2541), .A2(IR_REG_31__SCAN_IN), .ZN(n2540) );
  MUX2_X1 U3199 ( .A(IR_REG_31__SCAN_IN), .B(n2540), .S(IR_REG_9__SCAN_IN), 
        .Z(n2542) );
  MUX2_X1 U3200 ( .A(n4283), .B(DATAI_9_), .S(n3787), .Z(n3365) );
  NAND2_X1 U3201 ( .A1(n3365), .A2(n2816), .ZN(n2543) );
  NAND2_X1 U3202 ( .A1(n2544), .A2(n2543), .ZN(n2545) );
  XNOR2_X1 U3203 ( .A(n2545), .B(n2819), .ZN(n2546) );
  AOI22_X1 U3204 ( .A1(n3103), .A2(n2651), .B1(n2742), .B2(n3365), .ZN(n2547)
         );
  XNOR2_X1 U3205 ( .A(n2546), .B(n2547), .ZN(n3352) );
  INV_X1 U3206 ( .A(n2546), .ZN(n2548) );
  NAND2_X1 U3207 ( .A1(n2548), .A2(n2547), .ZN(n2549) );
  NOR2_X1 U3208 ( .A1(n2550), .A2(REG3_REG_10__SCAN_IN), .ZN(n2551) );
  OR2_X1 U3209 ( .A1(n2566), .A2(n2551), .ZN(n3397) );
  INV_X1 U32100 ( .A(n3397), .ZN(n3408) );
  NAND2_X1 U32110 ( .A1(n2773), .A2(n3408), .ZN(n2555) );
  NAND2_X1 U32120 ( .A1(n2877), .A2(REG0_REG_10__SCAN_IN), .ZN(n2554) );
  NAND2_X1 U32130 ( .A1(n3783), .A2(REG1_REG_10__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U32140 ( .A1(n2693), .A2(REG2_REG_10__SCAN_IN), .ZN(n2552) );
  NAND4_X1 U32150 ( .A1(n2555), .A2(n2554), .A3(n2553), .A4(n2552), .ZN(n3890)
         );
  NAND2_X1 U32160 ( .A1(n3890), .A2(n2815), .ZN(n2558) );
  NAND2_X1 U32170 ( .A1(n2608), .A2(IR_REG_31__SCAN_IN), .ZN(n2556) );
  XNOR2_X1 U32180 ( .A(n2556), .B(IR_REG_10__SCAN_IN), .ZN(n4285) );
  MUX2_X1 U32190 ( .A(n4285), .B(DATAI_10_), .S(n3787), .Z(n3390) );
  NAND2_X1 U32200 ( .A1(n3390), .A2(n2816), .ZN(n2557) );
  NAND2_X1 U32210 ( .A1(n2558), .A2(n2557), .ZN(n2559) );
  XNOR2_X1 U32220 ( .A(n2559), .B(n2832), .ZN(n2561) );
  AOI22_X1 U32230 ( .A1(n3890), .A2(n2651), .B1(n2742), .B2(n3390), .ZN(n2562)
         );
  XNOR2_X1 U32240 ( .A(n2561), .B(n2562), .ZN(n3406) );
  INV_X1 U32250 ( .A(n2561), .ZN(n2564) );
  INV_X1 U32260 ( .A(n2562), .ZN(n2563) );
  NAND2_X1 U32270 ( .A1(n2564), .A2(n2563), .ZN(n2565) );
  NAND2_X1 U32280 ( .A1(n3403), .A2(n2565), .ZN(n3382) );
  OR2_X1 U32290 ( .A1(n2566), .A2(REG3_REG_11__SCAN_IN), .ZN(n2567) );
  AND2_X1 U32300 ( .A1(n2580), .A2(n2567), .ZN(n3432) );
  NAND2_X1 U32310 ( .A1(n2773), .A2(n3432), .ZN(n2571) );
  NAND2_X1 U32320 ( .A1(n2877), .A2(REG0_REG_11__SCAN_IN), .ZN(n2570) );
  NAND2_X1 U32330 ( .A1(n3783), .A2(REG1_REG_11__SCAN_IN), .ZN(n2569) );
  NAND2_X1 U32340 ( .A1(n2693), .A2(REG2_REG_11__SCAN_IN), .ZN(n2568) );
  NAND4_X1 U32350 ( .A1(n2571), .A2(n2570), .A3(n2569), .A4(n2568), .ZN(n3442)
         );
  NAND2_X1 U32360 ( .A1(n3442), .A2(n2651), .ZN(n2573) );
  OAI21_X1 U32370 ( .B1(n2608), .B2(IR_REG_10__SCAN_IN), .A(IR_REG_31__SCAN_IN), .ZN(n2587) );
  XNOR2_X1 U32380 ( .A(n2587), .B(IR_REG_11__SCAN_IN), .ZN(n4287) );
  MUX2_X1 U32390 ( .A(n4287), .B(DATAI_11_), .S(n3787), .Z(n3425) );
  NAND2_X1 U32400 ( .A1(n3425), .A2(n2815), .ZN(n2572) );
  NAND2_X1 U32410 ( .A1(n2573), .A2(n2572), .ZN(n3380) );
  NAND2_X1 U32420 ( .A1(n3442), .A2(n2804), .ZN(n2575) );
  NAND2_X1 U32430 ( .A1(n3425), .A2(n2816), .ZN(n2574) );
  NAND2_X1 U32440 ( .A1(n2575), .A2(n2574), .ZN(n2576) );
  XNOR2_X1 U32450 ( .A(n2576), .B(n2819), .ZN(n3379) );
  OAI21_X1 U32460 ( .B1(n3382), .B2(n3380), .A(n3379), .ZN(n2578) );
  NAND2_X1 U32470 ( .A1(n3382), .A2(n3380), .ZN(n2577) );
  NAND2_X1 U32480 ( .A1(n2578), .A2(n2577), .ZN(n3413) );
  NAND2_X1 U32490 ( .A1(n2580), .A2(n2579), .ZN(n2581) );
  AND2_X1 U32500 ( .A1(n2599), .A2(n2581), .ZN(n3452) );
  NAND2_X1 U32510 ( .A1(n2773), .A2(n3452), .ZN(n2585) );
  NAND2_X1 U32520 ( .A1(n2877), .A2(REG0_REG_12__SCAN_IN), .ZN(n2584) );
  NAND2_X1 U32530 ( .A1(n3783), .A2(REG1_REG_12__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U32540 ( .A1(n2693), .A2(REG2_REG_12__SCAN_IN), .ZN(n2582) );
  NAND4_X1 U32550 ( .A1(n2585), .A2(n2584), .A3(n2583), .A4(n2582), .ZN(n3889)
         );
  NAND2_X1 U32560 ( .A1(n3889), .A2(n2804), .ZN(n2591) );
  INV_X1 U32570 ( .A(IR_REG_11__SCAN_IN), .ZN(n2586) );
  NAND2_X1 U32580 ( .A1(n2587), .A2(n2586), .ZN(n2588) );
  NAND2_X1 U32590 ( .A1(n2588), .A2(IR_REG_31__SCAN_IN), .ZN(n2589) );
  XNOR2_X1 U32600 ( .A(n2589), .B(IR_REG_12__SCAN_IN), .ZN(n4288) );
  MUX2_X1 U32610 ( .A(n4288), .B(DATAI_12_), .S(n3787), .Z(n3449) );
  NAND2_X1 U32620 ( .A1(n3449), .A2(n2816), .ZN(n2590) );
  NAND2_X1 U32630 ( .A1(n2591), .A2(n2590), .ZN(n2592) );
  XNOR2_X1 U32640 ( .A(n2592), .B(n2819), .ZN(n2595) );
  NAND2_X1 U32650 ( .A1(n3889), .A2(n2651), .ZN(n2594) );
  NAND2_X1 U32660 ( .A1(n3449), .A2(n2804), .ZN(n2593) );
  NAND2_X1 U32670 ( .A1(n2594), .A2(n2593), .ZN(n2596) );
  AND2_X1 U32680 ( .A1(n2595), .A2(n2596), .ZN(n3415) );
  INV_X1 U32690 ( .A(n2595), .ZN(n2598) );
  INV_X1 U32700 ( .A(n2596), .ZN(n2597) );
  NAND2_X1 U32710 ( .A1(n2598), .A2(n2597), .ZN(n3414) );
  NAND2_X1 U32720 ( .A1(n2599), .A2(n3460), .ZN(n2600) );
  AND2_X1 U32730 ( .A1(n2617), .A2(n2600), .ZN(n3495) );
  NAND2_X1 U32740 ( .A1(n2773), .A2(n3495), .ZN(n2604) );
  NAND2_X1 U32750 ( .A1(n2877), .A2(REG0_REG_13__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U32760 ( .A1(n3783), .A2(REG1_REG_13__SCAN_IN), .ZN(n2602) );
  NAND2_X1 U32770 ( .A1(n2693), .A2(REG2_REG_13__SCAN_IN), .ZN(n2601) );
  NAND4_X1 U32780 ( .A1(n2604), .A2(n2603), .A3(n2602), .A4(n2601), .ZN(n3477)
         );
  NAND2_X1 U32790 ( .A1(n3477), .A2(n2804), .ZN(n2612) );
  INV_X1 U32800 ( .A(IR_REG_12__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U32810 ( .A1(n2605), .A2(n2606), .ZN(n2607) );
  NAND2_X1 U32820 ( .A1(n2623), .A2(IR_REG_31__SCAN_IN), .ZN(n2609) );
  XNOR2_X1 U32830 ( .A(n2609), .B(IR_REG_13__SCAN_IN), .ZN(n4292) );
  INV_X1 U32840 ( .A(DATAI_13_), .ZN(n2610) );
  MUX2_X1 U32850 ( .A(n4468), .B(n2610), .S(n3787), .Z(n3493) );
  NAND2_X1 U32860 ( .A1(n3485), .A2(n2816), .ZN(n2611) );
  NAND2_X1 U32870 ( .A1(n2612), .A2(n2611), .ZN(n2613) );
  XNOR2_X1 U32880 ( .A(n2613), .B(n2832), .ZN(n3456) );
  NAND2_X1 U32890 ( .A1(n3477), .A2(n2651), .ZN(n2615) );
  NAND2_X1 U32900 ( .A1(n3485), .A2(n2804), .ZN(n2614) );
  NAND2_X1 U32910 ( .A1(n2615), .A2(n2614), .ZN(n3457) );
  AND2_X1 U32920 ( .A1(n2617), .A2(n2616), .ZN(n2618) );
  NOR2_X1 U32930 ( .A1(n2632), .A2(n2618), .ZN(n3537) );
  NAND2_X1 U32940 ( .A1(n2773), .A2(n3537), .ZN(n2622) );
  NAND2_X1 U32950 ( .A1(n2877), .A2(REG0_REG_14__SCAN_IN), .ZN(n2621) );
  NAND2_X1 U32960 ( .A1(n3783), .A2(REG1_REG_14__SCAN_IN), .ZN(n2620) );
  NAND2_X1 U32970 ( .A1(n2693), .A2(REG2_REG_14__SCAN_IN), .ZN(n2619) );
  NAND4_X1 U32980 ( .A1(n2622), .A2(n2621), .A3(n2620), .A4(n2619), .ZN(n3888)
         );
  NAND2_X1 U32990 ( .A1(n3888), .A2(n2804), .ZN(n2626) );
  OR2_X1 U33000 ( .A1(n2639), .A2(n2373), .ZN(n2624) );
  XNOR2_X1 U33010 ( .A(n2624), .B(IR_REG_14__SCAN_IN), .ZN(n4396) );
  MUX2_X1 U33020 ( .A(n4396), .B(DATAI_14_), .S(n3787), .Z(n3511) );
  NAND2_X1 U33030 ( .A1(n3511), .A2(n2816), .ZN(n2625) );
  NAND2_X1 U33040 ( .A1(n2626), .A2(n2625), .ZN(n2627) );
  XNOR2_X1 U33050 ( .A(n2627), .B(n2832), .ZN(n2631) );
  INV_X1 U33060 ( .A(n2631), .ZN(n2629) );
  AOI22_X1 U33070 ( .A1(n3888), .A2(n2651), .B1(n2742), .B2(n3511), .ZN(n2630)
         );
  INV_X1 U33080 ( .A(n2630), .ZN(n2628) );
  NAND2_X1 U33090 ( .A1(n2629), .A2(n2628), .ZN(n3530) );
  AND2_X1 U33100 ( .A1(n2631), .A2(n2630), .ZN(n3529) );
  AOI21_X1 U33110 ( .B1(n3528), .B2(n3530), .A(n3529), .ZN(n2660) );
  OR2_X1 U33120 ( .A1(n2632), .A2(REG3_REG_15__SCAN_IN), .ZN(n2633) );
  AND2_X1 U33130 ( .A1(n2633), .A2(n2670), .ZN(n3718) );
  NAND2_X1 U33140 ( .A1(n2773), .A2(n3718), .ZN(n2637) );
  NAND2_X1 U33150 ( .A1(n2877), .A2(REG0_REG_15__SCAN_IN), .ZN(n2636) );
  NAND2_X1 U33160 ( .A1(n3783), .A2(REG1_REG_15__SCAN_IN), .ZN(n2635) );
  NAND2_X1 U33170 ( .A1(n2693), .A2(REG2_REG_15__SCAN_IN), .ZN(n2634) );
  NAND4_X1 U33180 ( .A1(n2637), .A2(n2636), .A3(n2635), .A4(n2634), .ZN(n3551)
         );
  NAND2_X1 U33190 ( .A1(n3551), .A2(n2804), .ZN(n2645) );
  INV_X1 U33200 ( .A(IR_REG_14__SCAN_IN), .ZN(n2638) );
  NAND2_X1 U33210 ( .A1(n2639), .A2(n2638), .ZN(n2640) );
  NAND2_X1 U33220 ( .A1(n2640), .A2(IR_REG_31__SCAN_IN), .ZN(n2642) );
  INV_X1 U33230 ( .A(IR_REG_15__SCAN_IN), .ZN(n2641) );
  NAND2_X1 U33240 ( .A1(n2642), .A2(n2641), .ZN(n2652) );
  OR2_X1 U33250 ( .A1(n2642), .A2(n2641), .ZN(n2643) );
  MUX2_X1 U33260 ( .A(n4296), .B(DATAI_15_), .S(n2401), .Z(n3713) );
  NAND2_X1 U33270 ( .A1(n3713), .A2(n2816), .ZN(n2644) );
  NAND2_X1 U33280 ( .A1(n2645), .A2(n2644), .ZN(n2646) );
  XNOR2_X1 U33290 ( .A(n2646), .B(n2819), .ZN(n2659) );
  NAND2_X1 U33300 ( .A1(n2660), .A2(n2659), .ZN(n3708) );
  XNOR2_X1 U33310 ( .A(n2670), .B(REG3_REG_16__SCAN_IN), .ZN(n3646) );
  NAND2_X1 U33320 ( .A1(n2773), .A2(n3646), .ZN(n2650) );
  NAND2_X1 U33330 ( .A1(n2877), .A2(REG0_REG_16__SCAN_IN), .ZN(n2649) );
  NAND2_X1 U33340 ( .A1(n3783), .A2(REG1_REG_16__SCAN_IN), .ZN(n2648) );
  NAND2_X1 U33350 ( .A1(n2693), .A2(REG2_REG_16__SCAN_IN), .ZN(n2647) );
  NAND4_X1 U33360 ( .A1(n2650), .A2(n2649), .A3(n2648), .A4(n2647), .ZN(n4136)
         );
  INV_X1 U33370 ( .A(n4136), .ZN(n3653) );
  INV_X1 U33380 ( .A(n2651), .ZN(n2834) );
  NAND2_X1 U33390 ( .A1(n2652), .A2(IR_REG_31__SCAN_IN), .ZN(n2654) );
  INV_X1 U33400 ( .A(IR_REG_16__SCAN_IN), .ZN(n2653) );
  INV_X1 U33410 ( .A(n4465), .ZN(n2655) );
  MUX2_X1 U33420 ( .A(n2655), .B(DATAI_16_), .S(n2401), .Z(n3556) );
  INV_X1 U33430 ( .A(n3556), .ZN(n3643) );
  OAI22_X1 U33440 ( .A1(n3653), .A2(n2834), .B1(n3879), .B2(n3643), .ZN(n2663)
         );
  NAND2_X1 U33450 ( .A1(n4136), .A2(n2815), .ZN(n2657) );
  NAND2_X1 U33460 ( .A1(n3556), .A2(n2816), .ZN(n2656) );
  NAND2_X1 U33470 ( .A1(n2657), .A2(n2656), .ZN(n2658) );
  XNOR2_X1 U33480 ( .A(n2658), .B(n2819), .ZN(n2662) );
  XOR2_X1 U33490 ( .A(n2663), .B(n2662), .Z(n3640) );
  AND2_X1 U33500 ( .A1(n3713), .A2(n2804), .ZN(n2661) );
  AOI21_X1 U33510 ( .B1(n3551), .B2(n2651), .A(n2661), .ZN(n3710) );
  INV_X1 U33520 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2668) );
  INV_X1 U3353 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2667) );
  OAI21_X1 U33540 ( .B1(n2670), .B2(n2668), .A(n2667), .ZN(n2671) );
  NAND2_X1 U3355 ( .A1(REG3_REG_16__SCAN_IN), .A2(REG3_REG_17__SCAN_IN), .ZN(
        n2669) );
  AND2_X1 U3356 ( .A1(n2671), .A2(n2691), .ZN(n4144) );
  NAND2_X1 U3357 ( .A1(n2773), .A2(n4144), .ZN(n2676) );
  NAND2_X1 U3358 ( .A1(n2877), .A2(REG0_REG_17__SCAN_IN), .ZN(n2675) );
  NAND2_X1 U3359 ( .A1(n3783), .A2(REG1_REG_17__SCAN_IN), .ZN(n2674) );
  NAND2_X1 U3360 ( .A1(n2672), .A2(REG2_REG_17__SCAN_IN), .ZN(n2673) );
  NAND4_X1 U3361 ( .A1(n2676), .A2(n2675), .A3(n2674), .A4(n2673), .ZN(n3887)
         );
  INV_X1 U3362 ( .A(n2816), .ZN(n2831) );
  INV_X1 U3363 ( .A(n2677), .ZN(n2679) );
  AND2_X1 U3364 ( .A1(n2679), .A2(n2678), .ZN(n2680) );
  NAND2_X1 U3365 ( .A1(n2681), .A2(n2680), .ZN(n2682) );
  NAND2_X1 U3366 ( .A1(n2682), .A2(IR_REG_31__SCAN_IN), .ZN(n2683) );
  XNOR2_X1 U3367 ( .A(n2683), .B(IR_REG_17__SCAN_IN), .ZN(n4299) );
  INV_X1 U3368 ( .A(n4299), .ZN(n4463) );
  INV_X1 U3369 ( .A(DATAI_17_), .ZN(n2684) );
  MUX2_X1 U3370 ( .A(n4463), .B(n2684), .S(n2401), .Z(n4131) );
  OAI22_X1 U3371 ( .A1(n4113), .A2(n3879), .B1(n2831), .B2(n4131), .ZN(n2685)
         );
  XOR2_X1 U3372 ( .A(n2819), .B(n2685), .Z(n3651) );
  INV_X1 U3373 ( .A(n3651), .ZN(n2688) );
  NAND2_X1 U3374 ( .A1(n3887), .A2(n2651), .ZN(n2687) );
  NAND2_X1 U3375 ( .A1(n4141), .A2(n2804), .ZN(n2686) );
  NAND2_X1 U3376 ( .A1(n2687), .A2(n2686), .ZN(n2689) );
  NOR2_X1 U3377 ( .A1(n2688), .A2(n2689), .ZN(n2690) );
  INV_X1 U3378 ( .A(n2689), .ZN(n3650) );
  AND2_X1 U3379 ( .A1(n2691), .A2(n3689), .ZN(n2692) );
  NOR2_X1 U3380 ( .A1(n2709), .A2(n2692), .ZN(n4121) );
  NAND2_X1 U3381 ( .A1(n2429), .A2(n4121), .ZN(n2697) );
  NAND2_X1 U3382 ( .A1(n2877), .A2(REG0_REG_18__SCAN_IN), .ZN(n2696) );
  NAND2_X1 U3383 ( .A1(n3783), .A2(REG1_REG_18__SCAN_IN), .ZN(n2695) );
  NAND2_X1 U3384 ( .A1(n2693), .A2(REG2_REG_18__SCAN_IN), .ZN(n2694) );
  NAND4_X1 U3385 ( .A1(n2697), .A2(n2696), .A3(n2695), .A4(n2694), .ZN(n4092)
         );
  NAND2_X1 U3386 ( .A1(n4092), .A2(n2804), .ZN(n2701) );
  OR2_X1 U3387 ( .A1(n2698), .A2(n2373), .ZN(n2699) );
  XNOR2_X1 U3388 ( .A(n2699), .B(IR_REG_18__SCAN_IN), .ZN(n4300) );
  MUX2_X1 U3389 ( .A(n4300), .B(DATAI_18_), .S(n2401), .Z(n4108) );
  NAND2_X1 U3390 ( .A1(n4108), .A2(n2816), .ZN(n2700) );
  NAND2_X1 U3391 ( .A1(n2701), .A2(n2700), .ZN(n2702) );
  XNOR2_X1 U3392 ( .A(n2702), .B(n2819), .ZN(n2705) );
  NAND2_X1 U3393 ( .A1(n4092), .A2(n2651), .ZN(n2704) );
  NAND2_X1 U3394 ( .A1(n4108), .A2(n2804), .ZN(n2703) );
  NAND2_X1 U3395 ( .A1(n2704), .A2(n2703), .ZN(n2706) );
  AND2_X1 U3396 ( .A1(n2705), .A2(n2706), .ZN(n3685) );
  INV_X1 U3397 ( .A(n2705), .ZN(n2708) );
  INV_X1 U3398 ( .A(n2706), .ZN(n2707) );
  NAND2_X1 U3399 ( .A1(n2708), .A2(n2707), .ZN(n3684) );
  NOR2_X1 U3400 ( .A1(n2709), .A2(REG3_REG_19__SCAN_IN), .ZN(n2710) );
  OR2_X1 U3401 ( .A1(n2721), .A2(n2710), .ZN(n4097) );
  INV_X1 U3402 ( .A(n4097), .ZN(n3617) );
  NAND2_X1 U3403 ( .A1(n2429), .A2(n3617), .ZN(n2714) );
  NAND2_X1 U3404 ( .A1(n2877), .A2(REG0_REG_19__SCAN_IN), .ZN(n2713) );
  NAND2_X1 U3405 ( .A1(n3783), .A2(REG1_REG_19__SCAN_IN), .ZN(n2712) );
  NAND2_X1 U3406 ( .A1(n2672), .A2(REG2_REG_19__SCAN_IN), .ZN(n2711) );
  NAND2_X1 U3407 ( .A1(n4110), .A2(n2804), .ZN(n2716) );
  MUX2_X1 U3408 ( .A(n2961), .B(DATAI_19_), .S(n2401), .Z(n2951) );
  NAND2_X1 U3409 ( .A1(n2951), .A2(n2816), .ZN(n2715) );
  NAND2_X1 U3410 ( .A1(n2716), .A2(n2715), .ZN(n2717) );
  XNOR2_X1 U3411 ( .A(n2717), .B(n2819), .ZN(n2718) );
  AOI22_X1 U3412 ( .A1(n4110), .A2(n2651), .B1(n2742), .B2(n2951), .ZN(n2719)
         );
  XNOR2_X1 U3413 ( .A(n2718), .B(n2719), .ZN(n3614) );
  INV_X1 U3414 ( .A(n2718), .ZN(n2720) );
  OR2_X1 U3415 ( .A1(n2721), .A2(REG3_REG_20__SCAN_IN), .ZN(n2722) );
  AND2_X1 U3416 ( .A1(n2733), .A2(n2722), .ZN(n4074) );
  NAND2_X1 U3417 ( .A1(n2773), .A2(n4074), .ZN(n2726) );
  NAND2_X1 U3418 ( .A1(n2877), .A2(REG0_REG_20__SCAN_IN), .ZN(n2725) );
  NAND2_X1 U3419 ( .A1(n3783), .A2(REG1_REG_20__SCAN_IN), .ZN(n2724) );
  NAND2_X1 U3420 ( .A1(n2693), .A2(REG2_REG_20__SCAN_IN), .ZN(n2723) );
  NAND4_X1 U3421 ( .A1(n2726), .A2(n2725), .A3(n2724), .A4(n2723), .ZN(n4044)
         );
  NAND2_X1 U3422 ( .A1(n4044), .A2(n2804), .ZN(n2728) );
  NAND2_X1 U3423 ( .A1(n4075), .A2(n2816), .ZN(n2727) );
  NAND2_X1 U3424 ( .A1(n2728), .A2(n2727), .ZN(n2729) );
  XNOR2_X1 U3425 ( .A(n2729), .B(n2832), .ZN(n2732) );
  AND2_X1 U3426 ( .A1(n4075), .A2(n2742), .ZN(n2730) );
  AOI21_X1 U3427 ( .B1(n4044), .B2(n2651), .A(n2730), .ZN(n2731) );
  NOR2_X1 U3428 ( .A1(n2732), .A2(n2731), .ZN(n3667) );
  AND2_X1 U3429 ( .A1(n2732), .A2(n2731), .ZN(n3666) );
  NAND2_X1 U3430 ( .A1(n2733), .A2(n3623), .ZN(n2734) );
  AND2_X1 U3431 ( .A1(n2747), .A2(n2734), .ZN(n4050) );
  NAND2_X1 U3432 ( .A1(n2773), .A2(n4050), .ZN(n2738) );
  NAND2_X1 U3433 ( .A1(n2877), .A2(REG0_REG_21__SCAN_IN), .ZN(n2737) );
  NAND2_X1 U3434 ( .A1(n3783), .A2(REG1_REG_21__SCAN_IN), .ZN(n2736) );
  NAND2_X1 U3435 ( .A1(n2672), .A2(REG2_REG_21__SCAN_IN), .ZN(n2735) );
  NAND4_X1 U3436 ( .A1(n2738), .A2(n2737), .A3(n2736), .A4(n2735), .ZN(n4027)
         );
  NAND2_X1 U3437 ( .A1(n4027), .A2(n2804), .ZN(n2740) );
  NAND2_X1 U3438 ( .A1(n2974), .A2(n2816), .ZN(n2739) );
  NAND2_X1 U3439 ( .A1(n2740), .A2(n2739), .ZN(n2741) );
  XNOR2_X1 U3440 ( .A(n2741), .B(n2832), .ZN(n3621) );
  AND2_X1 U3441 ( .A1(n2974), .A2(n2742), .ZN(n2743) );
  AOI21_X1 U3442 ( .B1(n4027), .B2(n2651), .A(n2743), .ZN(n2744) );
  NAND2_X1 U3443 ( .A1(n3621), .A2(n2744), .ZN(n2746) );
  INV_X1 U3444 ( .A(n3621), .ZN(n2745) );
  INV_X1 U3445 ( .A(n2744), .ZN(n3620) );
  AND2_X1 U3446 ( .A1(n2747), .A2(n4850), .ZN(n2748) );
  NOR2_X1 U3447 ( .A1(n2756), .A2(n2748), .ZN(n4033) );
  NAND2_X1 U3448 ( .A1(n2429), .A2(n4033), .ZN(n2752) );
  NAND2_X1 U3449 ( .A1(n2877), .A2(REG0_REG_22__SCAN_IN), .ZN(n2751) );
  NAND2_X1 U3450 ( .A1(n3783), .A2(REG1_REG_22__SCAN_IN), .ZN(n2750) );
  NAND2_X1 U3451 ( .A1(n2693), .A2(REG2_REG_22__SCAN_IN), .ZN(n2749) );
  NAND4_X1 U3452 ( .A1(n2752), .A2(n2751), .A3(n2750), .A4(n2749), .ZN(n4010)
         );
  OAI22_X1 U3453 ( .A1(n4042), .A2(n2834), .B1(n3879), .B2(n4034), .ZN(n2767)
         );
  NAND2_X1 U3454 ( .A1(n4010), .A2(n2804), .ZN(n2754) );
  NAND2_X1 U3455 ( .A1(n2956), .A2(n2816), .ZN(n2753) );
  NAND2_X1 U3456 ( .A1(n2754), .A2(n2753), .ZN(n2755) );
  XNOR2_X1 U3457 ( .A(n2755), .B(n2819), .ZN(n2766) );
  XOR2_X1 U34580 ( .A(n2767), .B(n2766), .Z(n3677) );
  NAND2_X1 U34590 ( .A1(n3676), .A2(n3677), .ZN(n3605) );
  NOR2_X1 U3460 ( .A1(n2756), .A2(REG3_REG_23__SCAN_IN), .ZN(n2757) );
  NOR2_X1 U3461 ( .A1(n2771), .A2(n2757), .ZN(n4017) );
  NAND2_X1 U3462 ( .A1(n2429), .A2(n4017), .ZN(n2761) );
  NAND2_X1 U3463 ( .A1(n2877), .A2(REG0_REG_23__SCAN_IN), .ZN(n2760) );
  NAND2_X1 U3464 ( .A1(n3783), .A2(REG1_REG_23__SCAN_IN), .ZN(n2759) );
  NAND2_X1 U3465 ( .A1(n2693), .A2(REG2_REG_23__SCAN_IN), .ZN(n2758) );
  NAND2_X1 U3466 ( .A1(n4028), .A2(n2804), .ZN(n2763) );
  NAND2_X1 U34670 ( .A1(n4014), .A2(n2816), .ZN(n2762) );
  NAND2_X1 U3468 ( .A1(n2763), .A2(n2762), .ZN(n2764) );
  XNOR2_X1 U34690 ( .A(n2764), .B(n2819), .ZN(n2780) );
  NOR2_X1 U3470 ( .A1(n3803), .A2(n3879), .ZN(n2765) );
  AOI21_X1 U34710 ( .B1(n4028), .B2(n2651), .A(n2765), .ZN(n2781) );
  XNOR2_X1 U3472 ( .A(n2780), .B(n2781), .ZN(n3606) );
  INV_X1 U34730 ( .A(n2766), .ZN(n2769) );
  INV_X1 U3474 ( .A(n2767), .ZN(n2768) );
  NAND2_X1 U34750 ( .A1(n2769), .A2(n2768), .ZN(n3607) );
  NAND2_X1 U3476 ( .A1(n3605), .A2(n2770), .ZN(n3604) );
  OR2_X1 U34770 ( .A1(n2771), .A2(REG3_REG_24__SCAN_IN), .ZN(n2772) );
  AND2_X1 U3478 ( .A1(n2790), .A2(n2772), .ZN(n3997) );
  NAND2_X1 U34790 ( .A1(n2773), .A2(n3997), .ZN(n2777) );
  NAND2_X1 U3480 ( .A1(n2877), .A2(REG0_REG_24__SCAN_IN), .ZN(n2776) );
  NAND2_X1 U34810 ( .A1(n3783), .A2(REG1_REG_24__SCAN_IN), .ZN(n2775) );
  NAND2_X1 U3482 ( .A1(n2672), .A2(REG2_REG_24__SCAN_IN), .ZN(n2774) );
  NAND4_X1 U34830 ( .A1(n2777), .A2(n2776), .A3(n2775), .A4(n2774), .ZN(n4009)
         );
  NAND2_X1 U3484 ( .A1(n4009), .A2(n2651), .ZN(n2779) );
  NAND2_X1 U34850 ( .A1(n3989), .A2(n2804), .ZN(n2778) );
  NAND2_X1 U3486 ( .A1(n2779), .A2(n2778), .ZN(n2786) );
  INV_X1 U34870 ( .A(n2786), .ZN(n2784) );
  INV_X1 U3488 ( .A(n2780), .ZN(n2782) );
  NOR2_X1 U34890 ( .A1(n2782), .A2(n2781), .ZN(n2787) );
  INV_X1 U3490 ( .A(n2787), .ZN(n2783) );
  NAND3_X1 U34910 ( .A1(n3604), .A2(n2784), .A3(n2783), .ZN(n3658) );
  INV_X1 U3492 ( .A(n4009), .ZN(n3634) );
  OAI22_X1 U34930 ( .A1(n3634), .A2(n3879), .B1(n2831), .B2(n3995), .ZN(n2785)
         );
  XNOR2_X1 U3494 ( .A(n2785), .B(n2819), .ZN(n3661) );
  NAND2_X1 U34950 ( .A1(n3658), .A2(n3661), .ZN(n2789) );
  INV_X1 U3496 ( .A(n3604), .ZN(n2788) );
  NAND2_X1 U34970 ( .A1(n2789), .A2(n3659), .ZN(n3630) );
  AOI22_X1 U3498 ( .A1(n2877), .A2(REG0_REG_25__SCAN_IN), .B1(n3783), .B2(
        REG1_REG_25__SCAN_IN), .ZN(n2795) );
  INV_X1 U34990 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3633) );
  NAND2_X1 U3500 ( .A1(n2790), .A2(n3633), .ZN(n2791) );
  NAND2_X1 U35010 ( .A1(n2800), .A2(n2791), .ZN(n3632) );
  NAND2_X1 U3502 ( .A1(n2672), .A2(REG2_REG_25__SCAN_IN), .ZN(n2793) );
  OAI22_X1 U35030 ( .A1(n3699), .A2(n3879), .B1(n2831), .B2(n3975), .ZN(n2796)
         );
  XNOR2_X1 U3504 ( .A(n2796), .B(n2819), .ZN(n2798) );
  OAI22_X1 U35050 ( .A1(n3699), .A2(n2834), .B1(n3879), .B2(n3975), .ZN(n2797)
         );
  OR2_X1 U35060 ( .A1(n2798), .A2(n2797), .ZN(n3629) );
  NAND2_X1 U35070 ( .A1(n3630), .A2(n3629), .ZN(n2799) );
  NAND2_X1 U35080 ( .A1(n2798), .A2(n2797), .ZN(n3628) );
  INV_X1 U35090 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4844) );
  NAND2_X1 U35100 ( .A1(n2800), .A2(n4844), .ZN(n2801) );
  NAND2_X1 U35110 ( .A1(n2811), .A2(n2801), .ZN(n3958) );
  AOI22_X1 U35120 ( .A1(n2877), .A2(REG0_REG_26__SCAN_IN), .B1(n3783), .B2(
        REG1_REG_26__SCAN_IN), .ZN(n2803) );
  NAND2_X1 U35130 ( .A1(n2672), .A2(REG2_REG_26__SCAN_IN), .ZN(n2802) );
  NAND2_X1 U35140 ( .A1(n3969), .A2(n2804), .ZN(n2806) );
  INV_X1 U35150 ( .A(n3956), .ZN(n3949) );
  NAND2_X1 U35160 ( .A1(n3949), .A2(n2816), .ZN(n2805) );
  NAND2_X1 U35170 ( .A1(n2806), .A2(n2805), .ZN(n2807) );
  XNOR2_X1 U35180 ( .A(n2807), .B(n2832), .ZN(n2810) );
  NOR2_X1 U35190 ( .A1(n3956), .A2(n3879), .ZN(n2808) );
  AOI21_X1 U35200 ( .B1(n3969), .B2(n2651), .A(n2808), .ZN(n2809) );
  NOR2_X1 U35210 ( .A1(n2810), .A2(n2809), .ZN(n3696) );
  NAND2_X1 U35220 ( .A1(n2810), .A2(n2809), .ZN(n3694) );
  INV_X1 U35230 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4847) );
  AND2_X1 U35240 ( .A1(n2811), .A2(n4847), .ZN(n2812) );
  AOI22_X1 U35250 ( .A1(n2877), .A2(REG0_REG_27__SCAN_IN), .B1(n3783), .B2(
        REG1_REG_27__SCAN_IN), .ZN(n2814) );
  NAND2_X1 U35260 ( .A1(n2693), .A2(REG2_REG_27__SCAN_IN), .ZN(n2813) );
  NAND2_X1 U35270 ( .A1(n3950), .A2(n2815), .ZN(n2818) );
  INV_X1 U35280 ( .A(n3937), .ZN(n3928) );
  NAND2_X1 U35290 ( .A1(n3928), .A2(n2816), .ZN(n2817) );
  NAND2_X1 U35300 ( .A1(n2818), .A2(n2817), .ZN(n2820) );
  XNOR2_X1 U35310 ( .A(n2820), .B(n2819), .ZN(n2860) );
  NOR2_X1 U35320 ( .A1(n3937), .A2(n3879), .ZN(n2821) );
  AOI21_X1 U35330 ( .B1(n3950), .B2(n2651), .A(n2821), .ZN(n2858) );
  XNOR2_X1 U35340 ( .A(n2860), .B(n2858), .ZN(n3576) );
  NAND2_X1 U35350 ( .A1(n2822), .A2(REG3_REG_28__SCAN_IN), .ZN(n3600) );
  INV_X1 U35360 ( .A(n2822), .ZN(n2824) );
  INV_X1 U35370 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2823) );
  NAND2_X1 U35380 ( .A1(n2824), .A2(n2823), .ZN(n2825) );
  NAND2_X1 U35390 ( .A1(n3600), .A2(n2825), .ZN(n3920) );
  INV_X1 U35400 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4630) );
  NAND2_X1 U35410 ( .A1(n3783), .A2(REG1_REG_28__SCAN_IN), .ZN(n2827) );
  NAND2_X1 U35420 ( .A1(n2672), .A2(REG2_REG_28__SCAN_IN), .ZN(n2826) );
  OAI211_X1 U35430 ( .C1(n2395), .C2(n4630), .A(n2827), .B(n2826), .ZN(n2828)
         );
  INV_X1 U35440 ( .A(n2828), .ZN(n2829) );
  OAI22_X1 U35450 ( .A1(n3930), .A2(n3879), .B1(n2831), .B2(n3585), .ZN(n2833)
         );
  XNOR2_X1 U35460 ( .A(n2833), .B(n2832), .ZN(n2836) );
  OAI22_X1 U35470 ( .A1(n3930), .A2(n2834), .B1(n3879), .B2(n3585), .ZN(n2835)
         );
  XNOR2_X1 U35480 ( .A(n2836), .B(n2835), .ZN(n2865) );
  INV_X1 U35490 ( .A(n2865), .ZN(n2857) );
  INV_X1 U35500 ( .A(n2992), .ZN(n3000) );
  NAND2_X1 U35510 ( .A1(n2998), .A2(n3000), .ZN(n2837) );
  MUX2_X1 U35520 ( .A(n2998), .B(n2837), .S(B_REG_SCAN_IN), .Z(n2838) );
  OAI22_X1 U35530 ( .A1(n2997), .A2(D_REG_1__SCAN_IN), .B1(n4254), .B2(n2992), 
        .ZN(n2971) );
  INV_X1 U35540 ( .A(n2971), .ZN(n3212) );
  INV_X1 U35550 ( .A(D_REG_0__SCAN_IN), .ZN(n2999) );
  NAND2_X1 U35560 ( .A1(n2852), .A2(n2999), .ZN(n2841) );
  INV_X1 U35570 ( .A(n4254), .ZN(n2839) );
  NAND2_X1 U35580 ( .A1(n2839), .A2(n2998), .ZN(n2840) );
  NOR4_X1 U35590 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2850) );
  NOR4_X1 U35600 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2849) );
  INV_X1 U35610 ( .A(D_REG_17__SCAN_IN), .ZN(n4727) );
  INV_X1 U35620 ( .A(D_REG_4__SCAN_IN), .ZN(n4711) );
  INV_X1 U35630 ( .A(D_REG_8__SCAN_IN), .ZN(n4712) );
  INV_X1 U35640 ( .A(D_REG_7__SCAN_IN), .ZN(n4698) );
  NAND4_X1 U35650 ( .A1(n4727), .A2(n4711), .A3(n4712), .A4(n4698), .ZN(n2847)
         );
  NOR4_X1 U35660 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2845) );
  NOR4_X1 U35670 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_31__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2844) );
  NOR4_X1 U35680 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_29__SCAN_IN), .ZN(n2843) );
  NOR4_X1 U35690 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2842) );
  NAND4_X1 U35700 ( .A1(n2845), .A2(n2844), .A3(n2843), .A4(n2842), .ZN(n2846)
         );
  NOR4_X1 U35710 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(n2847), 
        .A4(n2846), .ZN(n2848) );
  NAND3_X1 U35720 ( .A1(n2850), .A2(n2849), .A3(n2848), .ZN(n2851) );
  NAND2_X1 U35730 ( .A1(n2852), .A2(n2851), .ZN(n2969) );
  NAND3_X1 U35740 ( .A1(n3212), .A2(n2979), .A3(n2969), .ZN(n2873) );
  OR2_X1 U35750 ( .A1(n2873), .A2(n3024), .ZN(n2883) );
  INV_X1 U35760 ( .A(n3021), .ZN(n2964) );
  NAND2_X1 U35770 ( .A1(n2884), .A2(n4305), .ZN(n2868) );
  NAND2_X1 U35780 ( .A1(n3132), .A2(n2868), .ZN(n2855) );
  NAND2_X1 U35790 ( .A1(n2964), .A2(n2855), .ZN(n2856) );
  NAND2_X1 U35800 ( .A1(n2857), .A2(n3678), .ZN(n2892) );
  INV_X1 U35810 ( .A(n2858), .ZN(n2859) );
  NAND2_X1 U3582 ( .A1(n2860), .A2(n2859), .ZN(n2864) );
  INV_X1 U3583 ( .A(n2864), .ZN(n2861) );
  AND2_X1 U3584 ( .A1(n2865), .A2(n2862), .ZN(n2863) );
  NOR3_X1 U3585 ( .A1(n2865), .A2(n4551), .A3(n2864), .ZN(n2889) );
  AND2_X1 U3586 ( .A1(n2884), .A2(n2961), .ZN(n4449) );
  NAND2_X1 U3587 ( .A1(n4517), .A2(n2867), .ZN(n2970) );
  NAND2_X1 U3588 ( .A1(n2873), .A2(n2970), .ZN(n3114) );
  AND2_X1 U3589 ( .A1(n3021), .A2(n2868), .ZN(n2968) );
  INV_X1 U3590 ( .A(n3023), .ZN(n2869) );
  NOR2_X1 U3591 ( .A1(n2968), .A2(n2869), .ZN(n2870) );
  AND2_X1 U3592 ( .A1(n2984), .A2(n2870), .ZN(n2871) );
  INV_X2 U3593 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3594 ( .A(n4547), .ZN(n3336) );
  OR2_X1 U3595 ( .A1(n3877), .A2(n3216), .ZN(n2872) );
  NOR2_X1 U3596 ( .A1(n2873), .A2(n2334), .ZN(n2882) );
  NAND2_X1 U3597 ( .A1(n2874), .A2(IR_REG_31__SCAN_IN), .ZN(n2875) );
  INV_X1 U3598 ( .A(n3715), .ZN(n4540) );
  AOI22_X1 U3599 ( .A1(n3950), .A2(n4540), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n2887) );
  INV_X1 U3600 ( .A(REG2_REG_29__SCAN_IN), .ZN(n2880) );
  OR2_X1 U3601 ( .A1(n3600), .A2(n2876), .ZN(n2879) );
  AOI22_X1 U3602 ( .A1(n2877), .A2(REG0_REG_29__SCAN_IN), .B1(n3783), .B2(
        REG1_REG_29__SCAN_IN), .ZN(n2878) );
  OAI211_X1 U3603 ( .C1(n2881), .C2(n2880), .A(n2879), .B(n2878), .ZN(n3790)
         );
  INV_X1 U3604 ( .A(n2883), .ZN(n2885) );
  INV_X1 U3605 ( .A(n2884), .ZN(n4257) );
  AOI21_X2 U3606 ( .B1(n2885), .B2(n4162), .A(n4453), .ZN(n3700) );
  AOI22_X1 U3607 ( .A1(n3790), .A2(n3712), .B1(n4542), .B2(n2975), .ZN(n2886)
         );
  OAI211_X1 U3608 ( .C1(n3336), .C2(n3920), .A(n2887), .B(n2886), .ZN(n2888)
         );
  NOR2_X1 U3609 ( .A1(n2889), .A2(n2888), .ZN(n2890) );
  OAI211_X1 U3610 ( .C1(n2893), .C2(n2892), .A(n2891), .B(n2890), .ZN(U3217)
         );
  INV_X1 U3611 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2973) );
  NAND2_X1 U3612 ( .A1(n3155), .A2(n3146), .ZN(n3725) );
  INV_X1 U3613 ( .A(n3193), .ZN(n2894) );
  NAND2_X1 U3614 ( .A1(n3173), .A2(n2894), .ZN(n3732) );
  NAND2_X1 U3615 ( .A1(n3732), .A2(n3729), .ZN(n2935) );
  NAND2_X1 U3616 ( .A1(n3155), .A2(n3122), .ZN(n3181) );
  NAND2_X1 U3617 ( .A1(n3222), .A2(n2894), .ZN(n2895) );
  NAND2_X1 U3618 ( .A1(n3894), .A2(n3220), .ZN(n2896) );
  INV_X1 U3619 ( .A(n3894), .ZN(n3163) );
  NAND2_X1 U3620 ( .A1(n3163), .A2(n3226), .ZN(n3241) );
  INV_X1 U3621 ( .A(n3893), .ZN(n3296) );
  INV_X1 U3622 ( .A(n3252), .ZN(n3165) );
  NAND2_X1 U3623 ( .A1(n3893), .A2(n3165), .ZN(n3738) );
  NAND2_X1 U3624 ( .A1(n3735), .A2(n3738), .ZN(n3239) );
  AND2_X1 U3625 ( .A1(n3241), .A2(n3239), .ZN(n2897) );
  NAND2_X1 U3626 ( .A1(n3242), .A2(n2897), .ZN(n2899) );
  NAND2_X1 U3627 ( .A1(n3893), .A2(n3252), .ZN(n2898) );
  NAND2_X1 U3628 ( .A1(n2899), .A2(n2898), .ZN(n3293) );
  INV_X1 U3629 ( .A(n3277), .ZN(n3164) );
  NAND2_X1 U3630 ( .A1(n3164), .A2(n2938), .ZN(n2900) );
  NAND2_X1 U3631 ( .A1(n3293), .A2(n2900), .ZN(n2902) );
  NAND2_X1 U3632 ( .A1(n3277), .A2(n3301), .ZN(n2901) );
  NAND2_X1 U3633 ( .A1(n2902), .A2(n2901), .ZN(n3281) );
  AND2_X1 U3634 ( .A1(n3892), .A2(n3276), .ZN(n2903) );
  OAI22_X1 U3635 ( .A1(n3281), .A2(n2903), .B1(n3276), .B2(n3892), .ZN(n3317)
         );
  INV_X1 U3636 ( .A(n3317), .ZN(n2905) );
  INV_X1 U3637 ( .A(n4539), .ZN(n3262) );
  NAND2_X1 U3638 ( .A1(n3262), .A2(n3331), .ZN(n2940) );
  NAND2_X1 U3639 ( .A1(n4539), .A2(n3310), .ZN(n3750) );
  NAND2_X1 U3640 ( .A1(n4539), .A2(n3331), .ZN(n2906) );
  INV_X1 U3641 ( .A(n3891), .ZN(n3353) );
  AND2_X1 U3642 ( .A1(n3103), .A2(n3365), .ZN(n2908) );
  INV_X1 U3643 ( .A(n3365), .ZN(n3360) );
  NAND2_X1 U3644 ( .A1(n4544), .A2(n3360), .ZN(n2907) );
  NOR2_X1 U3645 ( .A1(n3890), .A2(n3390), .ZN(n2909) );
  NAND2_X1 U3646 ( .A1(n3417), .A2(n3425), .ZN(n3437) );
  NAND2_X1 U3647 ( .A1(n3442), .A2(n3431), .ZN(n3440) );
  NAND2_X1 U3648 ( .A1(n3417), .A2(n3431), .ZN(n2910) );
  NAND2_X1 U3649 ( .A1(n3889), .A2(n3449), .ZN(n2911) );
  INV_X1 U3650 ( .A(n3477), .ZN(n3533) );
  NAND2_X1 U3651 ( .A1(n3533), .A2(n3493), .ZN(n2912) );
  INV_X1 U3652 ( .A(n3888), .ZN(n3716) );
  NAND2_X1 U3653 ( .A1(n3716), .A2(n3511), .ZN(n3766) );
  INV_X1 U3654 ( .A(n3511), .ZN(n3534) );
  NAND2_X1 U3655 ( .A1(n3888), .A2(n3534), .ZN(n3746) );
  NAND2_X1 U3656 ( .A1(n3766), .A2(n3746), .ZN(n3501) );
  NAND2_X1 U3657 ( .A1(n3502), .A2(n3501), .ZN(n3500) );
  NAND2_X1 U3658 ( .A1(n3716), .A2(n3534), .ZN(n2913) );
  NAND2_X1 U3659 ( .A1(n3500), .A2(n2913), .ZN(n3465) );
  NAND2_X1 U3660 ( .A1(n3551), .A2(n3713), .ZN(n2914) );
  INV_X1 U3661 ( .A(n3551), .ZN(n3642) );
  NAND2_X1 U3662 ( .A1(n3653), .A2(n3556), .ZN(n3844) );
  NAND2_X1 U3663 ( .A1(n4136), .A2(n3643), .ZN(n3847) );
  NAND2_X1 U3664 ( .A1(n3549), .A2(n2915), .ZN(n3548) );
  NAND2_X1 U3665 ( .A1(n4136), .A2(n3556), .ZN(n2916) );
  NAND2_X1 U3666 ( .A1(n3548), .A2(n2916), .ZN(n4128) );
  NAND2_X1 U3667 ( .A1(n4113), .A2(n4131), .ZN(n2917) );
  NAND2_X1 U3668 ( .A1(n4128), .A2(n2917), .ZN(n2919) );
  NAND2_X1 U3669 ( .A1(n3887), .A2(n4141), .ZN(n2918) );
  INV_X1 U3670 ( .A(n4092), .ZN(n4134) );
  NAND2_X1 U3671 ( .A1(n4134), .A2(n4108), .ZN(n4087) );
  NAND2_X1 U3672 ( .A1(n4092), .A2(n4117), .ZN(n4085) );
  NAND2_X1 U3673 ( .A1(n4134), .A2(n4117), .ZN(n2920) );
  NOR2_X1 U3674 ( .A1(n4110), .A2(n2951), .ZN(n4058) );
  NAND2_X1 U3675 ( .A1(n4044), .A2(n4075), .ZN(n3797) );
  NAND2_X1 U3676 ( .A1(n4110), .A2(n2951), .ZN(n4057) );
  OAI211_X1 U3677 ( .C1(n4081), .C2(n4058), .A(n3797), .B(n4057), .ZN(n2921)
         );
  INV_X1 U3678 ( .A(n4044), .ZN(n4090) );
  INV_X1 U3679 ( .A(n4075), .ZN(n4066) );
  NAND2_X1 U3680 ( .A1(n4090), .A2(n4066), .ZN(n3798) );
  NAND2_X1 U3681 ( .A1(n2921), .A2(n3798), .ZN(n4039) );
  NAND2_X1 U3682 ( .A1(n4027), .A2(n2974), .ZN(n2922) );
  INV_X1 U3683 ( .A(n4027), .ZN(n4067) );
  INV_X1 U3684 ( .A(n2974), .ZN(n4049) );
  NAND2_X1 U3685 ( .A1(n4067), .A2(n4049), .ZN(n2923) );
  XNOR2_X1 U3686 ( .A(n4010), .B(n2956), .ZN(n4023) );
  NAND2_X1 U3687 ( .A1(n4025), .A2(n2925), .ZN(n4002) );
  NAND2_X1 U3688 ( .A1(n3993), .A2(n3803), .ZN(n2926) );
  NAND2_X1 U3689 ( .A1(n4009), .A2(n3989), .ZN(n2927) );
  AOI22_X2 U3690 ( .A1(n3982), .A2(n2927), .B1(n3634), .B2(n3995), .ZN(n3963)
         );
  NAND2_X1 U3691 ( .A1(n3699), .A2(n3975), .ZN(n2928) );
  NAND2_X1 U3692 ( .A1(n3969), .A2(n3949), .ZN(n2929) );
  INV_X1 U3693 ( .A(n3969), .ZN(n3635) );
  INV_X1 U3694 ( .A(n3950), .ZN(n3701) );
  NAND2_X1 U3695 ( .A1(n3701), .A2(n3937), .ZN(n2930) );
  NAND2_X1 U3696 ( .A1(n3886), .A2(n3585), .ZN(n3723) );
  NAND2_X1 U3697 ( .A1(n3930), .A2(n2975), .ZN(n3782) );
  NAND2_X1 U3698 ( .A1(n3723), .A2(n3782), .ZN(n3584) );
  XNOR2_X1 U3699 ( .A(n3586), .B(n3584), .ZN(n3917) );
  XNOR2_X1 U3700 ( .A(n3216), .B(n3880), .ZN(n2931) );
  NAND2_X1 U3701 ( .A1(n2931), .A2(n4305), .ZN(n3508) );
  INV_X1 U3702 ( .A(n2932), .ZN(n3834) );
  INV_X1 U3703 ( .A(n3895), .ZN(n2933) );
  NAND2_X1 U3704 ( .A1(n2933), .A2(n3115), .ZN(n3724) );
  OR2_X1 U3705 ( .A1(n2932), .A2(n3724), .ZN(n3187) );
  NAND2_X1 U3706 ( .A1(n3187), .A2(n3728), .ZN(n2936) );
  NAND2_X1 U3707 ( .A1(n2936), .A2(n3832), .ZN(n3189) );
  NAND2_X1 U3708 ( .A1(n3189), .A2(n3729), .ZN(n3219) );
  NAND2_X1 U3709 ( .A1(n3163), .A2(n3220), .ZN(n3734) );
  NAND2_X1 U3710 ( .A1(n3894), .A2(n3226), .ZN(n3731) );
  INV_X1 U3711 ( .A(n3735), .ZN(n2937) );
  AND2_X1 U3712 ( .A1(n3277), .A2(n2938), .ZN(n3292) );
  NAND2_X1 U3713 ( .A1(n3164), .A2(n3301), .ZN(n3751) );
  OAI21_X1 U3714 ( .B1(n3294), .B2(n3292), .A(n3751), .ZN(n3275) );
  NAND2_X1 U3715 ( .A1(n3892), .A2(n3284), .ZN(n3752) );
  NAND2_X1 U3716 ( .A1(n3275), .A2(n3752), .ZN(n2939) );
  INV_X1 U3717 ( .A(n3892), .ZN(n3307) );
  NAND2_X1 U3718 ( .A1(n3307), .A2(n3276), .ZN(n3740) );
  NAND2_X1 U3719 ( .A1(n2939), .A2(n3740), .ZN(n3305) );
  INV_X1 U3720 ( .A(n2940), .ZN(n2941) );
  NAND2_X1 U3721 ( .A1(n3353), .A2(n4541), .ZN(n3743) );
  NAND2_X1 U3722 ( .A1(n3891), .A2(n3340), .ZN(n3753) );
  AND2_X1 U3723 ( .A1(n3103), .A2(n3360), .ZN(n3748) );
  OR2_X1 U3724 ( .A1(n3359), .A2(n3748), .ZN(n2942) );
  NAND2_X1 U3725 ( .A1(n4544), .A2(n3365), .ZN(n3744) );
  NAND2_X1 U3726 ( .A1(n2942), .A2(n3744), .ZN(n3389) );
  NAND2_X1 U3727 ( .A1(n3890), .A2(n3407), .ZN(n3760) );
  NAND2_X1 U3728 ( .A1(n3389), .A2(n3760), .ZN(n2943) );
  NAND2_X1 U3729 ( .A1(n3427), .A2(n3390), .ZN(n3758) );
  NAND2_X1 U3730 ( .A1(n2943), .A2(n3758), .ZN(n3439) );
  INV_X1 U3731 ( .A(n3449), .ZN(n3445) );
  NAND2_X1 U3732 ( .A1(n3889), .A2(n3445), .ZN(n3479) );
  NAND2_X1 U3733 ( .A1(n3477), .A2(n3493), .ZN(n2944) );
  NAND2_X1 U3734 ( .A1(n3479), .A2(n2944), .ZN(n2946) );
  INV_X1 U3735 ( .A(n3440), .ZN(n2945) );
  NOR2_X1 U3736 ( .A1(n2946), .A2(n2945), .ZN(n3761) );
  NAND2_X1 U3737 ( .A1(n3439), .A2(n3761), .ZN(n2950) );
  INV_X1 U3738 ( .A(n3889), .ZN(n3487) );
  NAND2_X1 U3739 ( .A1(n3487), .A2(n3449), .ZN(n3481) );
  NAND2_X1 U3740 ( .A1(n3437), .A2(n3481), .ZN(n2949) );
  INV_X1 U3741 ( .A(n2946), .ZN(n2948) );
  NOR2_X1 U3742 ( .A1(n3477), .A2(n3493), .ZN(n2947) );
  AOI21_X1 U3743 ( .B1(n2949), .B2(n2948), .A(n2947), .ZN(n3764) );
  NAND2_X1 U3744 ( .A1(n2950), .A2(n3764), .ZN(n3843) );
  INV_X1 U3745 ( .A(n3501), .ZN(n3833) );
  NAND2_X1 U3746 ( .A1(n3843), .A2(n3833), .ZN(n3503) );
  NAND2_X1 U3747 ( .A1(n3642), .A2(n3713), .ZN(n3765) );
  NAND2_X1 U3748 ( .A1(n3551), .A2(n3470), .ZN(n3747) );
  NAND2_X1 U3749 ( .A1(n3765), .A2(n3747), .ZN(n3809) );
  INV_X1 U3750 ( .A(n3847), .ZN(n3768) );
  NAND2_X1 U3751 ( .A1(n3887), .A2(n4131), .ZN(n3846) );
  AND2_X1 U3752 ( .A1(n4130), .A2(n3846), .ZN(n4084) );
  NAND2_X1 U3753 ( .A1(n4110), .A2(n4095), .ZN(n2952) );
  AND2_X1 U3754 ( .A1(n4085), .A2(n2952), .ZN(n3848) );
  NAND2_X1 U3755 ( .A1(n4084), .A2(n3848), .ZN(n4063) );
  NAND2_X1 U3756 ( .A1(n4113), .A2(n4141), .ZN(n4082) );
  NAND2_X1 U3757 ( .A1(n4087), .A2(n4082), .ZN(n2954) );
  NOR2_X1 U3758 ( .A1(n4110), .A2(n4095), .ZN(n2953) );
  AOI21_X1 U3759 ( .B1(n2954), .B2(n3848), .A(n2953), .ZN(n4062) );
  NAND2_X1 U3760 ( .A1(n4090), .A2(n4075), .ZN(n2955) );
  AND2_X1 U3761 ( .A1(n4044), .A2(n4066), .ZN(n3850) );
  NAND2_X1 U3762 ( .A1(n4067), .A2(n2974), .ZN(n4003) );
  NAND2_X1 U3763 ( .A1(n4042), .A2(n2956), .ZN(n4006) );
  NAND2_X1 U3764 ( .A1(n4003), .A2(n4006), .ZN(n3855) );
  AND2_X1 U3765 ( .A1(n4027), .A2(n4049), .ZN(n3796) );
  NAND2_X1 U3766 ( .A1(n4028), .A2(n3803), .ZN(n2958) );
  NAND2_X1 U3767 ( .A1(n4010), .A2(n4034), .ZN(n2957) );
  NAND2_X1 U3768 ( .A1(n2958), .A2(n2957), .ZN(n3775) );
  AOI21_X1 U3769 ( .B1(n3796), .B2(n4006), .A(n3775), .ZN(n3853) );
  NOR2_X1 U3770 ( .A1(n4009), .A2(n3995), .ZN(n3802) );
  NOR2_X1 U3771 ( .A1(n4028), .A2(n3803), .ZN(n3983) );
  NOR2_X1 U3772 ( .A1(n3802), .A2(n3983), .ZN(n3859) );
  NAND2_X1 U3773 ( .A1(n3990), .A2(n3975), .ZN(n3800) );
  NAND2_X1 U3774 ( .A1(n4009), .A2(n3995), .ZN(n3964) );
  AND2_X1 U3775 ( .A1(n3800), .A2(n3964), .ZN(n3856) );
  OR2_X1 U3776 ( .A1(n3969), .A2(n3956), .ZN(n3828) );
  NAND2_X1 U3777 ( .A1(n3699), .A2(n3968), .ZN(n3945) );
  NAND2_X1 U3778 ( .A1(n3828), .A2(n3945), .ZN(n3861) );
  INV_X1 U3779 ( .A(n3861), .ZN(n2959) );
  AND2_X1 U3780 ( .A1(n3969), .A2(n3956), .ZN(n3827) );
  AOI21_X1 U3781 ( .B1(n3946), .B2(n2959), .A(n3827), .ZN(n3927) );
  AND2_X1 U3782 ( .A1(n3950), .A2(n3937), .ZN(n3780) );
  INV_X1 U3783 ( .A(n3780), .ZN(n2960) );
  NAND2_X1 U3784 ( .A1(n3927), .A2(n3933), .ZN(n3926) );
  NAND2_X1 U3785 ( .A1(n3926), .A2(n3781), .ZN(n3590) );
  XNOR2_X1 U3786 ( .A(n3590), .B(n3584), .ZN(n2967) );
  NAND2_X1 U3787 ( .A1(n3880), .A2(n2961), .ZN(n2963) );
  NAND2_X1 U3788 ( .A1(n4257), .A2(n4256), .ZN(n2962) );
  AOI22_X1 U3789 ( .A1(n3790), .A2(n4109), .B1(n4162), .B2(n2975), .ZN(n2966)
         );
  NAND2_X1 U3790 ( .A1(n3950), .A2(n4137), .ZN(n2965) );
  OAI211_X1 U3791 ( .C1(n2967), .C2(n4139), .A(n2966), .B(n2965), .ZN(n3923)
         );
  AOI21_X1 U3792 ( .B1(n3917), .B2(n4496), .A(n3923), .ZN(n2981) );
  NAND2_X1 U3793 ( .A1(n2333), .A2(n2969), .ZN(n3213) );
  NAND2_X1 U3794 ( .A1(n2971), .A2(n2970), .ZN(n2972) );
  NAND2_X1 U3795 ( .A1(n3145), .A2(n3146), .ZN(n3194) );
  NAND2_X1 U3796 ( .A1(n3311), .A2(n3310), .ZN(n3345) );
  NAND2_X1 U3797 ( .A1(n3510), .A2(n3470), .ZN(n3557) );
  INV_X1 U3798 ( .A(n3936), .ZN(n2976) );
  OAI21_X1 U3799 ( .B1(n2976), .B2(n3585), .A(n3588), .ZN(n3918) );
  NAND2_X1 U3800 ( .A1(n2978), .A2(n2977), .ZN(U3546) );
  NAND2_X1 U3801 ( .A1(n2983), .A2(n2982), .ZN(U3514) );
  INV_X1 U3802 ( .A(n2154), .ZN(n3071) );
  INV_X1 U3803 ( .A(DATAI_1_), .ZN(n2985) );
  MUX2_X1 U3804 ( .A(n3071), .B(n2985), .S(U3149), .Z(n2986) );
  INV_X1 U3805 ( .A(n2986), .ZN(U3351) );
  INV_X1 U3806 ( .A(n3028), .ZN(n3906) );
  INV_X1 U3807 ( .A(DATAI_2_), .ZN(n2987) );
  MUX2_X1 U3808 ( .A(n3906), .B(n2987), .S(U3149), .Z(n2988) );
  INV_X1 U3809 ( .A(n2988), .ZN(U3350) );
  INV_X1 U3810 ( .A(DATAI_19_), .ZN(n2989) );
  MUX2_X1 U3811 ( .A(n2989), .B(n4305), .S(STATE_REG_SCAN_IN), .Z(n2990) );
  INV_X1 U3812 ( .A(n2990), .ZN(U3333) );
  INV_X1 U3813 ( .A(DATAI_22_), .ZN(n4639) );
  NAND2_X1 U3814 ( .A1(n3880), .A2(STATE_REG_SCAN_IN), .ZN(n2991) );
  OAI21_X1 U3815 ( .B1(STATE_REG_SCAN_IN), .B2(n4639), .A(n2991), .ZN(U3330)
         );
  INV_X1 U3816 ( .A(DATAI_25_), .ZN(n4729) );
  NAND2_X1 U3817 ( .A1(n2992), .A2(STATE_REG_SCAN_IN), .ZN(n2993) );
  OAI21_X1 U3818 ( .B1(STATE_REG_SCAN_IN), .B2(n4729), .A(n2993), .ZN(U3327)
         );
  INV_X1 U3819 ( .A(DATAI_27_), .ZN(n2995) );
  NAND2_X1 U3820 ( .A1(n4322), .A2(STATE_REG_SCAN_IN), .ZN(n2994) );
  OAI21_X1 U3821 ( .B1(STATE_REG_SCAN_IN), .B2(n2995), .A(n2994), .ZN(U3325)
         );
  INV_X1 U3822 ( .A(n3024), .ZN(n2996) );
  NOR2_X1 U3823 ( .A1(n4254), .A2(n3878), .ZN(n3001) );
  AOI22_X1 U3824 ( .A1(n4459), .A2(n2999), .B1(n3001), .B2(n2998), .ZN(U3458)
         );
  INV_X1 U3825 ( .A(D_REG_1__SCAN_IN), .ZN(n3002) );
  AOI22_X1 U3826 ( .A1(n4459), .A2(n3002), .B1(n3001), .B2(n3000), .ZN(U3459)
         );
  INV_X1 U3827 ( .A(DATAI_31_), .ZN(n4832) );
  OR4_X1 U3828 ( .A1(n2348), .A2(IR_REG_30__SCAN_IN), .A3(U3149), .A4(n2373), 
        .ZN(n3003) );
  OAI21_X1 U3829 ( .B1(STATE_REG_SCAN_IN), .B2(n4832), .A(n3003), .ZN(U3321)
         );
  INV_X1 U3830 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n3005) );
  NAND2_X1 U3831 ( .A1(n3173), .A2(U4043), .ZN(n3004) );
  OAI21_X1 U3832 ( .B1(U4043), .B2(n3005), .A(n3004), .ZN(U3552) );
  INV_X1 U3833 ( .A(REG1_REG_1__SCAN_IN), .ZN(n3006) );
  XNOR2_X1 U3834 ( .A(n3064), .B(n3006), .ZN(n3062) );
  AND2_X1 U3835 ( .A1(REG1_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n3063)
         );
  NAND2_X1 U3836 ( .A1(n3062), .A2(n3063), .ZN(n3008) );
  NAND2_X1 U3837 ( .A1(n2154), .A2(REG1_REG_1__SCAN_IN), .ZN(n3007) );
  NAND2_X1 U3838 ( .A1(n3008), .A2(n3007), .ZN(n3905) );
  NAND2_X1 U3839 ( .A1(n3009), .A2(n3905), .ZN(n3011) );
  NAND2_X1 U3840 ( .A1(n3028), .A2(REG1_REG_2__SCAN_IN), .ZN(n3010) );
  NAND2_X1 U3841 ( .A1(n3011), .A2(n3010), .ZN(n3012) );
  INV_X1 U3842 ( .A(n4262), .ZN(n3049) );
  XNOR2_X1 U3843 ( .A(n3012), .B(n3049), .ZN(n3043) );
  NAND2_X1 U3844 ( .A1(n3043), .A2(REG1_REG_3__SCAN_IN), .ZN(n3014) );
  NAND2_X1 U3845 ( .A1(n3012), .A2(n4262), .ZN(n3013) );
  INV_X1 U3846 ( .A(REG1_REG_4__SCAN_IN), .ZN(n3015) );
  NAND2_X1 U3847 ( .A1(n3016), .A2(n4336), .ZN(n3017) );
  INV_X1 U3848 ( .A(REG1_REG_5__SCAN_IN), .ZN(n3019) );
  MUX2_X1 U3849 ( .A(n3019), .B(REG1_REG_5__SCAN_IN), .S(n3061), .Z(n3018) );
  NOR2_X1 U3850 ( .A1(n3061), .A2(n3019), .ZN(n3020) );
  INV_X1 U3851 ( .A(n4260), .ZN(n3038) );
  XNOR2_X1 U3852 ( .A(n3072), .B(REG1_REG_6__SCAN_IN), .ZN(n3042) );
  NAND2_X1 U3853 ( .A1(n3023), .A2(n3021), .ZN(n3022) );
  OR2_X1 U3854 ( .A1(n3023), .A2(U3149), .ZN(n3883) );
  NAND2_X1 U3855 ( .A1(n3024), .A2(n3883), .ZN(n3033) );
  NAND2_X1 U3856 ( .A1(n3034), .A2(n3033), .ZN(n4325) );
  INV_X1 U3857 ( .A(n3061), .ZN(n4261) );
  NAND2_X1 U3858 ( .A1(n2154), .A2(REG2_REG_1__SCAN_IN), .ZN(n3908) );
  INV_X1 U3859 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3025) );
  MUX2_X1 U3860 ( .A(REG2_REG_1__SCAN_IN), .B(n3025), .S(n2154), .Z(n3026) );
  INV_X1 U3861 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3027) );
  INV_X1 U3862 ( .A(n3029), .ZN(n3030) );
  AOI22_X1 U3863 ( .A1(n3044), .A2(REG2_REG_3__SCAN_IN), .B1(n4262), .B2(n3030), .ZN(n3031) );
  XNOR2_X1 U3864 ( .A(n3031), .B(n4336), .ZN(n4327) );
  INV_X1 U3865 ( .A(n3031), .ZN(n3032) );
  INV_X1 U3866 ( .A(REG2_REG_5__SCAN_IN), .ZN(n4868) );
  MUX2_X1 U3867 ( .A(REG2_REG_5__SCAN_IN), .B(n4868), .S(n3061), .Z(n3051) );
  NOR2_X1 U3868 ( .A1(n3052), .A2(n3051), .ZN(n3050) );
  AOI21_X1 U3869 ( .B1(n4261), .B2(REG2_REG_5__SCAN_IN), .A(n3050), .ZN(n3075)
         );
  XNOR2_X1 U3870 ( .A(n3077), .B(n2215), .ZN(n3040) );
  INV_X1 U3871 ( .A(n4322), .ZN(n3896) );
  OR2_X1 U3872 ( .A1(n4311), .A2(n3896), .ZN(n3904) );
  INV_X1 U3873 ( .A(n3033), .ZN(n3035) );
  NOR2_X1 U3874 ( .A1(STATE_REG_SCAN_IN), .A2(n3036), .ZN(n3264) );
  AOI21_X1 U3875 ( .B1(n4440), .B2(ADDR_REG_6__SCAN_IN), .A(n3264), .ZN(n3037)
         );
  OAI21_X1 U3876 ( .B1(n3038), .B2(n4448), .A(n3037), .ZN(n3039) );
  AOI21_X1 U3877 ( .B1(n3040), .B2(n4433), .A(n3039), .ZN(n3041) );
  OAI21_X1 U3878 ( .B1(n3042), .B2(n4436), .A(n3041), .ZN(U3246) );
  XOR2_X1 U3879 ( .A(n3043), .B(REG1_REG_3__SCAN_IN), .Z(n3046) );
  INV_X1 U3880 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3228) );
  XNOR2_X1 U3881 ( .A(n3044), .B(n3228), .ZN(n3045) );
  AOI22_X1 U3882 ( .A1(n4431), .A2(n3046), .B1(n4433), .B2(n3045), .ZN(n3048)
         );
  AOI22_X1 U3883 ( .A1(n4440), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3047) );
  OAI211_X1 U3884 ( .C1(n3049), .C2(n4448), .A(n3048), .B(n3047), .ZN(U3243)
         );
  AOI211_X1 U3885 ( .C1(n3052), .C2(n3051), .A(n3050), .B(n4441), .ZN(n3058)
         );
  INV_X1 U3886 ( .A(n3053), .ZN(n3056) );
  MUX2_X1 U3887 ( .A(REG1_REG_5__SCAN_IN), .B(n3019), .S(n3061), .Z(n3055) );
  AOI211_X1 U3888 ( .C1(n3056), .C2(n3055), .A(n3054), .B(n4436), .ZN(n3057)
         );
  NOR2_X1 U3889 ( .A1(n3058), .A2(n3057), .ZN(n3060) );
  AND2_X1 U3890 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3206) );
  AOI21_X1 U3891 ( .B1(n4440), .B2(ADDR_REG_5__SCAN_IN), .A(n3206), .ZN(n3059)
         );
  OAI211_X1 U3892 ( .C1(n3061), .C2(n4448), .A(n3060), .B(n3059), .ZN(U3245)
         );
  XOR2_X1 U3893 ( .A(n3063), .B(n3062), .Z(n3068) );
  INV_X1 U3894 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4744) );
  OR2_X1 U3895 ( .A1(n4830), .A2(n4744), .ZN(n3903) );
  MUX2_X1 U3896 ( .A(n3025), .B(REG2_REG_1__SCAN_IN), .S(n2154), .Z(n3066) );
  INV_X1 U3897 ( .A(n3907), .ZN(n3065) );
  AOI211_X1 U3898 ( .C1(n3903), .C2(n3066), .A(n3065), .B(n4441), .ZN(n3067)
         );
  AOI21_X1 U3899 ( .B1(n4431), .B2(n3068), .A(n3067), .ZN(n3070) );
  AOI22_X1 U3900 ( .A1(n4440), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3069) );
  OAI211_X1 U3901 ( .C1(n3071), .C2(n4448), .A(n3070), .B(n3069), .ZN(U3241)
         );
  INV_X1 U3902 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4525) );
  XOR2_X1 U3903 ( .A(n4525), .B(n4259), .Z(n3073) );
  XNOR2_X1 U3904 ( .A(n3087), .B(n3073), .ZN(n3083) );
  INV_X1 U3905 ( .A(n4448), .ZN(n4397) );
  AND2_X1 U3906 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3332) );
  AOI21_X1 U3907 ( .B1(n4440), .B2(ADDR_REG_7__SCAN_IN), .A(n3332), .ZN(n3074)
         );
  INV_X1 U3908 ( .A(n3074), .ZN(n3081) );
  INV_X1 U3909 ( .A(n3075), .ZN(n3076) );
  INV_X1 U3910 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3313) );
  MUX2_X1 U3911 ( .A(n3313), .B(REG2_REG_7__SCAN_IN), .S(n4259), .Z(n3078) );
  AOI211_X1 U3912 ( .C1(n3079), .C2(n3078), .A(n4441), .B(n3084), .ZN(n3080)
         );
  AOI211_X1 U3913 ( .C1(n4397), .C2(n4259), .A(n3081), .B(n3080), .ZN(n3082)
         );
  OAI21_X1 U3914 ( .B1(n4436), .B2(n3083), .A(n3082), .ZN(U3247) );
  XNOR2_X1 U3915 ( .A(n4265), .B(n4280), .ZN(n4267) );
  XOR2_X1 U3916 ( .A(REG2_REG_8__SCAN_IN), .B(n4267), .Z(n3094) );
  NOR2_X1 U3917 ( .A1(STATE_REG_SCAN_IN), .A2(n3085), .ZN(n4546) );
  NOR2_X1 U3918 ( .A1(n4448), .A2(n4280), .ZN(n3086) );
  AOI211_X1 U3919 ( .C1(n4440), .C2(ADDR_REG_8__SCAN_IN), .A(n4546), .B(n3086), 
        .ZN(n3093) );
  OR2_X1 U3920 ( .A1(n4259), .A2(REG1_REG_7__SCAN_IN), .ZN(n3088) );
  NAND2_X1 U3921 ( .A1(n3089), .A2(n3088), .ZN(n4281) );
  XNOR2_X1 U3922 ( .A(n4281), .B(n4280), .ZN(n3090) );
  INV_X1 U3923 ( .A(n3090), .ZN(n3091) );
  INV_X1 U3924 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3374) );
  OAI211_X1 U3925 ( .C1(n3091), .C2(REG1_REG_8__SCAN_IN), .A(n4279), .B(n4431), 
        .ZN(n3092) );
  OAI211_X1 U3926 ( .C1(n3094), .C2(n4441), .A(n3093), .B(n3092), .ZN(U3248)
         );
  NOR2_X1 U3927 ( .A1(n4440), .A2(U4043), .ZN(U3148) );
  INV_X1 U3928 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n3096) );
  NAND2_X1 U3929 ( .A1(n3277), .A2(U4043), .ZN(n3095) );
  OAI21_X1 U3930 ( .B1(U4043), .B2(n3096), .A(n3095), .ZN(U3555) );
  INV_X1 U3931 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n3098) );
  NAND2_X1 U3932 ( .A1(n3442), .A2(U4043), .ZN(n3097) );
  OAI21_X1 U3933 ( .B1(U4043), .B2(n3098), .A(n3097), .ZN(U3561) );
  INV_X1 U3934 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n3100) );
  NAND2_X1 U3935 ( .A1(n3155), .A2(U4043), .ZN(n3099) );
  OAI21_X1 U3936 ( .B1(U4043), .B2(n3100), .A(n3099), .ZN(U3551) );
  INV_X1 U3937 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n3102) );
  NAND2_X1 U3938 ( .A1(n4110), .A2(U4043), .ZN(n3101) );
  OAI21_X1 U3939 ( .B1(U4043), .B2(n3102), .A(n3101), .ZN(U3569) );
  INV_X1 U3940 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n3105) );
  NAND2_X1 U3941 ( .A1(n3103), .A2(U4043), .ZN(n3104) );
  OAI21_X1 U3942 ( .B1(U4043), .B2(n3105), .A(n3104), .ZN(U3559) );
  INV_X1 U3943 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n3107) );
  NAND2_X1 U3944 ( .A1(n4539), .A2(U4043), .ZN(n3106) );
  OAI21_X1 U3945 ( .B1(U4043), .B2(n3107), .A(n3106), .ZN(U3557) );
  INV_X1 U3946 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n3109) );
  NAND2_X1 U3947 ( .A1(n4044), .A2(U4043), .ZN(n3108) );
  OAI21_X1 U3948 ( .B1(U4043), .B2(n3109), .A(n3108), .ZN(U3570) );
  INV_X1 U3949 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n3111) );
  NAND2_X1 U3950 ( .A1(n4010), .A2(U4043), .ZN(n3110) );
  OAI21_X1 U3951 ( .B1(U4043), .B2(n3111), .A(n3110), .ZN(U3572) );
  XNOR2_X1 U3952 ( .A(n3113), .B(n3112), .ZN(n3898) );
  NAND2_X1 U3953 ( .A1(n3114), .A2(n2333), .ZN(n3154) );
  AOI22_X1 U3954 ( .A1(n3712), .A2(n3155), .B1(REG3_REG_0__SCAN_IN), .B2(n3154), .ZN(n3117) );
  NAND2_X1 U3955 ( .A1(n4542), .A2(n3115), .ZN(n3116) );
  OAI211_X1 U3956 ( .C1(n3898), .C2(n4551), .A(n3117), .B(n3116), .ZN(U3229)
         );
  INV_X1 U3957 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n3119) );
  NAND2_X1 U3958 ( .A1(n4009), .A2(U4043), .ZN(n3118) );
  OAI21_X1 U3959 ( .B1(U4043), .B2(n3119), .A(n3118), .ZN(U3574) );
  XNOR2_X1 U3960 ( .A(n3121), .B(n3120), .ZN(n3125) );
  AOI22_X1 U3961 ( .A1(n3712), .A2(n3173), .B1(REG3_REG_1__SCAN_IN), .B2(n3154), .ZN(n3124) );
  AOI22_X1 U3962 ( .A1(n4542), .A2(n3122), .B1(n4540), .B2(n3895), .ZN(n3123)
         );
  OAI211_X1 U3963 ( .C1(n3125), .C2(n4551), .A(n3124), .B(n3123), .ZN(U3219)
         );
  INV_X1 U3964 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n3127) );
  NAND2_X1 U3965 ( .A1(n3551), .A2(U4043), .ZN(n3126) );
  OAI21_X1 U3966 ( .B1(U4043), .B2(n3127), .A(n3126), .ZN(U3565) );
  INV_X1 U3967 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n3129) );
  NAND2_X1 U3968 ( .A1(n3477), .A2(U4043), .ZN(n3128) );
  OAI21_X1 U3969 ( .B1(U4043), .B2(n3129), .A(n3128), .ZN(U3563) );
  INV_X1 U3970 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n3131) );
  NAND2_X1 U3971 ( .A1(n3990), .A2(U4043), .ZN(n3130) );
  OAI21_X1 U3972 ( .B1(U4043), .B2(n3131), .A(n3130), .ZN(U3575) );
  NAND2_X1 U3973 ( .A1(n3895), .A2(n3145), .ZN(n3726) );
  NAND2_X1 U3974 ( .A1(n3724), .A2(n3726), .ZN(n4455) );
  INV_X1 U3975 ( .A(n3132), .ZN(n3133) );
  NOR2_X1 U3976 ( .A1(n3145), .A2(n3133), .ZN(n4452) );
  INV_X1 U3977 ( .A(n3508), .ZN(n4072) );
  OAI21_X1 U3978 ( .B1(n4072), .B2(n4115), .A(n4455), .ZN(n3134) );
  OAI21_X1 U3979 ( .B1(n3186), .B2(n4133), .A(n3134), .ZN(n4450) );
  AOI211_X1 U3980 ( .C1(n4517), .C2(n4455), .A(n4452), .B(n4450), .ZN(n4477)
         );
  NAND2_X1 U3981 ( .A1(n4530), .A2(REG1_REG_0__SCAN_IN), .ZN(n3135) );
  OAI21_X1 U3982 ( .B1(n4477), .B2(n4530), .A(n3135), .ZN(U3518) );
  NAND2_X1 U3983 ( .A1(n2932), .A2(n3724), .ZN(n3136) );
  NAND2_X1 U3984 ( .A1(n3187), .A2(n3136), .ZN(n3140) );
  NAND2_X1 U3985 ( .A1(n3895), .A2(n4137), .ZN(n3138) );
  NAND2_X1 U3986 ( .A1(n3173), .A2(n4109), .ZN(n3137) );
  OAI211_X1 U3987 ( .C1(n4132), .C2(n3146), .A(n3138), .B(n3137), .ZN(n3139)
         );
  AOI21_X1 U3988 ( .B1(n3140), .B2(n4115), .A(n3139), .ZN(n3144) );
  INV_X1 U3989 ( .A(n3141), .ZN(n3142) );
  XNOR2_X1 U3990 ( .A(n2932), .B(n3142), .ZN(n3273) );
  NAND2_X1 U3991 ( .A1(n3273), .A2(n4072), .ZN(n3143) );
  NAND2_X1 U3992 ( .A1(n3144), .A2(n3143), .ZN(n3270) );
  INV_X1 U3993 ( .A(n3273), .ZN(n3147) );
  OAI21_X1 U3994 ( .B1(n3146), .B2(n3145), .A(n3194), .ZN(n3269) );
  OAI22_X1 U3995 ( .A1(n3147), .A2(n4480), .B1(n4512), .B2(n3269), .ZN(n3148)
         );
  NOR2_X1 U3996 ( .A1(n3270), .A2(n3148), .ZN(n4478) );
  NAND2_X1 U3997 ( .A1(n4530), .A2(REG1_REG_1__SCAN_IN), .ZN(n3149) );
  OAI21_X1 U3998 ( .B1(n4478), .B2(n4530), .A(n3149), .ZN(U3519) );
  INV_X1 U3999 ( .A(n3151), .ZN(n3152) );
  AOI21_X1 U4000 ( .B1(n3150), .B2(n3153), .A(n3152), .ZN(n3158) );
  AOI22_X1 U4001 ( .A1(n3712), .A2(n3894), .B1(REG3_REG_2__SCAN_IN), .B2(n3154), .ZN(n3157) );
  AOI22_X1 U4002 ( .A1(n4542), .A2(n3193), .B1(n4540), .B2(n3155), .ZN(n3156)
         );
  OAI211_X1 U4003 ( .C1(n3158), .C2(n4551), .A(n3157), .B(n3156), .ZN(U3234)
         );
  NAND2_X1 U4004 ( .A1(n3159), .A2(n3678), .ZN(n3170) );
  AOI21_X1 U4005 ( .B1(n3160), .B2(n3162), .A(n3161), .ZN(n3169) );
  NAND2_X1 U4006 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4331) );
  OAI21_X1 U4007 ( .B1(n3163), .B2(n3715), .A(n4331), .ZN(n3167) );
  OAI22_X1 U4008 ( .A1(n3700), .A2(n3165), .B1(n3164), .B2(n4543), .ZN(n3166)
         );
  AOI211_X1 U4009 ( .C1(n3253), .C2(n4547), .A(n3167), .B(n3166), .ZN(n3168)
         );
  OAI21_X1 U4010 ( .B1(n3170), .B2(n3169), .A(n3168), .ZN(U3227) );
  OAI21_X1 U4011 ( .B1(n3172), .B2(n3171), .A(n3160), .ZN(n3177) );
  MUX2_X1 U4012 ( .A(n3336), .B(STATE_REG_SCAN_IN), .S(REG3_REG_3__SCAN_IN), 
        .Z(n3175) );
  AOI22_X1 U4013 ( .A1(n4540), .A2(n3173), .B1(n3712), .B2(n3893), .ZN(n3174)
         );
  OAI211_X1 U4014 ( .C1(n3700), .C2(n3226), .A(n3175), .B(n3174), .ZN(n3176)
         );
  AOI21_X1 U4015 ( .B1(n3177), .B2(n3678), .A(n3176), .ZN(n3178) );
  INV_X1 U4016 ( .A(n3178), .ZN(U3215) );
  INV_X1 U4017 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n3180) );
  NAND2_X1 U4018 ( .A1(n3790), .A2(U4043), .ZN(n3179) );
  OAI21_X1 U4019 ( .B1(U4043), .B2(n3180), .A(n3179), .ZN(U3579) );
  AND2_X1 U4020 ( .A1(n3182), .A2(n3181), .ZN(n3184) );
  OAI21_X1 U4021 ( .B1(n3184), .B2(n2935), .A(n3183), .ZN(n3233) );
  AOI22_X1 U4022 ( .A1(n3894), .A2(n4109), .B1(n3193), .B2(n4162), .ZN(n3185)
         );
  OAI21_X1 U4023 ( .B1(n3186), .B2(n4112), .A(n3185), .ZN(n3191) );
  NAND3_X1 U4024 ( .A1(n2935), .A2(n3728), .A3(n3187), .ZN(n3188) );
  AOI21_X1 U4025 ( .B1(n3189), .B2(n3188), .A(n4139), .ZN(n3190) );
  AOI211_X1 U4026 ( .C1(n4072), .C2(n3233), .A(n3191), .B(n3190), .ZN(n3234)
         );
  INV_X1 U4027 ( .A(n3234), .ZN(n3192) );
  AOI21_X1 U4028 ( .B1(n4517), .B2(n3233), .A(n3192), .ZN(n3202) );
  AND2_X1 U4029 ( .A1(n3194), .A2(n3193), .ZN(n3195) );
  NOR2_X1 U4030 ( .A1(n3227), .A2(n3195), .ZN(n3235) );
  INV_X1 U4031 ( .A(n4211), .ZN(n3196) );
  AOI22_X1 U4032 ( .A1(n3235), .A2(n3196), .B1(REG1_REG_2__SCAN_IN), .B2(n4530), .ZN(n3197) );
  OAI21_X1 U4033 ( .B1(n3202), .B2(n4530), .A(n3197), .ZN(U3520) );
  INV_X1 U4034 ( .A(n4249), .ZN(n3200) );
  INV_X1 U4035 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3198) );
  NOR2_X1 U4036 ( .A1(n4520), .A2(n3198), .ZN(n3199) );
  AOI21_X1 U4037 ( .B1(n3235), .B2(n3200), .A(n3199), .ZN(n3201) );
  OAI21_X1 U4038 ( .B1(n3202), .B2(n4518), .A(n3201), .ZN(U3471) );
  XNOR2_X1 U4039 ( .A(n3203), .B(n3204), .ZN(n3209) );
  AOI22_X1 U4040 ( .A1(n4542), .A2(n3301), .B1(n4540), .B2(n3893), .ZN(n3208)
         );
  NOR2_X1 U4041 ( .A1(n3307), .A2(n4543), .ZN(n3205) );
  AOI211_X1 U4042 ( .C1(n3302), .C2(n4547), .A(n3206), .B(n3205), .ZN(n3207)
         );
  OAI211_X1 U40430 ( .C1(n3209), .C2(n4551), .A(n3208), .B(n3207), .ZN(U3224)
         );
  XNOR2_X1 U4044 ( .A(n3210), .B(n3810), .ZN(n4481) );
  NAND2_X1 U4045 ( .A1(n3212), .A2(n3211), .ZN(n3214) );
  OR2_X1 U4046 ( .A1(n3216), .A2(n4305), .ZN(n3282) );
  INV_X1 U4047 ( .A(n3282), .ZN(n3217) );
  NAND2_X1 U4048 ( .A1(n4125), .A2(n3217), .ZN(n4078) );
  OAI21_X1 U4049 ( .B1(n3810), .B2(n3219), .A(n3218), .ZN(n3224) );
  AOI22_X1 U4050 ( .A1(n3893), .A2(n4109), .B1(n4162), .B2(n3220), .ZN(n3221)
         );
  OAI21_X1 U4051 ( .B1(n3222), .B2(n4112), .A(n3221), .ZN(n3223) );
  AOI21_X1 U4052 ( .B1(n3224), .B2(n4115), .A(n3223), .ZN(n3225) );
  OAI21_X1 U4053 ( .B1(n4481), .B2(n3508), .A(n3225), .ZN(n4483) );
  NAND2_X1 U4054 ( .A1(n4483), .A2(n4125), .ZN(n3232) );
  OAI21_X1 U4055 ( .B1(n3227), .B2(n3226), .A(n3251), .ZN(n4479) );
  INV_X1 U4056 ( .A(n4479), .ZN(n3230) );
  OAI22_X1 U4057 ( .A1(n4125), .A2(n3228), .B1(REG3_REG_3__SCAN_IN), .B2(n4096), .ZN(n3229) );
  AOI21_X1 U4058 ( .B1(n3230), .B2(n4316), .A(n3229), .ZN(n3231) );
  OAI211_X1 U4059 ( .C1(n4481), .C2(n4078), .A(n3232), .B(n3231), .ZN(U3287)
         );
  INV_X1 U4060 ( .A(n3233), .ZN(n3238) );
  MUX2_X1 U4061 ( .A(n3027), .B(n3234), .S(n4125), .Z(n3237) );
  AOI22_X1 U4062 ( .A1(n3235), .A2(n4316), .B1(REG3_REG_2__SCAN_IN), .B2(n4453), .ZN(n3236) );
  OAI211_X1 U4063 ( .C1(n3238), .C2(n4078), .A(n3237), .B(n3236), .ZN(U3288)
         );
  XNOR2_X1 U4064 ( .A(n3240), .B(n3815), .ZN(n3249) );
  NAND2_X1 U4065 ( .A1(n3242), .A2(n3241), .ZN(n3243) );
  OR2_X1 U4066 ( .A1(n3243), .A2(n3815), .ZN(n3245) );
  NAND2_X1 U4067 ( .A1(n3243), .A2(n3815), .ZN(n3244) );
  NAND2_X1 U4068 ( .A1(n3245), .A2(n3244), .ZN(n3255) );
  AOI22_X1 U4069 ( .A1(n3894), .A2(n4137), .B1(n3252), .B2(n4162), .ZN(n3247)
         );
  NAND2_X1 U4070 ( .A1(n3277), .A2(n4109), .ZN(n3246) );
  OAI211_X1 U4071 ( .C1(n3255), .C2(n3508), .A(n3247), .B(n3246), .ZN(n3248)
         );
  AOI21_X1 U4072 ( .B1(n3249), .B2(n4115), .A(n3248), .ZN(n4485) );
  INV_X1 U4073 ( .A(n3300), .ZN(n3250) );
  AOI211_X1 U4074 ( .C1(n3252), .C2(n3251), .A(n4512), .B(n3250), .ZN(n4487)
         );
  AOI22_X1 U4075 ( .A1(n4487), .A2(n4305), .B1(n4453), .B2(n3253), .ZN(n3254)
         );
  AND2_X1 U4076 ( .A1(n4485), .A2(n3254), .ZN(n3257) );
  INV_X1 U4077 ( .A(n3255), .ZN(n4488) );
  INV_X1 U4078 ( .A(n4078), .ZN(n4454) );
  AOI22_X1 U4079 ( .A1(n4488), .A2(n4454), .B1(REG2_REG_4__SCAN_IN), .B2(n4315), .ZN(n3256) );
  OAI21_X1 U4080 ( .B1(n3257), .B2(n4315), .A(n3256), .ZN(U3286) );
  NOR2_X1 U4081 ( .A1(n2239), .A2(n3260), .ZN(n3261) );
  XNOR2_X1 U4082 ( .A(n3258), .B(n3261), .ZN(n3267) );
  AOI22_X1 U4083 ( .A1(n4542), .A2(n3276), .B1(n4540), .B2(n3277), .ZN(n3266)
         );
  NOR2_X1 U4084 ( .A1(n3262), .A2(n4543), .ZN(n3263) );
  AOI211_X1 U4085 ( .C1(n3286), .C2(n4547), .A(n3264), .B(n3263), .ZN(n3265)
         );
  OAI211_X1 U4086 ( .C1(n3267), .C2(n4551), .A(n3266), .B(n3265), .ZN(U3236)
         );
  INV_X1 U4087 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3268) );
  OAI22_X1 U4088 ( .A1(n4146), .A2(n3269), .B1(n3268), .B2(n4096), .ZN(n3272)
         );
  MUX2_X1 U4089 ( .A(n3270), .B(REG2_REG_1__SCAN_IN), .S(n4458), .Z(n3271) );
  AOI211_X1 U4090 ( .C1(n4454), .C2(n3273), .A(n3272), .B(n3271), .ZN(n3274)
         );
  INV_X1 U4091 ( .A(n3274), .ZN(U3289) );
  NAND2_X1 U4092 ( .A1(n3740), .A2(n3752), .ZN(n3808) );
  XNOR2_X1 U4093 ( .A(n3275), .B(n3808), .ZN(n3280) );
  AOI22_X1 U4094 ( .A1(n4539), .A2(n4109), .B1(n4162), .B2(n3276), .ZN(n3279)
         );
  NAND2_X1 U4095 ( .A1(n3277), .A2(n4137), .ZN(n3278) );
  OAI211_X1 U4096 ( .C1(n3280), .C2(n4139), .A(n3279), .B(n3278), .ZN(n3320)
         );
  INV_X1 U4097 ( .A(n3320), .ZN(n3291) );
  XOR2_X1 U4098 ( .A(n3281), .B(n3808), .Z(n3321) );
  NAND2_X1 U4099 ( .A1(n3508), .A2(n3282), .ZN(n3283) );
  INV_X1 U4100 ( .A(n4149), .ZN(n3935) );
  NOR2_X1 U4101 ( .A1(n3299), .A2(n3284), .ZN(n3285) );
  OR2_X1 U4102 ( .A1(n3311), .A2(n3285), .ZN(n3325) );
  NOR2_X1 U4103 ( .A1(n3325), .A2(n4146), .ZN(n3289) );
  INV_X1 U4104 ( .A(n3286), .ZN(n3287) );
  OAI22_X1 U4105 ( .A1(n4125), .A2(n2215), .B1(n3287), .B2(n4096), .ZN(n3288)
         );
  AOI211_X1 U4106 ( .C1(n3321), .C2(n3935), .A(n3289), .B(n3288), .ZN(n3290)
         );
  OAI21_X1 U4107 ( .B1(n3291), .B2(n4315), .A(n3290), .ZN(U3284) );
  INV_X1 U4108 ( .A(n3292), .ZN(n3737) );
  NAND2_X1 U4109 ( .A1(n3737), .A2(n3751), .ZN(n3814) );
  XNOR2_X1 U4110 ( .A(n3293), .B(n3814), .ZN(n4490) );
  XNOR2_X1 U4111 ( .A(n3294), .B(n3814), .ZN(n3298) );
  AOI22_X1 U4112 ( .A1(n3892), .A2(n4109), .B1(n4162), .B2(n3301), .ZN(n3295)
         );
  OAI21_X1 U4113 ( .B1(n3296), .B2(n4112), .A(n3295), .ZN(n3297) );
  AOI21_X1 U4114 ( .B1(n3298), .B2(n4115), .A(n3297), .ZN(n4491) );
  MUX2_X1 U4115 ( .A(n4491), .B(n4868), .S(n4458), .Z(n3304) );
  AOI21_X1 U4116 ( .B1(n3301), .B2(n3300), .A(n3299), .ZN(n4494) );
  AOI22_X1 U4117 ( .A1(n4494), .A2(n4316), .B1(n3302), .B2(n4453), .ZN(n3303)
         );
  OAI211_X1 U4118 ( .C1(n4149), .C2(n4490), .A(n3304), .B(n3303), .ZN(U3285)
         );
  XNOR2_X1 U4119 ( .A(n3305), .B(n3807), .ZN(n3309) );
  AOI22_X1 U4120 ( .A1(n3891), .A2(n4109), .B1(n4162), .B2(n3331), .ZN(n3306)
         );
  OAI21_X1 U4121 ( .B1(n3307), .B2(n4112), .A(n3306), .ZN(n3308) );
  AOI21_X1 U4122 ( .B1(n3309), .B2(n4115), .A(n3308), .ZN(n4500) );
  OAI211_X1 U4123 ( .C1(n3311), .C2(n3310), .A(n4506), .B(n3345), .ZN(n4499)
         );
  INV_X1 U4124 ( .A(n4499), .ZN(n3315) );
  INV_X1 U4125 ( .A(n3312), .ZN(n3335) );
  OAI22_X1 U4126 ( .A1(n4125), .A2(n3313), .B1(n3335), .B2(n4096), .ZN(n3314)
         );
  AOI21_X1 U4127 ( .B1(n3315), .B2(n4120), .A(n3314), .ZN(n3319) );
  NAND2_X1 U4128 ( .A1(n3317), .A2(n3807), .ZN(n4497) );
  NAND3_X1 U4129 ( .A1(n3316), .A2(n4497), .A3(n3935), .ZN(n3318) );
  OAI211_X1 U4130 ( .C1(n4500), .C2(n4315), .A(n3319), .B(n3318), .ZN(U3283)
         );
  AOI21_X1 U4131 ( .B1(n3321), .B2(n4496), .A(n3320), .ZN(n3328) );
  INV_X1 U4132 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3322) );
  OAI22_X1 U4133 ( .A1(n3325), .A2(n4249), .B1(n4520), .B2(n3322), .ZN(n3323)
         );
  INV_X1 U4134 ( .A(n3323), .ZN(n3324) );
  OAI21_X1 U4135 ( .B1(n3328), .B2(n4518), .A(n3324), .ZN(U3479) );
  OAI22_X1 U4136 ( .A1(n3325), .A2(n4211), .B1(n4533), .B2(n2270), .ZN(n3326)
         );
  INV_X1 U4137 ( .A(n3326), .ZN(n3327) );
  OAI21_X1 U4138 ( .B1(n3328), .B2(n4530), .A(n3327), .ZN(U3524) );
  AOI211_X1 U4139 ( .C1(n3330), .C2(n3329), .A(n4551), .B(n2185), .ZN(n3338)
         );
  AOI22_X1 U4140 ( .A1(n4542), .A2(n3331), .B1(n3712), .B2(n3891), .ZN(n3334)
         );
  AOI21_X1 U4141 ( .B1(n4540), .B2(n3892), .A(n3332), .ZN(n3333) );
  OAI211_X1 U4142 ( .C1(n3336), .C2(n3335), .A(n3334), .B(n3333), .ZN(n3337)
         );
  OR2_X1 U4143 ( .A1(n3338), .A2(n3337), .ZN(U3210) );
  NAND2_X1 U4144 ( .A1(n3743), .A2(n3753), .ZN(n3811) );
  XOR2_X1 U4145 ( .A(n3811), .B(n3339), .Z(n3343) );
  OAI22_X1 U4146 ( .A1(n4544), .A2(n4133), .B1(n3340), .B2(n4132), .ZN(n3341)
         );
  AOI21_X1 U4147 ( .B1(n4137), .B2(n4539), .A(n3341), .ZN(n3342) );
  OAI21_X1 U4148 ( .B1(n3343), .B2(n4139), .A(n3342), .ZN(n3372) );
  INV_X1 U4149 ( .A(n3372), .ZN(n3350) );
  XOR2_X1 U4150 ( .A(n3344), .B(n3811), .Z(n3373) );
  NAND2_X1 U4151 ( .A1(n3345), .A2(n4541), .ZN(n3346) );
  AOI22_X1 U4152 ( .A1(n4315), .A2(REG2_REG_8__SCAN_IN), .B1(n4548), .B2(n4453), .ZN(n3347) );
  OAI21_X1 U4153 ( .B1(n3378), .B2(n4146), .A(n3347), .ZN(n3348) );
  AOI21_X1 U4154 ( .B1(n3373), .B2(n3935), .A(n3348), .ZN(n3349) );
  OAI21_X1 U4155 ( .B1(n3350), .B2(n4315), .A(n3349), .ZN(U3282) );
  XOR2_X1 U4156 ( .A(n3351), .B(n3352), .Z(n3357) );
  AOI22_X1 U4157 ( .A1(n4542), .A2(n3365), .B1(n3712), .B2(n3890), .ZN(n3356)
         );
  AND2_X1 U4158 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4343) );
  NOR2_X1 U4159 ( .A1(n3353), .A2(n3715), .ZN(n3354) );
  AOI211_X1 U4160 ( .C1(n3366), .C2(n4547), .A(n4343), .B(n3354), .ZN(n3355)
         );
  OAI211_X1 U4161 ( .C1(n3357), .C2(n4551), .A(n3356), .B(n3355), .ZN(U3228)
         );
  INV_X1 U4162 ( .A(n3748), .ZN(n3754) );
  NAND2_X1 U4163 ( .A1(n3754), .A2(n3744), .ZN(n3812) );
  XNOR2_X1 U4164 ( .A(n3358), .B(n3812), .ZN(n4502) );
  XOR2_X1 U4165 ( .A(n3812), .B(n3359), .Z(n3363) );
  OAI22_X1 U4166 ( .A1(n3427), .A2(n4133), .B1(n4132), .B2(n3360), .ZN(n3361)
         );
  AOI21_X1 U4167 ( .B1(n4137), .B2(n3891), .A(n3361), .ZN(n3362) );
  OAI21_X1 U4168 ( .B1(n3363), .B2(n4139), .A(n3362), .ZN(n4503) );
  NAND2_X1 U4169 ( .A1(n4503), .A2(n4125), .ZN(n3371) );
  AOI21_X1 U4170 ( .B1(n3365), .B2(n3364), .A(n3396), .ZN(n4505) );
  INV_X1 U4171 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3368) );
  INV_X1 U4172 ( .A(n3366), .ZN(n3367) );
  OAI22_X1 U4173 ( .A1(n4125), .A2(n3368), .B1(n3367), .B2(n4096), .ZN(n3369)
         );
  AOI21_X1 U4174 ( .B1(n4505), .B2(n4316), .A(n3369), .ZN(n3370) );
  OAI211_X1 U4175 ( .C1(n4502), .C2(n4149), .A(n3371), .B(n3370), .ZN(U3281)
         );
  AOI21_X1 U4176 ( .B1(n3373), .B2(n4496), .A(n3372), .ZN(n3376) );
  MUX2_X1 U4177 ( .A(n3374), .B(n3376), .S(n4533), .Z(n3375) );
  OAI21_X1 U4178 ( .B1(n3378), .B2(n4211), .A(n3375), .ZN(U3526) );
  INV_X1 U4179 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4714) );
  MUX2_X1 U4180 ( .A(n4714), .B(n3376), .S(n4520), .Z(n3377) );
  OAI21_X1 U4181 ( .B1(n3378), .B2(n4249), .A(n3377), .ZN(U3483) );
  XOR2_X1 U4182 ( .A(n3380), .B(n3379), .Z(n3381) );
  XNOR2_X1 U4183 ( .A(n3382), .B(n3381), .ZN(n3387) );
  AOI22_X1 U4184 ( .A1(n4542), .A2(n3425), .B1(n3712), .B2(n3889), .ZN(n3386)
         );
  INV_X1 U4185 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3383) );
  NOR2_X1 U4186 ( .A1(STATE_REG_SCAN_IN), .A2(n3383), .ZN(n4361) );
  NOR2_X1 U4187 ( .A1(n3427), .A2(n3715), .ZN(n3384) );
  AOI211_X1 U4188 ( .C1(n3432), .C2(n4547), .A(n4361), .B(n3384), .ZN(n3385)
         );
  OAI211_X1 U4189 ( .C1(n3387), .C2(n4551), .A(n3386), .B(n3385), .ZN(U3233)
         );
  NAND2_X1 U4190 ( .A1(n3758), .A2(n3760), .ZN(n3818) );
  XOR2_X1 U4191 ( .A(n3388), .B(n3818), .Z(n3395) );
  XOR2_X1 U4192 ( .A(n3818), .B(n3389), .Z(n3393) );
  AOI22_X1 U4193 ( .A1(n3442), .A2(n4109), .B1(n4162), .B2(n3390), .ZN(n3391)
         );
  OAI21_X1 U4194 ( .B1(n4544), .B2(n4112), .A(n3391), .ZN(n3392) );
  AOI21_X1 U4195 ( .B1(n3393), .B2(n4115), .A(n3392), .ZN(n3394) );
  OAI21_X1 U4196 ( .B1(n3395), .B2(n3508), .A(n3394), .ZN(n4509) );
  INV_X1 U4197 ( .A(n4509), .ZN(n3402) );
  INV_X1 U4198 ( .A(n3395), .ZN(n4511) );
  NOR2_X1 U4199 ( .A1(n3396), .A2(n3407), .ZN(n4508) );
  NOR3_X1 U4200 ( .A1(n4508), .A2(n4507), .A3(n4146), .ZN(n3400) );
  INV_X1 U4201 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3398) );
  OAI22_X1 U4202 ( .A1(n4125), .A2(n3398), .B1(n3397), .B2(n4096), .ZN(n3399)
         );
  AOI211_X1 U4203 ( .C1(n4511), .C2(n4454), .A(n3400), .B(n3399), .ZN(n3401)
         );
  OAI21_X1 U4204 ( .B1(n3402), .B2(n4315), .A(n3401), .ZN(U3280) );
  INV_X1 U4205 ( .A(n3403), .ZN(n3404) );
  AOI211_X1 U4206 ( .C1(n3406), .C2(n3405), .A(n4551), .B(n3404), .ZN(n3412)
         );
  OAI22_X1 U4207 ( .A1(n3700), .A2(n3407), .B1(n4544), .B2(n3715), .ZN(n3411)
         );
  NAND2_X1 U4208 ( .A1(n4547), .A2(n3408), .ZN(n3409) );
  NAND2_X1 U4209 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4351) );
  OAI211_X1 U4210 ( .C1(n3417), .C2(n4543), .A(n3409), .B(n4351), .ZN(n3410)
         );
  OR3_X1 U4211 ( .A1(n3412), .A2(n3411), .A3(n3410), .ZN(U3214) );
  NOR2_X1 U4212 ( .A1(n2252), .A2(n3415), .ZN(n3416) );
  XNOR2_X1 U4213 ( .A(n3413), .B(n3416), .ZN(n3421) );
  NAND2_X1 U4214 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4370) );
  OAI21_X1 U4215 ( .B1(n3533), .B2(n4543), .A(n4370), .ZN(n3419) );
  OAI22_X1 U4216 ( .A1(n3700), .A2(n3445), .B1(n3417), .B2(n3715), .ZN(n3418)
         );
  AOI211_X1 U4217 ( .C1(n3452), .C2(n4547), .A(n3419), .B(n3418), .ZN(n3420)
         );
  OAI21_X1 U4218 ( .B1(n3421), .B2(n4551), .A(n3420), .ZN(U3221) );
  XOR2_X1 U4219 ( .A(n3816), .B(n3439), .Z(n3430) );
  NAND2_X1 U4220 ( .A1(n3422), .A2(n3816), .ZN(n3423) );
  NAND2_X1 U4221 ( .A1(n3424), .A2(n3423), .ZN(n4516) );
  AOI22_X1 U4222 ( .A1(n3889), .A2(n4109), .B1(n4162), .B2(n3425), .ZN(n3426)
         );
  OAI21_X1 U4223 ( .B1(n3427), .B2(n4112), .A(n3426), .ZN(n3428) );
  AOI21_X1 U4224 ( .B1(n4516), .B2(n4072), .A(n3428), .ZN(n3429) );
  OAI21_X1 U4225 ( .B1(n4139), .B2(n3430), .A(n3429), .ZN(n4514) );
  INV_X1 U4226 ( .A(n4514), .ZN(n3436) );
  OAI21_X1 U4227 ( .B1(n4507), .B2(n3431), .A(n3450), .ZN(n4513) );
  AOI22_X1 U4228 ( .A1(n4458), .A2(REG2_REG_11__SCAN_IN), .B1(n3432), .B2(
        n4453), .ZN(n3433) );
  OAI21_X1 U4229 ( .B1(n4513), .B2(n4146), .A(n3433), .ZN(n3434) );
  AOI21_X1 U4230 ( .B1(n4516), .B2(n4454), .A(n3434), .ZN(n3435) );
  OAI21_X1 U4231 ( .B1(n3436), .B2(n4315), .A(n3435), .ZN(U3279) );
  INV_X1 U4232 ( .A(n3437), .ZN(n3438) );
  OR2_X1 U4233 ( .A1(n3439), .A2(n3438), .ZN(n3441) );
  NAND2_X1 U4234 ( .A1(n3441), .A2(n3440), .ZN(n3482) );
  NAND2_X1 U4235 ( .A1(n3481), .A2(n3479), .ZN(n3819) );
  XNOR2_X1 U4236 ( .A(n3482), .B(n3819), .ZN(n3447) );
  NAND2_X1 U4237 ( .A1(n3442), .A2(n4137), .ZN(n3444) );
  NAND2_X1 U4238 ( .A1(n3477), .A2(n4109), .ZN(n3443) );
  OAI211_X1 U4239 ( .C1(n4132), .C2(n3445), .A(n3444), .B(n3443), .ZN(n3446)
         );
  AOI21_X1 U4240 ( .B1(n3447), .B2(n4115), .A(n3446), .ZN(n3521) );
  XNOR2_X1 U4241 ( .A(n3448), .B(n3819), .ZN(n3519) );
  NAND2_X1 U4242 ( .A1(n3450), .A2(n3449), .ZN(n3451) );
  NAND2_X1 U4243 ( .A1(n3492), .A2(n3451), .ZN(n3527) );
  AOI22_X1 U4244 ( .A1(n4315), .A2(REG2_REG_12__SCAN_IN), .B1(n3452), .B2(
        n4453), .ZN(n3453) );
  OAI21_X1 U4245 ( .B1(n3527), .B2(n4146), .A(n3453), .ZN(n3454) );
  AOI21_X1 U4246 ( .B1(n3519), .B2(n3935), .A(n3454), .ZN(n3455) );
  OAI21_X1 U4247 ( .B1(n3521), .B2(n4315), .A(n3455), .ZN(U3278) );
  XOR2_X1 U4248 ( .A(n3457), .B(n3456), .Z(n3458) );
  XNOR2_X1 U4249 ( .A(n3459), .B(n3458), .ZN(n3464) );
  AOI22_X1 U4250 ( .A1(n4542), .A2(n3485), .B1(n3712), .B2(n3888), .ZN(n3463)
         );
  NOR2_X1 U4251 ( .A1(STATE_REG_SCAN_IN), .A2(n3460), .ZN(n4380) );
  NOR2_X1 U4252 ( .A1(n3487), .A2(n3715), .ZN(n3461) );
  AOI211_X1 U4253 ( .C1(n3495), .C2(n4547), .A(n4380), .B(n3461), .ZN(n3462)
         );
  OAI211_X1 U4254 ( .C1(n3464), .C2(n4551), .A(n3463), .B(n3462), .ZN(U3231)
         );
  XNOR2_X1 U4255 ( .A(n3465), .B(n3809), .ZN(n3541) );
  INV_X1 U4256 ( .A(n3541), .ZN(n3476) );
  XNOR2_X1 U4257 ( .A(n3466), .B(n3809), .ZN(n3469) );
  OAI22_X1 U4258 ( .A1(n3653), .A2(n4133), .B1(n3470), .B2(n4132), .ZN(n3467)
         );
  AOI21_X1 U4259 ( .B1(n4137), .B2(n3888), .A(n3467), .ZN(n3468) );
  OAI21_X1 U4260 ( .B1(n3469), .B2(n4139), .A(n3468), .ZN(n3540) );
  OAI21_X1 U4261 ( .B1(n3510), .B2(n3470), .A(n3557), .ZN(n3546) );
  NOR2_X1 U4262 ( .A1(n3546), .A2(n4146), .ZN(n3474) );
  INV_X1 U4263 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3472) );
  INV_X1 U4264 ( .A(n3718), .ZN(n3471) );
  OAI22_X1 U4265 ( .A1(n4125), .A2(n3472), .B1(n3471), .B2(n4096), .ZN(n3473)
         );
  AOI211_X1 U4266 ( .C1(n3540), .C2(n4125), .A(n3474), .B(n3473), .ZN(n3475)
         );
  OAI21_X1 U4267 ( .B1(n3476), .B2(n4149), .A(n3475), .ZN(U3275) );
  XNOR2_X1 U4268 ( .A(n3477), .B(n3493), .ZN(n3483) );
  XNOR2_X1 U4269 ( .A(n3478), .B(n3483), .ZN(n3491) );
  INV_X1 U4270 ( .A(n3479), .ZN(n3480) );
  AOI21_X1 U4271 ( .B1(n3482), .B2(n3481), .A(n3480), .ZN(n3484) );
  INV_X1 U4272 ( .A(n3483), .ZN(n3823) );
  XNOR2_X1 U4273 ( .A(n3484), .B(n3823), .ZN(n3489) );
  AOI22_X1 U4274 ( .A1(n3888), .A2(n4109), .B1(n4162), .B2(n3485), .ZN(n3486)
         );
  OAI21_X1 U4275 ( .B1(n3487), .B2(n4112), .A(n3486), .ZN(n3488) );
  AOI21_X1 U4276 ( .B1(n3489), .B2(n4115), .A(n3488), .ZN(n3490) );
  OAI21_X1 U4277 ( .B1(n3491), .B2(n3508), .A(n3490), .ZN(n3564) );
  INV_X1 U4278 ( .A(n3564), .ZN(n3499) );
  INV_X1 U4279 ( .A(n3491), .ZN(n3565) );
  INV_X1 U4280 ( .A(n3492), .ZN(n3494) );
  OAI21_X1 U4281 ( .B1(n3494), .B2(n3493), .A(n3512), .ZN(n3569) );
  AOI22_X1 U4282 ( .A1(n4315), .A2(REG2_REG_13__SCAN_IN), .B1(n3495), .B2(
        n4453), .ZN(n3496) );
  OAI21_X1 U4283 ( .B1(n3569), .B2(n4146), .A(n3496), .ZN(n3497) );
  AOI21_X1 U4284 ( .B1(n3565), .B2(n4454), .A(n3497), .ZN(n3498) );
  OAI21_X1 U4285 ( .B1(n3499), .B2(n4458), .A(n3498), .ZN(U3277) );
  OAI21_X1 U4286 ( .B1(n3502), .B2(n3501), .A(n3500), .ZN(n3571) );
  INV_X1 U4287 ( .A(n3571), .ZN(n3509) );
  OAI21_X1 U4288 ( .B1(n3833), .B2(n3843), .A(n3503), .ZN(n3506) );
  AOI22_X1 U4289 ( .A1(n3551), .A2(n4109), .B1(n4162), .B2(n3511), .ZN(n3504)
         );
  OAI21_X1 U4290 ( .B1(n3533), .B2(n4112), .A(n3504), .ZN(n3505) );
  AOI21_X1 U4291 ( .B1(n3506), .B2(n4115), .A(n3505), .ZN(n3507) );
  OAI21_X1 U4292 ( .B1(n3509), .B2(n3508), .A(n3507), .ZN(n3570) );
  INV_X1 U4293 ( .A(n3570), .ZN(n3518) );
  INV_X1 U4294 ( .A(n3510), .ZN(n3514) );
  NAND2_X1 U4295 ( .A1(n3512), .A2(n3511), .ZN(n3513) );
  NAND2_X1 U4296 ( .A1(n3514), .A2(n3513), .ZN(n3575) );
  AOI22_X1 U4297 ( .A1(n4315), .A2(REG2_REG_14__SCAN_IN), .B1(n3537), .B2(
        n4453), .ZN(n3515) );
  OAI21_X1 U4298 ( .B1(n3575), .B2(n4146), .A(n3515), .ZN(n3516) );
  AOI21_X1 U4299 ( .B1(n3571), .B2(n4454), .A(n3516), .ZN(n3517) );
  OAI21_X1 U4300 ( .B1(n3518), .B2(n4315), .A(n3517), .ZN(U3276) );
  NAND2_X1 U4301 ( .A1(n3519), .A2(n4496), .ZN(n3520) );
  NAND2_X1 U4302 ( .A1(n3521), .A2(n3520), .ZN(n3524) );
  MUX2_X1 U4303 ( .A(n3524), .B(REG0_REG_12__SCAN_IN), .S(n4518), .Z(n3522) );
  INV_X1 U4304 ( .A(n3522), .ZN(n3523) );
  OAI21_X1 U4305 ( .B1(n3527), .B2(n4249), .A(n3523), .ZN(U3491) );
  MUX2_X1 U4306 ( .A(n3524), .B(REG1_REG_12__SCAN_IN), .S(n4530), .Z(n3525) );
  INV_X1 U4307 ( .A(n3525), .ZN(n3526) );
  OAI21_X1 U4308 ( .B1(n4211), .B2(n3527), .A(n3526), .ZN(U3530) );
  INV_X1 U4309 ( .A(n3529), .ZN(n3531) );
  NAND2_X1 U4310 ( .A1(n3531), .A2(n3530), .ZN(n3532) );
  XNOR2_X1 U4311 ( .A(n3528), .B(n3532), .ZN(n3539) );
  NAND2_X1 U4312 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4398) );
  OAI21_X1 U4313 ( .B1(n3642), .B2(n4543), .A(n4398), .ZN(n3536) );
  OAI22_X1 U4314 ( .A1(n3700), .A2(n3534), .B1(n3533), .B2(n3715), .ZN(n3535)
         );
  AOI211_X1 U4315 ( .C1(n3537), .C2(n4547), .A(n3536), .B(n3535), .ZN(n3538)
         );
  OAI21_X1 U4316 ( .B1(n3539), .B2(n4551), .A(n3538), .ZN(U3212) );
  INV_X1 U4317 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3542) );
  AOI21_X1 U4318 ( .B1(n3541), .B2(n4496), .A(n3540), .ZN(n3544) );
  MUX2_X1 U4319 ( .A(n3542), .B(n3544), .S(n4520), .Z(n3543) );
  OAI21_X1 U4320 ( .B1(n3546), .B2(n4249), .A(n3543), .ZN(U3497) );
  INV_X1 U4321 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4295) );
  MUX2_X1 U4322 ( .A(n4295), .B(n3544), .S(n4533), .Z(n3545) );
  OAI21_X1 U4323 ( .B1(n4211), .B2(n3546), .A(n3545), .ZN(U3533) );
  OAI21_X1 U4324 ( .B1(n3549), .B2(n2915), .A(n3548), .ZN(n4216) );
  XNOR2_X1 U4325 ( .A(n3550), .B(n2915), .ZN(n3555) );
  NAND2_X1 U4326 ( .A1(n3551), .A2(n4137), .ZN(n3553) );
  NAND2_X1 U4327 ( .A1(n3887), .A2(n4109), .ZN(n3552) );
  OAI211_X1 U4328 ( .C1(n4132), .C2(n3643), .A(n3553), .B(n3552), .ZN(n3554)
         );
  AOI21_X1 U4329 ( .B1(n3555), .B2(n4115), .A(n3554), .ZN(n4215) );
  INV_X1 U4330 ( .A(n4215), .ZN(n3562) );
  NAND2_X1 U4331 ( .A1(n3557), .A2(n3556), .ZN(n4212) );
  NAND3_X1 U4332 ( .A1(n4213), .A2(n4316), .A3(n4212), .ZN(n3560) );
  NAND2_X1 U4333 ( .A1(n4453), .A2(n3646), .ZN(n3559) );
  NAND2_X1 U4334 ( .A1(n4458), .A2(REG2_REG_16__SCAN_IN), .ZN(n3558) );
  NAND3_X1 U4335 ( .A1(n3560), .A2(n3559), .A3(n3558), .ZN(n3561) );
  AOI21_X1 U4336 ( .B1(n3562), .B2(n4125), .A(n3561), .ZN(n3563) );
  OAI21_X1 U4337 ( .B1(n4216), .B2(n4149), .A(n3563), .ZN(U3274) );
  INV_X1 U4338 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4291) );
  AOI21_X1 U4339 ( .B1(n4517), .B2(n3565), .A(n3564), .ZN(n3567) );
  MUX2_X1 U4340 ( .A(n4291), .B(n3567), .S(n4533), .Z(n3566) );
  OAI21_X1 U4341 ( .B1(n4211), .B2(n3569), .A(n3566), .ZN(U3531) );
  INV_X1 U4342 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4785) );
  MUX2_X1 U4343 ( .A(n4785), .B(n3567), .S(n4520), .Z(n3568) );
  OAI21_X1 U4344 ( .B1(n3569), .B2(n4249), .A(n3568), .ZN(U3493) );
  INV_X1 U4345 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4794) );
  AOI21_X1 U4346 ( .B1(n4517), .B2(n3571), .A(n3570), .ZN(n3573) );
  MUX2_X1 U4347 ( .A(n4794), .B(n3573), .S(n4520), .Z(n3572) );
  OAI21_X1 U4348 ( .B1(n3575), .B2(n4249), .A(n3572), .ZN(U3495) );
  INV_X1 U4349 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4393) );
  MUX2_X1 U4350 ( .A(n4393), .B(n3573), .S(n4533), .Z(n3574) );
  OAI21_X1 U4351 ( .B1(n4211), .B2(n3575), .A(n3574), .ZN(U3532) );
  XNOR2_X1 U4352 ( .A(n3577), .B(n3576), .ZN(n3578) );
  NAND2_X1 U4353 ( .A1(n3578), .A2(n3678), .ZN(n3583) );
  INV_X1 U4354 ( .A(n3939), .ZN(n3581) );
  OAI22_X1 U4355 ( .A1(n3635), .A2(n3715), .B1(STATE_REG_SCAN_IN), .B2(n4847), 
        .ZN(n3580) );
  OAI22_X1 U4356 ( .A1(n3930), .A2(n4543), .B1(n3700), .B2(n3937), .ZN(n3579)
         );
  AOI211_X1 U4357 ( .C1(n3581), .C2(n4547), .A(n3580), .B(n3579), .ZN(n3582)
         );
  NAND2_X1 U4358 ( .A1(n3583), .A2(n3582), .ZN(U3211) );
  INV_X1 U4359 ( .A(n3584), .ZN(n3830) );
  NAND2_X1 U4360 ( .A1(n3787), .A2(DATAI_29_), .ZN(n3789) );
  XNOR2_X1 U4361 ( .A(n3790), .B(n3789), .ZN(n3836) );
  AOI21_X1 U4362 ( .B1(n3596), .B2(n3588), .A(n4157), .ZN(n4166) );
  AOI22_X1 U4363 ( .A1(n4166), .A2(n4316), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4315), .ZN(n3603) );
  INV_X1 U4364 ( .A(n3782), .ZN(n3589) );
  AOI21_X1 U4365 ( .B1(n3590), .B2(n3723), .A(n3589), .ZN(n3592) );
  INV_X1 U4366 ( .A(n3836), .ZN(n3591) );
  XNOR2_X1 U4367 ( .A(n3592), .B(n3591), .ZN(n3599) );
  INV_X1 U4368 ( .A(REG0_REG_30__SCAN_IN), .ZN(n3595) );
  NAND2_X1 U4369 ( .A1(n3783), .A2(REG1_REG_30__SCAN_IN), .ZN(n3594) );
  NAND2_X1 U4370 ( .A1(n2693), .A2(REG2_REG_30__SCAN_IN), .ZN(n3593) );
  OAI211_X1 U4371 ( .C1(n2395), .C2(n3595), .A(n3594), .B(n3593), .ZN(n3885)
         );
  AOI21_X1 U4372 ( .B1(n4322), .B2(B_REG_SCAN_IN), .A(n4133), .ZN(n4153) );
  AOI22_X1 U4373 ( .A1(n3885), .A2(n4153), .B1(n4162), .B2(n3596), .ZN(n3598)
         );
  NAND2_X1 U4374 ( .A1(n3886), .A2(n4137), .ZN(n3597) );
  NOR2_X1 U4375 ( .A1(n3600), .A2(n4096), .ZN(n3601) );
  OAI21_X1 U4376 ( .B1(n4165), .B2(n3601), .A(n4125), .ZN(n3602) );
  OAI211_X1 U4377 ( .C1(n4167), .C2(n4149), .A(n3603), .B(n3602), .ZN(U3354)
         );
  NAND2_X1 U4378 ( .A1(n3604), .A2(n3678), .ZN(n3612) );
  AOI21_X1 U4379 ( .B1(n3605), .B2(n3607), .A(n3606), .ZN(n3611) );
  INV_X1 U4380 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4843) );
  OAI22_X1 U4381 ( .A1(n4042), .A2(n3715), .B1(STATE_REG_SCAN_IN), .B2(n4843), 
        .ZN(n3609) );
  OAI22_X1 U4382 ( .A1(n3700), .A2(n3803), .B1(n3634), .B2(n4543), .ZN(n3608)
         );
  AOI211_X1 U4383 ( .C1(n4017), .C2(n4547), .A(n3609), .B(n3608), .ZN(n3610)
         );
  OAI21_X1 U4384 ( .B1(n3612), .B2(n3611), .A(n3610), .ZN(U3213) );
  XOR2_X1 U4385 ( .A(n3614), .B(n3613), .Z(n3619) );
  NAND2_X1 U4386 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4303) );
  OAI21_X1 U4387 ( .B1(n4134), .B2(n3715), .A(n4303), .ZN(n3616) );
  OAI22_X1 U4388 ( .A1(n3700), .A2(n4095), .B1(n4090), .B2(n4543), .ZN(n3615)
         );
  AOI211_X1 U4389 ( .C1(n3617), .C2(n4547), .A(n3616), .B(n3615), .ZN(n3618)
         );
  OAI21_X1 U4390 ( .B1(n3619), .B2(n4551), .A(n3618), .ZN(U3216) );
  XNOR2_X1 U4391 ( .A(n3621), .B(n3620), .ZN(n3622) );
  XNOR2_X1 U4392 ( .A(n2168), .B(n3622), .ZN(n3627) );
  OAI22_X1 U4393 ( .A1(n4090), .A2(n3715), .B1(STATE_REG_SCAN_IN), .B2(n3623), 
        .ZN(n3625) );
  OAI22_X1 U4394 ( .A1(n3700), .A2(n4049), .B1(n4042), .B2(n4543), .ZN(n3624)
         );
  AOI211_X1 U4395 ( .C1(n4050), .C2(n4547), .A(n3625), .B(n3624), .ZN(n3626)
         );
  OAI21_X1 U4396 ( .B1(n3627), .B2(n4551), .A(n3626), .ZN(U3220) );
  NAND2_X1 U4397 ( .A1(n3629), .A2(n3628), .ZN(n3631) );
  XOR2_X1 U4398 ( .A(n3631), .B(n3630), .Z(n3639) );
  INV_X1 U4399 ( .A(n3632), .ZN(n3977) );
  OAI22_X1 U4400 ( .A1(n3634), .A2(n3715), .B1(STATE_REG_SCAN_IN), .B2(n3633), 
        .ZN(n3637) );
  OAI22_X1 U4401 ( .A1(n3635), .A2(n4543), .B1(n3700), .B2(n3975), .ZN(n3636)
         );
  AOI211_X1 U4402 ( .C1(n3977), .C2(n4547), .A(n3637), .B(n3636), .ZN(n3638)
         );
  OAI21_X1 U4403 ( .B1(n3639), .B2(n4551), .A(n3638), .ZN(U3222) );
  AOI21_X1 U4404 ( .B1(n3710), .B2(n3708), .A(n3707), .ZN(n3641) );
  XNOR2_X1 U4405 ( .A(n3641), .B(n3640), .ZN(n3648) );
  NAND2_X1 U4406 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4412) );
  OAI21_X1 U4407 ( .B1(n3642), .B2(n3715), .A(n4412), .ZN(n3645) );
  OAI22_X1 U4408 ( .A1(n3700), .A2(n3643), .B1(n4113), .B2(n4543), .ZN(n3644)
         );
  AOI211_X1 U4409 ( .C1(n3646), .C2(n4547), .A(n3645), .B(n3644), .ZN(n3647)
         );
  OAI21_X1 U4410 ( .B1(n3648), .B2(n4551), .A(n3647), .ZN(U3223) );
  XNOR2_X1 U4411 ( .A(n3651), .B(n3650), .ZN(n3652) );
  XNOR2_X1 U4412 ( .A(n3649), .B(n3652), .ZN(n3657) );
  AOI22_X1 U4413 ( .A1(n4542), .A2(n4141), .B1(n3712), .B2(n4092), .ZN(n3656)
         );
  AND2_X1 U4414 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4423) );
  NOR2_X1 U4415 ( .A1(n3653), .A2(n3715), .ZN(n3654) );
  AOI211_X1 U4416 ( .C1(n4144), .C2(n4547), .A(n4423), .B(n3654), .ZN(n3655)
         );
  OAI211_X1 U4417 ( .C1(n3657), .C2(n4551), .A(n3656), .B(n3655), .ZN(U3225)
         );
  NAND2_X1 U4418 ( .A1(n3659), .A2(n3658), .ZN(n3660) );
  XOR2_X1 U4419 ( .A(n3661), .B(n3660), .Z(n3665) );
  INV_X1 U4420 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4853) );
  OAI22_X1 U4421 ( .A1(n3993), .A2(n3715), .B1(STATE_REG_SCAN_IN), .B2(n4853), 
        .ZN(n3663) );
  OAI22_X1 U4422 ( .A1(n3700), .A2(n3995), .B1(n3699), .B2(n4543), .ZN(n3662)
         );
  AOI211_X1 U4423 ( .C1(n3997), .C2(n4547), .A(n3663), .B(n3662), .ZN(n3664)
         );
  OAI21_X1 U4424 ( .B1(n3665), .B2(n4551), .A(n3664), .ZN(U3226) );
  OR2_X1 U4425 ( .A1(n3667), .A2(n3666), .ZN(n3668) );
  AOI22_X1 U4426 ( .A1(n3670), .A2(n2227), .B1(n3669), .B2(n3668), .ZN(n3675)
         );
  INV_X1 U4427 ( .A(n4110), .ZN(n3671) );
  INV_X1 U4428 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4852) );
  OAI22_X1 U4429 ( .A1(n3671), .A2(n3715), .B1(STATE_REG_SCAN_IN), .B2(n4852), 
        .ZN(n3673) );
  OAI22_X1 U4430 ( .A1(n3700), .A2(n4066), .B1(n4067), .B2(n4543), .ZN(n3672)
         );
  AOI211_X1 U4431 ( .C1(n4074), .C2(n4547), .A(n3673), .B(n3672), .ZN(n3674)
         );
  OAI21_X1 U4432 ( .B1(n3675), .B2(n4551), .A(n3674), .ZN(U3230) );
  OAI21_X1 U4433 ( .B1(n3677), .B2(n3676), .A(n3605), .ZN(n3679) );
  NAND2_X1 U4434 ( .A1(n3679), .A2(n3678), .ZN(n3683) );
  OAI22_X1 U4435 ( .A1(n4067), .A2(n3715), .B1(STATE_REG_SCAN_IN), .B2(n4850), 
        .ZN(n3681) );
  OAI22_X1 U4436 ( .A1(n3700), .A2(n4034), .B1(n3993), .B2(n4543), .ZN(n3680)
         );
  AOI211_X1 U4437 ( .C1(n4033), .C2(n4547), .A(n3681), .B(n3680), .ZN(n3682)
         );
  NAND2_X1 U4438 ( .A1(n3683), .A2(n3682), .ZN(U3232) );
  INV_X1 U4439 ( .A(n3684), .ZN(n3686) );
  NOR2_X1 U4440 ( .A1(n3686), .A2(n3685), .ZN(n3687) );
  XNOR2_X1 U4441 ( .A(n3688), .B(n3687), .ZN(n3693) );
  AOI22_X1 U4442 ( .A1(n4542), .A2(n4108), .B1(n3712), .B2(n4110), .ZN(n3692)
         );
  NOR2_X1 U4443 ( .A1(n3689), .A2(STATE_REG_SCAN_IN), .ZN(n4439) );
  NOR2_X1 U4444 ( .A1(n4113), .A2(n3715), .ZN(n3690) );
  AOI211_X1 U4445 ( .C1(n4121), .C2(n4547), .A(n4439), .B(n3690), .ZN(n3691)
         );
  OAI211_X1 U4446 ( .C1(n3693), .C2(n4551), .A(n3692), .B(n3691), .ZN(U3235)
         );
  INV_X1 U4447 ( .A(n3694), .ZN(n3695) );
  NOR2_X1 U4448 ( .A1(n3696), .A2(n3695), .ZN(n3697) );
  XNOR2_X1 U4449 ( .A(n3698), .B(n3697), .ZN(n3706) );
  INV_X1 U4450 ( .A(n3958), .ZN(n3704) );
  OAI22_X1 U4451 ( .A1(n3699), .A2(n3715), .B1(STATE_REG_SCAN_IN), .B2(n4844), 
        .ZN(n3703) );
  OAI22_X1 U4452 ( .A1(n3701), .A2(n4543), .B1(n3700), .B2(n3956), .ZN(n3702)
         );
  AOI211_X1 U4453 ( .C1(n3704), .C2(n4547), .A(n3703), .B(n3702), .ZN(n3705)
         );
  OAI21_X1 U4454 ( .B1(n3706), .B2(n4551), .A(n3705), .ZN(U3237) );
  INV_X1 U4455 ( .A(n3707), .ZN(n3709) );
  NAND2_X1 U4456 ( .A1(n3709), .A2(n3708), .ZN(n3711) );
  XNOR2_X1 U4457 ( .A(n3711), .B(n3710), .ZN(n3721) );
  AOI22_X1 U4458 ( .A1(n4542), .A2(n3713), .B1(n3712), .B2(n4136), .ZN(n3720)
         );
  INV_X1 U4459 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3714) );
  NOR2_X1 U4460 ( .A1(STATE_REG_SCAN_IN), .A2(n3714), .ZN(n4405) );
  NOR2_X1 U4461 ( .A1(n3716), .A2(n3715), .ZN(n3717) );
  AOI211_X1 U4462 ( .C1(n3718), .C2(n4547), .A(n4405), .B(n3717), .ZN(n3719)
         );
  OAI211_X1 U4463 ( .C1(n3721), .C2(n4551), .A(n3720), .B(n3719), .ZN(U3238)
         );
  NAND2_X1 U4464 ( .A1(n3790), .A2(n3789), .ZN(n3722) );
  AND2_X1 U4465 ( .A1(n3723), .A2(n3722), .ZN(n3840) );
  INV_X1 U4466 ( .A(n3840), .ZN(n3779) );
  INV_X1 U4467 ( .A(n3724), .ZN(n3727) );
  OAI211_X1 U4468 ( .C1(n3727), .C2(n4256), .A(n3726), .B(n3725), .ZN(n3730)
         );
  NAND3_X1 U4469 ( .A1(n3730), .A2(n3729), .A3(n3728), .ZN(n3733) );
  NAND3_X1 U4470 ( .A1(n3733), .A2(n3732), .A3(n3731), .ZN(n3736) );
  NAND3_X1 U4471 ( .A1(n3736), .A2(n3735), .A3(n3734), .ZN(n3739) );
  NAND4_X1 U4472 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3752), .ZN(n3741)
         );
  NAND3_X1 U4473 ( .A1(n3741), .A2(n3807), .A3(n3740), .ZN(n3742) );
  NAND3_X1 U4474 ( .A1(n3742), .A2(n3750), .A3(n3753), .ZN(n3745) );
  AND3_X1 U4475 ( .A1(n3745), .A2(n3744), .A3(n3743), .ZN(n3749) );
  NAND2_X1 U4476 ( .A1(n3747), .A2(n3746), .ZN(n3756) );
  NOR3_X1 U4477 ( .A1(n3749), .A2(n3748), .A3(n3756), .ZN(n3763) );
  NOR2_X1 U4478 ( .A1(n2195), .A2(n3751), .ZN(n3755) );
  NAND4_X1 U4479 ( .A1(n3755), .A2(n3754), .A3(n3753), .A4(n3752), .ZN(n3759)
         );
  NAND2_X1 U4480 ( .A1(n3756), .A2(n3765), .ZN(n3841) );
  INV_X1 U4481 ( .A(n3841), .ZN(n3757) );
  AOI21_X1 U4482 ( .B1(n3759), .B2(n3758), .A(n3757), .ZN(n3762) );
  OAI211_X1 U4483 ( .C1(n3763), .C2(n3762), .A(n3761), .B(n3760), .ZN(n3770)
         );
  INV_X1 U4484 ( .A(n3764), .ZN(n3767) );
  NAND2_X1 U4485 ( .A1(n3766), .A2(n3765), .ZN(n3842) );
  OAI21_X1 U4486 ( .B1(n3767), .B2(n3842), .A(n3841), .ZN(n3769) );
  AOI21_X1 U4487 ( .B1(n3770), .B2(n3769), .A(n3768), .ZN(n3772) );
  INV_X1 U4488 ( .A(n3844), .ZN(n3771) );
  OAI211_X1 U4489 ( .C1(n3772), .C2(n3771), .A(n3848), .B(n3846), .ZN(n3773)
         );
  AOI211_X1 U4490 ( .C1(n3773), .C2(n3851), .A(n3850), .B(n3796), .ZN(n3774)
         );
  NOR2_X1 U4491 ( .A1(n3774), .A2(n3855), .ZN(n3776) );
  OAI21_X1 U4492 ( .B1(n3776), .B2(n3775), .A(n3859), .ZN(n3777) );
  AOI21_X1 U4493 ( .B1(n3856), .B2(n3777), .A(n3861), .ZN(n3778) );
  NOR4_X1 U4494 ( .A1(n3827), .A2(n3780), .A3(n3779), .A4(n3778), .ZN(n3795)
         );
  NAND2_X1 U4495 ( .A1(n3782), .A2(n3781), .ZN(n3862) );
  INV_X1 U4496 ( .A(n4163), .ZN(n4151) );
  INV_X1 U4497 ( .A(REG0_REG_31__SCAN_IN), .ZN(n3786) );
  NAND2_X1 U4498 ( .A1(n3783), .A2(REG1_REG_31__SCAN_IN), .ZN(n3785) );
  NAND2_X1 U4499 ( .A1(n2693), .A2(REG2_REG_31__SCAN_IN), .ZN(n3784) );
  OAI211_X1 U4500 ( .C1(n2395), .C2(n3786), .A(n3785), .B(n3784), .ZN(n4154)
         );
  AND2_X1 U4501 ( .A1(n3787), .A2(DATAI_31_), .ZN(n4155) );
  INV_X1 U4502 ( .A(n4155), .ZN(n4152) );
  NAND2_X1 U4503 ( .A1(n4154), .A2(n4152), .ZN(n3791) );
  OAI21_X1 U4504 ( .B1(n3885), .B2(n4151), .A(n3791), .ZN(n3788) );
  INV_X1 U4505 ( .A(n3788), .ZN(n3831) );
  OAI21_X1 U4506 ( .B1(n3790), .B2(n3789), .A(n3831), .ZN(n3860) );
  AOI21_X1 U4507 ( .B1(n3862), .B2(n3840), .A(n3860), .ZN(n3866) );
  INV_X1 U4508 ( .A(n3866), .ZN(n3794) );
  INV_X1 U4509 ( .A(n3791), .ZN(n3793) );
  INV_X1 U4510 ( .A(n4154), .ZN(n3867) );
  INV_X1 U4511 ( .A(n3885), .ZN(n3792) );
  NOR2_X1 U4512 ( .A1(n3792), .A2(n4163), .ZN(n3868) );
  AOI21_X1 U4513 ( .B1(n4155), .B2(n3867), .A(n3868), .ZN(n3804) );
  OAI22_X1 U4514 ( .A1(n3795), .A2(n3794), .B1(n3793), .B2(n3804), .ZN(n3875)
         );
  INV_X1 U4515 ( .A(n3796), .ZN(n4005) );
  AND2_X1 U4516 ( .A1(n3798), .A2(n3797), .ZN(n4064) );
  INV_X1 U4517 ( .A(n4057), .ZN(n3799) );
  NOR2_X1 U4518 ( .A1(n3799), .A2(n4058), .ZN(n4088) );
  INV_X1 U4519 ( .A(n3964), .ZN(n3801) );
  NOR2_X1 U4520 ( .A1(n3802), .A2(n3801), .ZN(n3986) );
  XNOR2_X1 U4521 ( .A(n4028), .B(n3803), .ZN(n4007) );
  INV_X1 U4522 ( .A(n4007), .ZN(n3805) );
  NAND4_X1 U4523 ( .A1(n3966), .A2(n3986), .A3(n3805), .A4(n3804), .ZN(n3806)
         );
  NOR3_X1 U4524 ( .A1(n4064), .A2(n4088), .A3(n3806), .ZN(n3826) );
  NOR4_X1 U4525 ( .A1(n2915), .A2(n2904), .A3(n3809), .A4(n3808), .ZN(n3824)
         );
  INV_X1 U4526 ( .A(n3810), .ZN(n3813) );
  NAND2_X1 U4527 ( .A1(n4082), .A2(n3846), .ZN(n4129) );
  NOR4_X1 U4528 ( .A1(n3813), .A2(n3812), .A3(n4129), .A4(n3811), .ZN(n3822)
         );
  INV_X1 U4529 ( .A(n3814), .ZN(n3817) );
  NAND4_X1 U4530 ( .A1(n3817), .A2(n4107), .A3(n3816), .A4(n3815), .ZN(n3820)
         );
  NOR4_X1 U4531 ( .A1(n3820), .A2(n3819), .A3(n4455), .A4(n3818), .ZN(n3821)
         );
  AND4_X1 U4532 ( .A1(n3824), .A2(n3823), .A3(n3822), .A4(n3821), .ZN(n3825)
         );
  NAND4_X1 U4533 ( .A1(n4023), .A2(n4041), .A3(n3826), .A4(n3825), .ZN(n3838)
         );
  INV_X1 U4534 ( .A(n3827), .ZN(n3839) );
  NAND2_X1 U4535 ( .A1(n3839), .A2(n3828), .ZN(n3947) );
  INV_X1 U4536 ( .A(n3947), .ZN(n3829) );
  NAND3_X1 U4537 ( .A1(n3933), .A2(n3830), .A3(n3829), .ZN(n3837) );
  NAND4_X1 U4538 ( .A1(n3834), .A2(n3833), .A3(n3832), .A4(n3831), .ZN(n3835)
         );
  OR4_X1 U4539 ( .A1(n3838), .A2(n3837), .A3(n3836), .A4(n3835), .ZN(n3873) );
  NAND3_X1 U4540 ( .A1(n3933), .A2(n3840), .A3(n3839), .ZN(n3865) );
  OAI21_X1 U4541 ( .B1(n3843), .B2(n3842), .A(n3841), .ZN(n3845) );
  NAND2_X1 U4542 ( .A1(n3845), .A2(n3844), .ZN(n3849) );
  NAND4_X1 U4543 ( .A1(n3849), .A2(n3848), .A3(n3847), .A4(n3846), .ZN(n3852)
         );
  AOI21_X1 U4544 ( .B1(n3852), .B2(n3851), .A(n3850), .ZN(n3854) );
  OAI21_X1 U4545 ( .B1(n3855), .B2(n3854), .A(n3853), .ZN(n3858) );
  INV_X1 U4546 ( .A(n3856), .ZN(n3857) );
  AOI21_X1 U4547 ( .B1(n3859), .B2(n3858), .A(n3857), .ZN(n3863) );
  NOR4_X1 U4548 ( .A1(n3863), .A2(n3862), .A3(n3861), .A4(n3860), .ZN(n3864)
         );
  AOI21_X1 U4549 ( .B1(n3866), .B2(n3865), .A(n3864), .ZN(n3871) );
  NOR2_X1 U4550 ( .A1(n4154), .A2(n4151), .ZN(n3870) );
  OAI21_X1 U4551 ( .B1(n3868), .B2(n3867), .A(n4155), .ZN(n3869) );
  OAI21_X1 U4552 ( .B1(n3871), .B2(n3870), .A(n3869), .ZN(n3872) );
  MUX2_X1 U4553 ( .A(n3873), .B(n3872), .S(n4256), .Z(n3874) );
  MUX2_X1 U4554 ( .A(n3875), .B(n3874), .S(n4257), .Z(n3876) );
  XNOR2_X1 U4555 ( .A(n3876), .B(n4305), .ZN(n3884) );
  NOR4_X1 U4556 ( .A1(n3904), .A2(n3879), .A3(n3878), .A4(n3877), .ZN(n3882)
         );
  OAI21_X1 U4557 ( .B1(n3883), .B2(n3880), .A(B_REG_SCAN_IN), .ZN(n3881) );
  OAI22_X1 U4558 ( .A1(n3884), .A2(n3883), .B1(n3882), .B2(n3881), .ZN(U3239)
         );
  MUX2_X1 U4559 ( .A(n4154), .B(DATAO_REG_31__SCAN_IN), .S(n3900), .Z(U3581)
         );
  MUX2_X1 U4560 ( .A(n3885), .B(DATAO_REG_30__SCAN_IN), .S(n3900), .Z(U3580)
         );
  MUX2_X1 U4561 ( .A(n3886), .B(DATAO_REG_28__SCAN_IN), .S(n3900), .Z(U3578)
         );
  MUX2_X1 U4562 ( .A(n3950), .B(DATAO_REG_27__SCAN_IN), .S(n3900), .Z(U3577)
         );
  MUX2_X1 U4563 ( .A(n3969), .B(DATAO_REG_26__SCAN_IN), .S(n3900), .Z(U3576)
         );
  MUX2_X1 U4564 ( .A(n4028), .B(DATAO_REG_23__SCAN_IN), .S(n3900), .Z(U3573)
         );
  MUX2_X1 U4565 ( .A(n4027), .B(DATAO_REG_21__SCAN_IN), .S(n3900), .Z(U3571)
         );
  MUX2_X1 U4566 ( .A(n4092), .B(DATAO_REG_18__SCAN_IN), .S(n3900), .Z(U3568)
         );
  MUX2_X1 U4567 ( .A(n3887), .B(DATAO_REG_17__SCAN_IN), .S(n3900), .Z(U3567)
         );
  MUX2_X1 U4568 ( .A(n4136), .B(DATAO_REG_16__SCAN_IN), .S(n3900), .Z(U3566)
         );
  MUX2_X1 U4569 ( .A(n3888), .B(DATAO_REG_14__SCAN_IN), .S(n3900), .Z(U3564)
         );
  MUX2_X1 U4570 ( .A(n3889), .B(DATAO_REG_12__SCAN_IN), .S(n3900), .Z(U3562)
         );
  MUX2_X1 U4571 ( .A(n3890), .B(DATAO_REG_10__SCAN_IN), .S(n3900), .Z(U3560)
         );
  MUX2_X1 U4572 ( .A(n3891), .B(DATAO_REG_8__SCAN_IN), .S(n3900), .Z(U3558) );
  MUX2_X1 U4573 ( .A(n3892), .B(DATAO_REG_6__SCAN_IN), .S(n3900), .Z(U3556) );
  MUX2_X1 U4574 ( .A(n3893), .B(DATAO_REG_4__SCAN_IN), .S(n3900), .Z(U3554) );
  MUX2_X1 U4575 ( .A(n3894), .B(DATAO_REG_3__SCAN_IN), .S(n3900), .Z(U3553) );
  MUX2_X1 U4576 ( .A(n3895), .B(DATAO_REG_0__SCAN_IN), .S(n3900), .Z(U3550) );
  NAND3_X1 U4577 ( .A1(n3898), .A2(n3897), .A3(n3896), .ZN(n3902) );
  AND2_X1 U4578 ( .A1(n4322), .A2(n4744), .ZN(n3899) );
  OR2_X1 U4579 ( .A1(n3899), .A2(n4311), .ZN(n4320) );
  AOI21_X1 U4580 ( .B1(n4320), .B2(n4830), .A(n3900), .ZN(n3901) );
  OAI211_X1 U4581 ( .C1(n3904), .C2(n3903), .A(n3902), .B(n3901), .ZN(n4337)
         );
  AOI22_X1 U4582 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4440), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3916) );
  NOR2_X1 U4583 ( .A1(n4448), .A2(n3906), .ZN(n3913) );
  AND3_X1 U4584 ( .A1(n3909), .A2(n3908), .A3(n3907), .ZN(n3910) );
  NOR3_X1 U4585 ( .A1(n4441), .A2(n3911), .A3(n3910), .ZN(n3912) );
  AOI211_X1 U4586 ( .C1(n4431), .C2(n3914), .A(n3913), .B(n3912), .ZN(n3915)
         );
  NAND3_X1 U4587 ( .A1(n4337), .A2(n3916), .A3(n3915), .ZN(U3242) );
  INV_X1 U4588 ( .A(n3917), .ZN(n3925) );
  NOR2_X1 U4589 ( .A1(n3918), .A2(n4146), .ZN(n3922) );
  INV_X1 U4590 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3919) );
  OAI22_X1 U4591 ( .A1(n3920), .A2(n4096), .B1(n3919), .B2(n4125), .ZN(n3921)
         );
  AOI211_X1 U4592 ( .C1(n3923), .C2(n4125), .A(n3922), .B(n3921), .ZN(n3924)
         );
  OAI21_X1 U4593 ( .B1(n3925), .B2(n4149), .A(n3924), .ZN(U3262) );
  OAI21_X1 U4594 ( .B1(n3927), .B2(n3933), .A(n3926), .ZN(n3932) );
  AOI22_X1 U4595 ( .A1(n3969), .A2(n4137), .B1(n3928), .B2(n4162), .ZN(n3929)
         );
  OAI21_X1 U4596 ( .B1(n3930), .B2(n4133), .A(n3929), .ZN(n3931) );
  AOI21_X1 U4597 ( .B1(n3932), .B2(n4115), .A(n3931), .ZN(n4169) );
  XNOR2_X1 U4598 ( .A(n3934), .B(n3933), .ZN(n4168) );
  NAND2_X1 U4599 ( .A1(n4168), .A2(n3935), .ZN(n3943) );
  OAI21_X1 U4600 ( .B1(n3954), .B2(n3937), .A(n3936), .ZN(n4171) );
  INV_X1 U4601 ( .A(n4171), .ZN(n3941) );
  INV_X1 U4602 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3938) );
  OAI22_X1 U4603 ( .A1(n3939), .A2(n4096), .B1(n3938), .B2(n4125), .ZN(n3940)
         );
  AOI21_X1 U4604 ( .B1(n3941), .B2(n4316), .A(n3940), .ZN(n3942) );
  OAI211_X1 U4605 ( .C1(n4169), .C2(n4315), .A(n3943), .B(n3942), .ZN(U3263)
         );
  XNOR2_X1 U4606 ( .A(n3944), .B(n3947), .ZN(n4173) );
  INV_X1 U4607 ( .A(n4173), .ZN(n3962) );
  NAND2_X1 U4608 ( .A1(n3946), .A2(n3945), .ZN(n3948) );
  XNOR2_X1 U4609 ( .A(n3948), .B(n3947), .ZN(n3953) );
  AOI22_X1 U4610 ( .A1(n3990), .A2(n4137), .B1(n3949), .B2(n4162), .ZN(n3952)
         );
  NAND2_X1 U4611 ( .A1(n3950), .A2(n4109), .ZN(n3951) );
  OAI211_X1 U4612 ( .C1(n3953), .C2(n4139), .A(n3952), .B(n3951), .ZN(n4172)
         );
  INV_X1 U4613 ( .A(n3954), .ZN(n3955) );
  OAI21_X1 U4614 ( .B1(n3973), .B2(n3956), .A(n3955), .ZN(n4226) );
  NOR2_X1 U4615 ( .A1(n4226), .A2(n4146), .ZN(n3960) );
  INV_X1 U4616 ( .A(REG2_REG_26__SCAN_IN), .ZN(n3957) );
  OAI22_X1 U4617 ( .A1(n3958), .A2(n4096), .B1(n4125), .B2(n3957), .ZN(n3959)
         );
  AOI211_X1 U4618 ( .C1(n4172), .C2(n4125), .A(n3960), .B(n3959), .ZN(n3961)
         );
  OAI21_X1 U4619 ( .B1(n3962), .B2(n4149), .A(n3961), .ZN(U3264) );
  XNOR2_X1 U4620 ( .A(n3963), .B(n3966), .ZN(n4176) );
  INV_X1 U4621 ( .A(n4176), .ZN(n3981) );
  NAND2_X1 U4622 ( .A1(n3965), .A2(n3964), .ZN(n3967) );
  XNOR2_X1 U4623 ( .A(n3967), .B(n3966), .ZN(n3972) );
  AOI22_X1 U4624 ( .A1(n3969), .A2(n4109), .B1(n4162), .B2(n3968), .ZN(n3971)
         );
  NAND2_X1 U4625 ( .A1(n4009), .A2(n4137), .ZN(n3970) );
  OAI211_X1 U4626 ( .C1(n3972), .C2(n4139), .A(n3971), .B(n3970), .ZN(n4175)
         );
  INV_X1 U4627 ( .A(n3994), .ZN(n3976) );
  INV_X1 U4628 ( .A(n3973), .ZN(n3974) );
  OAI21_X1 U4629 ( .B1(n3976), .B2(n3975), .A(n3974), .ZN(n4230) );
  AOI22_X1 U4630 ( .A1(n4458), .A2(REG2_REG_25__SCAN_IN), .B1(n3977), .B2(
        n4453), .ZN(n3978) );
  OAI21_X1 U4631 ( .B1(n4230), .B2(n4146), .A(n3978), .ZN(n3979) );
  AOI21_X1 U4632 ( .B1(n4175), .B2(n4125), .A(n3979), .ZN(n3980) );
  OAI21_X1 U4633 ( .B1(n3981), .B2(n4149), .A(n3980), .ZN(U3265) );
  XOR2_X1 U4634 ( .A(n3986), .B(n3982), .Z(n4180) );
  INV_X1 U4635 ( .A(n4180), .ZN(n4001) );
  INV_X1 U4636 ( .A(n3983), .ZN(n3984) );
  NAND2_X1 U4637 ( .A1(n3985), .A2(n3984), .ZN(n3987) );
  XNOR2_X1 U4638 ( .A(n3987), .B(n3986), .ZN(n3988) );
  NAND2_X1 U4639 ( .A1(n3988), .A2(n4115), .ZN(n3992) );
  AOI22_X1 U4640 ( .A1(n3990), .A2(n4109), .B1(n4162), .B2(n3989), .ZN(n3991)
         );
  OAI211_X1 U4641 ( .C1(n3993), .C2(n4112), .A(n3992), .B(n3991), .ZN(n4179)
         );
  INV_X1 U4642 ( .A(n4016), .ZN(n3996) );
  OAI21_X1 U4643 ( .B1(n3996), .B2(n3995), .A(n3994), .ZN(n4233) );
  AOI22_X1 U4644 ( .A1(n4458), .A2(REG2_REG_24__SCAN_IN), .B1(n3997), .B2(
        n4453), .ZN(n3998) );
  OAI21_X1 U4645 ( .B1(n4233), .B2(n4146), .A(n3998), .ZN(n3999) );
  AOI21_X1 U4646 ( .B1(n4179), .B2(n4125), .A(n3999), .ZN(n4000) );
  OAI21_X1 U4647 ( .B1(n4001), .B2(n4149), .A(n4000), .ZN(U3266) );
  XOR2_X1 U4648 ( .A(n4007), .B(n4002), .Z(n4183) );
  INV_X1 U4649 ( .A(n4183), .ZN(n4021) );
  INV_X1 U4650 ( .A(n4003), .ZN(n4004) );
  AOI21_X1 U4651 ( .B1(n4040), .B2(n4005), .A(n4004), .ZN(n4026) );
  OAI21_X1 U4652 ( .B1(n4026), .B2(n2924), .A(n4006), .ZN(n4008) );
  XNOR2_X1 U4653 ( .A(n4008), .B(n4007), .ZN(n4013) );
  AOI22_X1 U4654 ( .A1(n4009), .A2(n4109), .B1(n4014), .B2(n4162), .ZN(n4012)
         );
  NAND2_X1 U4655 ( .A1(n4010), .A2(n4137), .ZN(n4011) );
  OAI211_X1 U4656 ( .C1(n4013), .C2(n4139), .A(n4012), .B(n4011), .ZN(n4182)
         );
  NAND2_X1 U4657 ( .A1(n4188), .A2(n4014), .ZN(n4015) );
  NAND2_X1 U4658 ( .A1(n4016), .A2(n4015), .ZN(n4237) );
  AOI22_X1 U4659 ( .A1(n4458), .A2(REG2_REG_23__SCAN_IN), .B1(n4017), .B2(
        n4453), .ZN(n4018) );
  OAI21_X1 U4660 ( .B1(n4237), .B2(n4146), .A(n4018), .ZN(n4019) );
  AOI21_X1 U4661 ( .B1(n4182), .B2(n4125), .A(n4019), .ZN(n4020) );
  OAI21_X1 U4662 ( .B1(n4021), .B2(n4149), .A(n4020), .ZN(U3267) );
  NAND2_X1 U4663 ( .A1(n4022), .A2(n4023), .ZN(n4024) );
  NAND2_X1 U4664 ( .A1(n4025), .A2(n4024), .ZN(n4186) );
  XNOR2_X1 U4665 ( .A(n4026), .B(n2924), .ZN(n4032) );
  NAND2_X1 U4666 ( .A1(n4027), .A2(n4137), .ZN(n4030) );
  NAND2_X1 U4667 ( .A1(n4028), .A2(n4109), .ZN(n4029) );
  OAI211_X1 U4668 ( .C1(n4132), .C2(n4034), .A(n4030), .B(n4029), .ZN(n4031)
         );
  AOI21_X1 U4669 ( .B1(n4032), .B2(n4115), .A(n4031), .ZN(n4190) );
  AOI22_X1 U4670 ( .A1(n4458), .A2(REG2_REG_22__SCAN_IN), .B1(n4033), .B2(
        n4453), .ZN(n4036) );
  OR2_X1 U4671 ( .A1(n4047), .A2(n4034), .ZN(n4187) );
  NAND3_X1 U4672 ( .A1(n4188), .A2(n4187), .A3(n4316), .ZN(n4035) );
  OAI211_X1 U4673 ( .C1(n4190), .C2(n4315), .A(n4036), .B(n4035), .ZN(n4037)
         );
  INV_X1 U4674 ( .A(n4037), .ZN(n4038) );
  OAI21_X1 U4675 ( .B1(n4186), .B2(n4149), .A(n4038), .ZN(U3268) );
  XOR2_X1 U4676 ( .A(n4041), .B(n4039), .Z(n4194) );
  INV_X1 U4677 ( .A(n4194), .ZN(n4056) );
  XOR2_X1 U4678 ( .A(n4041), .B(n4040), .Z(n4046) );
  OAI22_X1 U4679 ( .A1(n4042), .A2(n4133), .B1(n4132), .B2(n4049), .ZN(n4043)
         );
  AOI21_X1 U4680 ( .B1(n4137), .B2(n4044), .A(n4043), .ZN(n4045) );
  OAI21_X1 U4681 ( .B1(n4046), .B2(n4139), .A(n4045), .ZN(n4193) );
  INV_X1 U4682 ( .A(n4047), .ZN(n4048) );
  OAI21_X1 U4683 ( .B1(n2206), .B2(n4049), .A(n4048), .ZN(n4241) );
  NOR2_X1 U4684 ( .A1(n4241), .A2(n4146), .ZN(n4054) );
  INV_X1 U4685 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4052) );
  INV_X1 U4686 ( .A(n4050), .ZN(n4051) );
  OAI22_X1 U4687 ( .A1(n4125), .A2(n4052), .B1(n4051), .B2(n4096), .ZN(n4053)
         );
  AOI211_X1 U4688 ( .C1(n4193), .C2(n4125), .A(n4054), .B(n4053), .ZN(n4055)
         );
  OAI21_X1 U4689 ( .B1(n4056), .B2(n4149), .A(n4055), .ZN(U3269) );
  NAND2_X1 U4690 ( .A1(n4081), .A2(n4057), .ZN(n4060) );
  INV_X1 U4691 ( .A(n4058), .ZN(n4059) );
  NAND2_X1 U4692 ( .A1(n4060), .A2(n4059), .ZN(n4061) );
  XNOR2_X1 U4693 ( .A(n4061), .B(n4064), .ZN(n4073) );
  NAND2_X1 U4694 ( .A1(n4063), .A2(n4062), .ZN(n4065) );
  XNOR2_X1 U4695 ( .A(n4065), .B(n4064), .ZN(n4070) );
  OAI22_X1 U4696 ( .A1(n4067), .A2(n4133), .B1(n4132), .B2(n4066), .ZN(n4068)
         );
  AOI21_X1 U4697 ( .B1(n4137), .B2(n4110), .A(n4068), .ZN(n4069) );
  OAI21_X1 U4698 ( .B1(n4070), .B2(n4139), .A(n4069), .ZN(n4071) );
  AOI21_X1 U4699 ( .B1(n4073), .B2(n4072), .A(n4071), .ZN(n4199) );
  INV_X1 U4700 ( .A(n4073), .ZN(n4200) );
  AOI22_X1 U4701 ( .A1(n4458), .A2(REG2_REG_20__SCAN_IN), .B1(n4074), .B2(
        n4453), .ZN(n4077) );
  NAND2_X1 U4702 ( .A1(n2164), .A2(n4075), .ZN(n4196) );
  NAND3_X1 U4703 ( .A1(n4197), .A2(n4316), .A3(n4196), .ZN(n4076) );
  OAI211_X1 U4704 ( .C1(n4200), .C2(n4078), .A(n4077), .B(n4076), .ZN(n4079)
         );
  INV_X1 U4705 ( .A(n4079), .ZN(n4080) );
  OAI21_X1 U4706 ( .B1(n4458), .B2(n4199), .A(n4080), .ZN(U3270) );
  XNOR2_X1 U4707 ( .A(n4081), .B(n4088), .ZN(n4202) );
  INV_X1 U4708 ( .A(n4202), .ZN(n4102) );
  INV_X1 U4709 ( .A(n4082), .ZN(n4083) );
  NOR2_X1 U4710 ( .A1(n4084), .A2(n4083), .ZN(n4106) );
  INV_X1 U4711 ( .A(n4085), .ZN(n4086) );
  AOI21_X1 U4712 ( .B1(n4106), .B2(n4087), .A(n4086), .ZN(n4089) );
  XNOR2_X1 U4713 ( .A(n4089), .B(n4088), .ZN(n4094) );
  OAI22_X1 U4714 ( .A1(n4090), .A2(n4133), .B1(n4132), .B2(n4095), .ZN(n4091)
         );
  AOI21_X1 U4715 ( .B1(n4137), .B2(n4092), .A(n4091), .ZN(n4093) );
  OAI21_X1 U4716 ( .B1(n4094), .B2(n4139), .A(n4093), .ZN(n4201) );
  OAI21_X1 U4717 ( .B1(n4118), .B2(n4095), .A(n2164), .ZN(n4245) );
  NOR2_X1 U4718 ( .A1(n4245), .A2(n4146), .ZN(n4100) );
  INV_X1 U4719 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4098) );
  OAI22_X1 U4720 ( .A1(n4125), .A2(n4098), .B1(n4097), .B2(n4096), .ZN(n4099)
         );
  AOI211_X1 U4721 ( .C1(n4201), .C2(n4125), .A(n4100), .B(n4099), .ZN(n4101)
         );
  OAI21_X1 U4722 ( .B1(n4102), .B2(n4149), .A(n4101), .ZN(U3271) );
  INV_X1 U4723 ( .A(n4103), .ZN(n4104) );
  AOI21_X1 U4724 ( .B1(n4107), .B2(n4105), .A(n4104), .ZN(n4207) );
  XOR2_X1 U4725 ( .A(n4107), .B(n4106), .Z(n4116) );
  AOI22_X1 U4726 ( .A1(n4110), .A2(n4109), .B1(n4108), .B2(n4162), .ZN(n4111)
         );
  OAI21_X1 U4727 ( .B1(n4113), .B2(n4112), .A(n4111), .ZN(n4114) );
  AOI21_X1 U4728 ( .B1(n4116), .B2(n4115), .A(n4114), .ZN(n4206) );
  INV_X1 U4729 ( .A(n4206), .ZN(n4126) );
  OAI21_X1 U4730 ( .B1(n4142), .B2(n4117), .A(n4506), .ZN(n4119) );
  OR2_X1 U4731 ( .A1(n4119), .A2(n4118), .ZN(n4205) );
  INV_X1 U4732 ( .A(n4120), .ZN(n4123) );
  AOI22_X1 U4733 ( .A1(n4315), .A2(REG2_REG_18__SCAN_IN), .B1(n4121), .B2(
        n4453), .ZN(n4122) );
  OAI21_X1 U4734 ( .B1(n4205), .B2(n4123), .A(n4122), .ZN(n4124) );
  AOI21_X1 U4735 ( .B1(n4126), .B2(n4125), .A(n4124), .ZN(n4127) );
  OAI21_X1 U4736 ( .B1(n4207), .B2(n4149), .A(n4127), .ZN(U3272) );
  XOR2_X1 U4737 ( .A(n4129), .B(n4128), .Z(n4209) );
  INV_X1 U4738 ( .A(n4209), .ZN(n4150) );
  XNOR2_X1 U4739 ( .A(n4130), .B(n4129), .ZN(n4140) );
  OAI22_X1 U4740 ( .A1(n4134), .A2(n4133), .B1(n4132), .B2(n4131), .ZN(n4135)
         );
  AOI21_X1 U4741 ( .B1(n4137), .B2(n4136), .A(n4135), .ZN(n4138) );
  OAI21_X1 U4742 ( .B1(n4140), .B2(n4139), .A(n4138), .ZN(n4208) );
  AND2_X1 U4743 ( .A1(n4213), .A2(n4141), .ZN(n4143) );
  OR2_X1 U4744 ( .A1(n4143), .A2(n4142), .ZN(n4250) );
  AOI22_X1 U4745 ( .A1(n4315), .A2(REG2_REG_17__SCAN_IN), .B1(n4144), .B2(
        n4453), .ZN(n4145) );
  OAI21_X1 U4746 ( .B1(n4250), .B2(n4146), .A(n4145), .ZN(n4147) );
  AOI21_X1 U4747 ( .B1(n4208), .B2(n4125), .A(n4147), .ZN(n4148) );
  OAI21_X1 U4748 ( .B1(n4150), .B2(n4149), .A(n4148), .ZN(U3273) );
  NAND2_X1 U4749 ( .A1(n4157), .A2(n4151), .ZN(n4158) );
  XNOR2_X1 U4750 ( .A(n4158), .B(n4152), .ZN(n4312) );
  INV_X1 U4751 ( .A(n4312), .ZN(n4218) );
  INV_X1 U4752 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4636) );
  AND2_X1 U4753 ( .A1(n4154), .A2(n4153), .ZN(n4161) );
  AOI21_X1 U4754 ( .B1(n4155), .B2(n4162), .A(n4161), .ZN(n4314) );
  MUX2_X1 U4755 ( .A(n4636), .B(n4314), .S(n4533), .Z(n4156) );
  OAI21_X1 U4756 ( .B1(n4218), .B2(n4211), .A(n4156), .ZN(U3549) );
  INV_X1 U4757 ( .A(n4157), .ZN(n4160) );
  INV_X1 U4758 ( .A(n4158), .ZN(n4159) );
  AOI21_X1 U4759 ( .B1(n4163), .B2(n4160), .A(n4159), .ZN(n4317) );
  INV_X1 U4760 ( .A(n4317), .ZN(n4220) );
  INV_X1 U4761 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4637) );
  AOI21_X1 U4762 ( .B1(n4163), .B2(n4162), .A(n4161), .ZN(n4319) );
  MUX2_X1 U4763 ( .A(n4637), .B(n4319), .S(n4533), .Z(n4164) );
  OAI21_X1 U4764 ( .B1(n4220), .B2(n4211), .A(n4164), .ZN(U3548) );
  NAND2_X1 U4765 ( .A1(n4168), .A2(n4496), .ZN(n4170) );
  OAI211_X1 U4766 ( .C1(n4512), .C2(n4171), .A(n4170), .B(n4169), .ZN(n4222)
         );
  MUX2_X1 U4767 ( .A(REG1_REG_27__SCAN_IN), .B(n4222), .S(n4533), .Z(U3545) );
  INV_X1 U4768 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4631) );
  AOI21_X1 U4769 ( .B1(n4173), .B2(n4496), .A(n4172), .ZN(n4223) );
  MUX2_X1 U4770 ( .A(n4631), .B(n4223), .S(n4533), .Z(n4174) );
  OAI21_X1 U4771 ( .B1(n4211), .B2(n4226), .A(n4174), .ZN(U3544) );
  INV_X1 U4772 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4177) );
  AOI21_X1 U4773 ( .B1(n4176), .B2(n4496), .A(n4175), .ZN(n4227) );
  MUX2_X1 U4774 ( .A(n4177), .B(n4227), .S(n4533), .Z(n4178) );
  OAI21_X1 U4775 ( .B1(n4211), .B2(n4230), .A(n4178), .ZN(U3543) );
  INV_X1 U4776 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4621) );
  AOI21_X1 U4777 ( .B1(n4180), .B2(n4496), .A(n4179), .ZN(n4231) );
  MUX2_X1 U4778 ( .A(n4621), .B(n4231), .S(n4533), .Z(n4181) );
  OAI21_X1 U4779 ( .B1(n4211), .B2(n4233), .A(n4181), .ZN(U3542) );
  INV_X1 U4780 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4184) );
  AOI21_X1 U4781 ( .B1(n4183), .B2(n4496), .A(n4182), .ZN(n4234) );
  MUX2_X1 U4782 ( .A(n4184), .B(n4234), .S(n4533), .Z(n4185) );
  OAI21_X1 U4783 ( .B1(n4211), .B2(n4237), .A(n4185), .ZN(U3541) );
  OR2_X1 U4784 ( .A1(n4186), .A2(n4501), .ZN(n4192) );
  NAND3_X1 U4785 ( .A1(n4188), .A2(n4187), .A3(n4506), .ZN(n4189) );
  AND2_X1 U4786 ( .A1(n4190), .A2(n4189), .ZN(n4191) );
  NAND2_X1 U4787 ( .A1(n4192), .A2(n4191), .ZN(n4238) );
  MUX2_X1 U4788 ( .A(REG1_REG_22__SCAN_IN), .B(n4238), .S(n4533), .Z(U3540) );
  INV_X1 U4789 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4775) );
  AOI21_X1 U4790 ( .B1(n4194), .B2(n4496), .A(n4193), .ZN(n4239) );
  MUX2_X1 U4791 ( .A(n4775), .B(n4239), .S(n4533), .Z(n4195) );
  OAI21_X1 U4792 ( .B1(n4211), .B2(n4241), .A(n4195), .ZN(U3539) );
  NAND3_X1 U4793 ( .A1(n4197), .A2(n4506), .A3(n4196), .ZN(n4198) );
  OAI211_X1 U4794 ( .C1(n4200), .C2(n4480), .A(n4199), .B(n4198), .ZN(n4242)
         );
  MUX2_X1 U4795 ( .A(REG1_REG_20__SCAN_IN), .B(n4242), .S(n4533), .Z(U3538) );
  INV_X1 U4796 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4203) );
  AOI21_X1 U4797 ( .B1(n4202), .B2(n4496), .A(n4201), .ZN(n4243) );
  MUX2_X1 U4798 ( .A(n4203), .B(n4243), .S(n4533), .Z(n4204) );
  OAI21_X1 U4799 ( .B1(n4211), .B2(n4245), .A(n4204), .ZN(U3537) );
  OAI211_X1 U4800 ( .C1(n4207), .C2(n4501), .A(n4206), .B(n4205), .ZN(n4246)
         );
  MUX2_X1 U4801 ( .A(REG1_REG_18__SCAN_IN), .B(n4246), .S(n4533), .Z(U3536) );
  INV_X1 U4802 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4278) );
  AOI21_X1 U4803 ( .B1(n4209), .B2(n4496), .A(n4208), .ZN(n4247) );
  MUX2_X1 U4804 ( .A(n4278), .B(n4247), .S(n4533), .Z(n4210) );
  OAI21_X1 U4805 ( .B1(n4211), .B2(n4250), .A(n4210), .ZN(U3535) );
  NAND3_X1 U4806 ( .A1(n4213), .A2(n4506), .A3(n4212), .ZN(n4214) );
  OAI211_X1 U4807 ( .C1(n4216), .C2(n4501), .A(n4215), .B(n4214), .ZN(n4251)
         );
  MUX2_X1 U4808 ( .A(REG1_REG_16__SCAN_IN), .B(n4251), .S(n4533), .Z(U3534) );
  MUX2_X1 U4809 ( .A(n3786), .B(n4314), .S(n4520), .Z(n4217) );
  OAI21_X1 U4810 ( .B1(n4218), .B2(n4249), .A(n4217), .ZN(U3517) );
  MUX2_X1 U4811 ( .A(n3595), .B(n4319), .S(n4520), .Z(n4219) );
  OAI21_X1 U4812 ( .B1(n4220), .B2(n4249), .A(n4219), .ZN(U3516) );
  MUX2_X1 U4813 ( .A(REG0_REG_29__SCAN_IN), .B(n4221), .S(n4520), .Z(U3515) );
  MUX2_X1 U4814 ( .A(REG0_REG_27__SCAN_IN), .B(n4222), .S(n4520), .Z(U3513) );
  INV_X1 U4815 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4224) );
  MUX2_X1 U4816 ( .A(n4224), .B(n4223), .S(n4520), .Z(n4225) );
  OAI21_X1 U4817 ( .B1(n4226), .B2(n4249), .A(n4225), .ZN(U3512) );
  INV_X1 U4818 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4228) );
  MUX2_X1 U4819 ( .A(n4228), .B(n4227), .S(n4520), .Z(n4229) );
  OAI21_X1 U4820 ( .B1(n4230), .B2(n4249), .A(n4229), .ZN(U3511) );
  INV_X1 U4821 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4624) );
  MUX2_X1 U4822 ( .A(n4624), .B(n4231), .S(n4520), .Z(n4232) );
  OAI21_X1 U4823 ( .B1(n4233), .B2(n4249), .A(n4232), .ZN(U3510) );
  INV_X1 U4824 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4235) );
  MUX2_X1 U4825 ( .A(n4235), .B(n4234), .S(n4520), .Z(n4236) );
  OAI21_X1 U4826 ( .B1(n4237), .B2(n4249), .A(n4236), .ZN(U3509) );
  MUX2_X1 U4827 ( .A(REG0_REG_22__SCAN_IN), .B(n4238), .S(n4520), .Z(U3508) );
  INV_X1 U4828 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4615) );
  MUX2_X1 U4829 ( .A(n4615), .B(n4239), .S(n4520), .Z(n4240) );
  OAI21_X1 U4830 ( .B1(n4241), .B2(n4249), .A(n4240), .ZN(U3507) );
  MUX2_X1 U4831 ( .A(REG0_REG_20__SCAN_IN), .B(n4242), .S(n4520), .Z(U3506) );
  INV_X1 U4832 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4770) );
  MUX2_X1 U4833 ( .A(n4770), .B(n4243), .S(n4520), .Z(n4244) );
  OAI21_X1 U4834 ( .B1(n4245), .B2(n4249), .A(n4244), .ZN(U3505) );
  MUX2_X1 U4835 ( .A(REG0_REG_18__SCAN_IN), .B(n4246), .S(n4520), .Z(U3503) );
  INV_X1 U4836 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4773) );
  MUX2_X1 U4837 ( .A(n4773), .B(n4247), .S(n4520), .Z(n4248) );
  OAI21_X1 U4838 ( .B1(n4250), .B2(n4249), .A(n4248), .ZN(U3501) );
  MUX2_X1 U4839 ( .A(REG0_REG_16__SCAN_IN), .B(n4251), .S(n4520), .Z(U3499) );
  MUX2_X1 U4840 ( .A(n4252), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U4841 ( .A(n4253), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U4842 ( .A(n4254), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4843 ( .A(DATAI_24_), .B(n4255), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U4844 ( .A(n4256), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U4845 ( .A(DATAI_20_), .B(n4257), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  INV_X1 U4846 ( .A(n4280), .ZN(n4258) );
  MUX2_X1 U4847 ( .A(DATAI_8_), .B(n4258), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U4848 ( .A(n4259), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4849 ( .A(n4260), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4850 ( .A(n4261), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4851 ( .A(DATAI_4_), .B(n4336), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4852 ( .A(n4262), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4853 ( .A(n4098), .B(REG2_REG_19__SCAN_IN), .S(n4305), .Z(n4277) );
  NAND2_X1 U4854 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4300), .ZN(n4263) );
  OAI21_X1 U4855 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4300), .A(n4263), .ZN(n4444) );
  NOR2_X1 U4856 ( .A1(n4299), .A2(REG2_REG_17__SCAN_IN), .ZN(n4264) );
  AOI21_X1 U4857 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4299), .A(n4264), .ZN(n4426) );
  INV_X1 U4858 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4382) );
  NOR2_X1 U4859 ( .A1(n4382), .A2(n4468), .ZN(n4381) );
  NAND2_X1 U4860 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4287), .ZN(n4270) );
  INV_X1 U4861 ( .A(n4287), .ZN(n4471) );
  INV_X1 U4862 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4745) );
  AOI22_X1 U4863 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4287), .B1(n4471), .B2(
        n4745), .ZN(n4365) );
  AOI22_X1 U4864 ( .A1(n4283), .A2(REG2_REG_9__SCAN_IN), .B1(n3368), .B2(n4475), .ZN(n4346) );
  INV_X1 U4865 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4266) );
  OAI22_X1 U4866 ( .A1(n4267), .A2(n4266), .B1(n4265), .B2(n4280), .ZN(n4345)
         );
  NAND2_X1 U4867 ( .A1(n4346), .A2(n4345), .ZN(n4344) );
  OAI21_X1 U4868 ( .B1(n3368), .B2(n4475), .A(n4344), .ZN(n4268) );
  NAND2_X1 U4869 ( .A1(n4285), .A2(n4268), .ZN(n4269) );
  XNOR2_X1 U4870 ( .A(n2262), .B(n4268), .ZN(n4355) );
  NAND2_X1 U4871 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4355), .ZN(n4354) );
  NAND2_X1 U4872 ( .A1(n4288), .A2(n4271), .ZN(n4272) );
  NAND2_X1 U4873 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4374), .ZN(n4373) );
  NOR2_X1 U4874 ( .A1(n2223), .A2(n4273), .ZN(n4274) );
  INV_X1 U4875 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4390) );
  INV_X1 U4876 ( .A(n4296), .ZN(n4467) );
  AOI22_X1 U4877 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4467), .B1(n4296), .B2(
        n3472), .ZN(n4408) );
  NAND2_X1 U4878 ( .A1(n4275), .A2(n4465), .ZN(n4276) );
  INV_X1 U4879 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4415) );
  NAND2_X1 U4880 ( .A1(n4276), .A2(n4414), .ZN(n4425) );
  NAND2_X1 U4881 ( .A1(n4426), .A2(n4425), .ZN(n4424) );
  INV_X1 U4882 ( .A(n4300), .ZN(n4462) );
  INV_X1 U4883 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4821) );
  AOI22_X1 U4884 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4462), .B1(n4300), .B2(
        n4821), .ZN(n4438) );
  AOI22_X1 U4885 ( .A1(n4299), .A2(REG1_REG_17__SCAN_IN), .B1(n4278), .B2(
        n4463), .ZN(n4429) );
  OAI21_X1 U4886 ( .B1(n4281), .B2(n4280), .A(n4279), .ZN(n4282) );
  INV_X1 U4887 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4527) );
  AOI22_X1 U4888 ( .A1(n4283), .A2(n4527), .B1(REG1_REG_9__SCAN_IN), .B2(n4475), .ZN(n4340) );
  NOR2_X1 U4889 ( .A1(n4284), .A2(n2262), .ZN(n4286) );
  INV_X1 U4890 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4788) );
  NOR2_X1 U4891 ( .A1(n4788), .A2(n4350), .ZN(n4349) );
  INV_X1 U4892 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4531) );
  AOI22_X1 U4893 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4471), .B1(n4287), .B2(
        n4531), .ZN(n4359) );
  NOR2_X1 U4894 ( .A1(n4360), .A2(n4359), .ZN(n4358) );
  INV_X1 U4895 ( .A(n4288), .ZN(n4469) );
  NOR2_X1 U4896 ( .A1(n4289), .A2(n4469), .ZN(n4290) );
  INV_X1 U4897 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4743) );
  AOI22_X1 U4898 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4468), .B1(n4292), .B2(
        n4291), .ZN(n4378) );
  NOR2_X1 U4899 ( .A1(n4293), .A2(n2223), .ZN(n4294) );
  XOR2_X1 U4900 ( .A(n4396), .B(n4293), .Z(n4392) );
  NOR2_X1 U4901 ( .A1(n4393), .A2(n4392), .ZN(n4391) );
  AOI22_X1 U4902 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4467), .B1(n4296), .B2(
        n4295), .ZN(n4402) );
  NOR2_X1 U4903 ( .A1(n4403), .A2(n4402), .ZN(n4401) );
  NAND2_X1 U4904 ( .A1(n4297), .A2(n4465), .ZN(n4298) );
  INV_X1 U4905 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4792) );
  NAND2_X1 U4906 ( .A1(n4429), .A2(n4428), .ZN(n4427) );
  AOI21_X1 U4907 ( .B1(n4300), .B2(REG1_REG_18__SCAN_IN), .A(n4437), .ZN(n4302) );
  XNOR2_X1 U4908 ( .A(n4305), .B(REG1_REG_19__SCAN_IN), .ZN(n4301) );
  XNOR2_X1 U4909 ( .A(n4302), .B(n4301), .ZN(n4307) );
  NAND2_X1 U4910 ( .A1(n4440), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4304) );
  OAI211_X1 U4911 ( .C1(n4448), .C2(n4305), .A(n4304), .B(n4303), .ZN(n4306)
         );
  AOI21_X1 U4912 ( .B1(n4307), .B2(n4431), .A(n4306), .ZN(n4308) );
  OAI21_X1 U4913 ( .B1(n4309), .B2(n4441), .A(n4308), .ZN(U3259) );
  INV_X1 U4914 ( .A(DATAI_28_), .ZN(n4310) );
  AOI22_X1 U4915 ( .A1(STATE_REG_SCAN_IN), .A2(n4311), .B1(n4310), .B2(U3149), 
        .ZN(U3324) );
  AOI22_X1 U4916 ( .A1(n4312), .A2(n4316), .B1(n4315), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4313) );
  OAI21_X1 U4917 ( .B1(n4458), .B2(n4314), .A(n4313), .ZN(U3260) );
  AOI22_X1 U4918 ( .A1(n4317), .A2(n4316), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4315), .ZN(n4318) );
  OAI21_X1 U4919 ( .B1(n4458), .B2(n4319), .A(n4318), .ZN(U3261) );
  INV_X1 U4920 ( .A(n4320), .ZN(n4321) );
  OAI21_X1 U4921 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4322), .A(n4321), .ZN(n4323)
         );
  XOR2_X1 U4922 ( .A(n4323), .B(IR_REG_0__SCAN_IN), .Z(n4326) );
  AOI22_X1 U4923 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4440), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4324) );
  OAI21_X1 U4924 ( .B1(n4326), .B2(n4325), .A(n4324), .ZN(U3240) );
  XNOR2_X1 U4925 ( .A(n4327), .B(REG2_REG_4__SCAN_IN), .ZN(n4330) );
  XOR2_X1 U4926 ( .A(n4328), .B(REG1_REG_4__SCAN_IN), .Z(n4329) );
  OAI22_X1 U4927 ( .A1(n4330), .A2(n4441), .B1(n4436), .B2(n4329), .ZN(n4335)
         );
  INV_X1 U4928 ( .A(n4440), .ZN(n4333) );
  INV_X1 U4929 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4332) );
  OAI21_X1 U4930 ( .B1(n4333), .B2(n4332), .A(n4331), .ZN(n4334) );
  AOI211_X1 U4931 ( .C1(n4336), .C2(n4397), .A(n4335), .B(n4334), .ZN(n4338)
         );
  NAND2_X1 U4932 ( .A1(n4338), .A2(n4337), .ZN(U3244) );
  AOI211_X1 U4933 ( .C1(n4341), .C2(n4340), .A(n4339), .B(n4436), .ZN(n4342)
         );
  AOI211_X1 U4934 ( .C1(n4440), .C2(ADDR_REG_9__SCAN_IN), .A(n4343), .B(n4342), 
        .ZN(n4348) );
  OAI211_X1 U4935 ( .C1(n4346), .C2(n4345), .A(n4433), .B(n4344), .ZN(n4347)
         );
  OAI211_X1 U4936 ( .C1(n4448), .C2(n4475), .A(n4348), .B(n4347), .ZN(U3249)
         );
  AOI211_X1 U4937 ( .C1(n4788), .C2(n4350), .A(n4349), .B(n4436), .ZN(n4353)
         );
  INV_X1 U4938 ( .A(n4351), .ZN(n4352) );
  AOI211_X1 U4939 ( .C1(n4440), .C2(ADDR_REG_10__SCAN_IN), .A(n4353), .B(n4352), .ZN(n4357) );
  OAI211_X1 U4940 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4355), .A(n4433), .B(n4354), .ZN(n4356) );
  OAI211_X1 U4941 ( .C1(n4448), .C2(n2262), .A(n4357), .B(n4356), .ZN(U3250)
         );
  AOI211_X1 U4942 ( .C1(n4360), .C2(n4359), .A(n4358), .B(n4436), .ZN(n4362)
         );
  AOI211_X1 U4943 ( .C1(n4440), .C2(ADDR_REG_11__SCAN_IN), .A(n4362), .B(n4361), .ZN(n4367) );
  OAI211_X1 U4944 ( .C1(n4365), .C2(n4364), .A(n4433), .B(n4363), .ZN(n4366)
         );
  OAI211_X1 U4945 ( .C1(n4448), .C2(n4471), .A(n4367), .B(n4366), .ZN(U3251)
         );
  AOI211_X1 U4946 ( .C1(n4743), .C2(n4369), .A(n4368), .B(n4436), .ZN(n4372)
         );
  INV_X1 U4947 ( .A(n4370), .ZN(n4371) );
  AOI211_X1 U4948 ( .C1(n4440), .C2(ADDR_REG_12__SCAN_IN), .A(n4372), .B(n4371), .ZN(n4376) );
  OAI211_X1 U4949 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4374), .A(n4433), .B(n4373), .ZN(n4375) );
  OAI211_X1 U4950 ( .C1(n4448), .C2(n4469), .A(n4376), .B(n4375), .ZN(U3252)
         );
  AOI211_X1 U4951 ( .C1(n2179), .C2(n4378), .A(n4377), .B(n4436), .ZN(n4379)
         );
  AOI211_X1 U4952 ( .C1(n4440), .C2(ADDR_REG_13__SCAN_IN), .A(n4380), .B(n4379), .ZN(n4387) );
  AOI21_X1 U4953 ( .B1(n4382), .B2(n4468), .A(n4381), .ZN(n4385) );
  AOI21_X1 U4954 ( .B1(n4385), .B2(n4384), .A(n4441), .ZN(n4383) );
  OAI21_X1 U4955 ( .B1(n4385), .B2(n4384), .A(n4383), .ZN(n4386) );
  OAI211_X1 U4956 ( .C1(n4448), .C2(n4468), .A(n4387), .B(n4386), .ZN(U3253)
         );
  NAND2_X1 U4957 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4440), .ZN(n4400) );
  AOI211_X1 U4958 ( .C1(n4390), .C2(n4389), .A(n4388), .B(n4441), .ZN(n4395)
         );
  AOI211_X1 U4959 ( .C1(n4393), .C2(n4392), .A(n4391), .B(n4436), .ZN(n4394)
         );
  AOI211_X1 U4960 ( .C1(n4397), .C2(n4396), .A(n4395), .B(n4394), .ZN(n4399)
         );
  NAND3_X1 U4961 ( .A1(n4400), .A2(n4399), .A3(n4398), .ZN(U3254) );
  AOI211_X1 U4962 ( .C1(n4403), .C2(n4402), .A(n4401), .B(n4436), .ZN(n4404)
         );
  AOI211_X1 U4963 ( .C1(n4440), .C2(ADDR_REG_15__SCAN_IN), .A(n4405), .B(n4404), .ZN(n4411) );
  AOI21_X1 U4964 ( .B1(n4408), .B2(n4407), .A(n4406), .ZN(n4409) );
  NAND2_X1 U4965 ( .A1(n4433), .A2(n4409), .ZN(n4410) );
  OAI211_X1 U4966 ( .C1(n4448), .C2(n4467), .A(n4411), .B(n4410), .ZN(U3255)
         );
  INV_X1 U4967 ( .A(n4412), .ZN(n4413) );
  AOI21_X1 U4968 ( .B1(n4440), .B2(ADDR_REG_16__SCAN_IN), .A(n4413), .ZN(n4422) );
  OAI21_X1 U4969 ( .B1(n4416), .B2(n4415), .A(n4414), .ZN(n4420) );
  OAI21_X1 U4970 ( .B1(n4418), .B2(n4792), .A(n4417), .ZN(n4419) );
  AOI22_X1 U4971 ( .A1(n4433), .A2(n4420), .B1(n4431), .B2(n4419), .ZN(n4421)
         );
  OAI211_X1 U4972 ( .C1(n4465), .C2(n4448), .A(n4422), .B(n4421), .ZN(U3256)
         );
  AOI21_X1 U4973 ( .B1(n4440), .B2(ADDR_REG_17__SCAN_IN), .A(n4423), .ZN(n4435) );
  OAI21_X1 U4974 ( .B1(n4426), .B2(n4425), .A(n4424), .ZN(n4432) );
  OAI21_X1 U4975 ( .B1(n4429), .B2(n4428), .A(n4427), .ZN(n4430) );
  AOI22_X1 U4976 ( .A1(n4433), .A2(n4432), .B1(n4431), .B2(n4430), .ZN(n4434)
         );
  OAI211_X1 U4977 ( .C1(n4463), .C2(n4448), .A(n4435), .B(n4434), .ZN(U3257)
         );
  AOI211_X1 U4978 ( .C1(n4444), .C2(n4443), .A(n4442), .B(n4441), .ZN(n4445)
         );
  INV_X1 U4979 ( .A(n4445), .ZN(n4446) );
  OAI211_X1 U4980 ( .C1(n4448), .C2(n4462), .A(n4447), .B(n4446), .ZN(U3258)
         );
  INV_X1 U4981 ( .A(n4449), .ZN(n4451) );
  AOI21_X1 U4982 ( .B1(n4452), .B2(n4451), .A(n4450), .ZN(n4457) );
  AOI22_X1 U4983 ( .A1(n4455), .A2(n4454), .B1(REG3_REG_0__SCAN_IN), .B2(n4453), .ZN(n4456) );
  OAI221_X1 U4984 ( .B1(n4458), .B2(n4457), .C1(n4125), .C2(n4744), .A(n4456), 
        .ZN(U3290) );
  INV_X1 U4985 ( .A(D_REG_31__SCAN_IN), .ZN(n4648) );
  NOR2_X1 U4986 ( .A1(n4460), .A2(n4648), .ZN(U3291) );
  INV_X1 U4987 ( .A(D_REG_30__SCAN_IN), .ZN(n4652) );
  NOR2_X1 U4988 ( .A1(n4460), .A2(n4652), .ZN(U3292) );
  AND2_X1 U4989 ( .A1(D_REG_29__SCAN_IN), .A2(n4459), .ZN(U3293) );
  INV_X1 U4990 ( .A(D_REG_28__SCAN_IN), .ZN(n4662) );
  NOR2_X1 U4991 ( .A1(n4460), .A2(n4662), .ZN(U3294) );
  AND2_X1 U4992 ( .A1(D_REG_27__SCAN_IN), .A2(n4459), .ZN(U3295) );
  AND2_X1 U4993 ( .A1(D_REG_26__SCAN_IN), .A2(n4459), .ZN(U3296) );
  AND2_X1 U4994 ( .A1(D_REG_25__SCAN_IN), .A2(n4459), .ZN(U3297) );
  INV_X1 U4995 ( .A(D_REG_24__SCAN_IN), .ZN(n4696) );
  NOR2_X1 U4996 ( .A1(n4460), .A2(n4696), .ZN(U3298) );
  INV_X1 U4997 ( .A(D_REG_23__SCAN_IN), .ZN(n4649) );
  NOR2_X1 U4998 ( .A1(n4460), .A2(n4649), .ZN(U3299) );
  AND2_X1 U4999 ( .A1(D_REG_22__SCAN_IN), .A2(n4459), .ZN(U3300) );
  INV_X1 U5000 ( .A(D_REG_21__SCAN_IN), .ZN(n4661) );
  NOR2_X1 U5001 ( .A1(n4460), .A2(n4661), .ZN(U3301) );
  AND2_X1 U5002 ( .A1(D_REG_20__SCAN_IN), .A2(n4459), .ZN(U3302) );
  AND2_X1 U5003 ( .A1(D_REG_19__SCAN_IN), .A2(n4459), .ZN(U3303) );
  INV_X1 U5004 ( .A(D_REG_18__SCAN_IN), .ZN(n4669) );
  NOR2_X1 U5005 ( .A1(n4460), .A2(n4669), .ZN(U3304) );
  NOR2_X1 U5006 ( .A1(n4460), .A2(n4727), .ZN(U3305) );
  AND2_X1 U5007 ( .A1(D_REG_16__SCAN_IN), .A2(n4459), .ZN(U3306) );
  AND2_X1 U5008 ( .A1(D_REG_15__SCAN_IN), .A2(n4459), .ZN(U3307) );
  AND2_X1 U5009 ( .A1(D_REG_14__SCAN_IN), .A2(n4459), .ZN(U3308) );
  INV_X1 U5010 ( .A(D_REG_13__SCAN_IN), .ZN(n4684) );
  NOR2_X1 U5011 ( .A1(n4460), .A2(n4684), .ZN(U3309) );
  INV_X1 U5012 ( .A(D_REG_12__SCAN_IN), .ZN(n4694) );
  NOR2_X1 U5013 ( .A1(n4460), .A2(n4694), .ZN(U3310) );
  AND2_X1 U5014 ( .A1(D_REG_11__SCAN_IN), .A2(n4459), .ZN(U3311) );
  AND2_X1 U5015 ( .A1(D_REG_10__SCAN_IN), .A2(n4459), .ZN(U3312) );
  AND2_X1 U5016 ( .A1(D_REG_9__SCAN_IN), .A2(n4459), .ZN(U3313) );
  NOR2_X1 U5017 ( .A1(n4460), .A2(n4712), .ZN(U3314) );
  NOR2_X1 U5018 ( .A1(n4460), .A2(n4698), .ZN(U3315) );
  AND2_X1 U5019 ( .A1(D_REG_6__SCAN_IN), .A2(n4459), .ZN(U3316) );
  INV_X1 U5020 ( .A(D_REG_5__SCAN_IN), .ZN(n4681) );
  NOR2_X1 U5021 ( .A1(n4460), .A2(n4681), .ZN(U3317) );
  NOR2_X1 U5022 ( .A1(n4460), .A2(n4711), .ZN(U3318) );
  AND2_X1 U5023 ( .A1(D_REG_3__SCAN_IN), .A2(n4459), .ZN(U3319) );
  INV_X1 U5024 ( .A(D_REG_2__SCAN_IN), .ZN(n4672) );
  NOR2_X1 U5025 ( .A1(n4460), .A2(n4672), .ZN(U3320) );
  INV_X1 U5026 ( .A(DATAI_23_), .ZN(n4668) );
  AOI21_X1 U5027 ( .B1(U3149), .B2(n4668), .A(n4461), .ZN(U3329) );
  INV_X1 U5028 ( .A(DATAI_18_), .ZN(n4645) );
  AOI22_X1 U5029 ( .A1(STATE_REG_SCAN_IN), .A2(n4462), .B1(n4645), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5030 ( .A1(STATE_REG_SCAN_IN), .A2(n4463), .B1(n2684), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5031 ( .A(DATAI_16_), .ZN(n4464) );
  AOI22_X1 U5032 ( .A1(STATE_REG_SCAN_IN), .A2(n4465), .B1(n4464), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5033 ( .A(DATAI_15_), .ZN(n4466) );
  AOI22_X1 U5034 ( .A1(STATE_REG_SCAN_IN), .A2(n4467), .B1(n4466), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5035 ( .A(DATAI_14_), .ZN(n4724) );
  AOI22_X1 U5036 ( .A1(STATE_REG_SCAN_IN), .A2(n2223), .B1(n4724), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5037 ( .A1(STATE_REG_SCAN_IN), .A2(n4468), .B1(n2610), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5038 ( .A(DATAI_12_), .ZN(n4660) );
  AOI22_X1 U5039 ( .A1(STATE_REG_SCAN_IN), .A2(n4469), .B1(n4660), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5040 ( .A(DATAI_11_), .ZN(n4470) );
  AOI22_X1 U5041 ( .A1(STATE_REG_SCAN_IN), .A2(n4471), .B1(n4470), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5042 ( .A(DATAI_10_), .ZN(n4472) );
  AOI22_X1 U5043 ( .A1(STATE_REG_SCAN_IN), .A2(n2262), .B1(n4472), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5044 ( .A(DATAI_9_), .ZN(n4474) );
  AOI22_X1 U5045 ( .A1(STATE_REG_SCAN_IN), .A2(n4475), .B1(n4474), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5046 ( .A(DATAI_0_), .ZN(n4476) );
  AOI22_X1 U5047 ( .A1(STATE_REG_SCAN_IN), .A2(n4830), .B1(n4476), .B2(U3149), 
        .ZN(U3352) );
  AOI22_X1 U5048 ( .A1(n4520), .A2(n4477), .B1(n2353), .B2(n4518), .ZN(U3467)
         );
  INV_X1 U5049 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4728) );
  AOI22_X1 U5050 ( .A1(n4520), .A2(n4478), .B1(n4728), .B2(n4518), .ZN(U3469)
         );
  OAI22_X1 U5051 ( .A1(n4481), .A2(n4480), .B1(n4512), .B2(n4479), .ZN(n4482)
         );
  NOR2_X1 U5052 ( .A1(n4483), .A2(n4482), .ZN(n4522) );
  INV_X1 U5053 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4484) );
  AOI22_X1 U5054 ( .A1(n4520), .A2(n4522), .B1(n4484), .B2(n4518), .ZN(U3473)
         );
  INV_X1 U5055 ( .A(n4485), .ZN(n4486) );
  AOI211_X1 U5056 ( .C1(n4488), .C2(n4517), .A(n4487), .B(n4486), .ZN(n4523)
         );
  INV_X1 U5057 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4489) );
  AOI22_X1 U5058 ( .A1(n4520), .A2(n4523), .B1(n4489), .B2(n4518), .ZN(U3475)
         );
  NOR2_X1 U5059 ( .A1(n4490), .A2(n4501), .ZN(n4493) );
  INV_X1 U5060 ( .A(n4491), .ZN(n4492) );
  AOI211_X1 U5061 ( .C1(n4506), .C2(n4494), .A(n4493), .B(n4492), .ZN(n4524)
         );
  INV_X1 U5062 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4495) );
  AOI22_X1 U5063 ( .A1(n4520), .A2(n4524), .B1(n4495), .B2(n4518), .ZN(U3477)
         );
  NAND3_X1 U5064 ( .A1(n3316), .A2(n4497), .A3(n4496), .ZN(n4498) );
  AND3_X1 U5065 ( .A1(n4500), .A2(n4499), .A3(n4498), .ZN(n4526) );
  INV_X1 U5066 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4685) );
  AOI22_X1 U5067 ( .A1(n4520), .A2(n4526), .B1(n4685), .B2(n4518), .ZN(U3481)
         );
  NOR2_X1 U5068 ( .A1(n4502), .A2(n4501), .ZN(n4504) );
  AOI211_X1 U5069 ( .C1(n4506), .C2(n4505), .A(n4504), .B(n4503), .ZN(n4528)
         );
  INV_X1 U5070 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4683) );
  AOI22_X1 U5071 ( .A1(n4520), .A2(n4528), .B1(n4683), .B2(n4518), .ZN(U3485)
         );
  NOR3_X1 U5072 ( .A1(n4508), .A2(n4507), .A3(n4512), .ZN(n4510) );
  AOI211_X1 U5073 ( .C1(n4517), .C2(n4511), .A(n4510), .B(n4509), .ZN(n4529)
         );
  INV_X1 U5074 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4786) );
  AOI22_X1 U5075 ( .A1(n4520), .A2(n4529), .B1(n4786), .B2(n4518), .ZN(U3487)
         );
  NOR2_X1 U5076 ( .A1(n4513), .A2(n4512), .ZN(n4515) );
  AOI211_X1 U5077 ( .C1(n4517), .C2(n4516), .A(n4515), .B(n4514), .ZN(n4532)
         );
  INV_X1 U5078 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4519) );
  AOI22_X1 U5079 ( .A1(n4520), .A2(n4532), .B1(n4519), .B2(n4518), .ZN(U3489)
         );
  INV_X1 U5080 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4521) );
  AOI22_X1 U5081 ( .A1(n4533), .A2(n4522), .B1(n4521), .B2(n4530), .ZN(U3521)
         );
  AOI22_X1 U5082 ( .A1(n4533), .A2(n4523), .B1(n3015), .B2(n4530), .ZN(U3522)
         );
  AOI22_X1 U5083 ( .A1(n4533), .A2(n4524), .B1(n3019), .B2(n4530), .ZN(U3523)
         );
  AOI22_X1 U5084 ( .A1(n4533), .A2(n4526), .B1(n4525), .B2(n4530), .ZN(U3525)
         );
  AOI22_X1 U5085 ( .A1(n4533), .A2(n4528), .B1(n4527), .B2(n4530), .ZN(U3527)
         );
  AOI22_X1 U5086 ( .A1(n4533), .A2(n4529), .B1(n4788), .B2(n4530), .ZN(U3528)
         );
  AOI22_X1 U5087 ( .A1(n4533), .A2(n4532), .B1(n4531), .B2(n4530), .ZN(U3529)
         );
  INV_X1 U5088 ( .A(n4534), .ZN(n4536) );
  NOR2_X1 U5089 ( .A1(n4536), .A2(n4535), .ZN(n4537) );
  XNOR2_X1 U5090 ( .A(n4538), .B(n4537), .ZN(n4552) );
  AOI22_X1 U5091 ( .A1(n4542), .A2(n4541), .B1(n4540), .B2(n4539), .ZN(n4550)
         );
  NOR2_X1 U5092 ( .A1(n4544), .A2(n4543), .ZN(n4545) );
  AOI211_X1 U5093 ( .C1(n4548), .C2(n4547), .A(n4546), .B(n4545), .ZN(n4549)
         );
  OAI211_X1 U5094 ( .C1(n4552), .C2(n4551), .A(n4550), .B(n4549), .ZN(n4870)
         );
  INV_X1 U5095 ( .A(keyinput71), .ZN(n4553) );
  NOR4_X1 U5096 ( .A1(keyinput98), .A2(keyinput92), .A3(keyinput23), .A4(n4553), .ZN(n4554) );
  NAND3_X1 U5097 ( .A1(keyinput99), .A2(keyinput26), .A3(n4554), .ZN(n4566) );
  NOR2_X1 U5098 ( .A1(keyinput25), .A2(keyinput120), .ZN(n4555) );
  NAND3_X1 U5099 ( .A1(keyinput116), .A2(keyinput51), .A3(n4555), .ZN(n4556)
         );
  NOR3_X1 U5100 ( .A1(keyinput27), .A2(keyinput8), .A3(n4556), .ZN(n4564) );
  INV_X1 U5101 ( .A(keyinput66), .ZN(n4557) );
  NAND4_X1 U5102 ( .A1(keyinput37), .A2(keyinput85), .A3(keyinput123), .A4(
        n4557), .ZN(n4562) );
  NAND3_X1 U5103 ( .A1(keyinput126), .A2(keyinput64), .A3(keyinput32), .ZN(
        n4561) );
  NOR2_X1 U5104 ( .A1(keyinput18), .A2(keyinput56), .ZN(n4558) );
  NAND3_X1 U5105 ( .A1(keyinput17), .A2(keyinput79), .A3(n4558), .ZN(n4560) );
  NAND4_X1 U5106 ( .A1(keyinput59), .A2(keyinput106), .A3(keyinput60), .A4(
        keyinput103), .ZN(n4559) );
  NOR4_X1 U5107 ( .A1(n4562), .A2(n4561), .A3(n4560), .A4(n4559), .ZN(n4563)
         );
  NAND4_X1 U5108 ( .A1(keyinput114), .A2(keyinput29), .A3(n4564), .A4(n4563), 
        .ZN(n4565) );
  NOR4_X1 U5109 ( .A1(keyinput93), .A2(keyinput21), .A3(n4566), .A4(n4565), 
        .ZN(n4613) );
  NAND2_X1 U5110 ( .A1(keyinput57), .A2(keyinput95), .ZN(n4567) );
  NOR3_X1 U5111 ( .A1(keyinput70), .A2(keyinput118), .A3(n4567), .ZN(n4568) );
  NAND3_X1 U5112 ( .A1(keyinput33), .A2(keyinput9), .A3(n4568), .ZN(n4581) );
  INV_X1 U5113 ( .A(keyinput24), .ZN(n4756) );
  INV_X1 U5114 ( .A(keyinput30), .ZN(n4762) );
  INV_X1 U5115 ( .A(keyinput19), .ZN(n4759) );
  OR4_X1 U5116 ( .A1(n4756), .A2(n4762), .A3(n4759), .A4(keyinput81), .ZN(
        n4569) );
  NOR3_X1 U5117 ( .A1(keyinput125), .A2(keyinput5), .A3(n4569), .ZN(n4579) );
  NOR2_X1 U5118 ( .A1(keyinput45), .A2(keyinput73), .ZN(n4570) );
  NAND3_X1 U5119 ( .A1(keyinput22), .A2(keyinput11), .A3(n4570), .ZN(n4577) );
  NOR2_X1 U5120 ( .A1(keyinput7), .A2(keyinput104), .ZN(n4571) );
  NAND3_X1 U5121 ( .A1(keyinput117), .A2(keyinput14), .A3(n4571), .ZN(n4576)
         );
  NOR3_X1 U5122 ( .A1(keyinput2), .A2(keyinput44), .A3(keyinput38), .ZN(n4572)
         );
  NAND2_X1 U5123 ( .A1(keyinput15), .A2(n4572), .ZN(n4575) );
  INV_X1 U5124 ( .A(keyinput107), .ZN(n4573) );
  NAND4_X1 U5125 ( .A1(keyinput50), .A2(keyinput28), .A3(keyinput48), .A4(
        n4573), .ZN(n4574) );
  NOR4_X1 U5126 ( .A1(n4577), .A2(n4576), .A3(n4575), .A4(n4574), .ZN(n4578)
         );
  NAND4_X1 U5127 ( .A1(keyinput76), .A2(keyinput55), .A3(n4579), .A4(n4578), 
        .ZN(n4580) );
  NOR4_X1 U5128 ( .A1(keyinput61), .A2(keyinput52), .A3(n4581), .A4(n4580), 
        .ZN(n4612) );
  INV_X1 U5129 ( .A(keyinput77), .ZN(n4582) );
  NAND4_X1 U5130 ( .A1(keyinput41), .A2(keyinput100), .A3(keyinput83), .A4(
        n4582), .ZN(n4596) );
  NAND4_X1 U5131 ( .A1(keyinput119), .A2(keyinput112), .A3(keyinput115), .A4(
        keyinput89), .ZN(n4595) );
  INV_X1 U5132 ( .A(keyinput97), .ZN(n4583) );
  NOR2_X1 U5133 ( .A1(keyinput113), .A2(n4583), .ZN(n4585) );
  NOR4_X1 U5134 ( .A1(keyinput101), .A2(keyinput105), .A3(keyinput13), .A4(
        keyinput1), .ZN(n4584) );
  NAND4_X1 U5135 ( .A1(keyinput65), .A2(keyinput69), .A3(n4585), .A4(n4584), 
        .ZN(n4594) );
  NAND2_X1 U5136 ( .A1(keyinput109), .A2(keyinput102), .ZN(n4586) );
  NOR3_X1 U5137 ( .A1(keyinput43), .A2(keyinput47), .A3(n4586), .ZN(n4592) );
  INV_X1 U5138 ( .A(keyinput34), .ZN(n4587) );
  NOR4_X1 U5139 ( .A1(keyinput121), .A2(keyinput96), .A3(keyinput54), .A4(
        n4587), .ZN(n4591) );
  NOR4_X1 U5140 ( .A1(keyinput88), .A2(keyinput80), .A3(keyinput108), .A4(
        keyinput72), .ZN(n4590) );
  NAND3_X1 U5141 ( .A1(keyinput0), .A2(keyinput84), .A3(keyinput49), .ZN(n4588) );
  NOR2_X1 U5142 ( .A1(keyinput53), .A2(n4588), .ZN(n4589) );
  NAND4_X1 U5143 ( .A1(n4592), .A2(n4591), .A3(n4590), .A4(n4589), .ZN(n4593)
         );
  NOR4_X1 U5144 ( .A1(n4596), .A2(n4595), .A3(n4594), .A4(n4593), .ZN(n4611)
         );
  NOR2_X1 U5145 ( .A1(keyinput36), .A2(keyinput68), .ZN(n4597) );
  NAND3_X1 U5146 ( .A1(keyinput4), .A2(keyinput40), .A3(n4597), .ZN(n4609) );
  NAND4_X1 U5147 ( .A1(keyinput124), .A2(keyinput16), .A3(keyinput12), .A4(
        keyinput20), .ZN(n4608) );
  NOR2_X1 U5148 ( .A1(keyinput87), .A2(keyinput86), .ZN(n4599) );
  NOR4_X1 U5149 ( .A1(keyinput91), .A2(keyinput90), .A3(keyinput94), .A4(
        keyinput111), .ZN(n4598) );
  NAND4_X1 U5150 ( .A1(n4599), .A2(keyinput110), .A3(keyinput122), .A4(n4598), 
        .ZN(n4607) );
  NAND3_X1 U5151 ( .A1(keyinput46), .A2(keyinput42), .A3(keyinput10), .ZN(
        n4600) );
  NOR2_X1 U5152 ( .A1(keyinput31), .A2(n4600), .ZN(n4605) );
  NOR4_X1 U5153 ( .A1(keyinput3), .A2(keyinput6), .A3(keyinput35), .A4(
        keyinput39), .ZN(n4604) );
  NAND2_X1 U5154 ( .A1(keyinput75), .A2(keyinput62), .ZN(n4601) );
  NOR3_X1 U5155 ( .A1(keyinput74), .A2(keyinput67), .A3(n4601), .ZN(n4603) );
  NOR4_X1 U5156 ( .A1(keyinput58), .A2(keyinput63), .A3(keyinput78), .A4(
        keyinput82), .ZN(n4602) );
  NAND4_X1 U5157 ( .A1(n4605), .A2(n4604), .A3(n4603), .A4(n4602), .ZN(n4606)
         );
  NOR4_X1 U5158 ( .A1(n4609), .A2(n4608), .A3(n4607), .A4(n4606), .ZN(n4610)
         );
  NAND4_X1 U5159 ( .A1(n4613), .A2(n4612), .A3(n4611), .A4(n4610), .ZN(n4867)
         );
  AOI22_X1 U5160 ( .A1(n4615), .A2(keyinput112), .B1(keyinput115), .B2(n4052), 
        .ZN(n4614) );
  OAI221_X1 U5161 ( .B1(n4615), .B2(keyinput112), .C1(n4052), .C2(keyinput115), 
        .A(n4614), .ZN(n4628) );
  INV_X1 U5162 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4618) );
  INV_X1 U5163 ( .A(keyinput89), .ZN(n4617) );
  AOI22_X1 U5164 ( .A1(n4618), .A2(keyinput100), .B1(DATAO_REG_22__SCAN_IN), 
        .B2(n4617), .ZN(n4616) );
  OAI221_X1 U5165 ( .B1(n4618), .B2(keyinput100), .C1(n4617), .C2(
        DATAO_REG_22__SCAN_IN), .A(n4616), .ZN(n4627) );
  INV_X1 U5166 ( .A(keyinput41), .ZN(n4620) );
  AOI22_X1 U5167 ( .A1(n4621), .A2(keyinput77), .B1(DATAO_REG_24__SCAN_IN), 
        .B2(n4620), .ZN(n4619) );
  OAI221_X1 U5168 ( .B1(n4621), .B2(keyinput77), .C1(n4620), .C2(
        DATAO_REG_24__SCAN_IN), .A(n4619), .ZN(n4626) );
  INV_X1 U5169 ( .A(keyinput121), .ZN(n4623) );
  AOI22_X1 U5170 ( .A1(n4624), .A2(keyinput83), .B1(DATAO_REG_25__SCAN_IN), 
        .B2(n4623), .ZN(n4622) );
  OAI221_X1 U5171 ( .B1(n4624), .B2(keyinput83), .C1(n4623), .C2(
        DATAO_REG_25__SCAN_IN), .A(n4622), .ZN(n4625) );
  NOR4_X1 U5172 ( .A1(n4628), .A2(n4627), .A3(n4626), .A4(n4625), .ZN(n4679)
         );
  AOI22_X1 U5173 ( .A1(n4631), .A2(keyinput96), .B1(n4630), .B2(keyinput34), 
        .ZN(n4629) );
  OAI221_X1 U5174 ( .B1(n4631), .B2(keyinput96), .C1(n4630), .C2(keyinput34), 
        .A(n4629), .ZN(n4643) );
  INV_X1 U5175 ( .A(REG1_REG_29__SCAN_IN), .ZN(n4634) );
  INV_X1 U5176 ( .A(keyinput54), .ZN(n4633) );
  AOI22_X1 U5177 ( .A1(n4634), .A2(keyinput102), .B1(DATAO_REG_29__SCAN_IN), 
        .B2(n4633), .ZN(n4632) );
  OAI221_X1 U5178 ( .B1(n4634), .B2(keyinput102), .C1(n4633), .C2(
        DATAO_REG_29__SCAN_IN), .A(n4632), .ZN(n4642) );
  AOI22_X1 U5179 ( .A1(n4637), .A2(keyinput47), .B1(keyinput43), .B2(n4636), 
        .ZN(n4635) );
  OAI221_X1 U5180 ( .B1(n4637), .B2(keyinput47), .C1(n4636), .C2(keyinput43), 
        .A(n4635), .ZN(n4641) );
  AOI22_X1 U5181 ( .A1(n3786), .A2(keyinput109), .B1(n4639), .B2(keyinput65), 
        .ZN(n4638) );
  OAI221_X1 U5182 ( .B1(n3786), .B2(keyinput109), .C1(n4639), .C2(keyinput65), 
        .A(n4638), .ZN(n4640) );
  NOR4_X1 U5183 ( .A1(n4643), .A2(n4642), .A3(n4641), .A4(n4640), .ZN(n4678)
         );
  INV_X1 U5184 ( .A(DATAI_20_), .ZN(n4646) );
  AOI22_X1 U5185 ( .A1(n4646), .A2(keyinput105), .B1(keyinput13), .B2(n4645), 
        .ZN(n4644) );
  OAI221_X1 U5186 ( .B1(n4646), .B2(keyinput105), .C1(n4645), .C2(keyinput13), 
        .A(n4644), .ZN(n4658) );
  AOI22_X1 U5187 ( .A1(n4649), .A2(keyinput97), .B1(keyinput101), .B2(n4648), 
        .ZN(n4647) );
  OAI221_X1 U5188 ( .B1(n4649), .B2(keyinput97), .C1(n4648), .C2(keyinput101), 
        .A(n4647), .ZN(n4657) );
  INV_X1 U5189 ( .A(DATAI_6_), .ZN(n4651) );
  AOI22_X1 U5190 ( .A1(n4652), .A2(keyinput69), .B1(keyinput113), .B2(n4651), 
        .ZN(n4650) );
  OAI221_X1 U5191 ( .B1(n4652), .B2(keyinput69), .C1(n4651), .C2(keyinput113), 
        .A(n4650), .ZN(n4656) );
  XNOR2_X1 U5192 ( .A(IR_REG_22__SCAN_IN), .B(keyinput1), .ZN(n4654) );
  XNOR2_X1 U5193 ( .A(keyinput49), .B(DATAI_5_), .ZN(n4653) );
  NAND2_X1 U5194 ( .A1(n4654), .A2(n4653), .ZN(n4655) );
  NOR4_X1 U5195 ( .A1(n4658), .A2(n4657), .A3(n4656), .A4(n4655), .ZN(n4677)
         );
  AOI22_X1 U5196 ( .A1(n4661), .A2(keyinput72), .B1(keyinput84), .B2(n4660), 
        .ZN(n4659) );
  OAI221_X1 U5197 ( .B1(n4661), .B2(keyinput72), .C1(n4660), .C2(keyinput84), 
        .A(n4659), .ZN(n4666) );
  XNOR2_X1 U5198 ( .A(n4662), .B(keyinput108), .ZN(n4665) );
  XNOR2_X1 U5199 ( .A(n4663), .B(keyinput80), .ZN(n4664) );
  OR3_X1 U5200 ( .A1(n4666), .A2(n4665), .A3(n4664), .ZN(n4675) );
  AOI22_X1 U5201 ( .A1(n4669), .A2(keyinput0), .B1(keyinput124), .B2(n4668), 
        .ZN(n4667) );
  OAI221_X1 U5202 ( .B1(n4669), .B2(keyinput0), .C1(n4668), .C2(keyinput124), 
        .A(n4667), .ZN(n4674) );
  INV_X1 U5203 ( .A(DATAI_26_), .ZN(n4671) );
  AOI22_X1 U5204 ( .A1(n4672), .A2(keyinput53), .B1(keyinput88), .B2(n4671), 
        .ZN(n4670) );
  OAI221_X1 U5205 ( .B1(n4672), .B2(keyinput53), .C1(n4671), .C2(keyinput88), 
        .A(n4670), .ZN(n4673) );
  NOR3_X1 U5206 ( .A1(n4675), .A2(n4674), .A3(n4673), .ZN(n4676) );
  NAND4_X1 U5207 ( .A1(n4679), .A2(n4678), .A3(n4677), .A4(n4676), .ZN(n4865)
         );
  AOI22_X1 U5208 ( .A1(n2538), .A2(keyinput40), .B1(keyinput3), .B2(n4681), 
        .ZN(n4680) );
  OAI221_X1 U5209 ( .B1(n2538), .B2(keyinput40), .C1(n4681), .C2(keyinput3), 
        .A(n4680), .ZN(n4692) );
  AOI22_X1 U5210 ( .A1(n4684), .A2(keyinput16), .B1(keyinput36), .B2(n4683), 
        .ZN(n4682) );
  OAI221_X1 U5211 ( .B1(n4684), .B2(keyinput16), .C1(n4683), .C2(keyinput36), 
        .A(n4682), .ZN(n4691) );
  XOR2_X1 U5212 ( .A(n4685), .B(keyinput4), .Z(n4689) );
  XOR2_X1 U5213 ( .A(n2367), .B(keyinput68), .Z(n4688) );
  XNOR2_X1 U5214 ( .A(IR_REG_10__SCAN_IN), .B(keyinput12), .ZN(n4687) );
  XNOR2_X1 U5215 ( .A(IR_REG_24__SCAN_IN), .B(keyinput20), .ZN(n4686) );
  NAND4_X1 U5216 ( .A1(n4689), .A2(n4688), .A3(n4687), .A4(n4686), .ZN(n4690)
         );
  NOR3_X1 U5217 ( .A1(n4692), .A2(n4691), .A3(n4690), .ZN(n4740) );
  INV_X1 U5218 ( .A(keyinput42), .ZN(n4693) );
  XNOR2_X1 U5219 ( .A(n4694), .B(n4693), .ZN(n4709) );
  INV_X1 U5220 ( .A(keyinput10), .ZN(n4695) );
  XNOR2_X1 U5221 ( .A(n4696), .B(n4695), .ZN(n4708) );
  INV_X1 U5222 ( .A(keyinput58), .ZN(n4697) );
  XNOR2_X1 U5223 ( .A(n4698), .B(n4697), .ZN(n4707) );
  XNOR2_X1 U5224 ( .A(IR_REG_13__SCAN_IN), .B(keyinput35), .ZN(n4701) );
  XNOR2_X1 U5225 ( .A(DATAI_4_), .B(keyinput6), .ZN(n4700) );
  XNOR2_X1 U5226 ( .A(keyinput31), .B(REG0_REG_6__SCAN_IN), .ZN(n4699) );
  NAND3_X1 U5227 ( .A1(n4701), .A2(n4700), .A3(n4699), .ZN(n4705) );
  XNOR2_X1 U5228 ( .A(IR_REG_28__SCAN_IN), .B(keyinput46), .ZN(n4703) );
  XNOR2_X1 U5229 ( .A(IR_REG_5__SCAN_IN), .B(keyinput39), .ZN(n4702) );
  NAND2_X1 U5230 ( .A1(n4703), .A2(n4702), .ZN(n4704) );
  NOR2_X1 U5231 ( .A1(n4705), .A2(n4704), .ZN(n4706) );
  AND4_X1 U5232 ( .A1(n4709), .A2(n4708), .A3(n4707), .A4(n4706), .ZN(n4739)
         );
  AOI22_X1 U5233 ( .A1(n4712), .A2(keyinput67), .B1(n4711), .B2(keyinput74), 
        .ZN(n4710) );
  OAI221_X1 U5234 ( .B1(n4712), .B2(keyinput67), .C1(n4711), .C2(keyinput74), 
        .A(n4710), .ZN(n4722) );
  XNOR2_X1 U5235 ( .A(n4713), .B(keyinput82), .ZN(n4721) );
  XNOR2_X1 U5236 ( .A(keyinput63), .B(n4714), .ZN(n4720) );
  XNOR2_X1 U5237 ( .A(IR_REG_8__SCAN_IN), .B(keyinput78), .ZN(n4718) );
  XNOR2_X1 U5238 ( .A(IR_REG_18__SCAN_IN), .B(keyinput62), .ZN(n4717) );
  XNOR2_X1 U5239 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput87), .ZN(n4716) );
  XNOR2_X1 U5240 ( .A(IR_REG_23__SCAN_IN), .B(keyinput75), .ZN(n4715) );
  NAND4_X1 U5241 ( .A1(n4718), .A2(n4717), .A3(n4716), .A4(n4715), .ZN(n4719)
         );
  NOR4_X1 U5242 ( .A1(n4722), .A2(n4721), .A3(n4720), .A4(n4719), .ZN(n4738)
         );
  AOI22_X1 U5243 ( .A1(n4724), .A2(keyinput111), .B1(keyinput110), .B2(n2521), 
        .ZN(n4723) );
  OAI221_X1 U5244 ( .B1(n4724), .B2(keyinput111), .C1(n2521), .C2(keyinput110), 
        .A(n4723), .ZN(n4736) );
  INV_X1 U5245 ( .A(DATAI_21_), .ZN(n4726) );
  AOI22_X1 U5246 ( .A1(n4727), .A2(keyinput90), .B1(keyinput94), .B2(n4726), 
        .ZN(n4725) );
  OAI221_X1 U5247 ( .B1(n4727), .B2(keyinput90), .C1(n4726), .C2(keyinput94), 
        .A(n4725), .ZN(n4735) );
  XOR2_X1 U5248 ( .A(n4728), .B(keyinput91), .Z(n4733) );
  XOR2_X1 U5249 ( .A(n4729), .B(keyinput122), .Z(n4732) );
  XNOR2_X1 U5250 ( .A(IR_REG_21__SCAN_IN), .B(keyinput86), .ZN(n4731) );
  XNOR2_X1 U5251 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput126), .ZN(n4730) );
  NAND4_X1 U5252 ( .A1(n4733), .A2(n4732), .A3(n4731), .A4(n4730), .ZN(n4734)
         );
  NOR3_X1 U5253 ( .A1(n4736), .A2(n4735), .A3(n4734), .ZN(n4737) );
  NAND4_X1 U5254 ( .A1(n4740), .A2(n4739), .A3(n4738), .A4(n4737), .ZN(n4864)
         );
  AOI22_X1 U5255 ( .A1(n3025), .A2(keyinput104), .B1(n3368), .B2(keyinput45), 
        .ZN(n4741) );
  OAI221_X1 U5256 ( .B1(n3025), .B2(keyinput104), .C1(n3368), .C2(keyinput45), 
        .A(n4741), .ZN(n4752) );
  AOI22_X1 U5257 ( .A1(n2999), .A2(keyinput73), .B1(keyinput70), .B2(n4743), 
        .ZN(n4742) );
  OAI221_X1 U5258 ( .B1(n2999), .B2(keyinput73), .C1(n4743), .C2(keyinput70), 
        .A(n4742), .ZN(n4751) );
  XOR2_X1 U5259 ( .A(n4744), .B(keyinput14), .Z(n4749) );
  XOR2_X1 U5260 ( .A(n4745), .B(keyinput22), .Z(n4748) );
  XNOR2_X1 U5261 ( .A(REG1_REG_1__SCAN_IN), .B(keyinput117), .ZN(n4747) );
  XNOR2_X1 U5262 ( .A(IR_REG_27__SCAN_IN), .B(keyinput11), .ZN(n4746) );
  NAND4_X1 U5263 ( .A1(n4749), .A2(n4748), .A3(n4747), .A4(n4746), .ZN(n4750)
         );
  NOR3_X1 U5264 ( .A1(n4752), .A2(n4751), .A3(n4750), .ZN(n4802) );
  INV_X1 U5265 ( .A(keyinput125), .ZN(n4754) );
  AOI22_X1 U5266 ( .A1(n2215), .A2(keyinput81), .B1(ADDR_REG_9__SCAN_IN), .B2(
        n4754), .ZN(n4753) );
  OAI221_X1 U5267 ( .B1(n2215), .B2(keyinput81), .C1(n4754), .C2(
        ADDR_REG_9__SCAN_IN), .A(n4753), .ZN(n4767) );
  INV_X1 U5268 ( .A(REG2_REG_4__SCAN_IN), .ZN(n4757) );
  AOI22_X1 U5269 ( .A1(n4757), .A2(keyinput55), .B1(ADDR_REG_5__SCAN_IN), .B2(
        n4756), .ZN(n4755) );
  OAI221_X1 U5270 ( .B1(n4757), .B2(keyinput55), .C1(n4756), .C2(
        ADDR_REG_5__SCAN_IN), .A(n4755), .ZN(n4766) );
  INV_X1 U5271 ( .A(ADDR_REG_17__SCAN_IN), .ZN(n4760) );
  AOI22_X1 U5272 ( .A1(n4760), .A2(keyinput7), .B1(ADDR_REG_16__SCAN_IN), .B2(
        n4759), .ZN(n4758) );
  OAI221_X1 U5273 ( .B1(n4760), .B2(keyinput7), .C1(n4759), .C2(
        ADDR_REG_16__SCAN_IN), .A(n4758), .ZN(n4765) );
  INV_X1 U5274 ( .A(keyinput5), .ZN(n4763) );
  AOI22_X1 U5275 ( .A1(n4763), .A2(ADDR_REG_13__SCAN_IN), .B1(
        ADDR_REG_15__SCAN_IN), .B2(n4762), .ZN(n4761) );
  OAI221_X1 U5276 ( .B1(n4763), .B2(ADDR_REG_13__SCAN_IN), .C1(n4762), .C2(
        ADDR_REG_15__SCAN_IN), .A(n4761), .ZN(n4764) );
  NOR4_X1 U5277 ( .A1(n4767), .A2(n4766), .A3(n4765), .A4(n4764), .ZN(n4801)
         );
  INV_X1 U5278 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4769) );
  AOI22_X1 U5279 ( .A1(n4770), .A2(keyinput15), .B1(n4769), .B2(keyinput28), 
        .ZN(n4768) );
  OAI221_X1 U5280 ( .B1(n4770), .B2(keyinput15), .C1(n4769), .C2(keyinput28), 
        .A(n4768), .ZN(n4783) );
  INV_X1 U5281 ( .A(keyinput2), .ZN(n4772) );
  AOI22_X1 U5282 ( .A1(n4773), .A2(keyinput107), .B1(DATAO_REG_19__SCAN_IN), 
        .B2(n4772), .ZN(n4771) );
  OAI221_X1 U5283 ( .B1(n4773), .B2(keyinput107), .C1(n4772), .C2(
        DATAO_REG_19__SCAN_IN), .A(n4771), .ZN(n4782) );
  INV_X1 U5284 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4776) );
  AOI22_X1 U5285 ( .A1(n4776), .A2(keyinput44), .B1(n4775), .B2(keyinput119), 
        .ZN(n4774) );
  OAI221_X1 U5286 ( .B1(n4776), .B2(keyinput44), .C1(n4775), .C2(keyinput119), 
        .A(n4774), .ZN(n4781) );
  INV_X1 U5287 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4779) );
  INV_X1 U5288 ( .A(keyinput48), .ZN(n4778) );
  AOI22_X1 U5289 ( .A1(n4779), .A2(keyinput38), .B1(DATAO_REG_20__SCAN_IN), 
        .B2(n4778), .ZN(n4777) );
  OAI221_X1 U5290 ( .B1(n4779), .B2(keyinput38), .C1(n4778), .C2(
        DATAO_REG_20__SCAN_IN), .A(n4777), .ZN(n4780) );
  NOR4_X1 U5291 ( .A1(n4783), .A2(n4782), .A3(n4781), .A4(n4780), .ZN(n4800)
         );
  AOI22_X1 U5292 ( .A1(n4786), .A2(keyinput118), .B1(n4785), .B2(keyinput33), 
        .ZN(n4784) );
  OAI221_X1 U5293 ( .B1(n4786), .B2(keyinput118), .C1(n4785), .C2(keyinput33), 
        .A(n4784), .ZN(n4798) );
  INV_X1 U5294 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4789) );
  AOI22_X1 U5295 ( .A1(n4789), .A2(keyinput95), .B1(keyinput57), .B2(n4788), 
        .ZN(n4787) );
  OAI221_X1 U5296 ( .B1(n4789), .B2(keyinput95), .C1(n4788), .C2(keyinput57), 
        .A(n4787), .ZN(n4797) );
  INV_X1 U5297 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4791) );
  AOI22_X1 U5298 ( .A1(n4792), .A2(keyinput52), .B1(n4791), .B2(keyinput50), 
        .ZN(n4790) );
  OAI221_X1 U5299 ( .B1(n4792), .B2(keyinput52), .C1(n4791), .C2(keyinput50), 
        .A(n4790), .ZN(n4796) );
  AOI22_X1 U5300 ( .A1(n4794), .A2(keyinput9), .B1(n2586), .B2(keyinput61), 
        .ZN(n4793) );
  OAI221_X1 U5301 ( .B1(n4794), .B2(keyinput9), .C1(n2586), .C2(keyinput61), 
        .A(n4793), .ZN(n4795) );
  NOR4_X1 U5302 ( .A1(n4798), .A2(n4797), .A3(n4796), .A4(n4795), .ZN(n4799)
         );
  NAND4_X1 U5303 ( .A1(n4802), .A2(n4801), .A3(n4800), .A4(n4799), .ZN(n4863)
         );
  INV_X1 U5304 ( .A(keyinput120), .ZN(n4805) );
  INV_X1 U5305 ( .A(keyinput114), .ZN(n4804) );
  AOI22_X1 U5306 ( .A1(n4805), .A2(DATAO_REG_11__SCAN_IN), .B1(
        DATAO_REG_5__SCAN_IN), .B2(n4804), .ZN(n4803) );
  OAI221_X1 U5307 ( .B1(n4805), .B2(DATAO_REG_11__SCAN_IN), .C1(n4804), .C2(
        DATAO_REG_5__SCAN_IN), .A(n4803), .ZN(n4817) );
  INV_X1 U5308 ( .A(keyinput116), .ZN(n4807) );
  AOI22_X1 U5309 ( .A1(n3228), .A2(keyinput8), .B1(DATAO_REG_1__SCAN_IN), .B2(
        n4807), .ZN(n4806) );
  OAI221_X1 U5310 ( .B1(n3228), .B2(keyinput8), .C1(n4807), .C2(
        DATAO_REG_1__SCAN_IN), .A(n4806), .ZN(n4816) );
  INV_X1 U5311 ( .A(keyinput51), .ZN(n4810) );
  INV_X1 U5312 ( .A(keyinput93), .ZN(n4809) );
  AOI22_X1 U5313 ( .A1(n4810), .A2(DATAO_REG_9__SCAN_IN), .B1(
        DATAO_REG_15__SCAN_IN), .B2(n4809), .ZN(n4808) );
  OAI221_X1 U5314 ( .B1(n4810), .B2(DATAO_REG_9__SCAN_IN), .C1(n4809), .C2(
        DATAO_REG_15__SCAN_IN), .A(n4808), .ZN(n4815) );
  INV_X1 U5315 ( .A(keyinput29), .ZN(n4813) );
  INV_X1 U5316 ( .A(keyinput25), .ZN(n4812) );
  AOI22_X1 U5317 ( .A1(n4813), .A2(DATAO_REG_2__SCAN_IN), .B1(
        DATAO_REG_13__SCAN_IN), .B2(n4812), .ZN(n4811) );
  OAI221_X1 U5318 ( .B1(n4813), .B2(DATAO_REG_2__SCAN_IN), .C1(n4812), .C2(
        DATAO_REG_13__SCAN_IN), .A(n4811), .ZN(n4814) );
  NOR4_X1 U5319 ( .A1(n4817), .A2(n4816), .A3(n4815), .A4(n4814), .ZN(n4861)
         );
  AOI22_X1 U5320 ( .A1(keyinput66), .A2(n3633), .B1(keyinput127), .B2(n4868), 
        .ZN(n4818) );
  OAI21_X1 U5321 ( .B1(n3633), .B2(keyinput66), .A(n4818), .ZN(n4827) );
  AOI22_X1 U5322 ( .A1(n3919), .A2(keyinput64), .B1(keyinput32), .B2(n3938), 
        .ZN(n4819) );
  OAI221_X1 U5323 ( .B1(n3919), .B2(keyinput64), .C1(n3938), .C2(keyinput32), 
        .A(n4819), .ZN(n4826) );
  AOI22_X1 U5324 ( .A1(n4821), .A2(keyinput123), .B1(U3149), .B2(keyinput27), 
        .ZN(n4820) );
  OAI221_X1 U5325 ( .B1(n4821), .B2(keyinput123), .C1(U3149), .C2(keyinput27), 
        .A(n4820), .ZN(n4825) );
  INV_X1 U5326 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4823) );
  AOI22_X1 U5327 ( .A1(n4098), .A2(keyinput37), .B1(keyinput85), .B2(n4823), 
        .ZN(n4822) );
  OAI221_X1 U5328 ( .B1(n4098), .B2(keyinput37), .C1(n4823), .C2(keyinput85), 
        .A(n4822), .ZN(n4824) );
  NOR4_X1 U5329 ( .A1(n4827), .A2(n4826), .A3(n4825), .A4(n4824), .ZN(n4860)
         );
  INV_X1 U5330 ( .A(keyinput76), .ZN(n4829) );
  AOI22_X1 U5331 ( .A1(n4830), .A2(keyinput79), .B1(ADDR_REG_4__SCAN_IN), .B2(
        n4829), .ZN(n4828) );
  OAI221_X1 U5332 ( .B1(n4830), .B2(keyinput79), .C1(n4829), .C2(
        ADDR_REG_4__SCAN_IN), .A(n4828), .ZN(n4841) );
  INV_X1 U5333 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4833) );
  AOI22_X1 U5334 ( .A1(n4833), .A2(keyinput106), .B1(keyinput18), .B2(n4832), 
        .ZN(n4831) );
  OAI221_X1 U5335 ( .B1(n4833), .B2(keyinput106), .C1(n4832), .C2(keyinput18), 
        .A(n4831), .ZN(n4840) );
  INV_X1 U5336 ( .A(DATAI_30_), .ZN(n4835) );
  AOI22_X1 U5337 ( .A1(n4835), .A2(keyinput17), .B1(n2684), .B2(keyinput60), 
        .ZN(n4834) );
  OAI221_X1 U5338 ( .B1(n4835), .B2(keyinput17), .C1(n2684), .C2(keyinput60), 
        .A(n4834), .ZN(n4839) );
  XOR2_X1 U5339 ( .A(n3268), .B(keyinput103), .Z(n4837) );
  XNOR2_X1 U5340 ( .A(REG1_REG_0__SCAN_IN), .B(keyinput56), .ZN(n4836) );
  NAND2_X1 U5341 ( .A1(n4837), .A2(n4836), .ZN(n4838) );
  NOR4_X1 U5342 ( .A1(n4841), .A2(n4840), .A3(n4839), .A4(n4838), .ZN(n4859)
         );
  AOI22_X1 U5343 ( .A1(n4844), .A2(keyinput71), .B1(keyinput99), .B2(n4843), 
        .ZN(n4842) );
  OAI221_X1 U5344 ( .B1(n4844), .B2(keyinput71), .C1(n4843), .C2(keyinput99), 
        .A(n4842), .ZN(n4857) );
  INV_X1 U5345 ( .A(keyinput21), .ZN(n4846) );
  AOI22_X1 U5346 ( .A1(n4847), .A2(keyinput98), .B1(DATAO_REG_7__SCAN_IN), 
        .B2(n4846), .ZN(n4845) );
  OAI221_X1 U5347 ( .B1(n4847), .B2(keyinput98), .C1(n4846), .C2(
        DATAO_REG_7__SCAN_IN), .A(n4845), .ZN(n4856) );
  INV_X1 U5348 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4849) );
  AOI22_X1 U5349 ( .A1(n4850), .A2(keyinput23), .B1(keyinput59), .B2(n4849), 
        .ZN(n4848) );
  OAI221_X1 U5350 ( .B1(n4850), .B2(keyinput23), .C1(n4849), .C2(keyinput59), 
        .A(n4848), .ZN(n4855) );
  AOI22_X1 U5351 ( .A1(n4853), .A2(keyinput26), .B1(keyinput92), .B2(n4852), 
        .ZN(n4851) );
  OAI221_X1 U5352 ( .B1(n4853), .B2(keyinput26), .C1(n4852), .C2(keyinput92), 
        .A(n4851), .ZN(n4854) );
  NOR4_X1 U5353 ( .A1(n4857), .A2(n4856), .A3(n4855), .A4(n4854), .ZN(n4858)
         );
  NAND4_X1 U5354 ( .A1(n4861), .A2(n4860), .A3(n4859), .A4(n4858), .ZN(n4862)
         );
  NOR4_X1 U5355 ( .A1(n4865), .A2(n4864), .A3(n4863), .A4(n4862), .ZN(n4866)
         );
  OAI221_X1 U5356 ( .B1(n4868), .B2(keyinput127), .C1(n4868), .C2(n4867), .A(
        n4866), .ZN(n4869) );
  XNOR2_X1 U5357 ( .A(n4870), .B(n4869), .ZN(U3218) );
  CLKBUF_X2 U2404 ( .A(n2401), .Z(n3787) );
  CLKBUF_X1 U2426 ( .A(n3064), .Z(n2154) );
endmodule

