

module b21_C_AntiSAT_k_256_8 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, 
        keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, 
        keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, 
        keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, 
        keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, 
        keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, 
        keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, 
        keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, 
        keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, 
        keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, 
        keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, 
        keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, 
        keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, 
        keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, 
        keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, 
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, 
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, 
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, 
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, 
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, 
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, 
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, 
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, 
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, 
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249, 
        keyinput250, keyinput251, keyinput252, keyinput253, keyinput254, 
        keyinput255, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, 
        ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, 
        ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, 
        ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, 
        ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, 
        P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, 
        P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, 
        P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, 
        P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, 
        P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, 
        P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, 
        P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, 
        P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, 
        P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, 
        P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, 
        P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, 
        P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, 
        P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, 
        P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, 
        P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, 
        P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, 
        P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, 
        P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, 
        P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, 
        P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521;

  CLKBUF_X2 U4977 ( .A(n5268), .Z(n5852) );
  BUF_X2 U4978 ( .A(n6497), .Z(n4474) );
  NOR2_X1 U4979 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5951) );
  INV_X1 U4980 ( .A(n9089), .ZN(n5973) );
  NAND2_X1 U4981 ( .A1(n8587), .A2(n8622), .ZN(n6617) );
  INV_X1 U4982 ( .A(n10035), .ZN(n6028) );
  INV_X1 U4983 ( .A(n7257), .ZN(n5855) );
  NOR2_X1 U4984 ( .A1(n8812), .A2(n6606), .ZN(n8804) );
  NAND2_X1 U4985 ( .A1(n5919), .A2(n8345), .ZN(n5174) );
  INV_X1 U4986 ( .A(n7351), .ZN(n9945) );
  NAND2_X2 U4987 ( .A1(n6187), .A2(n6186), .ZN(n7616) );
  NAND2_X1 U4988 ( .A1(n6236), .A2(n6235), .ZN(n9051) );
  MUX2_X1 U4989 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5961), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5962) );
  OAI211_X1 U4990 ( .C1(n5622), .C2(n6635), .A(n5142), .B(n5141), .ZN(n7332)
         );
  INV_X1 U4991 ( .A(n5972), .ZN(n8640) );
  NAND2_X1 U4992 ( .A1(n7236), .A2(n8720), .ZN(n4472) );
  XNOR2_X2 U4993 ( .A(n6366), .B(n6367), .ZN(n8684) );
  OAI211_X2 U4994 ( .C1(n6097), .C2(n4978), .A(n4977), .B(n6126), .ZN(n7321)
         );
  NAND2_X1 U4995 ( .A1(n4983), .A2(n7075), .ZN(n4977) );
  XNOR2_X2 U4996 ( .A(n9934), .B(n7186), .ZN(n4867) );
  NAND4_X4 U4997 ( .A1(n5160), .A2(n5159), .A3(n5158), .A4(n5157), .ZN(n7186)
         );
  INV_X2 U4998 ( .A(n4481), .ZN(n4473) );
  INV_X1 U4999 ( .A(n5121), .ZN(n5131) );
  NAND2_X2 U5000 ( .A1(n4697), .A2(n4696), .ZN(n5121) );
  BUF_X4 U5001 ( .A(n5121), .Z(n4481) );
  XNOR2_X1 U5002 ( .A(n6179), .B(n6177), .ZN(n7516) );
  NAND2_X2 U5003 ( .A1(n5962), .A2(n5965), .ZN(n8627) );
  NAND2_X4 U5004 ( .A1(n8640), .A2(n5973), .ZN(n6022) );
  AND2_X4 U5005 ( .A1(n6621), .A2(n7199), .ZN(n4475) );
  AND2_X1 U5006 ( .A1(n6621), .A2(n7199), .ZN(n5196) );
  NAND2_X1 U5007 ( .A1(n9303), .A2(n8411), .ZN(n9302) );
  OAI21_X1 U5008 ( .B1(n9348), .B2(n4879), .A(n4877), .ZN(n8410) );
  NAND2_X1 U5009 ( .A1(n9350), .A2(n9349), .ZN(n9348) );
  NAND2_X1 U5010 ( .A1(n5557), .A2(n5558), .ZN(n9136) );
  OAI21_X1 U5011 ( .B1(n9330), .B2(n8388), .A(n8389), .ZN(n9309) );
  OAI22_X1 U5012 ( .A1(n9341), .A2(n8387), .B1(n9509), .B2(n9367), .ZN(n9330)
         );
  NAND2_X1 U5013 ( .A1(n9400), .A2(n8401), .ZN(n9376) );
  NAND2_X1 U5014 ( .A1(n4744), .A2(n5536), .ZN(n7920) );
  OAI21_X1 U5015 ( .B1(n7299), .B2(n7298), .A(n8307), .ZN(n8146) );
  INV_X2 U5016 ( .A(n8877), .ZN(n4476) );
  INV_X1 U5017 ( .A(n7332), .ZN(n7250) );
  CLKBUF_X2 U5018 ( .A(n5268), .Z(n5882) );
  INV_X1 U5019 ( .A(n5204), .ZN(n7344) );
  NAND2_X1 U5020 ( .A1(n8723), .A2(n10078), .ZN(n6032) );
  CLKBUF_X1 U5021 ( .A(n6512), .Z(n4480) );
  NAND4_X2 U5022 ( .A1(n6006), .A2(n6005), .A3(n6004), .A4(n6003), .ZN(n7157)
         );
  INV_X1 U5023 ( .A(n6933), .ZN(n9934) );
  CLKBUF_X2 U5024 ( .A(n5238), .Z(n8133) );
  INV_X2 U5025 ( .A(n6022), .ZN(n6062) );
  NAND2_X4 U5026 ( .A1(n4474), .A2(n8627), .ZN(n6692) );
  INV_X2 U5027 ( .A(n6037), .ZN(n6438) );
  CLKBUF_X2 U5028 ( .A(n5174), .Z(n9755) );
  OR2_X1 U5029 ( .A1(n9185), .A2(n5000), .ZN(n4998) );
  NAND2_X1 U5030 ( .A1(n4478), .A2(n4868), .ZN(n9256) );
  NAND2_X1 U5031 ( .A1(n9286), .A2(n4532), .ZN(n4478) );
  AND2_X2 U5032 ( .A1(n9302), .A2(n8412), .ZN(n9286) );
  NAND2_X1 U5033 ( .A1(n8649), .A2(n6381), .ZN(n6391) );
  NAND2_X1 U5034 ( .A1(n9311), .A2(n9318), .ZN(n9310) );
  NAND2_X1 U5035 ( .A1(n4479), .A2(n8404), .ZN(n9350) );
  NAND2_X1 U5036 ( .A1(n9376), .A2(n8403), .ZN(n4479) );
  NAND2_X1 U5037 ( .A1(n9395), .A2(n8400), .ZN(n9400) );
  NAND2_X1 U5038 ( .A1(n9421), .A2(n9433), .ZN(n9395) );
  NAND2_X1 U5039 ( .A1(n9441), .A2(n8399), .ZN(n9421) );
  AND2_X1 U5040 ( .A1(n5533), .A2(n5535), .ZN(n5530) );
  NAND2_X1 U5041 ( .A1(n5504), .A2(n5503), .ZN(n4579) );
  NAND2_X1 U5042 ( .A1(n4876), .A2(n4875), .ZN(n9441) );
  NAND2_X1 U5043 ( .A1(n5778), .A2(n5777), .ZN(n9313) );
  NAND2_X1 U5044 ( .A1(n4833), .A2(n4832), .ZN(n7934) );
  OR2_X1 U5045 ( .A1(n9519), .A2(n8078), .ZN(n8269) );
  AND2_X1 U5046 ( .A1(n6286), .A2(n6247), .ZN(n7982) );
  NAND2_X1 U5047 ( .A1(n4727), .A2(n4725), .ZN(n4994) );
  NAND2_X1 U5048 ( .A1(n7586), .A2(n8132), .ZN(n5669) );
  OR2_X1 U5049 ( .A1(n9471), .A2(n9452), .ZN(n9450) );
  AND2_X1 U5050 ( .A1(n7786), .A2(n4506), .ZN(n4740) );
  XNOR2_X1 U5051 ( .A(n4614), .B(n5695), .ZN(n7586) );
  NAND2_X1 U5052 ( .A1(n7178), .A2(n7173), .ZN(n5336) );
  NAND2_X1 U5053 ( .A1(n7732), .A2(n7856), .ZN(n7855) );
  NAND2_X1 U5054 ( .A1(n6307), .A2(n6306), .ZN(n9042) );
  NAND2_X1 U5055 ( .A1(n7376), .A2(n4987), .ZN(n7178) );
  NAND2_X1 U5056 ( .A1(n7709), .A2(n8173), .ZN(n7710) );
  AND2_X1 U5057 ( .A1(n4967), .A2(n7569), .ZN(n4966) );
  NAND2_X1 U5058 ( .A1(n5282), .A2(n5281), .ZN(n7376) );
  OAI21_X1 U5059 ( .B1(n4587), .B2(n5235), .A(n5234), .ZN(n7117) );
  NAND2_X1 U5060 ( .A1(n6195), .A2(n6196), .ZN(n7568) );
  NAND2_X1 U5061 ( .A1(n5468), .A2(n5467), .ZN(n9712) );
  NAND2_X1 U5062 ( .A1(n6201), .A2(n6200), .ZN(n9057) );
  NAND2_X1 U5063 ( .A1(n5441), .A2(n5440), .ZN(n7851) );
  OR2_X1 U5064 ( .A1(n7706), .A2(n9651), .ZN(n8173) );
  OAI21_X1 U5065 ( .B1(n5539), .B2(n5538), .A(n5537), .ZN(n5560) );
  NAND2_X1 U5066 ( .A1(n5380), .A2(n5379), .ZN(n7706) );
  NAND2_X1 U5067 ( .A1(n5410), .A2(n5409), .ZN(n9737) );
  OR2_X1 U5068 ( .A1(n7412), .A2(n10064), .ZN(n7478) );
  NAND2_X1 U5069 ( .A1(n6169), .A2(n6168), .ZN(n7632) );
  NAND2_X1 U5070 ( .A1(n4908), .A2(n5428), .ZN(n4698) );
  OAI21_X2 U5071 ( .B1(n6493), .B2(n6607), .A(n8907), .ZN(n6494) );
  NAND2_X2 U5072 ( .A1(n6605), .A2(n8907), .ZN(n8877) );
  NAND2_X2 U5073 ( .A1(n6101), .A2(n6100), .ZN(n7420) );
  NAND2_X1 U5074 ( .A1(n6917), .A2(n6012), .ZN(n6907) );
  INV_X1 U5075 ( .A(n7163), .ZN(n7069) );
  AND2_X1 U5076 ( .A1(n6061), .A2(n6060), .ZN(n7163) );
  NAND2_X1 U5077 ( .A1(n7284), .A2(n7194), .ZN(n8073) );
  NAND2_X1 U5078 ( .A1(n7283), .A2(n7285), .ZN(n7284) );
  AND2_X1 U5079 ( .A1(n7195), .A2(n8071), .ZN(n8273) );
  INV_X1 U5080 ( .A(n10037), .ZN(n7152) );
  NAND2_X2 U5081 ( .A1(n7200), .A2(n7199), .ZN(n7257) );
  NAND4_X1 U5082 ( .A1(n5200), .A2(n5199), .A3(n5198), .A4(n5197), .ZN(n5204)
         );
  BUF_X4 U5083 ( .A(n6028), .Z(n10078) );
  NOR2_X1 U5084 ( .A1(n6933), .A2(n7192), .ZN(n7314) );
  OAI211_X1 U5085 ( .C1(n6643), .C2(n5223), .A(n5222), .B(n5221), .ZN(n7351)
         );
  NAND4_X1 U5086 ( .A1(n6027), .A2(n6026), .A3(n6025), .A4(n6024), .ZN(n8723)
         );
  NAND2_X1 U5087 ( .A1(n6062), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6005) );
  INV_X2 U5088 ( .A(n5622), .ZN(n8131) );
  INV_X2 U5089 ( .A(n5223), .ZN(n8132) );
  INV_X1 U5090 ( .A(n5153), .ZN(n8334) );
  NAND2_X1 U5091 ( .A1(n5886), .A2(n5110), .ZN(n6621) );
  XNOR2_X1 U5092 ( .A(n5992), .B(n5991), .ZN(n8587) );
  NAND2_X1 U5093 ( .A1(n5081), .A2(n5080), .ZN(n5082) );
  AOI21_X1 U5094 ( .B1(n5270), .B2(n4701), .A(n4521), .ZN(n4700) );
  INV_X1 U5095 ( .A(n6487), .ZN(n6304) );
  NAND2_X1 U5096 ( .A1(n5148), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5100) );
  NAND2_X1 U5097 ( .A1(n5112), .A2(n5113), .ZN(n5919) );
  NAND2_X1 U5098 ( .A1(n5105), .A2(n5104), .ZN(n7892) );
  NAND2_X1 U5099 ( .A1(n5080), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5078) );
  XNOR2_X1 U5100 ( .A(n5980), .B(n10398), .ZN(n8443) );
  XNOR2_X1 U5101 ( .A(n6452), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8628) );
  XNOR2_X1 U5102 ( .A(n5960), .B(n5959), .ZN(n6497) );
  XNOR2_X1 U5103 ( .A(n5967), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5972) );
  MUX2_X1 U5104 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5111), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5112) );
  NAND2_X2 U5105 ( .A1(n4473), .A2(P1_U3084), .ZN(n9599) );
  NAND2_X1 U5106 ( .A1(n5116), .A2(n5115), .ZN(n8345) );
  NAND2_X1 U5107 ( .A1(n5965), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U5108 ( .A1(n4814), .A2(n4813), .ZN(n5080) );
  NAND2_X1 U5109 ( .A1(n9080), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U5110 ( .A1(n5108), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5103) );
  INV_X2 U5111 ( .A(n7781), .ZN(n4477) );
  INV_X1 U5112 ( .A(n5903), .ZN(n4814) );
  AND2_X1 U5113 ( .A1(n4507), .A2(n5076), .ZN(n4813) );
  NAND2_X1 U5114 ( .A1(n5487), .A2(n5071), .ZN(n5903) );
  AND2_X1 U5115 ( .A1(n5487), .A2(n5090), .ZN(n5092) );
  OR2_X1 U5116 ( .A1(n5106), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5108) );
  XNOR2_X1 U5117 ( .A(n5218), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6892) );
  NAND2_X1 U5118 ( .A1(n4592), .A2(n5119), .ZN(n4697) );
  AND4_X1 U5119 ( .A1(n5955), .A2(n5954), .A3(n10398), .A4(n6457), .ZN(n5956)
         );
  XNOR2_X1 U5120 ( .A(n4862), .B(n5996), .ZN(n6701) );
  AND4_X1 U5121 ( .A1(n5066), .A2(n5065), .A3(n5064), .A4(n5063), .ZN(n5067)
         );
  INV_X1 U5122 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5062) );
  NOR2_X1 U5123 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5061) );
  INV_X1 U5124 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6249) );
  INV_X1 U5125 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6250) );
  NOR2_X1 U5126 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n6182) );
  INV_X1 U5127 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n10398) );
  NOR2_X1 U5128 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5981) );
  AND2_X1 U5129 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5236) );
  INV_X1 U5130 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6248) );
  INV_X2 U5131 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U5132 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5985) );
  INV_X1 U5133 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5119) );
  INV_X1 U5134 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5117) );
  INV_X1 U5135 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5564) );
  INV_X1 U5136 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n10230) );
  INV_X1 U5137 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6069) );
  INV_X1 U5138 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5952) );
  INV_X1 U5139 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5096) );
  INV_X1 U5140 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5099) );
  NOR2_X1 U5141 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5193) );
  INV_X1 U5142 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6128) );
  AND2_X2 U5143 ( .A1(n5067), .A2(n5244), .ZN(n5487) );
  NOR2_X4 U5144 ( .A1(n5138), .A2(n4996), .ZN(n5244) );
  INV_X1 U5145 ( .A(n4867), .ZN(n7283) );
  INV_X2 U5146 ( .A(n5174), .ZN(n5594) );
  NAND2_X1 U5147 ( .A1(n5594), .A2(n9214), .ZN(n4780) );
  NAND2_X1 U5148 ( .A1(n5040), .A2(n7527), .ZN(n7709) );
  AOI21_X2 U5149 ( .B1(n7550), .B2(n8094), .A(n4605), .ZN(n5040) );
  NAND2_X1 U5150 ( .A1(n7435), .A2(n4871), .ZN(n7550) );
  OAI21_X2 U5151 ( .B1(n6096), .B2(n7010), .A(n4984), .ZN(n4983) );
  NAND2_X2 U5152 ( .A1(n7984), .A2(n6286), .ZN(n7910) );
  NOR2_X2 U5153 ( .A1(n9450), .A2(n9431), .ZN(n9419) );
  AND2_X4 U5154 ( .A1(n8057), .A2(n5082), .ZN(n5382) );
  XNOR2_X1 U5155 ( .A(n5078), .B(n5077), .ZN(n8057) );
  NAND2_X2 U5156 ( .A1(n4714), .A2(n4712), .ZN(n6625) );
  OAI22_X2 U5157 ( .A1(n6907), .A2(n6906), .B1(n6021), .B2(n6020), .ZN(n6973)
         );
  BUF_X4 U5158 ( .A(n6429), .Z(n4482) );
  NAND2_X1 U5159 ( .A1(n5972), .A2(n5973), .ZN(n6429) );
  NAND2_X1 U5160 ( .A1(n8145), .A2(n8144), .ZN(n8155) );
  NAND2_X1 U5161 ( .A1(n8146), .A2(n8258), .ZN(n8145) );
  NAND2_X1 U5162 ( .A1(n8872), .A2(n4922), .ZN(n4917) );
  NAND2_X1 U5163 ( .A1(n6692), .A2(n6633), .ZN(n6058) );
  OR2_X1 U5164 ( .A1(n9485), .A2(n8120), .ZN(n8264) );
  NAND2_X1 U5165 ( .A1(n5834), .A2(n5833), .ZN(n5863) );
  OR2_X1 U5166 ( .A1(n8769), .A2(n8774), .ZN(n4860) );
  NAND2_X1 U5167 ( .A1(n8769), .A2(n8774), .ZN(n4861) );
  CLKBUF_X3 U5168 ( .A(n6058), .Z(n8436) );
  OAI211_X1 U5169 ( .C1(n8155), .C2(n8148), .A(n8147), .B(n8308), .ZN(n8152)
         );
  NAND2_X1 U5170 ( .A1(n8223), .A2(n8258), .ZN(n4811) );
  INV_X1 U5171 ( .A(n5459), .ZN(n4905) );
  INV_X1 U5172 ( .A(n6180), .ZN(n4969) );
  INV_X1 U5173 ( .A(n4894), .ZN(n4893) );
  OAI21_X1 U5174 ( .B1(n4896), .B2(n4895), .A(n5615), .ZN(n4894) );
  INV_X1 U5175 ( .A(n5486), .ZN(n4901) );
  NAND2_X1 U5176 ( .A1(n5371), .A2(n10238), .ZN(n5397) );
  NAND2_X1 U5177 ( .A1(n5316), .A2(n5315), .ZN(n5338) );
  AOI21_X1 U5178 ( .B1(n8666), .B2(n8665), .A(n4723), .ZN(n4722) );
  INV_X1 U5179 ( .A(n6425), .ZN(n4723) );
  XNOR2_X1 U5180 ( .A(n7616), .B(n6428), .ZN(n6195) );
  OR2_X1 U5181 ( .A1(n9035), .A2(n8659), .ZN(n8537) );
  OR2_X1 U5182 ( .A1(n7841), .A2(n7807), .ZN(n8515) );
  INV_X1 U5183 ( .A(n7454), .ZN(n4770) );
  OR2_X1 U5184 ( .A1(n9113), .A2(n4993), .ZN(n4992) );
  OR2_X1 U5185 ( .A1(n9514), .A2(n9380), .ZN(n8404) );
  OR2_X1 U5186 ( .A1(n9383), .A2(n8383), .ZN(n8385) );
  OR2_X1 U5187 ( .A1(n9474), .A2(n8106), .ZN(n8398) );
  OAI21_X1 U5188 ( .B1(n5751), .B2(n4543), .A(n4941), .ZN(n5834) );
  INV_X1 U5189 ( .A(n4942), .ZN(n4941) );
  OAI21_X1 U5190 ( .B1(n4945), .B2(n4543), .A(n5806), .ZN(n4942) );
  INV_X1 U5191 ( .A(n5149), .ZN(n5094) );
  AND2_X1 U5192 ( .A1(n5561), .A2(n5543), .ZN(n5559) );
  NAND2_X1 U5193 ( .A1(n5998), .A2(n5999), .ZN(n4976) );
  INV_X1 U5194 ( .A(n8443), .ZN(n8622) );
  NAND2_X1 U5195 ( .A1(n4852), .A2(n4851), .ZN(n4850) );
  INV_X1 U5196 ( .A(n6744), .ZN(n4851) );
  NAND2_X1 U5197 ( .A1(n4860), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n4859) );
  INV_X1 U5198 ( .A(n8571), .ZN(n8614) );
  INV_X1 U5199 ( .A(n8706), .ZN(n8821) );
  NAND2_X1 U5200 ( .A1(n4644), .A2(n4915), .ZN(n4921) );
  NAND2_X1 U5201 ( .A1(n8865), .A2(n4922), .ZN(n4644) );
  OR2_X1 U5202 ( .A1(n8891), .A2(n8892), .ZN(n4646) );
  OAI21_X1 U5203 ( .B1(n8979), .B2(n4549), .A(n4647), .ZN(n4761) );
  NAND2_X1 U5204 ( .A1(n8978), .A2(n7986), .ZN(n4647) );
  AOI21_X1 U5205 ( .B1(n7875), .B2(n4938), .A(n4771), .ZN(n8979) );
  INV_X1 U5206 ( .A(n4937), .ZN(n4771) );
  AOI21_X1 U5207 ( .B1(n4938), .B2(n8522), .A(n4940), .ZN(n4937) );
  NOR2_X1 U5208 ( .A1(n9051), .A2(n8967), .ZN(n4940) );
  INV_X1 U5209 ( .A(n7805), .ZN(n6565) );
  AND2_X1 U5210 ( .A1(n6535), .A2(n8520), .ZN(n8519) );
  INV_X1 U5211 ( .A(n6533), .ZN(n4637) );
  NOR2_X1 U5212 ( .A1(n6564), .A2(n4763), .ZN(n4762) );
  INV_X1 U5213 ( .A(n4767), .ZN(n4763) );
  OR2_X1 U5214 ( .A1(n7616), .A2(n8714), .ZN(n4767) );
  NAND2_X1 U5215 ( .A1(n7625), .A2(n8601), .ZN(n6532) );
  INV_X1 U5216 ( .A(n8971), .ZN(n8953) );
  OAI21_X1 U5217 ( .B1(n7061), .B2(n6524), .A(n6523), .ZN(n7225) );
  OR2_X1 U5218 ( .A1(n6666), .A2(n6694), .ZN(n8958) );
  INV_X1 U5219 ( .A(n8956), .ZN(n8966) );
  NAND2_X1 U5220 ( .A1(n4953), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U5221 ( .A1(n5988), .A2(n5987), .ZN(n4953) );
  NAND2_X1 U5222 ( .A1(n5181), .A2(n4584), .ZN(n6867) );
  AND2_X1 U5223 ( .A1(n6868), .A2(n5180), .ZN(n4584) );
  NAND3_X1 U5224 ( .A1(n5071), .A2(n5487), .A3(n4525), .ZN(n5115) );
  INV_X1 U5225 ( .A(n5845), .ZN(n5928) );
  NAND2_X1 U5226 ( .A1(n4792), .A2(n4791), .ZN(n4789) );
  OAI21_X1 U5227 ( .B1(n9294), .B2(n4513), .A(n8391), .ZN(n9280) );
  NOR2_X2 U5228 ( .A1(n9313), .A2(n9333), .ZN(n9312) );
  NAND2_X1 U5229 ( .A1(n7190), .A2(n7341), .ZN(n4828) );
  AND2_X1 U5230 ( .A1(n5174), .A2(n4481), .ZN(n5192) );
  NAND2_X1 U5231 ( .A1(n8119), .A2(n8118), .ZN(n9485) );
  AND2_X1 U5232 ( .A1(n9674), .A2(n9963), .ZN(n9970) );
  NAND2_X1 U5233 ( .A1(n5094), .A2(n5093), .ZN(n5148) );
  NAND2_X1 U5234 ( .A1(n6427), .A2(n6426), .ZN(n8999) );
  INV_X1 U5235 ( .A(n8721), .ZN(n7229) );
  OR2_X1 U5236 ( .A1(n6666), .A2(n4474), .ZN(n8956) );
  OAI21_X1 U5237 ( .B1(n8795), .B2(n9612), .A(n4866), .ZN(n4865) );
  AOI21_X1 U5238 ( .B1(n8796), .B2(n10010), .A(n9618), .ZN(n4866) );
  INV_X1 U5239 ( .A(n8259), .ZN(n8339) );
  AOI21_X1 U5240 ( .B1(n9284), .B2(n8413), .A(n8414), .ZN(n8416) );
  NAND2_X1 U5241 ( .A1(n8499), .A2(n4680), .ZN(n4679) );
  OAI211_X1 U5242 ( .C1(n4510), .C2(n4799), .A(n4798), .B(n4796), .ZN(n4795)
         );
  NAND2_X1 U5243 ( .A1(n8194), .A2(n8213), .ZN(n4799) );
  INV_X1 U5244 ( .A(n4797), .ZN(n4796) );
  NAND2_X1 U5245 ( .A1(n8271), .A2(n8272), .ZN(n4794) );
  NOR2_X1 U5246 ( .A1(n4676), .A2(n4674), .ZN(n4673) );
  NOR2_X1 U5247 ( .A1(n4677), .A2(n8950), .ZN(n4674) );
  NAND2_X1 U5248 ( .A1(n8538), .A2(n8539), .ZN(n4676) );
  NAND2_X1 U5249 ( .A1(n4673), .A2(n4677), .ZN(n4672) );
  AOI21_X1 U5250 ( .B1(n8224), .B2(n8213), .A(n8225), .ZN(n4810) );
  NAND2_X1 U5251 ( .A1(n8229), .A2(n8258), .ZN(n8233) );
  INV_X1 U5252 ( .A(n8559), .ZN(n4693) );
  NAND2_X1 U5253 ( .A1(n4694), .A2(n4690), .ZN(n4689) );
  INV_X1 U5254 ( .A(n8551), .ZN(n4690) );
  NAND2_X1 U5255 ( .A1(n4687), .A2(n4688), .ZN(n4686) );
  NAND2_X1 U5256 ( .A1(n4692), .A2(n4694), .ZN(n4688) );
  NAND2_X1 U5257 ( .A1(n6517), .A2(n10037), .ZN(n8474) );
  OR2_X1 U5258 ( .A1(n5685), .A2(n9120), .ZN(n5687) );
  NAND2_X1 U5259 ( .A1(n4740), .A2(n4738), .ZN(n4737) );
  INV_X1 U5260 ( .A(n7638), .ZN(n4738) );
  NOR2_X1 U5261 ( .A1(n7794), .A2(n4986), .ZN(n4591) );
  INV_X1 U5262 ( .A(n5458), .ZN(n4986) );
  NAND2_X1 U5263 ( .A1(n7855), .A2(n8282), .ZN(n4874) );
  INV_X1 U5264 ( .A(n5589), .ZN(n4895) );
  NAND2_X1 U5265 ( .A1(n5515), .A2(n5514), .ZN(n5537) );
  OAI21_X1 U5266 ( .B1(n4906), .B2(n4905), .A(n5051), .ZN(n4904) );
  NOR2_X1 U5267 ( .A1(n4520), .A2(n4608), .ZN(n4607) );
  INV_X1 U5268 ( .A(n5397), .ZN(n4608) );
  NOR2_X1 U5269 ( .A1(n4901), .A2(n4905), .ZN(n4900) );
  NAND2_X1 U5270 ( .A1(n4702), .A2(n5053), .ZN(n4708) );
  INV_X1 U5271 ( .A(n4924), .ZN(n4702) );
  OAI211_X1 U5272 ( .C1(n4697), .C2(n4596), .A(n4594), .B(n4593), .ZN(n5250)
         );
  NAND2_X1 U5273 ( .A1(n4595), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n4594) );
  INV_X1 U5274 ( .A(n4696), .ZN(n4595) );
  AND2_X1 U5275 ( .A1(n4958), .A2(n8642), .ZN(n4957) );
  NAND2_X1 U5276 ( .A1(n4722), .A2(n4720), .ZN(n4719) );
  NAND2_X1 U5277 ( .A1(n8694), .A2(n6425), .ZN(n4958) );
  NAND2_X1 U5278 ( .A1(n6214), .A2(n6232), .ZN(n4715) );
  NAND2_X1 U5279 ( .A1(n8438), .A2(n8577), .ZN(n4888) );
  OR2_X1 U5280 ( .A1(n9005), .A2(n8837), .ZN(n8560) );
  OR2_X1 U5281 ( .A1(n9014), .A2(n8669), .ZN(n8553) );
  NAND2_X1 U5282 ( .A1(n4631), .A2(n8922), .ZN(n4627) );
  NOR2_X1 U5283 ( .A1(n9030), .A2(n9025), .ZN(n4656) );
  OR2_X1 U5284 ( .A1(n9025), .A2(n8660), .ZN(n8546) );
  NAND2_X1 U5285 ( .A1(n6309), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6327) );
  INV_X1 U5286 ( .A(n6310), .ZN(n6309) );
  NAND2_X1 U5287 ( .A1(n8521), .A2(n8520), .ZN(n5006) );
  AND2_X1 U5288 ( .A1(n5039), .A2(n8487), .ZN(n4573) );
  NAND2_X1 U5289 ( .A1(n6130), .A2(n4881), .ZN(n8497) );
  NOR2_X1 U5290 ( .A1(n7406), .A2(n4882), .ZN(n4881) );
  INV_X1 U5291 ( .A(n6129), .ZN(n4882) );
  NAND2_X1 U5292 ( .A1(n4884), .A2(n7406), .ZN(n8500) );
  NAND2_X1 U5293 ( .A1(n7101), .A2(n8486), .ZN(n4574) );
  NOR2_X1 U5294 ( .A1(n6558), .A2(n5010), .ZN(n5009) );
  INV_X1 U5295 ( .A(n8458), .ZN(n5010) );
  NAND2_X1 U5296 ( .A1(n7064), .A2(n8479), .ZN(n8457) );
  INV_X1 U5297 ( .A(n6518), .ZN(n4621) );
  NAND2_X1 U5298 ( .A1(n4649), .A2(n6991), .ZN(n8458) );
  AND2_X1 U5299 ( .A1(n8473), .A2(n8474), .ZN(n6555) );
  NAND2_X1 U5300 ( .A1(n8635), .A2(n6554), .ZN(n8464) );
  NAND2_X1 U5301 ( .A1(n4480), .A2(n6513), .ZN(n8471) );
  OR2_X1 U5302 ( .A1(n6586), .A2(n6908), .ZN(n6601) );
  INV_X1 U5303 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5957) );
  INV_X1 U5304 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6457) );
  INV_X1 U5305 ( .A(n8057), .ZN(n5083) );
  INV_X1 U5306 ( .A(n4870), .ZN(n4869) );
  NOR2_X1 U5307 ( .A1(n8415), .A2(n8234), .ZN(n4870) );
  NAND2_X1 U5308 ( .A1(n8408), .A2(n8407), .ZN(n4879) );
  OR2_X1 U5309 ( .A1(n9313), .A2(n9194), .ZN(n8409) );
  AND2_X1 U5310 ( .A1(n8406), .A2(n8405), .ZN(n4880) );
  NAND2_X1 U5311 ( .A1(n9461), .A2(n9467), .ZN(n4876) );
  NOR2_X1 U5312 ( .A1(n9712), .A2(n8082), .ZN(n4779) );
  INV_X1 U5313 ( .A(n4835), .ZN(n4834) );
  OAI21_X1 U5314 ( .B1(n7739), .B2(n4836), .A(n7854), .ZN(n4835) );
  INV_X1 U5315 ( .A(n7852), .ZN(n4836) );
  OR2_X1 U5316 ( .A1(n7851), .A2(n7799), .ZN(n8184) );
  INV_X1 U5317 ( .A(n7524), .ZN(n4826) );
  INV_X1 U5318 ( .A(n7430), .ZN(n4827) );
  AND2_X1 U5319 ( .A1(n5153), .A2(n9430), .ZN(n5918) );
  INV_X1 U5320 ( .A(n8130), .ZN(n4936) );
  AND2_X1 U5321 ( .A1(n8127), .A2(n4936), .ZN(n4934) );
  INV_X1 U5322 ( .A(n8127), .ZN(n4931) );
  XNOR2_X1 U5323 ( .A(n8126), .B(n8125), .ZN(n8123) );
  AND2_X1 U5324 ( .A1(n5861), .A2(n5812), .ZN(n5833) );
  NOR2_X1 U5325 ( .A1(n5768), .A2(n4946), .ZN(n4945) );
  INV_X1 U5326 ( .A(n5750), .ZN(n4946) );
  OAI21_X1 U5327 ( .B1(n5093), .B2(n4749), .A(n5099), .ZN(n4748) );
  NOR2_X1 U5328 ( .A1(n5590), .A2(n4897), .ZN(n4896) );
  INV_X1 U5329 ( .A(n5561), .ZN(n4897) );
  NAND2_X1 U5330 ( .A1(n5432), .A2(n5431), .ZN(n5459) );
  NOR2_X1 U5331 ( .A1(n5460), .A2(n4907), .ZN(n4906) );
  INV_X1 U5332 ( .A(n5428), .ZN(n4907) );
  OR2_X1 U5333 ( .A1(n5430), .A2(n5429), .ZN(n4908) );
  NAND2_X1 U5334 ( .A1(n5398), .A2(n5397), .ZN(n5430) );
  AOI21_X1 U5335 ( .B1(n4924), .B2(n4926), .A(n4711), .ZN(n4710) );
  NAND2_X1 U5336 ( .A1(n4708), .A2(n5368), .ZN(n4707) );
  AOI21_X1 U5337 ( .B1(n5310), .B2(n4927), .A(n4925), .ZN(n4924) );
  INV_X1 U5338 ( .A(n5338), .ZN(n4925) );
  INV_X1 U5339 ( .A(n4927), .ZN(n4926) );
  NAND2_X1 U5340 ( .A1(n4612), .A2(SI_8_), .ZN(n5317) );
  INV_X1 U5341 ( .A(n5316), .ZN(n4612) );
  INV_X1 U5342 ( .A(n5247), .ZN(n5248) );
  NAND2_X1 U5343 ( .A1(n5136), .A2(n5135), .ZN(n5249) );
  NOR2_X1 U5344 ( .A1(n7836), .A2(n4975), .ZN(n4974) );
  INV_X1 U5345 ( .A(n6215), .ZN(n4975) );
  INV_X1 U5346 ( .A(n4960), .ZN(n4959) );
  OAI21_X1 U5347 ( .B1(n4963), .B2(n4961), .A(n4966), .ZN(n4960) );
  NAND2_X1 U5348 ( .A1(n6342), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6358) );
  INV_X1 U5349 ( .A(n6343), .ZN(n6342) );
  INV_X1 U5350 ( .A(n6414), .ZN(n6412) );
  AOI21_X1 U5351 ( .B1(n8430), .B2(n8573), .A(n8429), .ZN(n8433) );
  INV_X1 U5352 ( .A(n4888), .ZN(n8616) );
  INV_X1 U5353 ( .A(n8625), .ZN(n4571) );
  NAND2_X1 U5354 ( .A1(n4885), .A2(n8587), .ZN(n8625) );
  NAND2_X1 U5355 ( .A1(n4889), .A2(n4886), .ZN(n4885) );
  INV_X1 U5356 ( .A(n8583), .ZN(n4889) );
  OAI211_X1 U5357 ( .C1(n8617), .C2(n8572), .A(n8579), .B(n4887), .ZN(n4886)
         );
  AND2_X1 U5358 ( .A1(n4848), .A2(n4847), .ZN(n8726) );
  NAND2_X1 U5359 ( .A1(n7589), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4847) );
  NAND2_X1 U5360 ( .A1(n9079), .A2(n6547), .ZN(n4932) );
  INV_X1 U5361 ( .A(n8707), .ZN(n8837) );
  NAND2_X1 U5362 ( .A1(n8852), .A2(n8837), .ZN(n4920) );
  AND2_X1 U5363 ( .A1(n8553), .A2(n8551), .ZN(n8892) );
  NOR2_X1 U5364 ( .A1(n5034), .A2(n5033), .ZN(n8881) );
  INV_X1 U5365 ( .A(n8549), .ZN(n5033) );
  INV_X1 U5366 ( .A(n8896), .ZN(n5034) );
  INV_X1 U5367 ( .A(n8883), .ZN(n8924) );
  NAND2_X1 U5368 ( .A1(n8936), .A2(n5025), .ZN(n8926) );
  AND2_X1 U5369 ( .A1(n5029), .A2(n8538), .ZN(n5025) );
  NAND2_X1 U5370 ( .A1(n8945), .A2(n4656), .ZN(n8915) );
  AOI21_X1 U5371 ( .B1(n4631), .B2(n4629), .A(n4508), .ZN(n4628) );
  INV_X1 U5372 ( .A(n8955), .ZN(n4629) );
  INV_X1 U5373 ( .A(n8537), .ZN(n5028) );
  NAND2_X1 U5374 ( .A1(n8952), .A2(n5027), .ZN(n8936) );
  NOR2_X1 U5375 ( .A1(n8611), .A2(n5028), .ZN(n5027) );
  OAI21_X1 U5376 ( .B1(n4761), .B2(n4760), .A(n4544), .ZN(n8944) );
  NOR2_X1 U5377 ( .A1(n9042), .A2(n8969), .ZN(n4760) );
  INV_X1 U5378 ( .A(n6539), .ZN(n4939) );
  NAND2_X1 U5379 ( .A1(n6538), .A2(n6537), .ZN(n7873) );
  INV_X1 U5380 ( .A(n7875), .ZN(n6538) );
  NAND2_X1 U5381 ( .A1(n7649), .A2(n5020), .ZN(n5019) );
  AOI21_X1 U5382 ( .B1(n5022), .B2(n5018), .A(n5021), .ZN(n5017) );
  NAND2_X1 U5383 ( .A1(n4634), .A2(n4515), .ZN(n7808) );
  NAND2_X1 U5384 ( .A1(n4484), .A2(n6534), .ZN(n4636) );
  NAND2_X1 U5385 ( .A1(n6532), .A2(n4765), .ZN(n4764) );
  NOR2_X1 U5386 ( .A1(n8603), .A2(n4766), .ZN(n4765) );
  INV_X1 U5387 ( .A(n6531), .ZN(n4766) );
  NAND2_X1 U5388 ( .A1(n5024), .A2(n6564), .ZN(n7652) );
  AND2_X1 U5389 ( .A1(n8511), .A2(n8510), .ZN(n8603) );
  AOI21_X1 U5390 ( .B1(n7453), .B2(n4768), .A(n4519), .ZN(n7625) );
  NOR2_X1 U5391 ( .A1(n4770), .A2(n4769), .ZN(n4768) );
  INV_X1 U5392 ( .A(n6530), .ZN(n4769) );
  OR2_X1 U5393 ( .A1(n7401), .A2(n4618), .ZN(n7453) );
  NAND2_X1 U5394 ( .A1(n7403), .A2(n6528), .ZN(n4618) );
  AND2_X1 U5395 ( .A1(n8487), .A2(n8486), .ZN(n8595) );
  NAND2_X1 U5396 ( .A1(n8460), .A2(n8457), .ZN(n5015) );
  INV_X1 U5397 ( .A(n8719), .ZN(n7407) );
  INV_X1 U5398 ( .A(n6648), .ZN(n4641) );
  INV_X1 U5399 ( .A(n6058), .ZN(n4643) );
  INV_X1 U5400 ( .A(n6692), .ZN(n4639) );
  INV_X1 U5401 ( .A(n8958), .ZN(n8968) );
  OR2_X1 U5402 ( .A1(n6030), .A2(n6637), .ZN(n4773) );
  NAND2_X1 U5403 ( .A1(n6549), .A2(n6548), .ZN(n6606) );
  AND2_X1 U5404 ( .A1(n6580), .A2(n6579), .ZN(n6604) );
  NAND2_X1 U5405 ( .A1(n6323), .A2(n6322), .ZN(n9035) );
  NAND2_X1 U5406 ( .A1(n6289), .A2(n6288), .ZN(n9045) );
  NOR2_X1 U5407 ( .A1(n4499), .A2(n4651), .ZN(n4650) );
  OR2_X1 U5408 ( .A1(n8436), .A2(n6644), .ZN(n6031) );
  NAND2_X1 U5409 ( .A1(n4952), .A2(n4951), .ZN(n5994) );
  AOI21_X1 U5410 ( .B1(n4954), .B2(n5968), .A(n5968), .ZN(n4951) );
  INV_X1 U5411 ( .A(n4955), .ZN(n4954) );
  AND2_X1 U5412 ( .A1(n6098), .A2(n6074), .ZN(n6844) );
  NAND2_X1 U5413 ( .A1(n9188), .A2(n5832), .ZN(n5859) );
  OR2_X1 U5414 ( .A1(n9187), .A2(n9091), .ZN(n5000) );
  NAND2_X1 U5415 ( .A1(n7637), .A2(n7638), .ZN(n4741) );
  NAND2_X1 U5416 ( .A1(n7504), .A2(n4729), .ZN(n4728) );
  NOR2_X1 U5417 ( .A1(n4729), .A2(n7504), .ZN(n4730) );
  NAND2_X1 U5418 ( .A1(n5651), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U5419 ( .A1(n9177), .A2(n4735), .ZN(n4734) );
  NOR2_X1 U5420 ( .A1(n4991), .A2(n4736), .ZN(n4735) );
  AND2_X1 U5421 ( .A1(n5922), .A2(n9931), .ZN(n7047) );
  XNOR2_X1 U5422 ( .A(n5203), .B(n7257), .ZN(n5205) );
  OR2_X1 U5423 ( .A1(n8262), .A2(n5918), .ZN(n5922) );
  OR2_X1 U5424 ( .A1(n5803), .A2(n5802), .ZN(n5804) );
  NAND2_X1 U5425 ( .A1(n8339), .A2(n8297), .ZN(n8262) );
  NAND2_X1 U5426 ( .A1(n8339), .A2(n9430), .ZN(n7200) );
  INV_X1 U5427 ( .A(n5382), .ZN(n5848) );
  INV_X1 U5428 ( .A(n5238), .ZN(n5784) );
  AND2_X1 U5429 ( .A1(n5083), .A2(n5082), .ZN(n5238) );
  NAND2_X1 U5430 ( .A1(n6803), .A2(n6780), .ZN(n6879) );
  NOR2_X1 U5431 ( .A1(n9890), .A2(n4754), .ZN(n9906) );
  AND2_X1 U5432 ( .A1(n9234), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4754) );
  NOR2_X1 U5433 ( .A1(n8420), .A2(n9485), .ZN(n4792) );
  NAND2_X1 U5434 ( .A1(n9310), .A2(n8390), .ZN(n9294) );
  NAND2_X1 U5435 ( .A1(n5753), .A2(n5752), .ZN(n9331) );
  NAND2_X1 U5436 ( .A1(n9348), .A2(n4880), .ZN(n9326) );
  NOR2_X1 U5437 ( .A1(n8385), .A2(n4824), .ZN(n4823) );
  INV_X1 U5438 ( .A(n8375), .ZN(n4824) );
  OAI21_X1 U5439 ( .B1(n8385), .B2(n4822), .A(n8384), .ZN(n4820) );
  NAND2_X1 U5440 ( .A1(n4501), .A2(n8375), .ZN(n4822) );
  NOR2_X1 U5441 ( .A1(n5044), .A2(n5060), .ZN(n8384) );
  INV_X1 U5442 ( .A(n8156), .ZN(n4605) );
  NAND2_X1 U5443 ( .A1(n4827), .A2(n7431), .ZN(n7523) );
  NAND2_X1 U5444 ( .A1(n7296), .A2(n4500), .ZN(n7384) );
  AND3_X1 U5445 ( .A1(n4604), .A2(n5253), .A3(n4603), .ZN(n7246) );
  NAND2_X1 U5446 ( .A1(n5594), .A2(n6784), .ZN(n4603) );
  NAND2_X1 U5447 ( .A1(n6640), .A2(n8132), .ZN(n4604) );
  NAND2_X1 U5448 ( .A1(n7245), .A2(n8304), .ZN(n7299) );
  NAND2_X1 U5449 ( .A1(n4486), .A2(n7191), .ZN(n4829) );
  INV_X1 U5450 ( .A(n8273), .ZN(n7188) );
  NAND2_X1 U5451 ( .A1(n4867), .A2(n7280), .ZN(n7279) );
  INV_X1 U5452 ( .A(n9668), .ZN(n9705) );
  INV_X1 U5453 ( .A(n9670), .ZN(n9702) );
  OR2_X1 U5454 ( .A1(n8262), .A2(n6876), .ZN(n9670) );
  AND2_X1 U5455 ( .A1(n4502), .A2(n9264), .ZN(n9486) );
  NAND2_X1 U5456 ( .A1(n5596), .A2(n5595), .ZN(n9452) );
  AND2_X1 U5457 ( .A1(n8258), .A2(n5153), .ZN(n9950) );
  XNOR2_X1 U5458 ( .A(n8123), .B(SI_30_), .ZN(n8432) );
  NAND2_X1 U5459 ( .A1(n5092), .A2(n5047), .ZN(n5149) );
  NAND2_X1 U5460 ( .A1(n7666), .A2(n6215), .ZN(n7835) );
  NAND2_X1 U5461 ( .A1(n6221), .A2(n6220), .ZN(n7841) );
  NAND2_X1 U5462 ( .A1(n6153), .A2(n6152), .ZN(n7462) );
  NAND2_X1 U5463 ( .A1(n4972), .A2(n4551), .ZN(n4971) );
  NAND2_X1 U5464 ( .A1(n8993), .A2(n6494), .ZN(n4972) );
  AOI21_X1 U5465 ( .B1(n4558), .B2(n7516), .A(n6180), .ZN(n7571) );
  NAND2_X1 U5466 ( .A1(n6811), .A2(n6547), .ZN(n6187) );
  NAND2_X1 U5467 ( .A1(n6255), .A2(n6254), .ZN(n9632) );
  NAND2_X1 U5468 ( .A1(n6986), .A2(n6057), .ZN(n7034) );
  AND2_X1 U5469 ( .A1(n6496), .A2(n6488), .ZN(n9628) );
  NAND4_X1 U5470 ( .A1(n6067), .A2(n5050), .A3(n6066), .A4(n6065), .ZN(n8721)
         );
  NOR2_X1 U5471 ( .A1(n6696), .A2(n6695), .ZN(n6713) );
  OR2_X1 U5472 ( .A1(n6716), .A2(n6715), .ZN(n4856) );
  NOR2_X1 U5473 ( .A1(n6713), .A2(n4857), .ZN(n6716) );
  AND2_X1 U5474 ( .A1(n6717), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4857) );
  OR2_X1 U5475 ( .A1(n6742), .A2(n4546), .ZN(n4852) );
  INV_X1 U5476 ( .A(n4850), .ZN(n6840) );
  AND2_X1 U5477 ( .A1(n4859), .A2(n4861), .ZN(n8789) );
  XNOR2_X1 U5478 ( .A(n8988), .B(n8987), .ZN(n8986) );
  NAND2_X1 U5479 ( .A1(n4910), .A2(n4909), .ZN(n6550) );
  NAND2_X1 U5480 ( .A1(n4912), .A2(n4492), .ZN(n4909) );
  NOR2_X1 U5481 ( .A1(n8834), .A2(n8564), .ZN(n8820) );
  OAI21_X1 U5482 ( .B1(n4921), .B2(n8563), .A(n4918), .ZN(n8811) );
  AND2_X1 U5483 ( .A1(n7963), .A2(n4649), .ZN(n4648) );
  AOI21_X1 U5484 ( .B1(n8986), .B2(n10035), .A(n4659), .ZN(n4658) );
  OAI21_X1 U5485 ( .B1(n8987), .B2(n10076), .A(n8990), .ZN(n4659) );
  NOR2_X1 U5486 ( .A1(n7175), .A2(n4988), .ZN(n4987) );
  INV_X1 U5487 ( .A(n5286), .ZN(n4988) );
  NAND2_X1 U5488 ( .A1(n5571), .A2(n5570), .ZN(n9474) );
  NAND2_X1 U5489 ( .A1(n6930), .A2(n5187), .ZN(n5188) );
  MUX2_X1 U5490 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5114), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5116) );
  NAND2_X1 U5491 ( .A1(n5823), .A2(n5822), .ZN(n9287) );
  OR2_X1 U5492 ( .A1(n9190), .A2(n5928), .ZN(n5823) );
  NOR2_X1 U5493 ( .A1(n9855), .A2(n9854), .ZN(n9853) );
  XNOR2_X1 U5494 ( .A(n4843), .B(n9255), .ZN(n9484) );
  NAND2_X1 U5495 ( .A1(n9252), .A2(n4548), .ZN(n4843) );
  NAND2_X1 U5496 ( .A1(n5625), .A2(n5624), .ZN(n9431) );
  INV_X1 U5497 ( .A(n9271), .ZN(n4602) );
  OR2_X1 U5498 ( .A1(n9279), .A2(n9970), .ZN(n8422) );
  INV_X1 U5499 ( .A(n9931), .ZN(n8337) );
  AOI21_X1 U5500 ( .B1(n5902), .B2(n9930), .A(n5901), .ZN(n9928) );
  XNOR2_X1 U5501 ( .A(n5147), .B(n5146), .ZN(n8259) );
  INV_X1 U5502 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4597) );
  INV_X1 U5503 ( .A(n8457), .ZN(n8478) );
  NAND2_X1 U5504 ( .A1(n8476), .A2(n8481), .ZN(n4668) );
  OAI21_X1 U5505 ( .B1(n4669), .B2(n4667), .A(n4666), .ZN(n8489) );
  AND2_X1 U5506 ( .A1(n8595), .A2(n4503), .ZN(n4666) );
  AOI21_X1 U5507 ( .B1(n8470), .B2(n8469), .A(n4668), .ZN(n4667) );
  INV_X1 U5508 ( .A(n8484), .ZN(n4669) );
  AOI211_X1 U5509 ( .C1(n8177), .C2(n8176), .A(n8175), .B(n8174), .ZN(n8182)
         );
  NOR2_X1 U5510 ( .A1(n4682), .A2(n4681), .ZN(n4680) );
  NAND2_X1 U5511 ( .A1(n8501), .A2(n8572), .ZN(n4681) );
  INV_X1 U5512 ( .A(n8498), .ZN(n4682) );
  OAI21_X1 U5513 ( .B1(n8195), .B2(n8213), .A(n9672), .ZN(n4797) );
  NAND2_X1 U5514 ( .A1(n4678), .A2(n4514), .ZN(n8513) );
  NAND2_X1 U5515 ( .A1(n4793), .A2(n8258), .ZN(n8216) );
  OAI21_X1 U5516 ( .B1(n8212), .B2(n4794), .A(n8400), .ZN(n4793) );
  AND2_X1 U5517 ( .A1(n8546), .A2(n8540), .ZN(n4675) );
  NAND2_X1 U5518 ( .A1(n4809), .A2(n5052), .ZN(n8241) );
  NAND2_X1 U5519 ( .A1(n4811), .A2(n4810), .ZN(n4809) );
  AOI21_X1 U5520 ( .B1(n4523), .B2(n4692), .A(n4691), .ZN(n4687) );
  AND2_X1 U5521 ( .A1(n4496), .A2(n4932), .ZN(n8581) );
  INV_X1 U5522 ( .A(n8429), .ZN(n8574) );
  OR2_X1 U5523 ( .A1(n5795), .A2(n9129), .ZN(n5797) );
  NAND2_X1 U5524 ( .A1(n9313), .A2(n9194), .ZN(n8265) );
  INV_X1 U5525 ( .A(n9387), .ZN(n8383) );
  OAI21_X1 U5526 ( .B1(n5865), .B2(n4949), .A(n4947), .ZN(n8126) );
  AND2_X1 U5527 ( .A1(n4948), .A2(n8055), .ZN(n4947) );
  OR2_X1 U5528 ( .A1(n4557), .A2(n4949), .ZN(n4948) );
  INV_X1 U5529 ( .A(n5772), .ZN(n4943) );
  NOR2_X1 U5530 ( .A1(n5339), .A2(n4928), .ZN(n4927) );
  INV_X1 U5531 ( .A(n5251), .ZN(n4701) );
  INV_X1 U5532 ( .A(n7516), .ZN(n4968) );
  INV_X1 U5533 ( .A(n7359), .ZN(n4961) );
  OR3_X1 U5534 ( .A1(n6586), .A2(n6599), .A3(n6598), .ZN(n6504) );
  OR2_X1 U5535 ( .A1(n6606), .A2(n8822), .ZN(n8573) );
  AND2_X1 U5536 ( .A1(n6606), .A2(n8822), .ZN(n8429) );
  NAND2_X1 U5537 ( .A1(n4888), .A2(n8572), .ZN(n4887) );
  AND2_X1 U5538 ( .A1(n8573), .A2(n8574), .ZN(n8571) );
  INV_X1 U5539 ( .A(n6292), .ZN(n6290) );
  INV_X1 U5540 ( .A(n6256), .ZN(n6237) );
  NAND2_X1 U5541 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(n6237), .ZN(n6292) );
  NAND2_X1 U5542 ( .A1(n4665), .A2(n9637), .ZN(n4664) );
  NOR2_X1 U5543 ( .A1(n7815), .A2(n7841), .ZN(n4665) );
  NOR2_X1 U5544 ( .A1(n6564), .A2(n5023), .ZN(n5022) );
  INV_X1 U5545 ( .A(n8515), .ZN(n5021) );
  NAND2_X1 U5546 ( .A1(n7612), .A2(n7675), .ZN(n7656) );
  NOR3_X1 U5547 ( .A1(n7478), .A2(n4660), .A3(n7616), .ZN(n7612) );
  NAND2_X1 U5548 ( .A1(n4661), .A2(n7725), .ZN(n4660) );
  INV_X1 U5549 ( .A(n4662), .ZN(n4661) );
  NAND2_X1 U5550 ( .A1(n10071), .A2(n7479), .ZN(n4662) );
  NAND2_X1 U5551 ( .A1(n8721), .A2(n7163), .ZN(n8479) );
  NAND2_X1 U5552 ( .A1(n7273), .A2(n7152), .ZN(n8473) );
  NAND2_X1 U5553 ( .A1(n8464), .A2(n8471), .ZN(n7143) );
  NAND2_X1 U5554 ( .A1(n8464), .A2(n5016), .ZN(n7145) );
  AND3_X1 U5555 ( .A1(n8473), .A2(n8471), .A3(n8474), .ZN(n5016) );
  OAI21_X1 U5556 ( .B1(n5987), .B2(n5968), .A(n5989), .ZN(n4955) );
  OR2_X1 U5557 ( .A1(n6184), .A2(n5968), .ZN(n6147) );
  AND2_X1 U5558 ( .A1(n6018), .A2(n5951), .ZN(n6047) );
  NAND2_X1 U5559 ( .A1(n9166), .A2(n5721), .ZN(n4581) );
  NOR2_X1 U5560 ( .A1(n9166), .A2(n5721), .ZN(n4582) );
  INV_X1 U5561 ( .A(n9175), .ZN(n4736) );
  NOR2_X1 U5562 ( .A1(n9176), .A2(n4991), .ZN(n4732) );
  INV_X1 U5563 ( .A(n4989), .ZN(n4733) );
  AOI21_X1 U5564 ( .B1(n4990), .B2(n4993), .A(n4516), .ZN(n4989) );
  INV_X1 U5565 ( .A(n4740), .ZN(n4739) );
  NOR2_X1 U5566 ( .A1(n8257), .A2(n8321), .ZN(n4803) );
  AOI21_X1 U5567 ( .B1(n8253), .B2(n8321), .A(n4505), .ZN(n4801) );
  OAI21_X1 U5568 ( .B1(n8254), .B2(n9201), .A(n8255), .ZN(n4808) );
  NOR2_X1 U5569 ( .A1(n8251), .A2(n8321), .ZN(n4805) );
  INV_X1 U5570 ( .A(n5907), .ZN(n8297) );
  INV_X1 U5571 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5073) );
  INV_X1 U5572 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5324) );
  NOR2_X1 U5573 ( .A1(n9811), .A2(n4756), .ZN(n9826) );
  NOR2_X1 U5574 ( .A1(n4758), .A2(n4757), .ZN(n4756) );
  INV_X1 U5575 ( .A(n9816), .ZN(n4758) );
  NOR2_X1 U5576 ( .A1(n9826), .A2(n9825), .ZN(n9824) );
  OR2_X1 U5577 ( .A1(n8420), .A2(n9253), .ZN(n8249) );
  OR2_X1 U5578 ( .A1(n5755), .A2(n5754), .ZN(n5780) );
  NOR2_X1 U5579 ( .A1(n9509), .A2(n4784), .ZN(n4782) );
  INV_X1 U5580 ( .A(n4819), .ZN(n4818) );
  NOR2_X1 U5581 ( .A1(n9384), .A2(n8383), .ZN(n5044) );
  NOR2_X1 U5582 ( .A1(n9519), .A2(n9408), .ZN(n4786) );
  AND2_X1 U5583 ( .A1(n8199), .A2(n8198), .ZN(n9672) );
  INV_X1 U5584 ( .A(n7383), .ZN(n4839) );
  OAI21_X1 U5585 ( .B1(n4500), .B2(n4839), .A(n8277), .ZN(n4838) );
  OR2_X1 U5586 ( .A1(n7392), .A2(n7427), .ZN(n7439) );
  INV_X1 U5587 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5261) );
  NAND2_X1 U5588 ( .A1(n9210), .A2(n7246), .ZN(n8305) );
  NAND2_X1 U5589 ( .A1(n7310), .A2(n7351), .ZN(n8303) );
  NAND2_X1 U5590 ( .A1(n8073), .A2(n8273), .ZN(n4812) );
  NAND2_X1 U5591 ( .A1(n8419), .A2(n9275), .ZN(n9263) );
  NAND2_X1 U5592 ( .A1(n4874), .A2(n8097), .ZN(n9697) );
  AOI21_X1 U5593 ( .B1(n4893), .B2(n4895), .A(n4552), .ZN(n4891) );
  NAND2_X1 U5594 ( .A1(n5537), .A2(n5517), .ZN(n5538) );
  NAND2_X1 U5595 ( .A1(n5398), .A2(n4607), .ZN(n4611) );
  INV_X1 U5596 ( .A(n4904), .ZN(n4903) );
  NAND2_X1 U5597 ( .A1(n4995), .A2(n5062), .ZN(n5137) );
  INV_X1 U5598 ( .A(n5138), .ZN(n4995) );
  NAND2_X1 U5599 ( .A1(n5161), .A2(n5125), .ZN(n4898) );
  INV_X1 U5600 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4598) );
  INV_X1 U5601 ( .A(n8900), .ZN(n8669) );
  AOI21_X1 U5602 ( .B1(n4488), .B2(n4721), .A(n4547), .ZN(n4718) );
  INV_X1 U5603 ( .A(n4722), .ZN(n4721) );
  NAND2_X1 U5604 ( .A1(n6325), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6343) );
  INV_X1 U5605 ( .A(n6327), .ZN(n6325) );
  NAND2_X1 U5606 ( .A1(n4713), .A2(n6232), .ZN(n4712) );
  INV_X1 U5607 ( .A(n4974), .ZN(n4713) );
  NAND2_X1 U5608 ( .A1(n8684), .A2(n8683), .ZN(n8682) );
  AND2_X1 U5609 ( .A1(n6154), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U5610 ( .A1(n6170), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6189) );
  INV_X1 U5611 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6077) );
  NOR2_X1 U5612 ( .A1(n6078), .A2(n6077), .ZN(n6102) );
  NOR2_X1 U5613 ( .A1(n6223), .A2(n6222), .ZN(n6265) );
  AND2_X1 U5614 ( .A1(n6265), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6267) );
  NAND2_X1 U5615 ( .A1(n6459), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6452) );
  OR2_X1 U5616 ( .A1(n4482), .A2(n7089), .ZN(n5977) );
  AOI21_X1 U5617 ( .B1(n9605), .B2(P2_REG2_REG_1__SCAN_IN), .A(n9601), .ZN(
        n9615) );
  OR2_X1 U5618 ( .A1(n7214), .A2(n7213), .ZN(n4848) );
  NAND2_X1 U5619 ( .A1(n8726), .A2(n8727), .ZN(n8725) );
  NOR2_X1 U5620 ( .A1(n7768), .A2(n4854), .ZN(n7771) );
  NOR2_X1 U5621 ( .A1(n7765), .A2(n7614), .ZN(n4854) );
  NAND2_X1 U5622 ( .A1(n7771), .A2(n7770), .ZN(n7825) );
  NAND2_X1 U5623 ( .A1(n7825), .A2(n4853), .ZN(n7827) );
  OR2_X1 U5624 ( .A1(n7826), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4853) );
  NAND2_X1 U5625 ( .A1(n7827), .A2(n7828), .ZN(n8005) );
  NOR2_X1 U5626 ( .A1(n4913), .A2(n4774), .ZN(n4911) );
  NAND2_X1 U5627 ( .A1(n8836), .A2(n8819), .ZN(n4914) );
  OAI21_X1 U5628 ( .B1(n8835), .B2(n5037), .A(n5036), .ZN(n8818) );
  OR2_X1 U5629 ( .A1(n8819), .A2(n8836), .ZN(n5037) );
  OR2_X1 U5630 ( .A1(n8819), .A2(n8565), .ZN(n5036) );
  INV_X1 U5631 ( .A(n4919), .ZN(n4918) );
  OAI21_X1 U5632 ( .B1(n8563), .B2(n4920), .A(n6540), .ZN(n4919) );
  OR2_X1 U5633 ( .A1(n8999), .A2(n8706), .ZN(n6540) );
  NAND2_X1 U5634 ( .A1(n8857), .A2(n8561), .ZN(n8835) );
  NOR2_X1 U5635 ( .A1(n8835), .A2(n8836), .ZN(n8834) );
  NOR2_X1 U5636 ( .A1(n8846), .A2(n8999), .ZN(n8829) );
  NAND2_X1 U5637 ( .A1(n8853), .A2(n6573), .ZN(n8857) );
  AND2_X1 U5638 ( .A1(n8844), .A2(n8556), .ZN(n6573) );
  INV_X1 U5639 ( .A(n8844), .ZN(n8854) );
  AND2_X1 U5640 ( .A1(n8560), .A2(n8561), .ZN(n8844) );
  OR2_X1 U5641 ( .A1(n6398), .A2(n6397), .ZN(n6414) );
  OAI21_X1 U5642 ( .B1(n6572), .B2(n5032), .A(n5030), .ZN(n8873) );
  AOI21_X1 U5643 ( .B1(n5035), .B2(n8903), .A(n5031), .ZN(n5030) );
  INV_X1 U5644 ( .A(n5035), .ZN(n5032) );
  INV_X1 U5645 ( .A(n8553), .ZN(n5031) );
  NAND2_X1 U5646 ( .A1(n8945), .A2(n4652), .ZN(n8867) );
  NOR2_X1 U5647 ( .A1(n9014), .A2(n4654), .ZN(n4652) );
  NOR2_X1 U5648 ( .A1(n8867), .A2(n9011), .ZN(n8866) );
  AND2_X1 U5649 ( .A1(n4646), .A2(n4645), .ZN(n8865) );
  NAND2_X1 U5650 ( .A1(n8889), .A2(n8669), .ZN(n4645) );
  NAND2_X1 U5651 ( .A1(n6356), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6372) );
  OR2_X1 U5652 ( .A1(n6372), .A2(n8651), .ZN(n6398) );
  AND2_X1 U5653 ( .A1(n4626), .A2(n4624), .ZN(n8904) );
  INV_X1 U5654 ( .A(n4625), .ZN(n4624) );
  OAI21_X1 U5655 ( .B1(n4628), .B2(n5029), .A(n4491), .ZN(n4625) );
  NOR2_X1 U5656 ( .A1(n9045), .A2(n4483), .ZN(n8973) );
  NAND2_X1 U5657 ( .A1(n4578), .A2(n8451), .ZN(n8965) );
  OAI21_X1 U5658 ( .B1(n7805), .B2(n5005), .A(n4489), .ZN(n4578) );
  NAND2_X1 U5659 ( .A1(n5004), .A2(n5007), .ZN(n5002) );
  OR2_X1 U5660 ( .A1(n6566), .A2(n5008), .ZN(n5007) );
  NAND2_X1 U5661 ( .A1(n7808), .A2(n6536), .ZN(n7875) );
  NOR2_X1 U5662 ( .A1(n7656), .A2(n4663), .ZN(n7876) );
  INV_X1 U5663 ( .A(n4665), .ZN(n4663) );
  NOR2_X1 U5664 ( .A1(n7656), .A2(n7841), .ZN(n7810) );
  OR2_X1 U5665 ( .A1(n6203), .A2(n7669), .ZN(n6223) );
  OR2_X1 U5666 ( .A1(n6189), .A2(n6188), .ZN(n6203) );
  AOI21_X1 U5667 ( .B1(n8506), .B2(n8601), .A(n4576), .ZN(n4575) );
  INV_X1 U5668 ( .A(n8511), .ZN(n4576) );
  NAND2_X1 U5669 ( .A1(n7627), .A2(n7628), .ZN(n7626) );
  NOR2_X1 U5670 ( .A1(n7478), .A2(n4662), .ZN(n7630) );
  OR2_X1 U5671 ( .A1(n6529), .A2(n7468), .ZN(n7454) );
  NAND2_X1 U5672 ( .A1(n4574), .A2(n4573), .ZN(n6562) );
  INV_X1 U5673 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6131) );
  AND2_X1 U5674 ( .A1(n8598), .A2(n7467), .ZN(n7468) );
  NOR2_X1 U5675 ( .A1(n7478), .A2(n4884), .ZN(n7477) );
  INV_X1 U5676 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6115) );
  OR2_X1 U5677 ( .A1(n6116), .A2(n6115), .ZN(n6132) );
  AND2_X1 U5678 ( .A1(n4616), .A2(n6527), .ZN(n4615) );
  AND2_X1 U5679 ( .A1(n4574), .A2(n8487), .ZN(n7405) );
  NAND2_X1 U5680 ( .A1(n5014), .A2(n5012), .ZN(n7101) );
  NAND2_X1 U5681 ( .A1(n5013), .A2(n8485), .ZN(n5012) );
  NAND2_X1 U5682 ( .A1(n5015), .A2(n8594), .ZN(n5013) );
  AND2_X1 U5683 ( .A1(n7230), .A2(n10057), .ZN(n7232) );
  NOR2_X1 U5684 ( .A1(n7133), .A2(n7069), .ZN(n7230) );
  AND2_X1 U5685 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6063) );
  NAND2_X1 U5686 ( .A1(n6063), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6078) );
  OR2_X1 U5687 ( .A1(n4670), .A2(n7136), .ZN(n7064) );
  AND2_X1 U5688 ( .A1(n4620), .A2(n6520), .ZN(n4619) );
  NAND2_X1 U5689 ( .A1(n8590), .A2(n4621), .ZN(n4620) );
  NAND2_X1 U5690 ( .A1(n8459), .A2(n7064), .ZN(n8591) );
  NAND2_X1 U5691 ( .A1(n8588), .A2(n7141), .ZN(n4622) );
  NAND2_X1 U5692 ( .A1(n7145), .A2(n8473), .ZN(n7272) );
  INV_X1 U5693 ( .A(n6555), .ZN(n8588) );
  NOR2_X1 U5694 ( .A1(n6601), .A2(n6588), .ZN(n6593) );
  NAND2_X1 U5695 ( .A1(n5958), .A2(n5957), .ZN(n5965) );
  INV_X1 U5696 ( .A(n5958), .ZN(n6464) );
  OR3_X1 U5697 ( .A1(n6459), .A2(P2_IR_REG_23__SCAN_IN), .A3(n6458), .ZN(n6462) );
  NOR2_X2 U5698 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6018) );
  NAND2_X1 U5699 ( .A1(n9102), .A2(n9101), .ZN(n9100) );
  AND2_X1 U5700 ( .A1(n5383), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U5701 ( .A1(n5336), .A2(n5337), .ZN(n7505) );
  NAND2_X1 U5702 ( .A1(n5412), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5443) );
  INV_X1 U5703 ( .A(n7967), .ZN(n4743) );
  NOR2_X1 U5704 ( .A1(n5352), .A2(n9810), .ZN(n5383) );
  OR2_X1 U5705 ( .A1(n5325), .A2(n5324), .ZN(n5352) );
  NAND2_X1 U5706 ( .A1(n9111), .A2(n5641), .ZN(n9153) );
  OR2_X1 U5707 ( .A1(n5443), .A2(n5442), .ZN(n5469) );
  NAND2_X1 U5708 ( .A1(n5706), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5735) );
  AOI21_X1 U5709 ( .B1(n4730), .B2(n4728), .A(n4726), .ZN(n4725) );
  NAND2_X1 U5710 ( .A1(n5336), .A2(n4728), .ZN(n4727) );
  INV_X1 U5711 ( .A(n9657), .ZN(n4726) );
  NAND2_X1 U5712 ( .A1(n5572), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5599) );
  OR2_X1 U5713 ( .A1(n6865), .A2(n8337), .ZN(n5938) );
  NOR2_X1 U5714 ( .A1(n8357), .A2(n8137), .ZN(n8326) );
  AOI21_X1 U5715 ( .B1(n4807), .B2(n4804), .A(n4800), .ZN(n8261) );
  AND2_X1 U5716 ( .A1(n4806), .A2(n4805), .ZN(n4804) );
  NAND2_X1 U5717 ( .A1(n4808), .A2(n8252), .ZN(n4807) );
  NAND2_X1 U5718 ( .A1(n4802), .A2(n4801), .ZN(n4800) );
  NAND2_X1 U5719 ( .A1(n5062), .A2(n4997), .ZN(n4996) );
  INV_X1 U5720 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4997) );
  OAI21_X1 U5721 ( .B1(n6879), .B2(n6878), .A(n6783), .ZN(n9765) );
  NAND2_X1 U5722 ( .A1(n9796), .A2(n9795), .ZN(n6830) );
  INV_X1 U5723 ( .A(n7493), .ZN(n7487) );
  NOR2_X1 U5724 ( .A1(n9824), .A2(n4755), .ZN(n6834) );
  AND2_X1 U5725 ( .A1(n9823), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4755) );
  NAND2_X1 U5726 ( .A1(n6834), .A2(n6835), .ZN(n7486) );
  NOR2_X1 U5727 ( .A1(n9853), .A2(n4759), .ZN(n9225) );
  AND2_X1 U5728 ( .A1(n9858), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4759) );
  INV_X1 U5729 ( .A(n5092), .ZN(n5489) );
  NOR2_X1 U5730 ( .A1(n9906), .A2(n9907), .ZN(n9908) );
  NAND2_X1 U5731 ( .A1(n4869), .A2(n9254), .ZN(n4868) );
  NAND2_X1 U5732 ( .A1(n9286), .A2(n9285), .ZN(n9284) );
  AND2_X1 U5733 ( .A1(n8413), .A2(n8245), .ZN(n9285) );
  INV_X1 U5734 ( .A(n4878), .ZN(n4877) );
  OAI21_X1 U5735 ( .B1(n4880), .B2(n4879), .A(n8409), .ZN(n4878) );
  OR2_X1 U5736 ( .A1(n9331), .A2(n9332), .ZN(n9333) );
  OR2_X1 U5737 ( .A1(n9509), .A2(n9147), .ZN(n8405) );
  NAND2_X1 U5738 ( .A1(n9419), .A2(n9568), .ZN(n9405) );
  NAND2_X1 U5739 ( .A1(n9419), .A2(n4786), .ZN(n9372) );
  AND2_X1 U5740 ( .A1(n8271), .A2(n9396), .ZN(n9433) );
  OR2_X1 U5741 ( .A1(n9382), .A2(n9449), .ZN(n9447) );
  AND2_X1 U5742 ( .A1(n9449), .A2(n8398), .ZN(n4875) );
  NAND2_X1 U5743 ( .A1(n4876), .A2(n8398), .ZN(n9439) );
  AND2_X1 U5744 ( .A1(n8398), .A2(n8202), .ZN(n9467) );
  AND2_X1 U5745 ( .A1(n9687), .A2(n4777), .ZN(n9470) );
  AND2_X1 U5746 ( .A1(n4487), .A2(n9584), .ZN(n4777) );
  NAND2_X1 U5747 ( .A1(n5494), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5522) );
  NOR2_X1 U5748 ( .A1(n7921), .A2(n5522), .ZN(n5547) );
  AOI21_X1 U5749 ( .B1(n4834), .B2(n4836), .A(n4512), .ZN(n4832) );
  NAND2_X1 U5750 ( .A1(n9699), .A2(n8191), .ZN(n7928) );
  NAND2_X1 U5751 ( .A1(n9687), .A2(n9723), .ZN(n9689) );
  AND2_X1 U5752 ( .A1(n7743), .A2(n9732), .ZN(n9687) );
  AND2_X1 U5753 ( .A1(n8184), .A2(n8179), .ZN(n8282) );
  OR2_X1 U5754 ( .A1(n7554), .A2(n7706), .ZN(n7715) );
  NOR2_X1 U5755 ( .A1(n7715), .A2(n9737), .ZN(n7743) );
  AND2_X1 U5756 ( .A1(n7856), .A2(n8083), .ZN(n8283) );
  AOI21_X1 U5757 ( .B1(n4827), .B2(n4490), .A(n4825), .ZN(n7525) );
  OAI21_X1 U5758 ( .B1(n7522), .B2(n4826), .A(n4517), .ZN(n4825) );
  NOR2_X1 U5759 ( .A1(n4873), .A2(n4872), .ZN(n4871) );
  INV_X1 U5760 ( .A(n8086), .ZN(n4873) );
  INV_X1 U5761 ( .A(n8147), .ZN(n4872) );
  NOR2_X1 U5762 ( .A1(n7439), .A2(n8165), .ZN(n7555) );
  NAND2_X1 U5763 ( .A1(n7434), .A2(n7433), .ZN(n7435) );
  NOR2_X1 U5764 ( .A1(n4776), .A2(n4775), .ZN(n7241) );
  NAND2_X1 U5765 ( .A1(n7250), .A2(n9945), .ZN(n4775) );
  NAND2_X1 U5766 ( .A1(n7350), .A2(n9945), .ZN(n7349) );
  NAND2_X1 U5767 ( .A1(n4812), .A2(n7195), .ZN(n8301) );
  NOR2_X1 U5768 ( .A1(n6854), .A2(n8067), .ZN(n7285) );
  NAND2_X1 U5769 ( .A1(n5814), .A2(n5813), .ZN(n9494) );
  NOR2_X1 U5770 ( .A1(n4841), .A2(n4840), .ZN(n7297) );
  INV_X1 U5771 ( .A(n7295), .ZN(n4840) );
  INV_X1 U5772 ( .A(n7296), .ZN(n4841) );
  OR2_X1 U5773 ( .A1(n7052), .A2(n8334), .ZN(n9986) );
  OR2_X1 U5774 ( .A1(n7052), .A2(n5918), .ZN(n9976) );
  AND3_X1 U5775 ( .A1(n6862), .A2(n7047), .A3(n6861), .ZN(n6980) );
  INV_X1 U5776 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5075) );
  OAI211_X1 U5777 ( .C1(n8128), .C2(n4936), .A(n4933), .B(n4935), .ZN(n9079)
         );
  NAND2_X1 U5778 ( .A1(n4950), .A2(n6545), .ZN(n8056) );
  NAND2_X1 U5779 ( .A1(n5865), .A2(n4557), .ZN(n4950) );
  XNOR2_X1 U5780 ( .A(n6542), .B(n6541), .ZN(n7950) );
  XNOR2_X1 U5781 ( .A(n5839), .B(n5838), .ZN(n7945) );
  XNOR2_X1 U5782 ( .A(n5808), .B(n5807), .ZN(n6393) );
  NAND2_X1 U5783 ( .A1(n4944), .A2(n5772), .ZN(n5808) );
  OAI21_X1 U5784 ( .B1(n5724), .B2(n5723), .A(n5722), .ZN(n5731) );
  AND2_X1 U5785 ( .A1(n5750), .A2(n5729), .ZN(n5730) );
  NAND2_X1 U5786 ( .A1(n4746), .A2(n4745), .ZN(n5097) );
  AOI21_X1 U5787 ( .B1(n4747), .B2(n4749), .A(n4749), .ZN(n4745) );
  INV_X1 U5788 ( .A(n4748), .ZN(n4747) );
  NAND2_X1 U5789 ( .A1(n4930), .A2(n5667), .ZN(n4614) );
  NAND2_X1 U5790 ( .A1(n4892), .A2(n5589), .ZN(n5616) );
  NAND2_X1 U5791 ( .A1(n5562), .A2(n4896), .ZN(n4892) );
  NAND2_X1 U5792 ( .A1(n5562), .A2(n5561), .ZN(n5591) );
  NAND2_X1 U5793 ( .A1(n4902), .A2(n5459), .ZN(n5485) );
  NAND2_X1 U5794 ( .A1(n4908), .A2(n4906), .ZN(n4902) );
  NAND2_X1 U5795 ( .A1(n4704), .A2(n4703), .ZN(n5396) );
  INV_X1 U5796 ( .A(n4707), .ZN(n4703) );
  XNOR2_X1 U5797 ( .A(n5367), .B(n5053), .ZN(n6127) );
  OAI21_X1 U5798 ( .B1(n5312), .B2(n4926), .A(n4924), .ZN(n5367) );
  NAND2_X1 U5799 ( .A1(n4929), .A2(n5314), .ZN(n5340) );
  NAND2_X1 U5800 ( .A1(n4606), .A2(n5251), .ZN(n5252) );
  NAND2_X1 U5801 ( .A1(n5248), .A2(n5249), .ZN(n4606) );
  NOR2_X1 U5802 ( .A1(n4981), .A2(n4980), .ZN(n7011) );
  INV_X1 U5803 ( .A(n6096), .ZN(n4980) );
  INV_X1 U5804 ( .A(n6097), .ZN(n4981) );
  INV_X1 U5805 ( .A(n4983), .ZN(n4982) );
  NAND2_X1 U5806 ( .A1(n4976), .A2(n6012), .ZN(n6914) );
  INV_X1 U5807 ( .A(n7136), .ZN(n10052) );
  NAND2_X1 U5808 ( .A1(n4956), .A2(n6036), .ZN(n6986) );
  INV_X1 U5809 ( .A(n6984), .ZN(n6056) );
  INV_X1 U5810 ( .A(n8723), .ZN(n6991) );
  NAND2_X1 U5811 ( .A1(n4716), .A2(n6214), .ZN(n7666) );
  NOR2_X1 U5812 ( .A1(n7360), .A2(n7359), .ZN(n4965) );
  AND2_X1 U5813 ( .A1(n7993), .A2(n6303), .ZN(n7911) );
  NAND2_X1 U5814 ( .A1(n6410), .A2(n6409), .ZN(n9005) );
  INV_X1 U5815 ( .A(n9628), .ZN(n8701) );
  INV_X1 U5816 ( .A(n9631), .ZN(n8698) );
  INV_X1 U5817 ( .A(n8712), .ZN(n7807) );
  OR2_X1 U5818 ( .A1(n9635), .A2(n8956), .ZN(n8686) );
  OR2_X1 U5819 ( .A1(n8441), .A2(n4567), .ZN(n4572) );
  AND2_X1 U5820 ( .A1(n4684), .A2(n4570), .ZN(n4569) );
  NAND2_X1 U5821 ( .A1(n8625), .A2(n8624), .ZN(n4684) );
  NAND2_X1 U5822 ( .A1(n4571), .A2(n4498), .ZN(n4570) );
  NAND2_X1 U5823 ( .A1(n6689), .A2(n10025), .ZN(n10019) );
  OR2_X1 U5824 ( .A1(n6037), .A2(n10008), .ZN(n6003) );
  OR2_X1 U5825 ( .A1(n4482), .A2(n7158), .ZN(n6006) );
  AND2_X1 U5826 ( .A1(n4856), .A2(n4855), .ZN(n6731) );
  NAND2_X1 U5827 ( .A1(n6732), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4855) );
  AND2_X1 U5828 ( .A1(n4850), .A2(n4849), .ZN(n6843) );
  NAND2_X1 U5829 ( .A1(n6844), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4849) );
  NOR2_X1 U5830 ( .A1(n6843), .A2(n6842), .ZN(n6949) );
  AOI21_X1 U5831 ( .B1(n7211), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7210), .ZN(
        n7214) );
  INV_X1 U5832 ( .A(n4848), .ZN(n7588) );
  NAND2_X1 U5833 ( .A1(n8725), .A2(n4844), .ZN(n7593) );
  NAND2_X1 U5834 ( .A1(n4846), .A2(n4845), .ZN(n4844) );
  INV_X1 U5835 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n4845) );
  INV_X1 U5836 ( .A(n8731), .ZN(n4846) );
  NOR2_X1 U5837 ( .A1(n8752), .A2(n8751), .ZN(n8755) );
  NOR2_X1 U5838 ( .A1(n8755), .A2(n8754), .ZN(n8766) );
  NAND2_X1 U5839 ( .A1(n4860), .A2(n4861), .ZN(n8770) );
  INV_X1 U5840 ( .A(n4859), .ZN(n4858) );
  OAI21_X1 U5841 ( .B1(n8799), .B2(n4597), .A(n8798), .ZN(n4864) );
  AND2_X1 U5842 ( .A1(n4932), .A2(n4565), .ZN(n8987) );
  AOI21_X1 U5843 ( .B1(n8432), .B2(n6547), .A(n8431), .ZN(n8992) );
  OR2_X1 U5844 ( .A1(n6604), .A2(n4476), .ZN(n6616) );
  AND2_X1 U5845 ( .A1(n4921), .A2(n4920), .ZN(n8828) );
  INV_X1 U5846 ( .A(n4646), .ZN(n8890) );
  NAND2_X1 U5847 ( .A1(n8896), .A2(n5035), .ZN(n8880) );
  AND2_X1 U5848 ( .A1(n8902), .A2(n8901), .ZN(n9023) );
  NAND2_X1 U5849 ( .A1(n8936), .A2(n8538), .ZN(n8923) );
  NAND2_X1 U5850 ( .A1(n8945), .A2(n8935), .ZN(n8917) );
  NAND2_X1 U5851 ( .A1(n4623), .A2(n4628), .ZN(n8914) );
  OR2_X1 U5852 ( .A1(n8944), .A2(n4630), .ZN(n4623) );
  NOR2_X1 U5853 ( .A1(n5026), .A2(n5028), .ZN(n8937) );
  AND2_X1 U5854 ( .A1(n4632), .A2(n4485), .ZN(n8931) );
  NAND2_X1 U5855 ( .A1(n8944), .A2(n8955), .ZN(n4632) );
  INV_X1 U5856 ( .A(n4761), .ZN(n8027) );
  AND2_X1 U5857 ( .A1(n7873), .A2(n4938), .ZN(n7955) );
  NAND2_X1 U5858 ( .A1(n7873), .A2(n6539), .ZN(n7953) );
  NAND2_X1 U5859 ( .A1(n5003), .A2(n8520), .ZN(n7869) );
  NAND2_X1 U5860 ( .A1(n6565), .A2(n6535), .ZN(n5003) );
  OAI211_X1 U5861 ( .C1(n4762), .C2(n4484), .A(n4635), .B(n6534), .ZN(n7809)
         );
  OR2_X1 U5862 ( .A1(n4764), .A2(n4484), .ZN(n4635) );
  NAND2_X1 U5863 ( .A1(n7652), .A2(n8454), .ZN(n7751) );
  NAND2_X1 U5864 ( .A1(n7648), .A2(n6533), .ZN(n7750) );
  NAND2_X1 U5865 ( .A1(n4764), .A2(n4767), .ZN(n7646) );
  NAND2_X1 U5866 ( .A1(n6532), .A2(n6531), .ZN(n7608) );
  AND2_X1 U5867 ( .A1(n4617), .A2(n4472), .ZN(n7100) );
  NAND2_X1 U5868 ( .A1(n7225), .A2(n7226), .ZN(n4617) );
  INV_X1 U5869 ( .A(n5011), .ZN(n7227) );
  OAI21_X1 U5870 ( .B1(n8456), .B2(n7062), .A(n5015), .ZN(n5011) );
  NAND2_X1 U5871 ( .A1(n4639), .A2(n9617), .ZN(n4638) );
  NAND2_X1 U5872 ( .A1(n4643), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4642) );
  NAND2_X1 U5873 ( .A1(n6068), .A2(n4641), .ZN(n4640) );
  NAND2_X1 U5874 ( .A1(n8877), .A2(n6608), .ZN(n8977) );
  NAND2_X1 U5875 ( .A1(n8877), .A2(n6618), .ZN(n8981) );
  INV_X1 U5876 ( .A(n8977), .ZN(n7963) );
  INV_X2 U5877 ( .A(n10096), .ZN(n10098) );
  OAI21_X1 U5878 ( .B1(n6619), .B2(n9054), .A(n6583), .ZN(n6594) );
  AND2_X1 U5879 ( .A1(n6604), .A2(n6582), .ZN(n6583) );
  AND2_X1 U5880 ( .A1(n8996), .A2(n8995), .ZN(n8997) );
  AOI21_X1 U5881 ( .B1(n7561), .B2(n10035), .A(n4566), .ZN(n7562) );
  AND2_X1 U5882 ( .A1(n6663), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10025) );
  AND2_X1 U5883 ( .A1(n4527), .A2(n5966), .ZN(n5038) );
  XNOR2_X1 U5884 ( .A(n6454), .B(P2_IR_REG_24__SCAN_IN), .ZN(n7844) );
  NAND2_X1 U5885 ( .A1(n5990), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5992) );
  CLKBUF_X1 U5886 ( .A(n6487), .Z(n8618) );
  INV_X1 U5887 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7002) );
  INV_X1 U5888 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6948) );
  INV_X1 U5889 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6905) );
  INV_X1 U5890 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6812) );
  AND2_X1 U5891 ( .A1(n6151), .A2(n6166), .ZN(n7589) );
  INV_X1 U5892 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6662) );
  NAND2_X1 U5893 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4862) );
  INV_X1 U5894 ( .A(n5859), .ZN(n9094) );
  NAND2_X1 U5895 ( .A1(n5493), .A2(n5492), .ZN(n8082) );
  NAND2_X1 U5896 ( .A1(n4994), .A2(n5366), .ZN(n7541) );
  NAND2_X1 U5897 ( .A1(n5859), .A2(n5858), .ZN(n5916) );
  OR2_X1 U5898 ( .A1(n5001), .A2(n9091), .ZN(n4999) );
  AND2_X1 U5899 ( .A1(n5832), .A2(n9092), .ZN(n5001) );
  OR2_X1 U5900 ( .A1(n5336), .A2(n5337), .ZN(n7507) );
  NAND2_X1 U5901 ( .A1(n6867), .A2(n5186), .ZN(n6930) );
  AND2_X1 U5902 ( .A1(n4741), .A2(n4506), .ZN(n7785) );
  NAND2_X1 U5903 ( .A1(n7916), .A2(n7920), .ZN(n7970) );
  NAND2_X1 U5904 ( .A1(n5546), .A2(n5545), .ZN(n8372) );
  OR2_X1 U5905 ( .A1(n5336), .A2(n4730), .ZN(n4724) );
  NAND2_X1 U5906 ( .A1(n7784), .A2(n5458), .ZN(n7797) );
  NAND2_X1 U5907 ( .A1(n4583), .A2(n5720), .ZN(n9163) );
  NAND2_X1 U5908 ( .A1(n4580), .A2(n5721), .ZN(n9164) );
  INV_X1 U5909 ( .A(n4583), .ZN(n4580) );
  INV_X1 U5910 ( .A(n9193), .ZN(n9655) );
  AND2_X1 U5911 ( .A1(n7374), .A2(n5280), .ZN(n5281) );
  OR2_X1 U5912 ( .A1(n7115), .A2(n7114), .ZN(n5280) );
  AND2_X1 U5913 ( .A1(n9659), .A2(n9959), .ZN(n9170) );
  NAND2_X1 U5914 ( .A1(n4586), .A2(n4585), .ZN(n9188) );
  INV_X1 U5915 ( .A(n9187), .ZN(n4585) );
  INV_X1 U5916 ( .A(n9185), .ZN(n4586) );
  NAND2_X1 U5917 ( .A1(n7919), .A2(n7918), .ZN(n7916) );
  INV_X1 U5918 ( .A(n9186), .ZN(n9660) );
  INV_X1 U5919 ( .A(n9665), .ZN(n9191) );
  NAND2_X1 U5920 ( .A1(n5851), .A2(n5850), .ZN(n9304) );
  OR2_X1 U5921 ( .A1(n9315), .A2(n5928), .ZN(n5787) );
  NAND4_X1 U5922 ( .A1(n5089), .A2(n5088), .A3(n5087), .A4(n5086), .ZN(n9212)
         );
  NAND2_X1 U5923 ( .A1(n5845), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5159) );
  NAND2_X1 U5924 ( .A1(n5210), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5158) );
  NAND2_X1 U5925 ( .A1(n9217), .A2(n9216), .ZN(n9215) );
  NAND2_X1 U5926 ( .A1(n6804), .A2(n6805), .ZN(n6803) );
  NOR2_X1 U5927 ( .A1(n9779), .A2(n4545), .ZN(n6790) );
  NAND2_X1 U5928 ( .A1(n6790), .A2(n6791), .ZN(n6828) );
  NAND2_X1 U5929 ( .A1(n6828), .A2(n4750), .ZN(n9796) );
  OR2_X1 U5930 ( .A1(n6829), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4750) );
  NOR2_X1 U5931 ( .A1(n9840), .A2(n4550), .ZN(n9855) );
  XNOR2_X1 U5932 ( .A(n9225), .B(n7496), .ZN(n7489) );
  XNOR2_X1 U5933 ( .A(n4752), .B(n9232), .ZN(n9247) );
  OR2_X1 U5934 ( .A1(n9908), .A2(n4753), .ZN(n4752) );
  AND2_X1 U5935 ( .A1(n9233), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4753) );
  NOR2_X1 U5936 ( .A1(n9295), .A2(n4790), .ZN(n8358) );
  NAND2_X1 U5937 ( .A1(n9326), .A2(n8407), .ZN(n9319) );
  AND2_X1 U5938 ( .A1(n9354), .A2(n9353), .ZN(n9512) );
  NAND2_X1 U5939 ( .A1(n4817), .A2(n4821), .ZN(n9359) );
  INV_X1 U5940 ( .A(n4820), .ZN(n4821) );
  NAND2_X1 U5941 ( .A1(n9468), .A2(n4823), .ZN(n4817) );
  NAND2_X1 U5942 ( .A1(n7853), .A2(n7852), .ZN(n9686) );
  NAND2_X1 U5943 ( .A1(n7523), .A2(n7522), .ZN(n7553) );
  NAND2_X1 U5944 ( .A1(n7384), .A2(n7383), .ZN(n7426) );
  INV_X1 U5945 ( .A(n7246), .ZN(n7294) );
  INV_X1 U5946 ( .A(n4828), .ZN(n4830) );
  NAND2_X1 U5947 ( .A1(n5192), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4781) );
  INV_X1 U5948 ( .A(n9475), .ZN(n9713) );
  AOI22_X1 U5949 ( .A1(n9079), .A2(n8132), .B1(n8131), .B2(
        P2_DATAO_REG_31__SCAN_IN), .ZN(n8369) );
  OAI21_X1 U5950 ( .B1(n9484), .B2(n9970), .A(n4842), .ZN(n9552) );
  AND2_X1 U5951 ( .A1(n9487), .A2(n9488), .ZN(n4842) );
  NAND2_X1 U5952 ( .A1(n5104), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5102) );
  OR2_X1 U5953 ( .A1(n5103), .A2(n5101), .ZN(n5105) );
  INV_X1 U5954 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7358) );
  NAND2_X1 U5955 ( .A1(n5148), .A2(n5151), .ZN(n9430) );
  AND2_X1 U5956 ( .A1(n5592), .A2(n5569), .ZN(n9234) );
  INV_X1 U5957 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7003) );
  INV_X1 U5958 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6946) );
  INV_X1 U5959 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6903) );
  INV_X1 U5960 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6813) );
  XNOR2_X1 U5961 ( .A(n4751), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9214) );
  NAND2_X1 U5962 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4751) );
  AND2_X1 U5963 ( .A1(n8993), .A2(n9628), .ZN(n4973) );
  INV_X1 U5964 ( .A(n4856), .ZN(n6728) );
  INV_X1 U5965 ( .A(n4852), .ZN(n6745) );
  OAI21_X1 U5966 ( .B1(n8797), .B2(n6304), .A(n4863), .ZN(P2_U3264) );
  AOI21_X1 U5967 ( .B1(n4865), .B2(n6304), .A(n4864), .ZN(n4863) );
  NOR2_X1 U5968 ( .A1(n7271), .A2(n4648), .ZN(n7278) );
  INV_X1 U5969 ( .A(n4658), .ZN(n9064) );
  NAND2_X1 U5970 ( .A1(n10084), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n4657) );
  MUX2_X1 U5971 ( .A(n8336), .B(n8335), .S(n8334), .Z(n8343) );
  NAND2_X1 U5972 ( .A1(n9990), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n4599) );
  NAND2_X1 U5973 ( .A1(n8423), .A2(n9992), .ZN(n4600) );
  NAND2_X1 U5974 ( .A1(n6130), .A2(n6129), .ZN(n4884) );
  OR3_X1 U5975 ( .A1(n7656), .A2(n4664), .A3(n9051), .ZN(n4483) );
  OAI21_X1 U5976 ( .B1(n9468), .B2(n4501), .A(n8375), .ZN(n9382) );
  NAND2_X1 U5977 ( .A1(n5118), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4696) );
  OR2_X1 U5978 ( .A1(n5018), .A2(n4637), .ZN(n4484) );
  NAND2_X1 U5979 ( .A1(n9035), .A2(n8939), .ZN(n4485) );
  INV_X1 U5980 ( .A(n7650), .ZN(n6564) );
  XNOR2_X1 U5981 ( .A(n8993), .B(n8838), .ZN(n8819) );
  INV_X1 U5982 ( .A(n8819), .ZN(n8810) );
  AND2_X1 U5983 ( .A1(n8303), .A2(n8074), .ZN(n4486) );
  AND2_X1 U5984 ( .A1(n4779), .A2(n4778), .ZN(n4487) );
  OAI21_X1 U5985 ( .B1(n8668), .B2(n8666), .A(n8665), .ZN(n8693) );
  AND2_X1 U5986 ( .A1(n4957), .A2(n4719), .ZN(n4488) );
  AOI21_X1 U5987 ( .B1(n9200), .B2(n8263), .A(n8369), .ZN(n8300) );
  INV_X1 U5988 ( .A(n8300), .ZN(n4806) );
  AND2_X1 U5989 ( .A1(n5002), .A2(n8607), .ZN(n4489) );
  AND2_X1 U5990 ( .A1(n7431), .A2(n7524), .ZN(n4490) );
  NAND2_X1 U5991 ( .A1(n5734), .A2(n5733), .ZN(n9509) );
  INV_X1 U5992 ( .A(n8590), .ZN(n8467) );
  INV_X1 U5993 ( .A(n9014), .ZN(n8889) );
  NAND2_X1 U5994 ( .A1(n6354), .A2(n6353), .ZN(n9025) );
  AND2_X1 U5995 ( .A1(n5246), .A2(n5245), .ZN(n6784) );
  OR2_X1 U5996 ( .A1(n8938), .A2(n9025), .ZN(n4491) );
  OR2_X1 U5997 ( .A1(n4914), .A2(n4916), .ZN(n4492) );
  NAND2_X1 U5998 ( .A1(n6526), .A2(n4472), .ZN(n4493) );
  AOI22_X1 U5999 ( .A1(n8432), .A2(n8132), .B1(n8131), .B2(
        P2_DATAO_REG_30__SCAN_IN), .ZN(n8356) );
  NOR2_X1 U6000 ( .A1(n8935), .A2(n8959), .ZN(n4494) );
  INV_X1 U6001 ( .A(n8705), .ZN(n8838) );
  NAND2_X1 U6002 ( .A1(n9687), .A2(n4487), .ZN(n4495) );
  NAND2_X1 U6003 ( .A1(n4562), .A2(n6545), .ZN(n4949) );
  AND2_X1 U6004 ( .A1(n8801), .A2(n4565), .ZN(n4496) );
  NOR2_X1 U6005 ( .A1(n7327), .A2(n4564), .ZN(n4497) );
  AND2_X1 U6006 ( .A1(n6491), .A2(n8620), .ZN(n4498) );
  NAND4_X1 U6007 ( .A1(n5173), .A2(n5172), .A3(n5171), .A4(n5170), .ZN(n6854)
         );
  INV_X1 U6008 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10015) );
  INV_X1 U6009 ( .A(n6517), .ZN(n7273) );
  NAND2_X1 U6010 ( .A1(n8873), .A2(n8872), .ZN(n8853) );
  NAND2_X2 U6011 ( .A1(n5972), .A2(n9089), .ZN(n6037) );
  INV_X1 U6012 ( .A(n4991), .ZN(n4990) );
  NAND2_X1 U6013 ( .A1(n5686), .A2(n4992), .ZN(n4991) );
  AND2_X1 U6014 ( .A1(n6031), .A2(n4650), .ZN(n6519) );
  INV_X1 U6015 ( .A(n8722), .ZN(n4670) );
  NOR2_X1 U6016 ( .A1(n6643), .A2(n6030), .ZN(n4499) );
  AND2_X1 U6017 ( .A1(n8143), .A2(n7295), .ZN(n4500) );
  AND2_X1 U6018 ( .A1(n9474), .A2(n9443), .ZN(n4501) );
  INV_X1 U6019 ( .A(n5425), .ZN(n5429) );
  XNOR2_X1 U6020 ( .A(n5426), .B(SI_11_), .ZN(n5425) );
  INV_X1 U6021 ( .A(n4884), .ZN(n7479) );
  NAND4_X1 U6022 ( .A1(n5977), .A2(n5976), .A3(n5975), .A4(n5974), .ZN(n6512)
         );
  XNOR2_X1 U6023 ( .A(n9011), .B(n8882), .ZN(n8872) );
  INV_X1 U6024 ( .A(n8520), .ZN(n5008) );
  OR2_X1 U6025 ( .A1(n9295), .A2(n4789), .ZN(n4502) );
  XNOR2_X1 U6026 ( .A(n8999), .B(n8821), .ZN(n8836) );
  INV_X1 U6027 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9081) );
  INV_X1 U6028 ( .A(n8454), .ZN(n5023) );
  NAND2_X1 U6029 ( .A1(n6341), .A2(n6340), .ZN(n9030) );
  OR2_X1 U6030 ( .A1(n8485), .A2(n8580), .ZN(n4503) );
  OR3_X1 U6031 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4504) );
  AND2_X1 U6032 ( .A1(n8300), .A2(n8258), .ZN(n4505) );
  NAND2_X1 U6033 ( .A1(n5424), .A2(n5423), .ZN(n4506) );
  AND2_X1 U6034 ( .A1(n4525), .A2(n5075), .ZN(n4507) );
  NAND2_X1 U6035 ( .A1(n8445), .A2(n8549), .ZN(n8903) );
  NOR2_X1 U6036 ( .A1(n8607), .A2(n4939), .ZN(n4938) );
  AND2_X1 U6037 ( .A1(n8505), .A2(n8498), .ZN(n7628) );
  INV_X1 U6038 ( .A(n7628), .ZN(n8601) );
  OR2_X1 U6039 ( .A1(n9489), .A2(n8065), .ZN(n8413) );
  INV_X1 U6040 ( .A(n8420), .ZN(n9275) );
  NAND2_X1 U6041 ( .A1(n5868), .A2(n5867), .ZN(n8420) );
  INV_X1 U6042 ( .A(n8993), .ZN(n8817) );
  NAND2_X1 U6043 ( .A1(n5964), .A2(n5963), .ZN(n8993) );
  AND2_X1 U6044 ( .A1(n8935), .A2(n8959), .ZN(n4508) );
  NAND2_X1 U6045 ( .A1(n6264), .A2(n6263), .ZN(n7815) );
  AND2_X1 U6046 ( .A1(n8272), .A2(n8399), .ZN(n9449) );
  INV_X1 U6047 ( .A(n8522), .ZN(n6537) );
  AND2_X1 U6048 ( .A1(n8453), .A2(n8452), .ZN(n8522) );
  AND2_X1 U6049 ( .A1(n9284), .A2(n4870), .ZN(n4509) );
  INV_X1 U6050 ( .A(n5053), .ZN(n4711) );
  AND3_X1 U6051 ( .A1(n8193), .A2(n8192), .A3(n8191), .ZN(n4510) );
  AND2_X1 U6052 ( .A1(n4600), .A2(n4599), .ZN(n4511) );
  AND2_X1 U6053 ( .A1(n9712), .A2(n9204), .ZN(n4512) );
  NOR2_X1 U6054 ( .A1(n9494), .A2(n9287), .ZN(n4513) );
  INV_X1 U6055 ( .A(n8419), .ZN(n9281) );
  NOR2_X1 U6056 ( .A1(n9295), .A2(n9489), .ZN(n8419) );
  AND2_X1 U6057 ( .A1(n6564), .A2(n8512), .ZN(n4514) );
  INV_X1 U6058 ( .A(n4913), .ZN(n4912) );
  OAI21_X1 U6059 ( .B1(n4918), .B2(n8810), .A(n4524), .ZN(n4913) );
  AND2_X1 U6060 ( .A1(n4636), .A2(n8606), .ZN(n4515) );
  NOR2_X1 U6061 ( .A1(n5694), .A2(n5693), .ZN(n4516) );
  NAND2_X1 U6062 ( .A1(n8166), .A2(n9207), .ZN(n4517) );
  INV_X1 U6063 ( .A(n5337), .ZN(n4729) );
  NAND2_X1 U6064 ( .A1(n6692), .A2(n4481), .ZN(n6030) );
  INV_X1 U6065 ( .A(n6030), .ZN(n6068) );
  AND2_X1 U6066 ( .A1(n4858), .A2(n4861), .ZN(n4518) );
  XNOR2_X1 U6067 ( .A(n5313), .B(SI_7_), .ZN(n5310) );
  INV_X1 U6068 ( .A(n5005), .ZN(n5004) );
  OAI21_X1 U6069 ( .B1(n6566), .B2(n5006), .A(n8453), .ZN(n5005) );
  AND2_X1 U6070 ( .A1(n6530), .A2(n7457), .ZN(n4519) );
  NAND2_X1 U6071 ( .A1(n5425), .A2(n4900), .ZN(n4520) );
  INV_X1 U6072 ( .A(n4654), .ZN(n4653) );
  NAND2_X1 U6073 ( .A1(n4656), .A2(n4655), .ZN(n4654) );
  INV_X1 U6074 ( .A(n4784), .ZN(n4783) );
  NAND2_X1 U6075 ( .A1(n4786), .A2(n4785), .ZN(n4784) );
  INV_X1 U6076 ( .A(n4916), .ZN(n4915) );
  NAND2_X1 U6077 ( .A1(n8854), .A2(n4917), .ZN(n4916) );
  AND2_X1 U6078 ( .A1(n5271), .A2(SI_5_), .ZN(n4521) );
  AND2_X1 U6079 ( .A1(n5048), .A2(n5049), .ZN(n4522) );
  AND2_X1 U6080 ( .A1(n8249), .A2(n9254), .ZN(n8414) );
  INV_X1 U6081 ( .A(n4631), .ZN(n4630) );
  NOR2_X1 U6082 ( .A1(n4494), .A2(n4633), .ZN(n4631) );
  NAND2_X1 U6083 ( .A1(n4693), .A2(n4689), .ZN(n4523) );
  OR2_X1 U6084 ( .A1(n8993), .A2(n8705), .ZN(n4524) );
  INV_X1 U6085 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4749) );
  INV_X1 U6086 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5968) );
  AND2_X1 U6087 ( .A1(n4522), .A2(n5074), .ZN(n4525) );
  AND2_X1 U6088 ( .A1(n8810), .A2(n8567), .ZN(n4526) );
  AND2_X1 U6089 ( .A1(n5957), .A2(n5959), .ZN(n4527) );
  INV_X1 U6090 ( .A(n8408), .ZN(n9318) );
  AND2_X1 U6091 ( .A1(n8409), .A2(n8265), .ZN(n8408) );
  AND2_X1 U6092 ( .A1(n9514), .A2(n9351), .ZN(n4528) );
  INV_X1 U6093 ( .A(n8506), .ZN(n4577) );
  OR2_X1 U6094 ( .A1(n6320), .A2(n7994), .ZN(n4529) );
  AND2_X1 U6095 ( .A1(n8481), .A2(n8485), .ZN(n8594) );
  AND2_X1 U6096 ( .A1(n7859), .A2(n8097), .ZN(n4530) );
  AND2_X1 U6097 ( .A1(n8303), .A2(n7195), .ZN(n4531) );
  AND2_X1 U6098 ( .A1(n9254), .A2(n9285), .ZN(n4532) );
  AND2_X1 U6099 ( .A1(n9348), .A2(n8405), .ZN(n4533) );
  AND2_X1 U6100 ( .A1(n4591), .A2(n4737), .ZN(n4534) );
  AND2_X1 U6101 ( .A1(n5057), .A2(n5366), .ZN(n4535) );
  AND2_X1 U6102 ( .A1(n4572), .A2(n4569), .ZN(n4536) );
  AND2_X1 U6103 ( .A1(n4526), .A2(n4686), .ZN(n4537) );
  AND2_X1 U6104 ( .A1(n4675), .A2(n4672), .ZN(n4538) );
  INV_X1 U6105 ( .A(n6165), .ZN(n4964) );
  OR2_X1 U6106 ( .A1(n4903), .A2(n4901), .ZN(n4539) );
  AND2_X1 U6107 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4540) );
  INV_X1 U6108 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5904) );
  INV_X1 U6109 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6660) );
  INV_X1 U6110 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5093) );
  AND2_X1 U6111 ( .A1(n8945), .A2(n4653), .ZN(n4541) );
  INV_X1 U6112 ( .A(n8708), .ZN(n8959) );
  NAND2_X1 U6113 ( .A1(n6371), .A2(n6370), .ZN(n9020) );
  INV_X1 U6114 ( .A(n9020), .ZN(n4655) );
  AND2_X1 U6115 ( .A1(n8892), .A2(n8549), .ZN(n5035) );
  AND2_X1 U6116 ( .A1(n9687), .A2(n4779), .ZN(n4542) );
  INV_X1 U6117 ( .A(n8938), .ZN(n8660) );
  OR2_X1 U6118 ( .A1(n5807), .A2(n4943), .ZN(n4543) );
  OR2_X1 U6119 ( .A1(n8039), .A2(n8957), .ZN(n4544) );
  XNOR2_X1 U6120 ( .A(n5102), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5886) );
  INV_X1 U6121 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4596) );
  AND2_X1 U6122 ( .A1(n6789), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4545) );
  NAND2_X1 U6123 ( .A1(n5841), .A2(n5840), .ZN(n9489) );
  INV_X1 U6124 ( .A(n9489), .ZN(n4791) );
  INV_X1 U6125 ( .A(n9329), .ZN(n8406) );
  INV_X1 U6126 ( .A(n8665), .ZN(n4720) );
  NAND2_X1 U6127 ( .A1(n6395), .A2(n6394), .ZN(n9011) );
  INV_X1 U6128 ( .A(n9011), .ZN(n4923) );
  AND2_X1 U6129 ( .A1(n6747), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4546) );
  OAI21_X1 U6130 ( .B1(n7627), .B2(n4577), .A(n4575), .ZN(n7649) );
  NAND2_X1 U6131 ( .A1(n8926), .A2(n8546), .ZN(n8897) );
  NAND2_X1 U6132 ( .A1(n8951), .A2(n6569), .ZN(n8952) );
  INV_X1 U6133 ( .A(n8952), .ZN(n5026) );
  AND2_X1 U6134 ( .A1(n6437), .A2(n6436), .ZN(n4547) );
  NAND2_X1 U6135 ( .A1(n6572), .A2(n6571), .ZN(n8896) );
  INV_X1 U6136 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5101) );
  OR2_X1 U6137 ( .A1(n9275), .A2(n9253), .ZN(n4548) );
  AND2_X1 U6138 ( .A1(n9045), .A2(n8709), .ZN(n4549) );
  NAND2_X1 U6139 ( .A1(n9419), .A2(n4783), .ZN(n4787) );
  NAND2_X1 U6140 ( .A1(n4923), .A2(n8695), .ZN(n4922) );
  INV_X1 U6141 ( .A(n4922), .ZN(n4774) );
  AND2_X1 U6142 ( .A1(n9845), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4550) );
  AND3_X1 U6143 ( .A1(n6510), .A2(n6509), .A3(n6508), .ZN(n4551) );
  AND2_X1 U6144 ( .A1(n5617), .A2(SI_18_), .ZN(n4552) );
  AND2_X1 U6145 ( .A1(n5695), .A2(n5667), .ZN(n4553) );
  OR2_X1 U6146 ( .A1(n9275), .A2(n9551), .ZN(n4554) );
  INV_X1 U6147 ( .A(n4485), .ZN(n4633) );
  NOR2_X1 U6148 ( .A1(n9709), .A2(n8139), .ZN(n4555) );
  NAND2_X1 U6149 ( .A1(n7740), .A2(n7739), .ZN(n7853) );
  INV_X1 U6150 ( .A(n9992), .ZN(n9990) );
  NAND2_X1 U6151 ( .A1(n6556), .A2(n8458), .ZN(n7062) );
  NOR2_X1 U6152 ( .A1(n7478), .A2(n4660), .ZN(n4556) );
  AND2_X1 U6153 ( .A1(n6541), .A2(n5864), .ZN(n4557) );
  OAI21_X1 U6154 ( .B1(n7388), .B2(n8275), .A(n8066), .ZN(n7434) );
  NAND2_X1 U6155 ( .A1(n4588), .A2(n5395), .ZN(n7637) );
  NAND2_X1 U6156 ( .A1(n4724), .A2(n4728), .ZN(n9656) );
  NAND2_X1 U6157 ( .A1(n7435), .A2(n8147), .ZN(n7526) );
  NAND2_X1 U6158 ( .A1(n4622), .A2(n6518), .ZN(n7266) );
  OR2_X1 U6159 ( .A1(n5490), .A2(n5092), .ZN(n9238) );
  NAND2_X1 U6160 ( .A1(n5705), .A2(n5704), .ZN(n9514) );
  INV_X1 U6161 ( .A(n9514), .ZN(n4785) );
  NAND2_X1 U6162 ( .A1(n5521), .A2(n5520), .ZN(n9682) );
  INV_X1 U6163 ( .A(n9682), .ZN(n4778) );
  OAI21_X1 U6164 ( .B1(n4962), .B2(n4963), .A(n4959), .ZN(n7664) );
  OR2_X1 U6165 ( .A1(n4965), .A2(n4964), .ZN(n4558) );
  NAND2_X1 U6166 ( .A1(n4741), .A2(n4740), .ZN(n7784) );
  NAND2_X1 U6167 ( .A1(n7376), .A2(n5286), .ZN(n7174) );
  AND2_X1 U6168 ( .A1(n7505), .A2(n7504), .ZN(n4559) );
  AND2_X1 U6169 ( .A1(n7666), .A2(n4974), .ZN(n4560) );
  OR2_X1 U6170 ( .A1(n7656), .A2(n4664), .ZN(n4561) );
  INV_X1 U6171 ( .A(n8456), .ZN(n6557) );
  OR2_X1 U6172 ( .A1(n8054), .A2(SI_29_), .ZN(n4562) );
  NOR2_X1 U6173 ( .A1(n4831), .A2(n4830), .ZN(n4563) );
  OR2_X1 U6174 ( .A1(n7328), .A2(n4883), .ZN(n4564) );
  INV_X2 U6175 ( .A(n10084), .ZN(n10086) );
  OR2_X1 U6176 ( .A1(n8436), .A2(n9082), .ZN(n4565) );
  AND2_X1 U6177 ( .A1(n4884), .A2(n9058), .ZN(n4566) );
  INV_X1 U6178 ( .A(n6581), .ZN(n6513) );
  OAI211_X1 U6179 ( .C1(n6058), .C2(n6632), .A(n4773), .B(n4772), .ZN(n6581)
         );
  NAND2_X1 U6180 ( .A1(n6036), .A2(n6035), .ZN(n6983) );
  INV_X1 U6181 ( .A(n4776), .ZN(n7350) );
  AND2_X1 U6182 ( .A1(n10078), .A2(n8442), .ZN(n4567) );
  AND2_X1 U6183 ( .A1(n5181), .A2(n5180), .ZN(n4568) );
  INV_X1 U6184 ( .A(n6491), .ZN(n10027) );
  NAND2_X1 U6185 ( .A1(n7622), .A2(n8443), .ZN(n6491) );
  INV_X1 U6186 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n4757) );
  NAND2_X1 U6187 ( .A1(n4609), .A2(n5512), .ZN(n5539) );
  NAND2_X4 U6188 ( .A1(n5669), .A2(n5668), .ZN(n9519) );
  NAND2_X1 U6189 ( .A1(n5666), .A2(n5665), .ZN(n4930) );
  MUX2_X2 U6190 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n8423), .S(n10004), .Z(n8424) );
  NAND2_X1 U6191 ( .A1(n4611), .A2(n4539), .ZN(n4610) );
  AOI21_X1 U6192 ( .B1(n4818), .B2(n4820), .A(n4528), .ZN(n4816) );
  NAND2_X1 U6193 ( .A1(n8422), .A2(n4602), .ZN(n4601) );
  NAND2_X1 U6194 ( .A1(n4597), .A2(n4598), .ZN(n4592) );
  INV_X1 U6195 ( .A(n5314), .ZN(n4928) );
  OAI21_X1 U6196 ( .B1(n4823), .B2(n4820), .A(n8386), .ZN(n4819) );
  INV_X1 U6197 ( .A(n7405), .ZN(n7404) );
  NAND2_X1 U6198 ( .A1(n4579), .A2(n7901), .ZN(n5534) );
  NAND2_X1 U6199 ( .A1(n5533), .A2(n4579), .ZN(n7900) );
  OAI21_X2 U6200 ( .B1(n4583), .B2(n4582), .A(n4581), .ZN(n5748) );
  NAND2_X1 U6201 ( .A1(n4731), .A2(n4734), .ZN(n4583) );
  OR2_X2 U6202 ( .A1(n5916), .A2(n5915), .ZN(n5943) );
  XNOR2_X1 U6203 ( .A(n4587), .B(n6967), .ZN(n6972) );
  NAND2_X1 U6204 ( .A1(n5231), .A2(n5230), .ZN(n4587) );
  NAND2_X2 U6205 ( .A1(n5613), .A2(n5612), .ZN(n9176) );
  OAI21_X2 U6206 ( .B1(n9136), .B2(n9135), .A(n5586), .ZN(n5613) );
  NAND2_X1 U6207 ( .A1(n4994), .A2(n4535), .ZN(n4588) );
  NAND2_X1 U6208 ( .A1(n4534), .A2(n7637), .ZN(n4590) );
  NAND3_X1 U6209 ( .A1(n4590), .A2(n7795), .A3(n4589), .ZN(n5508) );
  NAND3_X1 U6210 ( .A1(n4591), .A2(n4737), .A3(n4739), .ZN(n4589) );
  NAND4_X1 U6211 ( .A1(n5071), .A2(n5244), .A3(n5067), .A4(n5904), .ZN(n5106)
         );
  INV_X4 U6212 ( .A(n4481), .ZN(n6633) );
  NAND3_X1 U6213 ( .A1(n4697), .A2(n4696), .A3(P2_DATAO_REG_4__SCAN_IN), .ZN(
        n4593) );
  OR2_X2 U6214 ( .A1(n9277), .A2(n4601), .ZN(n8423) );
  NAND2_X1 U6215 ( .A1(n8418), .A2(n8417), .ZN(n9277) );
  OAI21_X2 U6216 ( .B1(n7928), .B2(n8285), .A(n8194), .ZN(n9667) );
  NAND2_X1 U6217 ( .A1(n8425), .A2(n4554), .ZN(P1_U3551) );
  NAND2_X2 U6218 ( .A1(n8269), .A2(n9364), .ZN(n9387) );
  NAND2_X2 U6219 ( .A1(n9519), .A2(n8078), .ZN(n9364) );
  INV_X1 U6220 ( .A(n4610), .ZN(n5513) );
  NAND2_X1 U6221 ( .A1(n4610), .A2(n5509), .ZN(n4609) );
  OAI21_X1 U6222 ( .B1(n4481), .B2(P2_DATAO_REG_8__SCAN_IN), .A(n4613), .ZN(
        n5316) );
  NAND2_X1 U6223 ( .A1(n4481), .A2(n6662), .ZN(n4613) );
  OAI21_X1 U6224 ( .B1(n4493), .B2(n7225), .A(n4615), .ZN(n7401) );
  NAND3_X1 U6225 ( .A1(n6526), .A2(n4472), .A3(n8594), .ZN(n4616) );
  OAI21_X1 U6226 ( .B1(n8467), .B2(n4622), .A(n4619), .ZN(n7137) );
  OR2_X1 U6227 ( .A1(n8944), .A2(n4627), .ZN(n4626) );
  NAND3_X1 U6228 ( .A1(n4764), .A2(n6534), .A3(n4762), .ZN(n4634) );
  NAND2_X1 U6229 ( .A1(n4764), .A2(n4762), .ZN(n7648) );
  AND3_X2 U6230 ( .A1(n4642), .A2(n4640), .A3(n4638), .ZN(n10037) );
  XNOR2_X1 U6231 ( .A(n6519), .B(n5997), .ZN(n6033) );
  INV_X1 U6232 ( .A(n6519), .ZN(n4649) );
  NOR2_X1 U6233 ( .A1(n6692), .A2(n6710), .ZN(n4651) );
  OAI21_X1 U6234 ( .B1(n4658), .B2(n10084), .A(n4657), .ZN(P2_U3519) );
  NAND2_X1 U6235 ( .A1(n4671), .A2(n4538), .ZN(n8542) );
  NAND2_X1 U6236 ( .A1(n8535), .A2(n4673), .ZN(n4671) );
  NAND2_X1 U6237 ( .A1(n8537), .A2(n8536), .ZN(n4677) );
  NAND3_X1 U6238 ( .A1(n4683), .A2(n4679), .A3(n8509), .ZN(n4678) );
  NAND4_X1 U6239 ( .A1(n8504), .A2(n8505), .A3(n8580), .A4(n8503), .ZN(n4683)
         );
  NAND2_X1 U6240 ( .A1(n4685), .A2(n4537), .ZN(n8569) );
  NAND2_X1 U6241 ( .A1(n8552), .A2(n4687), .ZN(n4685) );
  NAND2_X1 U6242 ( .A1(n8563), .A2(n8562), .ZN(n4691) );
  AND2_X1 U6243 ( .A1(n8558), .A2(n8557), .ZN(n4692) );
  INV_X1 U6244 ( .A(n8550), .ZN(n4694) );
  NAND2_X1 U6245 ( .A1(n8682), .A2(n6369), .ZN(n6380) );
  NAND2_X1 U6246 ( .A1(n8656), .A2(n6352), .ZN(n6366) );
  NAND2_X1 U6247 ( .A1(n8042), .A2(n6339), .ZN(n8658) );
  OR2_X2 U6248 ( .A1(n8044), .A2(n8045), .ZN(n8042) );
  AND2_X2 U6249 ( .A1(n4695), .A2(n4529), .ZN(n8044) );
  NAND2_X1 U6250 ( .A1(n7910), .A2(n6321), .ZN(n4695) );
  NAND3_X1 U6251 ( .A1(n4697), .A2(n4696), .A3(n4540), .ZN(n5122) );
  XNOR2_X2 U6252 ( .A(n4698), .B(n5460), .ZN(n6811) );
  NAND2_X1 U6253 ( .A1(n4700), .A2(n4699), .ZN(n5289) );
  NAND3_X1 U6254 ( .A1(n5249), .A2(n5248), .A3(n5270), .ZN(n4699) );
  NAND3_X1 U6255 ( .A1(n4969), .A2(n7568), .A3(n6165), .ZN(n4963) );
  OAI211_X2 U6256 ( .C1(n4709), .C2(n4707), .A(n5055), .B(n4705), .ZN(n5398)
         );
  INV_X1 U6257 ( .A(n5312), .ZN(n4709) );
  NAND2_X1 U6258 ( .A1(n4709), .A2(n4710), .ZN(n4704) );
  NAND3_X1 U6259 ( .A1(n4706), .A2(n4708), .A3(n5368), .ZN(n4705) );
  INV_X1 U6260 ( .A(n4710), .ZN(n4706) );
  OR2_X2 U6261 ( .A1(n7664), .A2(n4715), .ZN(n4714) );
  INV_X1 U6262 ( .A(n7664), .ZN(n4716) );
  NAND2_X1 U6263 ( .A1(n4717), .A2(n4718), .ZN(n6451) );
  NAND2_X1 U6264 ( .A1(n8668), .A2(n4488), .ZN(n4717) );
  NOR2_X1 U6265 ( .A1(n4732), .A2(n4733), .ZN(n4731) );
  NAND2_X1 U6266 ( .A1(n9174), .A2(n9176), .ZN(n9112) );
  NAND2_X1 U6267 ( .A1(n9177), .A2(n9175), .ZN(n9174) );
  NAND2_X1 U6268 ( .A1(n4742), .A2(n7968), .ZN(n5558) );
  NAND3_X1 U6269 ( .A1(n7916), .A2(n7920), .A3(n4743), .ZN(n4742) );
  NAND2_X1 U6270 ( .A1(n5534), .A2(n5533), .ZN(n4744) );
  NAND2_X1 U6271 ( .A1(n5534), .A2(n5530), .ZN(n7919) );
  NAND2_X1 U6272 ( .A1(n5094), .A2(n4747), .ZN(n4746) );
  NAND3_X1 U6273 ( .A1(n5916), .A2(n5909), .A3(n5910), .ZN(n5945) );
  MUX2_X1 U6274 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6775), .S(n9214), .Z(n9217)
         );
  AND2_X2 U6275 ( .A1(n4985), .A2(n5056), .ZN(n5958) );
  OR2_X1 U6276 ( .A1(n6692), .A2(n6701), .ZN(n4772) );
  NAND2_X1 U6277 ( .A1(n7314), .A2(n9939), .ZN(n4776) );
  NAND2_X1 U6278 ( .A1(n7246), .A2(n7241), .ZN(n7303) );
  INV_X2 U6279 ( .A(n5192), .ZN(n5622) );
  OAI211_X2 U6280 ( .C1(n6637), .C2(n5223), .A(n4781), .B(n4780), .ZN(n6933)
         );
  NAND2_X1 U6281 ( .A1(n9419), .A2(n4782), .ZN(n9332) );
  INV_X1 U6282 ( .A(n4787), .ZN(n9360) );
  NAND2_X1 U6283 ( .A1(n4788), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5114) );
  NAND4_X1 U6284 ( .A1(n5244), .A2(n5071), .A3(n5067), .A4(n4522), .ZN(n4788)
         );
  NAND3_X1 U6285 ( .A1(n4792), .A2(n4791), .A3(n8356), .ZN(n4790) );
  AOI21_X1 U6286 ( .B1(n4795), .B2(n5043), .A(n8206), .ZN(n8207) );
  OR2_X1 U6287 ( .A1(n8196), .A2(n8197), .ZN(n4798) );
  NAND3_X1 U6288 ( .A1(n8254), .A2(n4803), .A3(n4806), .ZN(n4802) );
  NAND2_X1 U6289 ( .A1(n4812), .A2(n4531), .ZN(n7196) );
  NAND2_X1 U6290 ( .A1(n4814), .A2(n4507), .ZN(n5113) );
  OAI21_X1 U6291 ( .B1(n8221), .B2(n8220), .A(n8288), .ZN(n8222) );
  NOR2_X1 U6292 ( .A1(n8260), .A2(n8326), .ZN(n8333) );
  OAI211_X1 U6293 ( .C1(n8248), .C2(n8247), .A(n8414), .B(n8246), .ZN(n8254)
         );
  NOR2_X1 U6294 ( .A1(n8208), .A2(n8207), .ZN(n8212) );
  NAND2_X1 U6295 ( .A1(n8216), .A2(n8215), .ZN(n8219) );
  MUX2_X1 U6296 ( .A(n8244), .B(n8243), .S(n8258), .Z(n8247) );
  AOI21_X1 U6297 ( .B1(n8219), .B2(n9375), .A(n8402), .ZN(n8221) );
  AOI21_X1 U6298 ( .B1(n8297), .B2(n8259), .A(n8261), .ZN(n8260) );
  NOR2_X2 U6299 ( .A1(n7153), .A2(n7152), .ZN(n10039) );
  NAND2_X1 U6300 ( .A1(n9468), .A2(n4818), .ZN(n4815) );
  NAND2_X1 U6301 ( .A1(n4815), .A2(n4816), .ZN(n9341) );
  NAND3_X1 U6302 ( .A1(n4828), .A2(n7249), .A3(n4829), .ZN(n7252) );
  NAND2_X1 U6303 ( .A1(n7189), .A2(n7188), .ZN(n7341) );
  INV_X1 U6304 ( .A(n4829), .ZN(n4831) );
  NAND2_X1 U6305 ( .A1(n7740), .A2(n4834), .ZN(n4833) );
  OAI21_X1 U6306 ( .B1(n7296), .B2(n4839), .A(n4837), .ZN(n7429) );
  INV_X1 U6307 ( .A(n4838), .ZN(n4837) );
  NAND2_X1 U6308 ( .A1(n5115), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5111) );
  MUX2_X1 U6309 ( .A(n6686), .B(P2_REG2_REG_1__SCAN_IN), .S(n6701), .Z(n6687)
         );
  OAI21_X1 U6310 ( .B1(n7280), .B2(n4867), .A(n7279), .ZN(n9932) );
  NAND2_X1 U6311 ( .A1(n4874), .A2(n4530), .ZN(n9699) );
  NAND2_X1 U6312 ( .A1(n7479), .A2(n7406), .ZN(n6528) );
  XNOR2_X1 U6313 ( .A(n4884), .B(n6448), .ZN(n6138) );
  AND2_X1 U6314 ( .A1(n6494), .A2(n4884), .ZN(n4883) );
  AOI21_X1 U6315 ( .B1(n7478), .B2(n4884), .A(n7477), .ZN(n7561) );
  NAND2_X1 U6316 ( .A1(n5562), .A2(n4893), .ZN(n4890) );
  NAND2_X1 U6317 ( .A1(n4890), .A2(n4891), .ZN(n5644) );
  NAND2_X1 U6318 ( .A1(n5162), .A2(n5125), .ZN(n4899) );
  NAND3_X1 U6319 ( .A1(n4899), .A2(n5191), .A3(n4898), .ZN(n5130) );
  XNOR2_X1 U6320 ( .A(n5127), .B(SI_2_), .ZN(n5191) );
  OAI21_X1 U6321 ( .B1(n5162), .B2(n5161), .A(n5125), .ZN(n5190) );
  MUX2_X1 U6322 ( .A(n5126), .B(n6649), .S(n5121), .Z(n5127) );
  NAND2_X1 U6323 ( .A1(n4911), .A2(n8865), .ZN(n4910) );
  OAI21_X1 U6324 ( .B1(n8865), .B2(n8872), .A(n4922), .ZN(n8845) );
  NAND2_X1 U6325 ( .A1(n5312), .A2(n5311), .ZN(n4929) );
  NAND2_X1 U6326 ( .A1(n4930), .A2(n4553), .ZN(n5699) );
  NAND2_X1 U6327 ( .A1(n8128), .A2(n4934), .ZN(n4933) );
  NAND2_X1 U6328 ( .A1(n4931), .A2(n8130), .ZN(n4935) );
  NAND2_X1 U6329 ( .A1(n5751), .A2(n4945), .ZN(n4944) );
  NAND2_X1 U6330 ( .A1(n5751), .A2(n5750), .ZN(n5769) );
  AND2_X1 U6331 ( .A1(n5865), .A2(n5864), .ZN(n6542) );
  NAND2_X1 U6332 ( .A1(n5988), .A2(n4954), .ZN(n4952) );
  AND2_X1 U6333 ( .A1(n6056), .A2(n6035), .ZN(n4956) );
  OAI21_X1 U6334 ( .B1(n8693), .B2(n8694), .A(n6425), .ZN(n8643) );
  INV_X1 U6335 ( .A(n7360), .ZN(n4962) );
  NAND3_X1 U6336 ( .A1(n4968), .A2(n7568), .A3(n4969), .ZN(n4967) );
  OAI21_X1 U6337 ( .B1(n6511), .B2(n8993), .A(n4970), .ZN(P2_U3222) );
  AOI21_X1 U6338 ( .B1(n6490), .B2(n4973), .A(n4971), .ZN(n4970) );
  NAND3_X1 U6339 ( .A1(n4976), .A2(n6011), .A3(n6012), .ZN(n6917) );
  NAND2_X1 U6340 ( .A1(n6000), .A2(n6001), .ZN(n6012) );
  OAI21_X1 U6341 ( .B1(n6097), .B2(n7010), .A(n4982), .ZN(n7076) );
  NAND2_X1 U6342 ( .A1(n7075), .A2(n4979), .ZN(n4978) );
  INV_X1 U6343 ( .A(n7010), .ZN(n4979) );
  OR2_X1 U6344 ( .A1(n6110), .A2(n6109), .ZN(n4984) );
  AND2_X1 U6345 ( .A1(n6111), .A2(n5956), .ZN(n4985) );
  AND2_X1 U6346 ( .A1(n5056), .A2(n6111), .ZN(n5978) );
  NAND2_X1 U6347 ( .A1(n6464), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5961) );
  INV_X1 U6348 ( .A(n5641), .ZN(n4993) );
  NAND2_X1 U6349 ( .A1(n9112), .A2(n9113), .ZN(n9111) );
  NAND2_X1 U6350 ( .A1(n4998), .A2(n4999), .ZN(n5914) );
  OAI21_X1 U6351 ( .B1(n6565), .B2(n5007), .A(n5004), .ZN(n7956) );
  NAND3_X1 U6352 ( .A1(n6557), .A2(n5009), .A3(n6556), .ZN(n5014) );
  NAND3_X1 U6353 ( .A1(n6018), .A2(n5951), .A3(n5952), .ZN(n6059) );
  INV_X1 U6354 ( .A(n7649), .ZN(n5024) );
  NAND2_X1 U6355 ( .A1(n5019), .A2(n5017), .ZN(n7805) );
  INV_X1 U6356 ( .A(n8605), .ZN(n5018) );
  NOR2_X1 U6357 ( .A1(n8605), .A2(n5023), .ZN(n5020) );
  INV_X1 U6358 ( .A(n8922), .ZN(n5029) );
  NOR2_X1 U6359 ( .A1(n8818), .A2(n5045), .ZN(n8430) );
  AND2_X1 U6360 ( .A1(n5958), .A2(n4527), .ZN(n5969) );
  NAND2_X1 U6361 ( .A1(n5958), .A2(n5038), .ZN(n9080) );
  NAND2_X1 U6362 ( .A1(n6522), .A2(n6521), .ZN(n7061) );
  NAND2_X1 U6363 ( .A1(n6574), .A2(n8971), .ZN(n6580) );
  INV_X2 U6364 ( .A(n6058), .ZN(n6305) );
  AND2_X1 U6365 ( .A1(n6705), .A2(n8627), .ZN(n10010) );
  XNOR2_X1 U6366 ( .A(n8056), .B(n6546), .ZN(n9086) );
  INV_X1 U6367 ( .A(n7308), .ZN(n7189) );
  NAND2_X1 U6368 ( .A1(n6594), .A2(n10098), .ZN(n6592) );
  NAND2_X1 U6369 ( .A1(n7157), .A2(n10026), .ZN(n7087) );
  NAND2_X1 U6370 ( .A1(n5914), .A2(n5913), .ZN(n5944) );
  OAI22_X1 U6371 ( .A1(n7087), .A2(n10035), .B1(n10026), .B2(n6428), .ZN(n6915) );
  OR2_X1 U6372 ( .A1(n5969), .A2(n5968), .ZN(n5970) );
  INV_X1 U6373 ( .A(n6361), .ZN(n6498) );
  OR2_X1 U6374 ( .A1(n6361), .A2(n5971), .ZN(n5976) );
  INV_X1 U6375 ( .A(n5082), .ZN(n5085) );
  NOR2_X1 U6376 ( .A1(n7403), .A2(n6560), .ZN(n5039) );
  OR2_X1 U6377 ( .A1(n9262), .A2(n9693), .ZN(n5041) );
  NOR2_X1 U6378 ( .A1(n6284), .A2(n6283), .ZN(n5042) );
  AND2_X1 U6379 ( .A1(n8201), .A2(n8200), .ZN(n5043) );
  AND2_X1 U6380 ( .A1(n8817), .A2(n8705), .ZN(n5045) );
  OR2_X1 U6381 ( .A1(n6619), .A2(n8981), .ZN(n5046) );
  AND4_X1 U6382 ( .A1(n5567), .A2(n10230), .A3(n5091), .A4(n5564), .ZN(n5047)
         );
  AND2_X1 U6383 ( .A1(n5101), .A2(n5904), .ZN(n5048) );
  AND2_X1 U6384 ( .A1(n5073), .A2(n5072), .ZN(n5049) );
  INV_X1 U6385 ( .A(n9288), .ZN(n9253) );
  NAND2_X1 U6386 ( .A1(n6062), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5050) );
  AND2_X1 U6387 ( .A1(n5486), .A2(n5464), .ZN(n5051) );
  AND2_X1 U6388 ( .A1(n8233), .A2(n8232), .ZN(n5052) );
  AND2_X1 U6389 ( .A1(n5368), .A2(n5345), .ZN(n5053) );
  AND2_X1 U6390 ( .A1(n8800), .A2(n8703), .ZN(n5054) );
  AND2_X1 U6391 ( .A1(n5397), .A2(n5373), .ZN(n5055) );
  AND4_X1 U6392 ( .A1(n5984), .A2(n5950), .A3(n5949), .A4(n5948), .ZN(n5056)
         );
  NAND2_X1 U6393 ( .A1(n7539), .A2(n7538), .ZN(n5057) );
  XOR2_X1 U6394 ( .A(n9256), .B(n9255), .Z(n5058) );
  AND2_X1 U6395 ( .A1(n6616), .A2(n6615), .ZN(n5059) );
  AND2_X1 U6396 ( .A1(n9519), .A2(n9402), .ZN(n5060) );
  NAND2_X1 U6397 ( .A1(n7198), .A2(n7197), .ZN(n9700) );
  INV_X1 U6398 ( .A(n9700), .ZN(n9426) );
  INV_X1 U6399 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5179) );
  NAND2_X1 U6400 ( .A1(n9467), .A2(n8205), .ZN(n8206) );
  INV_X1 U6401 ( .A(n8258), .ZN(n8213) );
  NAND2_X1 U6402 ( .A1(n8214), .A2(n8213), .ZN(n8215) );
  NAND2_X1 U6403 ( .A1(n8231), .A2(n8213), .ZN(n8232) );
  INV_X1 U6404 ( .A(n8241), .ZN(n8239) );
  INV_X1 U6405 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5072) );
  INV_X1 U6406 ( .A(n9696), .ZN(n7859) );
  INV_X1 U6407 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5091) );
  OAI22_X1 U6408 ( .A1(n8433), .A2(n8444), .B1(n8443), .B2(n8801), .ZN(n8434)
         );
  INV_X1 U6409 ( .A(n6358), .ZN(n6356) );
  INV_X1 U6410 ( .A(n8903), .ZN(n6571) );
  AOI21_X1 U6411 ( .B1(n8705), .B2(n8966), .A(n5054), .ZN(n6579) );
  INV_X1 U6412 ( .A(n8611), .ZN(n6570) );
  AND2_X1 U6413 ( .A1(n6182), .A2(n6249), .ZN(n5984) );
  NAND2_X1 U6414 ( .A1(n5202), .A2(n5201), .ZN(n5203) );
  INV_X1 U6415 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5074) );
  INV_X1 U6416 ( .A(n5708), .ZN(n5706) );
  INV_X1 U6417 ( .A(n5599), .ZN(n5597) );
  INV_X1 U6418 ( .A(n9301), .ZN(n8411) );
  INV_X1 U6419 ( .A(n7436), .ZN(n7431) );
  NOR2_X1 U6420 ( .A1(n5070), .A2(n5069), .ZN(n5071) );
  INV_X1 U6421 ( .A(n5614), .ZN(n5615) );
  INV_X1 U6422 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5090) );
  INV_X1 U6423 ( .A(SI_10_), .ZN(n10238) );
  INV_X1 U6424 ( .A(n5310), .ZN(n5311) );
  INV_X1 U6425 ( .A(n7324), .ZN(n6143) );
  NAND2_X1 U6426 ( .A1(n6412), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6441) );
  NAND2_X1 U6427 ( .A1(n6290), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6310) );
  NOR2_X1 U6428 ( .A1(n6132), .A2(n6131), .ZN(n6154) );
  NAND2_X1 U6429 ( .A1(n6102), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6116) );
  OR2_X1 U6430 ( .A1(n6199), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6252) );
  INV_X1 U6431 ( .A(n5720), .ZN(n5721) );
  OR2_X1 U6432 ( .A1(n5843), .A2(n5842), .ZN(n5871) );
  INV_X1 U6433 ( .A(n5210), .ZN(n5932) );
  NOR2_X1 U6434 ( .A1(n5262), .A2(n5261), .ZN(n5299) );
  OR2_X2 U6435 ( .A1(n5671), .A2(n5670), .ZN(n5708) );
  NAND2_X1 U6436 ( .A1(n5597), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5627) );
  NOR2_X1 U6437 ( .A1(n5469), .A2(n7798), .ZN(n5494) );
  INV_X1 U6438 ( .A(n7256), .ZN(n7253) );
  INV_X1 U6439 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5076) );
  NAND2_X1 U6440 ( .A1(n5619), .A2(n5618), .ZN(n5642) );
  INV_X1 U6441 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5567) );
  NAND2_X1 U6442 ( .A1(n5462), .A2(n5461), .ZN(n5486) );
  OR3_X1 U6443 ( .A1(n5377), .A2(P1_IR_REG_8__SCAN_IN), .A3(n5376), .ZN(n5400)
         );
  AND2_X1 U6444 ( .A1(n6405), .A2(n6406), .ZN(n8666) );
  AND2_X1 U6445 ( .A1(n7982), .A2(n6275), .ZN(n6285) );
  OR3_X1 U6446 ( .A1(n6441), .A2(n10322), .A3(n6440), .ZN(n6609) );
  NAND2_X1 U6447 ( .A1(n6267), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6256) );
  OR2_X1 U6448 ( .A1(n6022), .A2(n10352), .ZN(n5974) );
  AND2_X1 U6449 ( .A1(n8757), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8751) );
  INV_X1 U6450 ( .A(n8519), .ZN(n8606) );
  OR2_X1 U6451 ( .A1(n10019), .A2(n6587), .ZN(n8907) );
  INV_X1 U6452 ( .A(n10076), .ZN(n9058) );
  INV_X1 U6453 ( .A(n8600), .ZN(n7457) );
  OR2_X1 U6454 ( .A1(n5627), .A2(n5626), .ZN(n5653) );
  AND2_X1 U6455 ( .A1(n5911), .A2(n9660), .ZN(n5909) );
  OR2_X1 U6456 ( .A1(n5938), .A2(n5920), .ZN(n9193) );
  OR2_X1 U6457 ( .A1(n5938), .A2(n5937), .ZN(n9652) );
  AND2_X1 U6458 ( .A1(n5871), .A2(n5844), .ZN(n9282) );
  NAND2_X1 U6459 ( .A1(n5547), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U6460 ( .A1(n5238), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5157) );
  INV_X1 U6461 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9810) );
  INV_X1 U6462 ( .A(n9430), .ZN(n8139) );
  INV_X1 U6463 ( .A(n9986), .ZN(n9960) );
  NAND2_X1 U6464 ( .A1(n9755), .A2(n9600), .ZN(n5178) );
  AND2_X1 U6465 ( .A1(n5667), .A2(n5648), .ZN(n5665) );
  AND2_X1 U6466 ( .A1(n6506), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9631) );
  INV_X1 U6467 ( .A(n6495), .ZN(n8626) );
  OR2_X1 U6468 ( .A1(n4482), .A2(n8849), .ZN(n6418) );
  OR2_X1 U6469 ( .A1(n6022), .A2(n6720), .ZN(n6045) );
  AOI21_X1 U6470 ( .B1(n6950), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6949), .ZN(
        n6954) );
  AND2_X1 U6471 ( .A1(n7648), .A2(n7647), .ZN(n9056) );
  INV_X1 U6472 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6595) );
  AND2_X1 U6473 ( .A1(n9063), .A2(n7961), .ZN(n9054) );
  AND2_X1 U6474 ( .A1(n6492), .A2(n8587), .ZN(n10070) );
  INV_X1 U6475 ( .A(n9054), .ZN(n10082) );
  AND2_X1 U6476 ( .A1(n6466), .A2(n6478), .ZN(n10018) );
  AND2_X1 U6477 ( .A1(n6261), .A2(n6219), .ZN(n8006) );
  INV_X1 U6478 ( .A(n9652), .ZN(n9196) );
  OR2_X1 U6479 ( .A1(n5921), .A2(n5928), .ZN(n5877) );
  NAND2_X1 U6480 ( .A1(n5382), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5089) );
  AND2_X1 U6481 ( .A1(n9751), .A2(n6773), .ZN(n9911) );
  INV_X1 U6482 ( .A(n9914), .ZN(n9883) );
  NAND2_X1 U6483 ( .A1(n8264), .A2(n8322), .ZN(n9255) );
  INV_X1 U6484 ( .A(n9415), .ZN(n9469) );
  NAND2_X1 U6485 ( .A1(n9950), .A2(n7050), .ZN(n9693) );
  INV_X1 U6486 ( .A(n9266), .ZN(n9691) );
  INV_X1 U6487 ( .A(n9976), .ZN(n9959) );
  INV_X1 U6488 ( .A(n9970), .ZN(n9988) );
  XNOR2_X1 U6489 ( .A(n5100), .B(n5099), .ZN(n5153) );
  INV_X1 U6490 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10365) );
  INV_X1 U6491 ( .A(n8799), .ZN(n10013) );
  INV_X1 U6492 ( .A(n9042), .ZN(n8039) );
  OR2_X1 U6493 ( .A1(n9635), .A2(n8958), .ZN(n8687) );
  INV_X1 U6494 ( .A(n6494), .ZN(n8692) );
  INV_X1 U6495 ( .A(n9618), .ZN(n10005) );
  AND2_X1 U6496 ( .A1(n8885), .A2(n8884), .ZN(n9017) );
  OR2_X1 U6497 ( .A1(n10098), .A2(n6590), .ZN(n6591) );
  NAND2_X1 U6498 ( .A1(n6593), .A2(n6589), .ZN(n10096) );
  NAND2_X1 U6499 ( .A1(n6593), .A2(n6599), .ZN(n10084) );
  NOR2_X1 U6500 ( .A1(n10019), .A2(n10018), .ZN(n10020) );
  INV_X1 U6501 ( .A(n10020), .ZN(n10128) );
  INV_X1 U6502 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n10341) );
  INV_X1 U6503 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10383) );
  INV_X1 U6504 ( .A(n7006), .ZN(n9087) );
  AND2_X1 U6505 ( .A1(n5927), .A2(n5926), .ZN(n9665) );
  OR2_X1 U6506 ( .A1(n5938), .A2(n5908), .ZN(n9186) );
  NAND2_X1 U6507 ( .A1(n5877), .A2(n5876), .ZN(n9288) );
  INV_X1 U6508 ( .A(P1_U4006), .ZN(n9211) );
  OR2_X1 U6509 ( .A1(P1_U3083), .A2(n6792), .ZN(n9924) );
  OR2_X1 U6510 ( .A1(n9709), .A2(n7053), .ZN(n9475) );
  INV_X1 U6511 ( .A(n9478), .ZN(n9678) );
  OR2_X1 U6512 ( .A1(n9709), .A2(n7258), .ZN(n9415) );
  AND2_X1 U6513 ( .A1(n7051), .A2(n9693), .ZN(n9709) );
  AND2_X2 U6514 ( .A1(n6980), .A2(n9928), .ZN(n10004) );
  INV_X1 U6515 ( .A(n10004), .ZN(n10002) );
  INV_X1 U6516 ( .A(n9408), .ZN(n9568) );
  AND2_X2 U6517 ( .A1(n6980), .A2(n7049), .ZN(n9992) );
  AND2_X1 U6518 ( .A1(n9931), .A2(n9925), .ZN(n9926) );
  INV_X1 U6519 ( .A(n9926), .ZN(n9927) );
  AND2_X1 U6520 ( .A1(n6621), .A2(n5906), .ZN(n9931) );
  INV_X1 U6521 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7008) );
  INV_X1 U6522 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6684) );
  NAND2_X1 U6523 ( .A1(n5059), .A2(n5046), .ZN(P2_U3267) );
  NAND2_X1 U6524 ( .A1(n5193), .A2(n5061), .ZN(n5138) );
  NOR2_X1 U6525 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5066) );
  NOR2_X1 U6526 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5065) );
  NOR2_X1 U6527 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5064) );
  NOR2_X1 U6528 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5063) );
  NOR2_X1 U6529 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5068) );
  NAND4_X1 U6530 ( .A1(n5068), .A2(n5564), .A3(n10230), .A4(n5096), .ZN(n5070)
         );
  NAND4_X1 U6531 ( .A1(n5093), .A2(n5090), .A3(n5091), .A4(n5099), .ZN(n5069)
         );
  INV_X1 U6532 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5077) );
  NAND2_X1 U6533 ( .A1(n5113), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5079) );
  MUX2_X1 U6534 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5079), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5081) );
  INV_X1 U6535 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6782) );
  OR2_X1 U6536 ( .A1(n5784), .A2(n6782), .ZN(n5088) );
  AND2_X4 U6537 ( .A1(n5083), .A2(n5085), .ZN(n5845) );
  NOR2_X1 U6538 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5084) );
  NOR2_X1 U6539 ( .A1(n5236), .A2(n5084), .ZN(n7331) );
  NAND2_X1 U6540 ( .A1(n5845), .A2(n7331), .ZN(n5087) );
  AND2_X4 U6541 ( .A1(n8057), .A2(n5085), .ZN(n5210) );
  NAND2_X1 U6542 ( .A1(n5210), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5086) );
  INV_X1 U6543 ( .A(n5097), .ZN(n5095) );
  NAND2_X1 U6544 ( .A1(n5095), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n5098) );
  NAND2_X1 U6545 ( .A1(n5097), .A2(n5096), .ZN(n5145) );
  NAND2_X1 U6546 ( .A1(n5098), .A2(n5145), .ZN(n5907) );
  OR2_X2 U6547 ( .A1(n5907), .A2(n8334), .ZN(n7199) );
  INV_X1 U6548 ( .A(n7199), .ZN(n7281) );
  NAND2_X1 U6549 ( .A1(n5103), .A2(n5101), .ZN(n5104) );
  NAND2_X1 U6550 ( .A1(n5106), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5107) );
  MUX2_X1 U6551 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5107), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5109) );
  NAND2_X1 U6552 ( .A1(n5109), .A2(n5108), .ZN(n7850) );
  NOR2_X1 U6553 ( .A1(n7892), .A2(n7850), .ZN(n5110) );
  AND2_X2 U6554 ( .A1(n7281), .A2(n6621), .ZN(n5268) );
  NAND2_X1 U6555 ( .A1(n9212), .A2(n5882), .ZN(n5144) );
  NAND2_X1 U6556 ( .A1(n5117), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5118) );
  INV_X1 U6557 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6635) );
  NAND2_X2 U6558 ( .A1(n5174), .A2(n6633), .ZN(n5223) );
  AND2_X1 U6559 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5120) );
  NAND2_X1 U6560 ( .A1(n5121), .A2(n5120), .ZN(n6009) );
  NAND2_X1 U6561 ( .A1(n5122), .A2(n6009), .ZN(n5124) );
  XNOR2_X1 U6562 ( .A(n5124), .B(SI_1_), .ZN(n5162) );
  INV_X1 U6563 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6632) );
  INV_X1 U6564 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5123) );
  MUX2_X1 U6565 ( .A(n6632), .B(n5123), .S(n5131), .Z(n5161) );
  NAND2_X1 U6566 ( .A1(n5124), .A2(SI_1_), .ZN(n5125) );
  INV_X1 U6567 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6649) );
  INV_X1 U6568 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5126) );
  INV_X1 U6569 ( .A(n5127), .ZN(n5128) );
  NAND2_X1 U6570 ( .A1(n5128), .A2(SI_2_), .ZN(n5129) );
  NAND2_X1 U6571 ( .A1(n5130), .A2(n5129), .ZN(n5216) );
  INV_X1 U6572 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6644) );
  INV_X1 U6573 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5132) );
  MUX2_X1 U6574 ( .A(n6644), .B(n5132), .S(n5131), .Z(n5133) );
  XNOR2_X1 U6575 ( .A(n5133), .B(SI_3_), .ZN(n5215) );
  NAND2_X1 U6576 ( .A1(n5216), .A2(n5215), .ZN(n5136) );
  INV_X1 U6577 ( .A(n5133), .ZN(n5134) );
  NAND2_X1 U6578 ( .A1(n5134), .A2(SI_3_), .ZN(n5135) );
  XNOR2_X1 U6579 ( .A(n5250), .B(SI_4_), .ZN(n5247) );
  XNOR2_X1 U6580 ( .A(n5249), .B(n5247), .ZN(n6634) );
  NAND2_X1 U6581 ( .A1(n8132), .A2(n6634), .ZN(n5142) );
  NAND2_X1 U6582 ( .A1(n5138), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5139) );
  MUX2_X1 U6583 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5139), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5140) );
  AND2_X1 U6584 ( .A1(n5137), .A2(n5140), .ZN(n6781) );
  NAND2_X1 U6585 ( .A1(n5594), .A2(n6781), .ZN(n5141) );
  NAND2_X1 U6586 ( .A1(n7332), .A2(n4475), .ZN(n5143) );
  NAND2_X1 U6587 ( .A1(n5144), .A2(n5143), .ZN(n5152) );
  NAND2_X1 U6588 ( .A1(n5145), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5147) );
  INV_X1 U6589 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U6590 ( .A1(n5149), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5150) );
  MUX2_X1 U6591 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5150), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n5151) );
  XNOR2_X1 U6592 ( .A(n5152), .B(n5855), .ZN(n6966) );
  NAND2_X1 U6593 ( .A1(n8259), .A2(n5918), .ZN(n5154) );
  AND2_X4 U6594 ( .A1(n4475), .A2(n5154), .ZN(n5878) );
  NAND2_X1 U6595 ( .A1(n9212), .A2(n5878), .ZN(n5156) );
  NAND2_X1 U6596 ( .A1(n5882), .A2(n7332), .ZN(n5155) );
  AND2_X1 U6597 ( .A1(n5156), .A2(n5155), .ZN(n6965) );
  AND2_X1 U6598 ( .A1(n6966), .A2(n6965), .ZN(n5235) );
  NAND2_X1 U6599 ( .A1(n5382), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5160) );
  NAND2_X1 U6600 ( .A1(n7186), .A2(n5268), .ZN(n5164) );
  XNOR2_X1 U6601 ( .A(n5162), .B(n5161), .ZN(n6637) );
  NAND2_X1 U6602 ( .A1(n6933), .A2(n4475), .ZN(n5163) );
  NAND2_X1 U6603 ( .A1(n5164), .A2(n5163), .ZN(n5165) );
  XNOR2_X1 U6604 ( .A(n5165), .B(n7257), .ZN(n5169) );
  INV_X1 U6605 ( .A(n5169), .ZN(n6931) );
  NAND2_X1 U6606 ( .A1(n7186), .A2(n5878), .ZN(n5167) );
  NAND2_X1 U6607 ( .A1(n6933), .A2(n5268), .ZN(n5166) );
  NAND2_X1 U6608 ( .A1(n5167), .A2(n5166), .ZN(n5168) );
  INV_X1 U6609 ( .A(n5168), .ZN(n6929) );
  NAND2_X1 U6610 ( .A1(n6931), .A2(n6929), .ZN(n5189) );
  NAND2_X1 U6611 ( .A1(n5169), .A2(n5168), .ZN(n5187) );
  NAND2_X1 U6612 ( .A1(n5210), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5173) );
  NAND2_X1 U6613 ( .A1(n5845), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U6614 ( .A1(n5382), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5171) );
  NAND2_X1 U6615 ( .A1(n5238), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6616 ( .A1(n6854), .A2(n5878), .ZN(n5181) );
  INV_X1 U6617 ( .A(SI_0_), .ZN(n5175) );
  NOR2_X1 U6618 ( .A1(n4481), .A2(n5175), .ZN(n5177) );
  INV_X1 U6619 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5176) );
  XNOR2_X1 U6620 ( .A(n5177), .B(n5176), .ZN(n9600) );
  OAI21_X2 U6621 ( .B1(n9755), .B2(n5179), .A(n5178), .ZN(n7192) );
  INV_X1 U6622 ( .A(n6621), .ZN(n5182) );
  AOI22_X1 U6623 ( .A1(n5268), .A2(n7192), .B1(n5182), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5180) );
  NAND2_X1 U6624 ( .A1(n6854), .A2(n5268), .ZN(n5184) );
  AOI22_X1 U6625 ( .A1(n7192), .A2(n5196), .B1(n5182), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6626 ( .A1(n5184), .A2(n5183), .ZN(n6868) );
  INV_X1 U6627 ( .A(n6868), .ZN(n5185) );
  NAND2_X1 U6628 ( .A1(n5185), .A2(n7257), .ZN(n5186) );
  NAND2_X1 U6629 ( .A1(n5189), .A2(n5188), .ZN(n6939) );
  XNOR2_X1 U6630 ( .A(n5190), .B(n5191), .ZN(n6648) );
  NAND2_X1 U6631 ( .A1(n5192), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5195) );
  INV_X1 U6632 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9590) );
  OR2_X1 U6633 ( .A1(n5193), .A2(n9590), .ZN(n5218) );
  NAND2_X1 U6634 ( .A1(n5594), .A2(n6892), .ZN(n5194) );
  OAI211_X1 U6635 ( .C1(n6648), .C2(n5223), .A(n5195), .B(n5194), .ZN(n7315)
         );
  NAND2_X1 U6636 ( .A1(n7315), .A2(n4475), .ZN(n5202) );
  NAND2_X1 U6637 ( .A1(n5210), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U6638 ( .A1(n5845), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5199) );
  NAND2_X1 U6639 ( .A1(n5382), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6640 ( .A1(n5238), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6641 ( .A1(n5204), .A2(n5268), .ZN(n5201) );
  AOI22_X1 U6642 ( .A1(n5204), .A2(n5878), .B1(n5268), .B2(n7315), .ZN(n5206)
         );
  XNOR2_X1 U6643 ( .A(n5205), .B(n5206), .ZN(n6938) );
  NAND2_X1 U6644 ( .A1(n6939), .A2(n6938), .ZN(n5209) );
  INV_X1 U6645 ( .A(n5205), .ZN(n5207) );
  NAND2_X1 U6646 ( .A1(n5207), .A2(n5206), .ZN(n5208) );
  NAND2_X1 U6647 ( .A1(n5209), .A2(n5208), .ZN(n6921) );
  INV_X1 U6648 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6925) );
  NAND2_X1 U6649 ( .A1(n5845), .A2(n6925), .ZN(n5214) );
  NAND2_X1 U6650 ( .A1(n5238), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U6651 ( .A1(n5210), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5212) );
  NAND2_X1 U6652 ( .A1(n5382), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5211) );
  NAND4_X1 U6653 ( .A1(n5214), .A2(n5213), .A3(n5212), .A4(n5211), .ZN(n9213)
         );
  NAND2_X1 U6654 ( .A1(n9213), .A2(n5268), .ZN(n5225) );
  XNOR2_X1 U6655 ( .A(n5216), .B(n5215), .ZN(n6643) );
  NAND2_X1 U6656 ( .A1(n5192), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5222) );
  INV_X1 U6657 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U6658 ( .A1(n5218), .A2(n5217), .ZN(n5219) );
  NAND2_X1 U6659 ( .A1(n5219), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5220) );
  XNOR2_X1 U6660 ( .A(n5220), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6809) );
  NAND2_X1 U6661 ( .A1(n5594), .A2(n6809), .ZN(n5221) );
  NAND2_X1 U6662 ( .A1(n7351), .A2(n4475), .ZN(n5224) );
  NAND2_X1 U6663 ( .A1(n5225), .A2(n5224), .ZN(n5226) );
  XNOR2_X1 U6664 ( .A(n5226), .B(n7257), .ZN(n5227) );
  AOI22_X1 U6665 ( .A1(n9213), .A2(n5878), .B1(n5882), .B2(n7351), .ZN(n5228)
         );
  XNOR2_X1 U6666 ( .A(n5227), .B(n5228), .ZN(n6922) );
  NAND2_X1 U6667 ( .A1(n6921), .A2(n6922), .ZN(n5231) );
  INV_X1 U6668 ( .A(n5227), .ZN(n5229) );
  NAND2_X1 U6669 ( .A1(n5229), .A2(n5228), .ZN(n5230) );
  INV_X1 U6670 ( .A(n6966), .ZN(n5233) );
  INV_X1 U6671 ( .A(n6965), .ZN(n5232) );
  NAND2_X1 U6672 ( .A1(n5233), .A2(n5232), .ZN(n5234) );
  NAND2_X1 U6673 ( .A1(n5382), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5242) );
  NAND2_X1 U6674 ( .A1(n5210), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U6675 ( .A1(n5236), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5262) );
  OAI21_X1 U6676 ( .B1(n5236), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5262), .ZN(
        n7244) );
  INV_X1 U6677 ( .A(n7244), .ZN(n5237) );
  NAND2_X1 U6678 ( .A1(n5845), .A2(n5237), .ZN(n5240) );
  NAND2_X1 U6679 ( .A1(n8133), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5239) );
  NAND4_X1 U6680 ( .A1(n5242), .A2(n5241), .A3(n5240), .A4(n5239), .ZN(n9210)
         );
  NAND2_X1 U6681 ( .A1(n9210), .A2(n5882), .ZN(n5255) );
  NAND2_X1 U6682 ( .A1(n5137), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5243) );
  MUX2_X1 U6683 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5243), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5246) );
  INV_X1 U6684 ( .A(n5244), .ZN(n5245) );
  INV_X1 U6685 ( .A(n6784), .ZN(n9771) );
  NAND2_X1 U6686 ( .A1(n5250), .A2(SI_4_), .ZN(n5251) );
  MUX2_X1 U6687 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5131), .Z(n5271) );
  XNOR2_X1 U6688 ( .A(n5271), .B(SI_5_), .ZN(n5269) );
  XNOR2_X1 U6689 ( .A(n5252), .B(n5269), .ZN(n6640) );
  NAND2_X1 U6690 ( .A1(n8131), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5253) );
  NAND2_X1 U6691 ( .A1(n7294), .A2(n4475), .ZN(n5254) );
  NAND2_X1 U6692 ( .A1(n5255), .A2(n5254), .ZN(n5256) );
  XNOR2_X1 U6693 ( .A(n5256), .B(n5855), .ZN(n7115) );
  NAND2_X1 U6694 ( .A1(n9210), .A2(n5878), .ZN(n5258) );
  NAND2_X1 U6695 ( .A1(n7294), .A2(n5882), .ZN(n5257) );
  AND2_X1 U6696 ( .A1(n5258), .A2(n5257), .ZN(n7114) );
  NAND2_X1 U6697 ( .A1(n7115), .A2(n7114), .ZN(n5259) );
  NAND2_X1 U6698 ( .A1(n7117), .A2(n5259), .ZN(n5282) );
  INV_X1 U6699 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5260) );
  OR2_X1 U6700 ( .A1(n5784), .A2(n5260), .ZN(n5267) );
  NAND2_X1 U6701 ( .A1(n5382), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5266) );
  AND2_X1 U6702 ( .A1(n5262), .A2(n5261), .ZN(n5263) );
  NOR2_X1 U6703 ( .A1(n5299), .A2(n5263), .ZN(n7368) );
  NAND2_X1 U6704 ( .A1(n5845), .A2(n7368), .ZN(n5265) );
  NAND2_X1 U6705 ( .A1(n5210), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5264) );
  NAND4_X1 U6706 ( .A1(n5267), .A2(n5266), .A3(n5265), .A4(n5264), .ZN(n9209)
         );
  NAND2_X1 U6707 ( .A1(n9209), .A2(n5852), .ZN(n5276) );
  INV_X1 U6708 ( .A(n5269), .ZN(n5270) );
  MUX2_X1 U6709 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6633), .Z(n5290) );
  XNOR2_X1 U6710 ( .A(n5290), .B(SI_6_), .ZN(n5287) );
  XNOR2_X1 U6711 ( .A(n5289), .B(n5287), .ZN(n6650) );
  NAND2_X1 U6712 ( .A1(n6650), .A2(n8132), .ZN(n5274) );
  OR2_X1 U6713 ( .A1(n5244), .A2(n9590), .ZN(n5272) );
  XNOR2_X1 U6714 ( .A(n5272), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6789) );
  AOI22_X1 U6715 ( .A1(n8131), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5594), .B2(
        n6789), .ZN(n5273) );
  NAND2_X1 U6716 ( .A1(n5274), .A2(n5273), .ZN(n9958) );
  NAND2_X1 U6717 ( .A1(n9958), .A2(n4475), .ZN(n5275) );
  NAND2_X1 U6718 ( .A1(n5276), .A2(n5275), .ZN(n5277) );
  XNOR2_X1 U6719 ( .A(n5277), .B(n5855), .ZN(n5285) );
  NAND2_X1 U6720 ( .A1(n9209), .A2(n5878), .ZN(n5279) );
  NAND2_X1 U6721 ( .A1(n9958), .A2(n5882), .ZN(n5278) );
  NAND2_X1 U6722 ( .A1(n5279), .A2(n5278), .ZN(n5283) );
  XNOR2_X1 U6723 ( .A(n5285), .B(n5283), .ZN(n7374) );
  INV_X1 U6724 ( .A(n5283), .ZN(n5284) );
  NAND2_X1 U6725 ( .A1(n5285), .A2(n5284), .ZN(n5286) );
  INV_X1 U6726 ( .A(n5287), .ZN(n5288) );
  NAND2_X1 U6727 ( .A1(n5289), .A2(n5288), .ZN(n5292) );
  NAND2_X1 U6728 ( .A1(n5290), .A2(SI_6_), .ZN(n5291) );
  NAND2_X1 U6729 ( .A1(n5292), .A2(n5291), .ZN(n5312) );
  MUX2_X1 U6730 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4473), .Z(n5313) );
  XNOR2_X1 U6731 ( .A(n5312), .B(n5310), .ZN(n6655) );
  NAND2_X1 U6732 ( .A1(n6655), .A2(n8132), .ZN(n5296) );
  INV_X1 U6733 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6657) );
  INV_X1 U6734 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6735 ( .A1(n5244), .A2(n5293), .ZN(n5377) );
  NAND2_X1 U6736 ( .A1(n5377), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5318) );
  XNOR2_X1 U6737 ( .A(n5318), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6829) );
  INV_X1 U6738 ( .A(n6829), .ZN(n6774) );
  OAI22_X1 U6739 ( .A1(n5622), .A2(n6657), .B1(n9755), .B2(n6774), .ZN(n5294)
         );
  INV_X1 U6740 ( .A(n5294), .ZN(n5295) );
  NAND2_X1 U6741 ( .A1(n5296), .A2(n5295), .ZN(n7427) );
  NAND2_X1 U6742 ( .A1(n7427), .A2(n4475), .ZN(n5306) );
  INV_X1 U6743 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5297) );
  OR2_X1 U6744 ( .A1(n5784), .A2(n5297), .ZN(n5304) );
  INV_X1 U6745 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5298) );
  OR2_X1 U6746 ( .A1(n5848), .A2(n5298), .ZN(n5303) );
  NAND2_X1 U6747 ( .A1(n5299), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5325) );
  OR2_X1 U6748 ( .A1(n5299), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5300) );
  AND2_X1 U6749 ( .A1(n5325), .A2(n5300), .ZN(n7395) );
  NAND2_X1 U6750 ( .A1(n5845), .A2(n7395), .ZN(n5302) );
  NAND2_X1 U6751 ( .A1(n5210), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5301) );
  NAND4_X1 U6752 ( .A1(n5304), .A2(n5303), .A3(n5302), .A4(n5301), .ZN(n9208)
         );
  NAND2_X1 U6753 ( .A1(n9208), .A2(n5852), .ZN(n5305) );
  NAND2_X1 U6754 ( .A1(n5306), .A2(n5305), .ZN(n5307) );
  XNOR2_X1 U6755 ( .A(n5307), .B(n5855), .ZN(n5309) );
  AOI22_X1 U6756 ( .A1(n7427), .A2(n5882), .B1(n5878), .B2(n9208), .ZN(n5308)
         );
  AND2_X1 U6757 ( .A1(n5309), .A2(n5308), .ZN(n7175) );
  OR2_X1 U6758 ( .A1(n5309), .A2(n5308), .ZN(n7173) );
  NAND2_X1 U6759 ( .A1(n5313), .A2(SI_7_), .ZN(n5314) );
  INV_X1 U6760 ( .A(SI_8_), .ZN(n5315) );
  NAND2_X1 U6761 ( .A1(n5338), .A2(n5317), .ZN(n5339) );
  XNOR2_X1 U6762 ( .A(n5340), .B(n5339), .ZN(n6659) );
  NAND2_X1 U6763 ( .A1(n6659), .A2(n8132), .ZN(n5322) );
  INV_X1 U6764 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U6765 ( .A1(n5318), .A2(n5375), .ZN(n5319) );
  NAND2_X1 U6766 ( .A1(n5319), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5347) );
  XNOR2_X1 U6767 ( .A(n5347), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9803) );
  INV_X1 U6768 ( .A(n9803), .ZN(n6827) );
  OAI22_X1 U6769 ( .A1(n5622), .A2(n6660), .B1(n9755), .B2(n6827), .ZN(n5320)
         );
  INV_X1 U6770 ( .A(n5320), .ZN(n5321) );
  NAND2_X1 U6771 ( .A1(n5322), .A2(n5321), .ZN(n8165) );
  NAND2_X1 U6772 ( .A1(n8165), .A2(n5882), .ZN(n5332) );
  INV_X1 U6773 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5323) );
  OR2_X1 U6774 ( .A1(n5848), .A2(n5323), .ZN(n5330) );
  NAND2_X1 U6775 ( .A1(n5325), .A2(n5324), .ZN(n5326) );
  AND2_X1 U6776 ( .A1(n5352), .A2(n5326), .ZN(n7442) );
  NAND2_X1 U6777 ( .A1(n5845), .A2(n7442), .ZN(n5329) );
  INV_X1 U6778 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7443) );
  OR2_X1 U6779 ( .A1(n5784), .A2(n7443), .ZN(n5328) );
  NAND2_X1 U6780 ( .A1(n5210), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5327) );
  NAND4_X1 U6781 ( .A1(n5330), .A2(n5329), .A3(n5328), .A4(n5327), .ZN(n9654)
         );
  NAND2_X1 U6782 ( .A1(n9654), .A2(n5878), .ZN(n5331) );
  NAND2_X1 U6783 ( .A1(n5332), .A2(n5331), .ZN(n5337) );
  NAND2_X1 U6784 ( .A1(n8165), .A2(n4475), .ZN(n5334) );
  NAND2_X1 U6785 ( .A1(n9654), .A2(n5852), .ZN(n5333) );
  NAND2_X1 U6786 ( .A1(n5334), .A2(n5333), .ZN(n5335) );
  XNOR2_X1 U6787 ( .A(n5335), .B(n5855), .ZN(n7504) );
  INV_X1 U6788 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5341) );
  MUX2_X1 U6789 ( .A(n10383), .B(n5341), .S(n6633), .Z(n5343) );
  INV_X1 U6790 ( .A(SI_9_), .ZN(n5342) );
  NAND2_X1 U6791 ( .A1(n5343), .A2(n5342), .ZN(n5368) );
  INV_X1 U6792 ( .A(n5343), .ZN(n5344) );
  NAND2_X1 U6793 ( .A1(n5344), .A2(SI_9_), .ZN(n5345) );
  NAND2_X1 U6794 ( .A1(n6127), .A2(n8132), .ZN(n5351) );
  INV_X1 U6795 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6796 ( .A1(n5347), .A2(n5346), .ZN(n5348) );
  NAND2_X1 U6797 ( .A1(n5348), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5349) );
  XNOR2_X1 U6798 ( .A(n5349), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9816) );
  AOI22_X1 U6799 ( .A1(n8131), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5594), .B2(
        n9816), .ZN(n5350) );
  NAND2_X1 U6800 ( .A1(n5351), .A2(n5350), .ZN(n8166) );
  NAND2_X1 U6801 ( .A1(n8166), .A2(n4475), .ZN(n5360) );
  AND2_X1 U6802 ( .A1(n5352), .A2(n9810), .ZN(n5353) );
  OR2_X1 U6803 ( .A1(n5353), .A2(n5383), .ZN(n9664) );
  INV_X1 U6804 ( .A(n9664), .ZN(n5354) );
  NAND2_X1 U6805 ( .A1(n5845), .A2(n5354), .ZN(n5358) );
  NAND2_X1 U6806 ( .A1(n8133), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5357) );
  NAND2_X1 U6807 ( .A1(n5210), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6808 ( .A1(n5382), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5355) );
  NAND4_X1 U6809 ( .A1(n5358), .A2(n5357), .A3(n5356), .A4(n5355), .ZN(n9207)
         );
  NAND2_X1 U6810 ( .A1(n9207), .A2(n5852), .ZN(n5359) );
  NAND2_X1 U6811 ( .A1(n5360), .A2(n5359), .ZN(n5361) );
  XNOR2_X1 U6812 ( .A(n5361), .B(n7257), .ZN(n5363) );
  AND2_X1 U6813 ( .A1(n9207), .A2(n5878), .ZN(n5362) );
  AOI21_X1 U6814 ( .B1(n8166), .B2(n5852), .A(n5362), .ZN(n5364) );
  XNOR2_X1 U6815 ( .A(n5363), .B(n5364), .ZN(n9657) );
  INV_X1 U6816 ( .A(n5363), .ZN(n5365) );
  NAND2_X1 U6817 ( .A1(n5365), .A2(n5364), .ZN(n5366) );
  INV_X1 U6818 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5370) );
  INV_X1 U6819 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5369) );
  MUX2_X1 U6820 ( .A(n5370), .B(n5369), .S(n5131), .Z(n5371) );
  INV_X1 U6821 ( .A(n5371), .ZN(n5372) );
  NAND2_X1 U6822 ( .A1(n5372), .A2(SI_10_), .ZN(n5373) );
  XNOR2_X1 U6823 ( .A(n5396), .B(n5055), .ZN(n6678) );
  NAND2_X1 U6824 ( .A1(n6678), .A2(n8132), .ZN(n5380) );
  INV_X1 U6825 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6826 ( .A1(n5375), .A2(n5374), .ZN(n5376) );
  NAND2_X1 U6827 ( .A1(n5400), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5378) );
  XNOR2_X1 U6828 ( .A(n5378), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9823) );
  AOI22_X1 U6829 ( .A1(n8131), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5594), .B2(
        n9823), .ZN(n5379) );
  NAND2_X1 U6830 ( .A1(n7706), .A2(n4475), .ZN(n5390) );
  INV_X1 U6831 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5381) );
  OR2_X1 U6832 ( .A1(n5784), .A2(n5381), .ZN(n5388) );
  NAND2_X1 U6833 ( .A1(n5382), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5387) );
  NOR2_X1 U6834 ( .A1(n5383), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5384) );
  OR2_X1 U6835 ( .A1(n5412), .A2(n5384), .ZN(n7544) );
  INV_X1 U6836 ( .A(n7544), .ZN(n7531) );
  NAND2_X1 U6837 ( .A1(n5845), .A2(n7531), .ZN(n5386) );
  NAND2_X1 U6838 ( .A1(n5210), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5385) );
  NAND4_X1 U6839 ( .A1(n5388), .A2(n5387), .A3(n5386), .A4(n5385), .ZN(n9206)
         );
  NAND2_X1 U6840 ( .A1(n9206), .A2(n5852), .ZN(n5389) );
  NAND2_X1 U6841 ( .A1(n5390), .A2(n5389), .ZN(n5391) );
  XNOR2_X1 U6842 ( .A(n5391), .B(n5855), .ZN(n7539) );
  AND2_X1 U6843 ( .A1(n9206), .A2(n5878), .ZN(n5392) );
  AOI21_X1 U6844 ( .B1(n7706), .B2(n5852), .A(n5392), .ZN(n7538) );
  INV_X1 U6845 ( .A(n7539), .ZN(n5394) );
  INV_X1 U6846 ( .A(n7538), .ZN(n5393) );
  NAND2_X1 U6847 ( .A1(n5394), .A2(n5393), .ZN(n5395) );
  INV_X1 U6848 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5399) );
  MUX2_X1 U6849 ( .A(n5399), .B(n6684), .S(n6633), .Z(n5426) );
  XNOR2_X1 U6850 ( .A(n5430), .B(n5425), .ZN(n6682) );
  NAND2_X1 U6851 ( .A1(n6682), .A2(n8132), .ZN(n5410) );
  INV_X1 U6852 ( .A(n5400), .ZN(n5402) );
  INV_X1 U6853 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6854 ( .A1(n5402), .A2(n5401), .ZN(n5404) );
  NAND2_X1 U6855 ( .A1(n5404), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5403) );
  MUX2_X1 U6856 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5403), .S(
        P1_IR_REG_11__SCAN_IN), .Z(n5407) );
  INV_X1 U6857 ( .A(n5404), .ZN(n5406) );
  INV_X1 U6858 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6859 ( .A1(n5406), .A2(n5405), .ZN(n5435) );
  NAND2_X1 U6860 ( .A1(n5407), .A2(n5435), .ZN(n7493) );
  OAI22_X1 U6861 ( .A1(n5622), .A2(n6684), .B1(n9755), .B2(n7493), .ZN(n5408)
         );
  INV_X1 U6862 ( .A(n5408), .ZN(n5409) );
  NAND2_X1 U6863 ( .A1(n9737), .A2(n4475), .ZN(n5419) );
  INV_X1 U6864 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5411) );
  OR2_X1 U6865 ( .A1(n5848), .A2(n5411), .ZN(n5417) );
  NAND2_X1 U6866 ( .A1(n5210), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5416) );
  INV_X1 U6867 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7714) );
  OR2_X1 U6868 ( .A1(n5784), .A2(n7714), .ZN(n5415) );
  OR2_X1 U6869 ( .A1(n5412), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5413) );
  AND2_X1 U6870 ( .A1(n5443), .A2(n5413), .ZN(n7639) );
  NAND2_X1 U6871 ( .A1(n5845), .A2(n7639), .ZN(n5414) );
  NAND4_X1 U6872 ( .A1(n5417), .A2(n5416), .A3(n5415), .A4(n5414), .ZN(n9205)
         );
  NAND2_X1 U6873 ( .A1(n9205), .A2(n5882), .ZN(n5418) );
  NAND2_X1 U6874 ( .A1(n5419), .A2(n5418), .ZN(n5420) );
  XNOR2_X1 U6875 ( .A(n5420), .B(n7257), .ZN(n5424) );
  AND2_X1 U6876 ( .A1(n9205), .A2(n5878), .ZN(n5421) );
  AOI21_X1 U6877 ( .B1(n9737), .B2(n5882), .A(n5421), .ZN(n5422) );
  XNOR2_X1 U6878 ( .A(n5424), .B(n5422), .ZN(n7638) );
  INV_X1 U6879 ( .A(n5422), .ZN(n5423) );
  INV_X1 U6880 ( .A(n5426), .ZN(n5427) );
  NAND2_X1 U6881 ( .A1(n5427), .A2(SI_11_), .ZN(n5428) );
  MUX2_X1 U6882 ( .A(n6812), .B(n6813), .S(n6633), .Z(n5432) );
  INV_X1 U6883 ( .A(SI_12_), .ZN(n5431) );
  INV_X1 U6884 ( .A(n5432), .ZN(n5433) );
  NAND2_X1 U6885 ( .A1(n5433), .A2(SI_12_), .ZN(n5434) );
  NAND2_X1 U6886 ( .A1(n5459), .A2(n5434), .ZN(n5460) );
  NAND2_X1 U6887 ( .A1(n6811), .A2(n8132), .ZN(n5441) );
  NAND2_X1 U6888 ( .A1(n5435), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5437) );
  INV_X1 U6889 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U6890 ( .A1(n5437), .A2(n5436), .ZN(n5465) );
  OR2_X1 U6891 ( .A1(n5437), .A2(n5436), .ZN(n5438) );
  NAND2_X1 U6892 ( .A1(n5465), .A2(n5438), .ZN(n7494) );
  OAI22_X1 U6893 ( .A1(n5622), .A2(n6813), .B1(n9755), .B2(n7494), .ZN(n5439)
         );
  INV_X1 U6894 ( .A(n5439), .ZN(n5440) );
  NAND2_X1 U6895 ( .A1(n7851), .A2(n4475), .ZN(n5450) );
  NAND2_X1 U6896 ( .A1(n5382), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U6897 ( .A1(n5210), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5447) );
  INV_X1 U6898 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U6899 ( .A1(n5443), .A2(n5442), .ZN(n5444) );
  AND2_X1 U6900 ( .A1(n5469), .A2(n5444), .ZN(n7791) );
  NAND2_X1 U6901 ( .A1(n5845), .A2(n7791), .ZN(n5446) );
  NAND2_X1 U6902 ( .A1(n8133), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5445) );
  NAND4_X1 U6903 ( .A1(n5448), .A2(n5447), .A3(n5446), .A4(n5445), .ZN(n9704)
         );
  NAND2_X1 U6904 ( .A1(n9704), .A2(n5852), .ZN(n5449) );
  NAND2_X1 U6905 ( .A1(n5450), .A2(n5449), .ZN(n5451) );
  XNOR2_X1 U6906 ( .A(n5451), .B(n5855), .ZN(n5453) );
  AND2_X1 U6907 ( .A1(n9704), .A2(n5878), .ZN(n5452) );
  AOI21_X1 U6908 ( .B1(n7851), .B2(n5852), .A(n5452), .ZN(n5454) );
  NAND2_X1 U6909 ( .A1(n5453), .A2(n5454), .ZN(n5458) );
  INV_X1 U6910 ( .A(n5453), .ZN(n5456) );
  INV_X1 U6911 ( .A(n5454), .ZN(n5455) );
  NAND2_X1 U6912 ( .A1(n5456), .A2(n5455), .ZN(n5457) );
  AND2_X1 U6913 ( .A1(n5458), .A2(n5457), .ZN(n7786) );
  MUX2_X1 U6914 ( .A(n6905), .B(n6903), .S(n6633), .Z(n5462) );
  INV_X1 U6915 ( .A(SI_13_), .ZN(n5461) );
  INV_X1 U6916 ( .A(n5462), .ZN(n5463) );
  NAND2_X1 U6917 ( .A1(n5463), .A2(SI_13_), .ZN(n5464) );
  XNOR2_X1 U6918 ( .A(n5485), .B(n5051), .ZN(n6902) );
  NAND2_X1 U6919 ( .A1(n6902), .A2(n8132), .ZN(n5468) );
  NAND2_X1 U6920 ( .A1(n5465), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5466) );
  XNOR2_X1 U6921 ( .A(n5466), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9858) );
  AOI22_X1 U6922 ( .A1(n8131), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5594), .B2(
        n9858), .ZN(n5467) );
  NAND2_X1 U6923 ( .A1(n9712), .A2(n4475), .ZN(n5477) );
  NAND2_X1 U6924 ( .A1(n8133), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U6925 ( .A1(n5382), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5474) );
  INV_X1 U6926 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7798) );
  AND2_X1 U6927 ( .A1(n5469), .A2(n7798), .ZN(n5470) );
  OR2_X1 U6928 ( .A1(n5494), .A2(n5470), .ZN(n9694) );
  INV_X1 U6929 ( .A(n9694), .ZN(n5471) );
  NAND2_X1 U6930 ( .A1(n5845), .A2(n5471), .ZN(n5473) );
  NAND2_X1 U6931 ( .A1(n5210), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5472) );
  NAND4_X1 U6932 ( .A1(n5475), .A2(n5474), .A3(n5473), .A4(n5472), .ZN(n9204)
         );
  NAND2_X1 U6933 ( .A1(n9204), .A2(n5852), .ZN(n5476) );
  NAND2_X1 U6934 ( .A1(n5477), .A2(n5476), .ZN(n5478) );
  XNOR2_X1 U6935 ( .A(n5478), .B(n5855), .ZN(n5481) );
  AND2_X1 U6936 ( .A1(n9204), .A2(n5878), .ZN(n5479) );
  AOI21_X1 U6937 ( .B1(n9712), .B2(n5882), .A(n5479), .ZN(n5482) );
  AND2_X1 U6938 ( .A1(n5481), .A2(n5482), .ZN(n7794) );
  INV_X1 U6939 ( .A(n7794), .ZN(n5480) );
  INV_X1 U6940 ( .A(n5481), .ZN(n5484) );
  INV_X1 U6941 ( .A(n5482), .ZN(n5483) );
  NAND2_X1 U6942 ( .A1(n5484), .A2(n5483), .ZN(n7795) );
  INV_X1 U6943 ( .A(n5508), .ZN(n5504) );
  MUX2_X1 U6944 ( .A(n6948), .B(n6946), .S(n6633), .Z(n5510) );
  XNOR2_X1 U6945 ( .A(n5510), .B(SI_14_), .ZN(n5509) );
  XNOR2_X1 U6946 ( .A(n5513), .B(n5509), .ZN(n6945) );
  NAND2_X1 U6947 ( .A1(n6945), .A2(n8132), .ZN(n5493) );
  NOR2_X1 U6948 ( .A1(n5487), .A2(n9590), .ZN(n5488) );
  MUX2_X1 U6949 ( .A(n9590), .B(n5488), .S(P1_IR_REG_14__SCAN_IN), .Z(n5490)
         );
  OAI22_X1 U6950 ( .A1(n5622), .A2(n6946), .B1(n9755), .B2(n9238), .ZN(n5491)
         );
  INV_X1 U6951 ( .A(n5491), .ZN(n5492) );
  NAND2_X1 U6952 ( .A1(n8082), .A2(n4475), .ZN(n5501) );
  NAND2_X1 U6953 ( .A1(n5382), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U6954 ( .A1(n5210), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5498) );
  OR2_X1 U6955 ( .A1(n5494), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5495) );
  AND2_X1 U6956 ( .A1(n5495), .A2(n5522), .ZN(n7902) );
  NAND2_X1 U6957 ( .A1(n5845), .A2(n7902), .ZN(n5497) );
  NAND2_X1 U6958 ( .A1(n8133), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5496) );
  NAND4_X1 U6959 ( .A1(n5499), .A2(n5498), .A3(n5497), .A4(n5496), .ZN(n9703)
         );
  NAND2_X1 U6960 ( .A1(n9703), .A2(n5852), .ZN(n5500) );
  NAND2_X1 U6961 ( .A1(n5501), .A2(n5500), .ZN(n5502) );
  XNOR2_X1 U6962 ( .A(n5502), .B(n7257), .ZN(n5507) );
  INV_X1 U6963 ( .A(n5507), .ZN(n5503) );
  NAND2_X1 U6964 ( .A1(n8082), .A2(n5852), .ZN(n5506) );
  NAND2_X1 U6965 ( .A1(n9703), .A2(n5878), .ZN(n5505) );
  NAND2_X1 U6966 ( .A1(n5506), .A2(n5505), .ZN(n7901) );
  NAND2_X1 U6967 ( .A1(n5508), .A2(n5507), .ZN(n5533) );
  INV_X1 U6968 ( .A(n5510), .ZN(n5511) );
  NAND2_X1 U6969 ( .A1(n5511), .A2(SI_14_), .ZN(n5512) );
  MUX2_X1 U6970 ( .A(n7002), .B(n7003), .S(n6633), .Z(n5515) );
  INV_X1 U6971 ( .A(SI_15_), .ZN(n5514) );
  INV_X1 U6972 ( .A(n5515), .ZN(n5516) );
  NAND2_X1 U6973 ( .A1(n5516), .A2(SI_15_), .ZN(n5517) );
  XNOR2_X1 U6974 ( .A(n5539), .B(n5538), .ZN(n7001) );
  NAND2_X1 U6975 ( .A1(n7001), .A2(n8132), .ZN(n5521) );
  NAND2_X1 U6976 ( .A1(n5489), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5518) );
  XNOR2_X1 U6977 ( .A(n5518), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9870) );
  INV_X1 U6978 ( .A(n9870), .ZN(n9240) );
  OAI22_X1 U6979 ( .A1(n5622), .A2(n7003), .B1(n9755), .B2(n9240), .ZN(n5519)
         );
  INV_X1 U6980 ( .A(n5519), .ZN(n5520) );
  NAND2_X1 U6981 ( .A1(n9682), .A2(n4475), .ZN(n5528) );
  NAND2_X1 U6982 ( .A1(n5210), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U6983 ( .A1(n8133), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5525) );
  INV_X1 U6984 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7921) );
  AOI21_X1 U6985 ( .B1(n7921), .B2(n5522), .A(n5547), .ZN(n9680) );
  NAND2_X1 U6986 ( .A1(n5845), .A2(n9680), .ZN(n5524) );
  NAND2_X1 U6987 ( .A1(n5382), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5523) );
  NAND4_X1 U6988 ( .A1(n5526), .A2(n5525), .A3(n5524), .A4(n5523), .ZN(n9203)
         );
  NAND2_X1 U6989 ( .A1(n9203), .A2(n5852), .ZN(n5527) );
  NAND2_X1 U6990 ( .A1(n5528), .A2(n5527), .ZN(n5529) );
  XNOR2_X1 U6991 ( .A(n5529), .B(n5855), .ZN(n5535) );
  NAND2_X1 U6992 ( .A1(n9682), .A2(n5852), .ZN(n5532) );
  NAND2_X1 U6993 ( .A1(n9203), .A2(n5878), .ZN(n5531) );
  NAND2_X1 U6994 ( .A1(n5532), .A2(n5531), .ZN(n7918) );
  INV_X1 U6995 ( .A(n5535), .ZN(n5536) );
  INV_X1 U6996 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5540) );
  MUX2_X1 U6997 ( .A(n5540), .B(n7008), .S(n6633), .Z(n5541) );
  INV_X1 U6998 ( .A(SI_16_), .ZN(n10338) );
  NAND2_X1 U6999 ( .A1(n5541), .A2(n10338), .ZN(n5561) );
  INV_X1 U7000 ( .A(n5541), .ZN(n5542) );
  NAND2_X1 U7001 ( .A1(n5542), .A2(SI_16_), .ZN(n5543) );
  XNOR2_X1 U7002 ( .A(n5560), .B(n5559), .ZN(n7005) );
  NAND2_X1 U7003 ( .A1(n7005), .A2(n8132), .ZN(n5546) );
  OR2_X1 U7004 ( .A1(n5489), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7005 ( .A1(n5544), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5565) );
  XNOR2_X1 U7006 ( .A(n5565), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9882) );
  AOI22_X1 U7007 ( .A1(n8131), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5594), .B2(
        n9882), .ZN(n5545) );
  NAND2_X1 U7008 ( .A1(n8372), .A2(n4475), .ZN(n5553) );
  OAI21_X1 U7009 ( .B1(n5547), .B2(P1_REG3_REG_16__SCAN_IN), .A(n5573), .ZN(
        n7974) );
  INV_X1 U7010 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9235) );
  NAND2_X1 U7011 ( .A1(n8133), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U7012 ( .A1(n5382), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5548) );
  OAI211_X1 U7013 ( .C1(n5932), .C2(n9235), .A(n5549), .B(n5548), .ZN(n5550)
         );
  INV_X1 U7014 ( .A(n5550), .ZN(n5551) );
  OAI21_X1 U7015 ( .B1(n7974), .B2(n5928), .A(n5551), .ZN(n9463) );
  NAND2_X1 U7016 ( .A1(n9463), .A2(n5882), .ZN(n5552) );
  NAND2_X1 U7017 ( .A1(n5553), .A2(n5552), .ZN(n5554) );
  XNOR2_X1 U7018 ( .A(n5554), .B(n7257), .ZN(n7967) );
  NAND2_X1 U7019 ( .A1(n8372), .A2(n5852), .ZN(n5556) );
  NAND2_X1 U7020 ( .A1(n9463), .A2(n5878), .ZN(n5555) );
  NAND2_X1 U7021 ( .A1(n5556), .A2(n5555), .ZN(n7968) );
  NAND2_X1 U7022 ( .A1(n7970), .A2(n7967), .ZN(n5557) );
  NAND2_X1 U7023 ( .A1(n5560), .A2(n5559), .ZN(n5562) );
  MUX2_X1 U7024 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n4473), .Z(n5588) );
  INV_X1 U7025 ( .A(SI_17_), .ZN(n5563) );
  XNOR2_X1 U7026 ( .A(n5588), .B(n5563), .ZN(n5587) );
  XNOR2_X1 U7027 ( .A(n5591), .B(n5587), .ZN(n7059) );
  NAND2_X1 U7028 ( .A1(n7059), .A2(n8132), .ZN(n5571) );
  NAND2_X1 U7029 ( .A1(n5565), .A2(n5564), .ZN(n5566) );
  NAND2_X1 U7030 ( .A1(n5566), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U7031 ( .A1(n5568), .A2(n5567), .ZN(n5592) );
  OR2_X1 U7032 ( .A1(n5568), .A2(n5567), .ZN(n5569) );
  AOI22_X1 U7033 ( .A1(n8131), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5594), .B2(
        n9234), .ZN(n5570) );
  NAND2_X1 U7034 ( .A1(n9474), .A2(n5196), .ZN(n5581) );
  INV_X1 U7035 ( .A(n5573), .ZN(n5572) );
  INV_X1 U7036 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9137) );
  NAND2_X1 U7037 ( .A1(n5573), .A2(n9137), .ZN(n5574) );
  NAND2_X1 U7038 ( .A1(n5599), .A2(n5574), .ZN(n9476) );
  OR2_X1 U7039 ( .A1(n9476), .A2(n5928), .ZN(n5579) );
  INV_X1 U7040 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10394) );
  NAND2_X1 U7041 ( .A1(n5382), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7042 ( .A1(n8133), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5575) );
  OAI211_X1 U7043 ( .C1(n5932), .C2(n10394), .A(n5576), .B(n5575), .ZN(n5577)
         );
  INV_X1 U7044 ( .A(n5577), .ZN(n5578) );
  NAND2_X1 U7045 ( .A1(n5579), .A2(n5578), .ZN(n9443) );
  NAND2_X1 U7046 ( .A1(n9443), .A2(n5852), .ZN(n5580) );
  NAND2_X1 U7047 ( .A1(n5581), .A2(n5580), .ZN(n5582) );
  XNOR2_X1 U7048 ( .A(n5582), .B(n5855), .ZN(n5585) );
  AND2_X1 U7049 ( .A1(n9443), .A2(n5878), .ZN(n5583) );
  AOI21_X1 U7050 ( .B1(n9474), .B2(n5852), .A(n5583), .ZN(n5584) );
  XNOR2_X1 U7051 ( .A(n5585), .B(n5584), .ZN(n9135) );
  NAND2_X1 U7052 ( .A1(n5585), .A2(n5584), .ZN(n5586) );
  INV_X1 U7053 ( .A(n5613), .ZN(n5610) );
  INV_X1 U7054 ( .A(n5587), .ZN(n5590) );
  NAND2_X1 U7055 ( .A1(n5588), .A2(SI_17_), .ZN(n5589) );
  MUX2_X1 U7056 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5131), .Z(n5617) );
  XNOR2_X1 U7057 ( .A(n5617), .B(SI_18_), .ZN(n5614) );
  XNOR2_X1 U7058 ( .A(n5616), .B(n5614), .ZN(n7262) );
  NAND2_X1 U7059 ( .A1(n7262), .A2(n8132), .ZN(n5596) );
  NAND2_X1 U7060 ( .A1(n5592), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5593) );
  XNOR2_X1 U7061 ( .A(n5593), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9233) );
  AOI22_X1 U7062 ( .A1(n8131), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9233), .B2(
        n5594), .ZN(n5595) );
  NAND2_X1 U7063 ( .A1(n9452), .A2(n4475), .ZN(n5607) );
  INV_X1 U7064 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U7065 ( .A1(n5599), .A2(n5598), .ZN(n5600) );
  NAND2_X1 U7066 ( .A1(n5627), .A2(n5600), .ZN(n9453) );
  OR2_X1 U7067 ( .A1(n9453), .A2(n5928), .ZN(n5605) );
  INV_X1 U7068 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9454) );
  NAND2_X1 U7069 ( .A1(n5210), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5602) );
  NAND2_X1 U7070 ( .A1(n5382), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5601) );
  OAI211_X1 U7071 ( .C1(n5784), .C2(n9454), .A(n5602), .B(n5601), .ZN(n5603)
         );
  INV_X1 U7072 ( .A(n5603), .ZN(n5604) );
  NAND2_X1 U7073 ( .A1(n5605), .A2(n5604), .ZN(n9464) );
  NAND2_X1 U7074 ( .A1(n9464), .A2(n5882), .ZN(n5606) );
  NAND2_X1 U7075 ( .A1(n5607), .A2(n5606), .ZN(n5608) );
  XNOR2_X1 U7076 ( .A(n5608), .B(n5855), .ZN(n5612) );
  INV_X1 U7077 ( .A(n5612), .ZN(n5609) );
  NAND2_X1 U7078 ( .A1(n5610), .A2(n5609), .ZN(n9177) );
  AND2_X1 U7079 ( .A1(n9464), .A2(n5878), .ZN(n5611) );
  AOI21_X1 U7080 ( .B1(n9452), .B2(n5852), .A(n5611), .ZN(n9175) );
  INV_X1 U7081 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8427) );
  MUX2_X1 U7082 ( .A(n8427), .B(n7358), .S(n4473), .Z(n5619) );
  INV_X1 U7083 ( .A(SI_19_), .ZN(n5618) );
  INV_X1 U7084 ( .A(n5619), .ZN(n5620) );
  NAND2_X1 U7085 ( .A1(n5620), .A2(SI_19_), .ZN(n5621) );
  NAND2_X1 U7086 ( .A1(n5642), .A2(n5621), .ZN(n5643) );
  XNOR2_X1 U7087 ( .A(n5644), .B(n5643), .ZN(n7357) );
  NAND2_X1 U7088 ( .A1(n7357), .A2(n8132), .ZN(n5625) );
  OAI22_X1 U7089 ( .A1(n5622), .A2(n7358), .B1(n9430), .B2(n9755), .ZN(n5623)
         );
  INV_X1 U7090 ( .A(n5623), .ZN(n5624) );
  NAND2_X1 U7091 ( .A1(n9431), .A2(n5196), .ZN(n5635) );
  INV_X1 U7092 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U7093 ( .A1(n5627), .A2(n5626), .ZN(n5628) );
  AND2_X1 U7094 ( .A1(n5653), .A2(n5628), .ZN(n9420) );
  NAND2_X1 U7095 ( .A1(n9420), .A2(n5845), .ZN(n5633) );
  INV_X1 U7096 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9232) );
  NAND2_X1 U7097 ( .A1(n5382), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U7098 ( .A1(n5210), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5629) );
  OAI211_X1 U7099 ( .C1(n5784), .C2(n9232), .A(n5630), .B(n5629), .ZN(n5631)
         );
  INV_X1 U7100 ( .A(n5631), .ZN(n5632) );
  NAND2_X1 U7101 ( .A1(n5633), .A2(n5632), .ZN(n9444) );
  NAND2_X1 U7102 ( .A1(n9444), .A2(n5852), .ZN(n5634) );
  NAND2_X1 U7103 ( .A1(n5635), .A2(n5634), .ZN(n5636) );
  XNOR2_X1 U7104 ( .A(n5636), .B(n7257), .ZN(n5638) );
  AND2_X1 U7105 ( .A1(n9444), .A2(n5878), .ZN(n5637) );
  AOI21_X1 U7106 ( .B1(n9431), .B2(n5852), .A(n5637), .ZN(n5639) );
  XNOR2_X1 U7107 ( .A(n5638), .B(n5639), .ZN(n9113) );
  INV_X1 U7108 ( .A(n5638), .ZN(n5640) );
  NAND2_X1 U7109 ( .A1(n5640), .A2(n5639), .ZN(n5641) );
  OAI21_X2 U7110 ( .B1(n5644), .B2(n5643), .A(n5642), .ZN(n5666) );
  INV_X1 U7111 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7549) );
  INV_X1 U7112 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7515) );
  MUX2_X1 U7113 ( .A(n7549), .B(n7515), .S(n6633), .Z(n5646) );
  INV_X1 U7114 ( .A(SI_20_), .ZN(n5645) );
  NAND2_X1 U7115 ( .A1(n5646), .A2(n5645), .ZN(n5667) );
  INV_X1 U7116 ( .A(n5646), .ZN(n5647) );
  NAND2_X1 U7117 ( .A1(n5647), .A2(SI_20_), .ZN(n5648) );
  XNOR2_X1 U7118 ( .A(n5666), .B(n5665), .ZN(n7514) );
  NAND2_X1 U7119 ( .A1(n7514), .A2(n8132), .ZN(n5650) );
  NAND2_X1 U7120 ( .A1(n8131), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5649) );
  NAND2_X2 U7121 ( .A1(n5650), .A2(n5649), .ZN(n9408) );
  NAND2_X1 U7122 ( .A1(n9408), .A2(n5196), .ZN(n5661) );
  INV_X1 U7123 ( .A(n5653), .ZN(n5651) );
  INV_X1 U7124 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U7125 ( .A1(n5653), .A2(n5652), .ZN(n5654) );
  NAND2_X1 U7126 ( .A1(n5671), .A2(n5654), .ZN(n9409) );
  OR2_X1 U7127 ( .A1(n9409), .A2(n5928), .ZN(n5659) );
  INV_X1 U7128 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9527) );
  NAND2_X1 U7129 ( .A1(n5382), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U7130 ( .A1(n8133), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5655) );
  OAI211_X1 U7131 ( .C1(n5932), .C2(n9527), .A(n5656), .B(n5655), .ZN(n5657)
         );
  INV_X1 U7132 ( .A(n5657), .ZN(n5658) );
  NAND2_X1 U7133 ( .A1(n5659), .A2(n5658), .ZN(n9202) );
  NAND2_X1 U7134 ( .A1(n9202), .A2(n5852), .ZN(n5660) );
  NAND2_X1 U7135 ( .A1(n5661), .A2(n5660), .ZN(n5662) );
  XNOR2_X1 U7136 ( .A(n5662), .B(n7257), .ZN(n5688) );
  NAND2_X1 U7137 ( .A1(n9408), .A2(n5852), .ZN(n5664) );
  NAND2_X1 U7138 ( .A1(n9202), .A2(n5878), .ZN(n5663) );
  NAND2_X1 U7139 ( .A1(n5664), .A2(n5663), .ZN(n5689) );
  NAND2_X1 U7140 ( .A1(n5688), .A2(n5689), .ZN(n9154) );
  INV_X1 U7141 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7587) );
  INV_X1 U7142 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8060) );
  MUX2_X1 U7143 ( .A(n7587), .B(n8060), .S(n6633), .Z(n5696) );
  XNOR2_X1 U7144 ( .A(n5696), .B(SI_21_), .ZN(n5695) );
  NAND2_X1 U7145 ( .A1(n8131), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U7146 ( .A1(n9519), .A2(n4475), .ZN(n5679) );
  INV_X1 U7147 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U7148 ( .A1(n5671), .A2(n5670), .ZN(n5672) );
  AND2_X1 U7149 ( .A1(n5708), .A2(n5672), .ZN(n9374) );
  NAND2_X1 U7150 ( .A1(n9374), .A2(n5845), .ZN(n5677) );
  INV_X1 U7151 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10404) );
  NAND2_X1 U7152 ( .A1(n5210), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U7153 ( .A1(n8133), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5673) );
  OAI211_X1 U7154 ( .C1(n5848), .C2(n10404), .A(n5674), .B(n5673), .ZN(n5675)
         );
  INV_X1 U7155 ( .A(n5675), .ZN(n5676) );
  NAND2_X1 U7156 ( .A1(n5677), .A2(n5676), .ZN(n9402) );
  NAND2_X1 U7157 ( .A1(n9402), .A2(n5852), .ZN(n5678) );
  NAND2_X1 U7158 ( .A1(n5679), .A2(n5678), .ZN(n5680) );
  XNOR2_X1 U7159 ( .A(n5680), .B(n7257), .ZN(n5684) );
  INV_X1 U7160 ( .A(n5684), .ZN(n5682) );
  AND2_X1 U7161 ( .A1(n9402), .A2(n5878), .ZN(n5681) );
  AOI21_X1 U7162 ( .B1(n9519), .B2(n5882), .A(n5681), .ZN(n5683) );
  NAND2_X1 U7163 ( .A1(n5682), .A2(n5683), .ZN(n5692) );
  INV_X1 U7164 ( .A(n5692), .ZN(n5685) );
  XNOR2_X1 U7165 ( .A(n5684), .B(n5683), .ZN(n9120) );
  AND2_X1 U7166 ( .A1(n9154), .A2(n5687), .ZN(n5686) );
  INV_X1 U7167 ( .A(n5687), .ZN(n5694) );
  INV_X1 U7168 ( .A(n5688), .ZN(n5691) );
  INV_X1 U7169 ( .A(n5689), .ZN(n5690) );
  NAND2_X1 U7170 ( .A1(n5691), .A2(n5690), .ZN(n9156) );
  AND2_X1 U7171 ( .A1(n9156), .A2(n5692), .ZN(n5693) );
  INV_X1 U7172 ( .A(n5696), .ZN(n5697) );
  NAND2_X1 U7173 ( .A1(n5697), .A2(SI_21_), .ZN(n5698) );
  NAND2_X1 U7174 ( .A1(n5699), .A2(n5698), .ZN(n5724) );
  INV_X1 U7175 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7623) );
  MUX2_X1 U7176 ( .A(n10341), .B(n7623), .S(n6633), .Z(n5701) );
  INV_X1 U7177 ( .A(SI_22_), .ZN(n5700) );
  NAND2_X1 U7178 ( .A1(n5701), .A2(n5700), .ZN(n5722) );
  INV_X1 U7179 ( .A(n5701), .ZN(n5702) );
  NAND2_X1 U7180 ( .A1(n5702), .A2(SI_22_), .ZN(n5703) );
  NAND2_X1 U7181 ( .A1(n5722), .A2(n5703), .ZN(n5723) );
  XNOR2_X1 U7182 ( .A(n5724), .B(n5723), .ZN(n7621) );
  NAND2_X1 U7183 ( .A1(n7621), .A2(n8132), .ZN(n5705) );
  NAND2_X1 U7184 ( .A1(n8131), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5704) );
  INV_X1 U7185 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U7186 ( .A1(n5708), .A2(n5707), .ZN(n5709) );
  NAND2_X1 U7187 ( .A1(n5735), .A2(n5709), .ZN(n9361) );
  OR2_X1 U7188 ( .A1(n9361), .A2(n5928), .ZN(n5715) );
  INV_X1 U7189 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U7190 ( .A1(n8133), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U7191 ( .A1(n5382), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5710) );
  OAI211_X1 U7192 ( .C1(n5712), .C2(n5932), .A(n5711), .B(n5710), .ZN(n5713)
         );
  INV_X1 U7193 ( .A(n5713), .ZN(n5714) );
  NAND2_X1 U7194 ( .A1(n5715), .A2(n5714), .ZN(n9351) );
  AND2_X1 U7195 ( .A1(n9351), .A2(n5878), .ZN(n5716) );
  AOI21_X1 U7196 ( .B1(n9514), .B2(n5852), .A(n5716), .ZN(n5720) );
  NAND2_X1 U7197 ( .A1(n9514), .A2(n5196), .ZN(n5718) );
  NAND2_X1 U7198 ( .A1(n9351), .A2(n5882), .ZN(n5717) );
  NAND2_X1 U7199 ( .A1(n5718), .A2(n5717), .ZN(n5719) );
  XNOR2_X1 U7200 ( .A(n5719), .B(n7257), .ZN(n9166) );
  INV_X1 U7201 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n10218) );
  INV_X1 U7202 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5725) );
  MUX2_X1 U7203 ( .A(n10218), .B(n5725), .S(n6633), .Z(n5727) );
  INV_X1 U7204 ( .A(SI_23_), .ZN(n5726) );
  NAND2_X1 U7205 ( .A1(n5727), .A2(n5726), .ZN(n5750) );
  INV_X1 U7206 ( .A(n5727), .ZN(n5728) );
  NAND2_X1 U7207 ( .A1(n5728), .A2(SI_23_), .ZN(n5729) );
  NAND2_X1 U7208 ( .A1(n5731), .A2(n5730), .ZN(n5751) );
  OR2_X1 U7209 ( .A1(n5731), .A2(n5730), .ZN(n5732) );
  NAND2_X1 U7210 ( .A1(n5751), .A2(n5732), .ZN(n7782) );
  NAND2_X1 U7211 ( .A1(n7782), .A2(n8132), .ZN(n5734) );
  NAND2_X1 U7212 ( .A1(n8131), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U7213 ( .A1(n9509), .A2(n5196), .ZN(n5744) );
  INV_X1 U7214 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9106) );
  OR2_X2 U7215 ( .A1(n5735), .A2(n9106), .ZN(n5755) );
  NAND2_X1 U7216 ( .A1(n5735), .A2(n9106), .ZN(n5736) );
  NAND2_X1 U7217 ( .A1(n5755), .A2(n5736), .ZN(n9344) );
  OR2_X1 U7218 ( .A1(n9344), .A2(n5928), .ZN(n5742) );
  INV_X1 U7219 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U7220 ( .A1(n5382), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U7221 ( .A1(n5210), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5737) );
  OAI211_X1 U7222 ( .C1(n5784), .C2(n5739), .A(n5738), .B(n5737), .ZN(n5740)
         );
  INV_X1 U7223 ( .A(n5740), .ZN(n5741) );
  NAND2_X1 U7224 ( .A1(n5742), .A2(n5741), .ZN(n9367) );
  NAND2_X1 U7225 ( .A1(n9367), .A2(n5852), .ZN(n5743) );
  NAND2_X1 U7226 ( .A1(n5744), .A2(n5743), .ZN(n5745) );
  XNOR2_X1 U7227 ( .A(n5745), .B(n7257), .ZN(n5747) );
  NAND2_X1 U7228 ( .A1(n5748), .A2(n5747), .ZN(n9102) );
  AND2_X1 U7229 ( .A1(n9367), .A2(n5878), .ZN(n5746) );
  AOI21_X1 U7230 ( .B1(n9509), .B2(n5852), .A(n5746), .ZN(n9101) );
  NOR2_X1 U7231 ( .A1(n5748), .A2(n5747), .ZN(n5749) );
  INV_X1 U7232 ( .A(n5749), .ZN(n9103) );
  NAND2_X1 U7233 ( .A1(n9100), .A2(n9103), .ZN(n9126) );
  INV_X1 U7234 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7846) );
  INV_X1 U7235 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7848) );
  MUX2_X1 U7236 ( .A(n7846), .B(n7848), .S(n4473), .Z(n5770) );
  XNOR2_X1 U7237 ( .A(n5770), .B(SI_24_), .ZN(n5767) );
  XNOR2_X1 U7238 ( .A(n5769), .B(n5767), .ZN(n7845) );
  NAND2_X1 U7239 ( .A1(n7845), .A2(n8132), .ZN(n5753) );
  NAND2_X1 U7240 ( .A1(n8131), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U7241 ( .A1(n9331), .A2(n4475), .ZN(n5764) );
  INV_X1 U7242 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U7243 ( .A1(n5755), .A2(n5754), .ZN(n5756) );
  AND2_X1 U7244 ( .A1(n5780), .A2(n5756), .ZN(n9334) );
  NAND2_X1 U7245 ( .A1(n9334), .A2(n5845), .ZN(n5762) );
  INV_X1 U7246 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5759) );
  NAND2_X1 U7247 ( .A1(n5382), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U7248 ( .A1(n8133), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5757) );
  OAI211_X1 U7249 ( .C1(n5932), .C2(n5759), .A(n5758), .B(n5757), .ZN(n5760)
         );
  INV_X1 U7250 ( .A(n5760), .ZN(n5761) );
  NAND2_X1 U7251 ( .A1(n5762), .A2(n5761), .ZN(n9352) );
  NAND2_X1 U7252 ( .A1(n9352), .A2(n5852), .ZN(n5763) );
  NAND2_X1 U7253 ( .A1(n5764), .A2(n5763), .ZN(n5765) );
  XNOR2_X1 U7254 ( .A(n5765), .B(n7257), .ZN(n5798) );
  AND2_X1 U7255 ( .A1(n9352), .A2(n5878), .ZN(n5766) );
  AOI21_X1 U7256 ( .B1(n9331), .B2(n5882), .A(n5766), .ZN(n5799) );
  XNOR2_X1 U7257 ( .A(n5798), .B(n5799), .ZN(n9144) );
  INV_X1 U7258 ( .A(n5767), .ZN(n5768) );
  INV_X1 U7259 ( .A(n5770), .ZN(n5771) );
  NAND2_X1 U7260 ( .A1(n5771), .A2(SI_24_), .ZN(n5772) );
  INV_X1 U7261 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7895) );
  INV_X1 U7262 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10217) );
  MUX2_X1 U7263 ( .A(n7895), .B(n10217), .S(n6633), .Z(n5774) );
  INV_X1 U7264 ( .A(SI_25_), .ZN(n5773) );
  NAND2_X1 U7265 ( .A1(n5774), .A2(n5773), .ZN(n5806) );
  INV_X1 U7266 ( .A(n5774), .ZN(n5775) );
  NAND2_X1 U7267 ( .A1(n5775), .A2(SI_25_), .ZN(n5776) );
  NAND2_X1 U7268 ( .A1(n5806), .A2(n5776), .ZN(n5807) );
  NAND2_X1 U7269 ( .A1(n6393), .A2(n8132), .ZN(n5778) );
  NAND2_X1 U7270 ( .A1(n8131), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U7271 ( .A1(n9313), .A2(n5196), .ZN(n5789) );
  INV_X1 U7272 ( .A(n5780), .ZN(n5779) );
  NAND2_X1 U7273 ( .A1(n5779), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5817) );
  INV_X1 U7274 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10310) );
  NAND2_X1 U7275 ( .A1(n5780), .A2(n10310), .ZN(n5781) );
  NAND2_X1 U7276 ( .A1(n5817), .A2(n5781), .ZN(n9315) );
  INV_X1 U7277 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9314) );
  NAND2_X1 U7278 ( .A1(n5210), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U7279 ( .A1(n5382), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5782) );
  OAI211_X1 U7280 ( .C1(n5784), .C2(n9314), .A(n5783), .B(n5782), .ZN(n5785)
         );
  INV_X1 U7281 ( .A(n5785), .ZN(n5786) );
  NAND2_X1 U7282 ( .A1(n5787), .A2(n5786), .ZN(n9327) );
  NAND2_X1 U7283 ( .A1(n9327), .A2(n5882), .ZN(n5788) );
  NAND2_X1 U7284 ( .A1(n5789), .A2(n5788), .ZN(n5790) );
  XNOR2_X1 U7285 ( .A(n5790), .B(n7257), .ZN(n5794) );
  INV_X1 U7286 ( .A(n5794), .ZN(n5792) );
  AND2_X1 U7287 ( .A1(n9327), .A2(n5878), .ZN(n5791) );
  AOI21_X1 U7288 ( .B1(n9313), .B2(n5882), .A(n5791), .ZN(n5793) );
  NAND2_X1 U7289 ( .A1(n5792), .A2(n5793), .ZN(n5801) );
  INV_X1 U7290 ( .A(n5801), .ZN(n5795) );
  XNOR2_X1 U7291 ( .A(n5794), .B(n5793), .ZN(n9129) );
  AND2_X1 U7292 ( .A1(n9144), .A2(n5797), .ZN(n5796) );
  NAND2_X1 U7293 ( .A1(n9126), .A2(n5796), .ZN(n5805) );
  INV_X1 U7294 ( .A(n5797), .ZN(n5803) );
  INV_X1 U7295 ( .A(n5798), .ZN(n5800) );
  NAND2_X1 U7296 ( .A1(n5800), .A2(n5799), .ZN(n9127) );
  AND2_X1 U7297 ( .A1(n9127), .A2(n5801), .ZN(n5802) );
  NAND2_X1 U7298 ( .A1(n5805), .A2(n5804), .ZN(n9185) );
  INV_X1 U7299 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n10335) );
  INV_X1 U7300 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10321) );
  MUX2_X1 U7301 ( .A(n10335), .B(n10321), .S(n6633), .Z(n5810) );
  INV_X1 U7302 ( .A(SI_26_), .ZN(n5809) );
  NAND2_X1 U7303 ( .A1(n5810), .A2(n5809), .ZN(n5861) );
  INV_X1 U7304 ( .A(n5810), .ZN(n5811) );
  NAND2_X1 U7305 ( .A1(n5811), .A2(SI_26_), .ZN(n5812) );
  XNOR2_X1 U7306 ( .A(n5834), .B(n5833), .ZN(n7896) );
  NAND2_X1 U7307 ( .A1(n7896), .A2(n8132), .ZN(n5814) );
  NAND2_X1 U7308 ( .A1(n8131), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7309 ( .A1(n9494), .A2(n4475), .ZN(n5825) );
  INV_X1 U7310 ( .A(n5817), .ZN(n5815) );
  NAND2_X1 U7311 ( .A1(n5815), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5843) );
  INV_X1 U7312 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U7313 ( .A1(n5817), .A2(n5816), .ZN(n5818) );
  NAND2_X1 U7314 ( .A1(n5843), .A2(n5818), .ZN(n9190) );
  INV_X1 U7315 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10333) );
  NAND2_X1 U7316 ( .A1(n8133), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U7317 ( .A1(n5382), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5819) );
  OAI211_X1 U7318 ( .C1(n10333), .C2(n5932), .A(n5820), .B(n5819), .ZN(n5821)
         );
  INV_X1 U7319 ( .A(n5821), .ZN(n5822) );
  NAND2_X1 U7320 ( .A1(n9287), .A2(n5882), .ZN(n5824) );
  NAND2_X1 U7321 ( .A1(n5825), .A2(n5824), .ZN(n5826) );
  XNOR2_X1 U7322 ( .A(n5826), .B(n5855), .ZN(n5828) );
  AND2_X1 U7323 ( .A1(n9287), .A2(n5878), .ZN(n5827) );
  AOI21_X1 U7324 ( .B1(n9494), .B2(n5852), .A(n5827), .ZN(n5829) );
  XNOR2_X1 U7325 ( .A(n5828), .B(n5829), .ZN(n9187) );
  INV_X1 U7326 ( .A(n5828), .ZN(n5831) );
  INV_X1 U7327 ( .A(n5829), .ZN(n5830) );
  NAND2_X1 U7328 ( .A1(n5831), .A2(n5830), .ZN(n5832) );
  NAND2_X1 U7329 ( .A1(n5863), .A2(n5861), .ZN(n5839) );
  INV_X1 U7330 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7949) );
  INV_X1 U7331 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5835) );
  MUX2_X1 U7332 ( .A(n7949), .B(n5835), .S(n4473), .Z(n5836) );
  INV_X1 U7333 ( .A(SI_27_), .ZN(n10267) );
  NAND2_X1 U7334 ( .A1(n5836), .A2(n10267), .ZN(n5860) );
  INV_X1 U7335 ( .A(n5836), .ZN(n5837) );
  NAND2_X1 U7336 ( .A1(n5837), .A2(SI_27_), .ZN(n5864) );
  AND2_X1 U7337 ( .A1(n5860), .A2(n5864), .ZN(n5838) );
  NAND2_X1 U7338 ( .A1(n7945), .A2(n8132), .ZN(n5841) );
  NAND2_X1 U7339 ( .A1(n8131), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U7340 ( .A1(n9489), .A2(n5196), .ZN(n5854) );
  INV_X1 U7341 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5842) );
  NAND2_X1 U7342 ( .A1(n5843), .A2(n5842), .ZN(n5844) );
  NAND2_X1 U7343 ( .A1(n9282), .A2(n5845), .ZN(n5851) );
  INV_X1 U7344 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10405) );
  NAND2_X1 U7345 ( .A1(n8133), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U7346 ( .A1(n5210), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5846) );
  OAI211_X1 U7347 ( .C1(n5848), .C2(n10405), .A(n5847), .B(n5846), .ZN(n5849)
         );
  INV_X1 U7348 ( .A(n5849), .ZN(n5850) );
  NAND2_X1 U7349 ( .A1(n9304), .A2(n5852), .ZN(n5853) );
  NAND2_X1 U7350 ( .A1(n5854), .A2(n5853), .ZN(n5856) );
  XNOR2_X1 U7351 ( .A(n5856), .B(n5855), .ZN(n9092) );
  AND2_X1 U7352 ( .A1(n9304), .A2(n5878), .ZN(n5857) );
  AOI21_X1 U7353 ( .B1(n9489), .B2(n5882), .A(n5857), .ZN(n9091) );
  INV_X1 U7354 ( .A(n5914), .ZN(n5910) );
  INV_X1 U7355 ( .A(n9092), .ZN(n5858) );
  AND2_X1 U7356 ( .A1(n5861), .A2(n5860), .ZN(n5862) );
  NAND2_X1 U7357 ( .A1(n5863), .A2(n5862), .ZN(n5865) );
  INV_X1 U7358 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10290) );
  INV_X1 U7359 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5866) );
  MUX2_X1 U7360 ( .A(n10290), .B(n5866), .S(n4473), .Z(n6544) );
  XNOR2_X1 U7361 ( .A(n6544), .B(SI_28_), .ZN(n6541) );
  NAND2_X1 U7362 ( .A1(n7950), .A2(n8132), .ZN(n5868) );
  NAND2_X1 U7363 ( .A1(n8131), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U7364 ( .A1(n8420), .A2(n5852), .ZN(n5880) );
  INV_X1 U7365 ( .A(n5871), .ZN(n5869) );
  NAND2_X1 U7366 ( .A1(n5869), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9262) );
  INV_X1 U7367 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U7368 ( .A1(n5871), .A2(n5870), .ZN(n5872) );
  NAND2_X1 U7369 ( .A1(n9262), .A2(n5872), .ZN(n5921) );
  INV_X1 U7370 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10397) );
  NAND2_X1 U7371 ( .A1(n8133), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7372 ( .A1(n5382), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5873) );
  OAI211_X1 U7373 ( .C1(n10397), .C2(n5932), .A(n5874), .B(n5873), .ZN(n5875)
         );
  INV_X1 U7374 ( .A(n5875), .ZN(n5876) );
  NAND2_X1 U7375 ( .A1(n9288), .A2(n5878), .ZN(n5879) );
  NAND2_X1 U7376 ( .A1(n5880), .A2(n5879), .ZN(n5881) );
  XNOR2_X1 U7377 ( .A(n5881), .B(n7257), .ZN(n5884) );
  AOI22_X1 U7378 ( .A1(n8420), .A2(n5196), .B1(n5882), .B2(n9288), .ZN(n5883)
         );
  XNOR2_X1 U7379 ( .A(n5884), .B(n5883), .ZN(n5911) );
  NAND2_X1 U7380 ( .A1(n7892), .A2(P1_B_REG_SCAN_IN), .ZN(n5885) );
  MUX2_X1 U7381 ( .A(P1_B_REG_SCAN_IN), .B(n5885), .S(n7850), .Z(n5887) );
  NAND2_X1 U7382 ( .A1(n5887), .A2(n5886), .ZN(n9925) );
  INV_X1 U7383 ( .A(n7892), .ZN(n5888) );
  OAI22_X1 U7384 ( .A1(n9925), .A2(P1_D_REG_1__SCAN_IN), .B1(n5886), .B2(n5888), .ZN(n6859) );
  NOR4_X1 U7385 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5892) );
  NOR4_X1 U7386 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n5891) );
  NOR4_X1 U7387 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5890) );
  NOR4_X1 U7388 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5889) );
  NAND4_X1 U7389 ( .A1(n5892), .A2(n5891), .A3(n5890), .A4(n5889), .ZN(n5898)
         );
  NOR2_X1 U7390 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .ZN(
        n5896) );
  NOR4_X1 U7391 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5895) );
  NOR4_X1 U7392 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5894) );
  NOR4_X1 U7393 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n5893) );
  NAND4_X1 U7394 ( .A1(n5896), .A2(n5895), .A3(n5894), .A4(n5893), .ZN(n5897)
         );
  NOR2_X1 U7395 ( .A1(n5898), .A2(n5897), .ZN(n5899) );
  NOR2_X1 U7396 ( .A1(n9925), .A2(n5899), .ZN(n6858) );
  NOR2_X1 U7397 ( .A1(n6859), .A2(n6858), .ZN(n7048) );
  INV_X1 U7398 ( .A(n9925), .ZN(n5902) );
  INV_X1 U7399 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9930) );
  INV_X1 U7400 ( .A(n7850), .ZN(n5900) );
  NOR2_X1 U7401 ( .A1(n5886), .A2(n5900), .ZN(n5901) );
  NAND2_X1 U7402 ( .A1(n7048), .A2(n9928), .ZN(n6865) );
  NAND2_X1 U7403 ( .A1(n5903), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5905) );
  XNOR2_X1 U7404 ( .A(n5905), .B(n5904), .ZN(n7778) );
  AND2_X1 U7405 ( .A1(n7778), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7406 ( .A1(n8259), .A2(n5907), .ZN(n7052) );
  AND2_X1 U7407 ( .A1(n9976), .A2(n8262), .ZN(n5924) );
  INV_X1 U7408 ( .A(n5924), .ZN(n5908) );
  INV_X1 U7409 ( .A(n5911), .ZN(n5912) );
  NAND2_X1 U7410 ( .A1(n5912), .A2(n9660), .ZN(n5915) );
  INV_X1 U7411 ( .A(n5915), .ZN(n5913) );
  OR2_X1 U7412 ( .A1(n7199), .A2(n7200), .ZN(n8338) );
  OR2_X1 U7413 ( .A1(n7052), .A2(n5153), .ZN(n7053) );
  AOI21_X1 U7414 ( .B1(n8338), .B2(n7053), .A(n8337), .ZN(n5917) );
  NAND2_X1 U7415 ( .A1(n6865), .A2(n5917), .ZN(n5926) );
  AND2_X1 U7416 ( .A1(n5926), .A2(n7047), .ZN(n9659) );
  INV_X1 U7417 ( .A(n9304), .ZN(n8065) );
  INV_X1 U7418 ( .A(n8338), .ZN(n5936) );
  INV_X1 U7419 ( .A(n5919), .ZN(n6876) );
  NAND2_X1 U7420 ( .A1(n5936), .A2(n6876), .ZN(n5920) );
  INV_X1 U7421 ( .A(n5921), .ZN(n9272) );
  NAND3_X1 U7422 ( .A1(n5922), .A2(n6621), .A3(n7778), .ZN(n5923) );
  AOI21_X1 U7423 ( .B1(n6865), .B2(n5924), .A(n5923), .ZN(n5925) );
  OR2_X1 U7424 ( .A1(n5925), .A2(P1_U3084), .ZN(n5927) );
  AOI22_X1 U7425 ( .A1(n9272), .A2(n9191), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n5940) );
  OR2_X1 U7426 ( .A1(n9262), .A2(n5928), .ZN(n5935) );
  INV_X1 U7427 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7428 ( .A1(n5382), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5930) );
  NAND2_X1 U7429 ( .A1(n8133), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5929) );
  OAI211_X1 U7430 ( .C1(n5932), .C2(n5931), .A(n5930), .B(n5929), .ZN(n5933)
         );
  INV_X1 U7431 ( .A(n5933), .ZN(n5934) );
  NAND2_X1 U7432 ( .A1(n5935), .A2(n5934), .ZN(n9201) );
  NAND2_X1 U7433 ( .A1(n5936), .A2(n5919), .ZN(n5937) );
  NAND2_X1 U7434 ( .A1(n9201), .A2(n9196), .ZN(n5939) );
  OAI211_X1 U7435 ( .C1(n8065), .C2(n9193), .A(n5940), .B(n5939), .ZN(n5941)
         );
  AOI21_X1 U7436 ( .B1(n8420), .B2(n9170), .A(n5941), .ZN(n5942) );
  NAND4_X1 U7437 ( .A1(n5945), .A2(n5944), .A3(n5943), .A4(n5942), .ZN(
        P1_U3218) );
  INV_X1 U7438 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5946) );
  NAND4_X1 U7439 ( .A1(n6250), .A2(n5946), .A3(n6128), .A4(n6248), .ZN(n5982)
         );
  INV_X1 U7440 ( .A(n5982), .ZN(n5950) );
  NOR2_X1 U7441 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5947) );
  AND2_X1 U7442 ( .A1(n5981), .A2(n5947), .ZN(n5949) );
  NOR2_X1 U7443 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5948) );
  NAND2_X1 U7444 ( .A1(n5985), .A2(n6069), .ZN(n5953) );
  NOR2_X2 U7445 ( .A1(n6059), .A2(n5953), .ZN(n6111) );
  NOR2_X1 U7446 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5955) );
  NOR2_X1 U7447 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5954) );
  INV_X1 U7448 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7449 ( .A1(n7950), .A2(n6068), .ZN(n5964) );
  OR2_X1 U7450 ( .A1(n8436), .A2(n10290), .ZN(n5963) );
  INV_X1 U7451 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5966) );
  XNOR2_X2 U7452 ( .A(n5970), .B(n5966), .ZN(n9089) );
  INV_X1 U7453 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7089) );
  NAND2_X2 U7454 ( .A1(n8640), .A2(n9089), .ZN(n6361) );
  INV_X1 U7455 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U7456 ( .A1(n6438), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5975) );
  INV_X1 U7457 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10352) );
  NAND2_X1 U7458 ( .A1(n5978), .A2(n10398), .ZN(n6459) );
  INV_X1 U7459 ( .A(n8628), .ZN(n7622) );
  INV_X1 U7460 ( .A(n5978), .ZN(n5979) );
  NAND2_X1 U7461 ( .A1(n5979), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5980) );
  NAND3_X1 U7462 ( .A1(n5981), .A2(n6069), .A3(n5952), .ZN(n5983) );
  NOR2_X1 U7463 ( .A1(n5983), .A2(n5982), .ZN(n5986) );
  NAND4_X1 U7464 ( .A1(n6047), .A2(n5986), .A3(n5985), .A4(n5984), .ZN(n6233)
         );
  INV_X1 U7465 ( .A(n6233), .ZN(n5988) );
  INV_X1 U7466 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5987) );
  INV_X1 U7467 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5989) );
  INV_X1 U7468 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U7469 ( .A1(n5994), .A2(n5993), .ZN(n5990) );
  INV_X1 U7470 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5991) );
  AND2_X2 U7471 ( .A1(n10027), .A2(n8587), .ZN(n10035) );
  NAND2_X1 U7472 ( .A1(n6512), .A2(n6028), .ZN(n6001) );
  INV_X1 U7473 ( .A(n6001), .ZN(n5999) );
  XNOR2_X1 U7474 ( .A(n5994), .B(n5993), .ZN(n6487) );
  NAND2_X1 U7475 ( .A1(n8628), .A2(n6304), .ZN(n8620) );
  NAND3_X1 U7476 ( .A1(n6491), .A2(n8620), .A3(n8443), .ZN(n5995) );
  NAND2_X4 U7477 ( .A1(n5995), .A2(n6617), .ZN(n6428) );
  INV_X1 U7478 ( .A(n6428), .ZN(n5997) );
  INV_X1 U7479 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5996) );
  XNOR2_X1 U7480 ( .A(n5997), .B(n6581), .ZN(n6000) );
  INV_X1 U7481 ( .A(n6000), .ZN(n5998) );
  INV_X1 U7482 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7158) );
  INV_X1 U7483 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6002) );
  OR2_X1 U7484 ( .A1(n6361), .A2(n6002), .ZN(n6004) );
  INV_X1 U7485 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10008) );
  NAND2_X1 U7486 ( .A1(n4481), .A2(SI_0_), .ZN(n6008) );
  INV_X1 U7487 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7488 ( .A1(n6008), .A2(n6007), .ZN(n6010) );
  AND2_X1 U7489 ( .A1(n6010), .A2(n6009), .ZN(n9090) );
  MUX2_X1 U7490 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9090), .S(n6692), .Z(n10026)
         );
  INV_X1 U7491 ( .A(n6915), .ZN(n6011) );
  NAND2_X1 U7492 ( .A1(n6438), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6017) );
  INV_X1 U7493 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7149) );
  OR2_X1 U7494 ( .A1(n4482), .A2(n7149), .ZN(n6016) );
  INV_X1 U7495 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6700) );
  OR2_X1 U7496 ( .A1(n6022), .A2(n6700), .ZN(n6015) );
  INV_X1 U7497 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6013) );
  OR2_X1 U7498 ( .A1(n6361), .A2(n6013), .ZN(n6014) );
  NAND4_X1 U7499 ( .A1(n6017), .A2(n6016), .A3(n6015), .A4(n6014), .ZN(n6517)
         );
  NAND2_X1 U7500 ( .A1(n6517), .A2(n6028), .ZN(n6020) );
  OR2_X1 U7501 ( .A1(n6018), .A2(n5968), .ZN(n6019) );
  XNOR2_X1 U7502 ( .A(n6019), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9617) );
  INV_X1 U7503 ( .A(n9617), .ZN(n6647) );
  INV_X2 U7504 ( .A(n6428), .ZN(n6448) );
  XNOR2_X1 U7505 ( .A(n7152), .B(n6448), .ZN(n6021) );
  XNOR2_X1 U7506 ( .A(n6020), .B(n6021), .ZN(n6906) );
  NAND2_X1 U7507 ( .A1(n6498), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6027) );
  OR2_X1 U7508 ( .A1(n4482), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6026) );
  INV_X1 U7509 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6703) );
  OR2_X1 U7510 ( .A1(n6022), .A2(n6703), .ZN(n6025) );
  INV_X1 U7511 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6023) );
  OR2_X1 U7512 ( .A1(n6037), .A2(n6023), .ZN(n6024) );
  NAND2_X1 U7513 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4504), .ZN(n6029) );
  XNOR2_X1 U7514 ( .A(n6029), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6717) );
  INV_X1 U7515 ( .A(n6717), .ZN(n6710) );
  XNOR2_X1 U7516 ( .A(n6032), .B(n6033), .ZN(n6974) );
  NAND2_X1 U7517 ( .A1(n6973), .A2(n6974), .ZN(n6036) );
  INV_X1 U7518 ( .A(n6032), .ZN(n6034) );
  NAND2_X1 U7519 ( .A1(n6034), .A2(n6033), .ZN(n6035) );
  NAND2_X1 U7520 ( .A1(n6438), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6046) );
  INV_X1 U7521 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6720) );
  INV_X1 U7522 ( .A(n6063), .ZN(n6041) );
  INV_X1 U7523 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6039) );
  INV_X1 U7524 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U7525 ( .A1(n6039), .A2(n6038), .ZN(n6040) );
  NAND2_X1 U7526 ( .A1(n6041), .A2(n6040), .ZN(n7131) );
  OR2_X1 U7527 ( .A1(n4482), .A2(n7131), .ZN(n6044) );
  INV_X1 U7528 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6042) );
  OR2_X1 U7529 ( .A1(n6361), .A2(n6042), .ZN(n6043) );
  NAND4_X1 U7530 ( .A1(n6046), .A2(n6045), .A3(n6044), .A4(n6043), .ZN(n8722)
         );
  AND2_X1 U7531 ( .A1(n8722), .A2(n10078), .ZN(n6051) );
  OR2_X1 U7532 ( .A1(n6047), .A2(n5968), .ZN(n6048) );
  XNOR2_X1 U7533 ( .A(n6048), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6732) );
  INV_X1 U7534 ( .A(n6732), .ZN(n6725) );
  NAND2_X1 U7535 ( .A1(n6634), .A2(n6547), .ZN(n6050) );
  OR2_X1 U7536 ( .A1(n8436), .A2(n4596), .ZN(n6049) );
  OAI211_X1 U7537 ( .C1(n6692), .C2(n6725), .A(n6050), .B(n6049), .ZN(n7136)
         );
  XNOR2_X1 U7538 ( .A(n7136), .B(n6428), .ZN(n6052) );
  NAND2_X1 U7539 ( .A1(n6051), .A2(n6052), .ZN(n6055) );
  INV_X1 U7540 ( .A(n6051), .ZN(n6054) );
  INV_X1 U7541 ( .A(n6052), .ZN(n6053) );
  NAND2_X1 U7542 ( .A1(n6054), .A2(n6053), .ZN(n6057) );
  NAND2_X1 U7543 ( .A1(n6055), .A2(n6057), .ZN(n6984) );
  INV_X2 U7544 ( .A(n6692), .ZN(n6664) );
  NAND2_X1 U7545 ( .A1(n6059), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6070) );
  XNOR2_X1 U7546 ( .A(n6070), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6747) );
  AOI22_X1 U7547 ( .A1(n6305), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6664), .B2(
        n6747), .ZN(n6061) );
  NAND2_X1 U7548 ( .A1(n6640), .A2(n6547), .ZN(n6060) );
  XNOR2_X1 U7549 ( .A(n7069), .B(n6448), .ZN(n6091) );
  NAND2_X1 U7550 ( .A1(n6438), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6067) );
  OAI21_X1 U7551 ( .B1(n6063), .B2(P2_REG3_REG_5__SCAN_IN), .A(n6078), .ZN(
        n7164) );
  OR2_X1 U7552 ( .A1(n4482), .A2(n7164), .ZN(n6066) );
  INV_X1 U7553 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6064) );
  OR2_X1 U7554 ( .A1(n6361), .A2(n6064), .ZN(n6065) );
  NAND2_X1 U7555 ( .A1(n8721), .A2(n10078), .ZN(n6092) );
  XNOR2_X1 U7556 ( .A(n6091), .B(n6092), .ZN(n7033) );
  BUF_X4 U7557 ( .A(n6068), .Z(n6547) );
  NAND2_X1 U7558 ( .A1(n6650), .A2(n6547), .ZN(n6076) );
  NAND2_X1 U7559 ( .A1(n6070), .A2(n6069), .ZN(n6071) );
  NAND2_X1 U7560 ( .A1(n6071), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6073) );
  INV_X1 U7561 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7562 ( .A1(n6073), .A2(n6072), .ZN(n6098) );
  OR2_X1 U7563 ( .A1(n6073), .A2(n6072), .ZN(n6074) );
  AOI22_X1 U7564 ( .A1(n6305), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6664), .B2(
        n6844), .ZN(n6075) );
  NAND2_X1 U7565 ( .A1(n6076), .A2(n6075), .ZN(n7236) );
  XNOR2_X1 U7566 ( .A(n7236), .B(n6448), .ZN(n6085) );
  NAND2_X1 U7567 ( .A1(n6498), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6083) );
  INV_X1 U7568 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6750) );
  OR2_X1 U7569 ( .A1(n6022), .A2(n6750), .ZN(n6082) );
  AND2_X1 U7570 ( .A1(n6078), .A2(n6077), .ZN(n6079) );
  OR2_X1 U7571 ( .A1(n6079), .A2(n6102), .ZN(n7233) );
  OR2_X1 U7572 ( .A1(n4482), .A2(n7233), .ZN(n6081) );
  INV_X1 U7573 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7234) );
  OR2_X1 U7574 ( .A1(n6037), .A2(n7234), .ZN(n6080) );
  NAND4_X1 U7575 ( .A1(n6083), .A2(n6082), .A3(n6081), .A4(n6080), .ZN(n8720)
         );
  NAND2_X1 U7576 ( .A1(n8720), .A2(n10078), .ZN(n6086) );
  NAND2_X1 U7577 ( .A1(n6085), .A2(n6086), .ZN(n6090) );
  INV_X1 U7578 ( .A(n6090), .ZN(n6095) );
  OR2_X1 U7579 ( .A1(n7033), .A2(n6095), .ZN(n6084) );
  OR2_X2 U7580 ( .A1(n7034), .A2(n6084), .ZN(n6097) );
  INV_X1 U7581 ( .A(n6085), .ZN(n6088) );
  INV_X1 U7582 ( .A(n6086), .ZN(n6087) );
  NAND2_X1 U7583 ( .A1(n6088), .A2(n6087), .ZN(n6089) );
  AND2_X1 U7584 ( .A1(n6090), .A2(n6089), .ZN(n7040) );
  INV_X1 U7585 ( .A(n6091), .ZN(n6094) );
  INV_X1 U7586 ( .A(n6092), .ZN(n6093) );
  NAND2_X1 U7587 ( .A1(n6094), .A2(n6093), .ZN(n7035) );
  AND2_X1 U7588 ( .A1(n7040), .A2(n7035), .ZN(n7036) );
  OR2_X1 U7589 ( .A1(n6095), .A2(n7036), .ZN(n6096) );
  NAND2_X1 U7590 ( .A1(n6655), .A2(n6547), .ZN(n6101) );
  NAND2_X1 U7591 ( .A1(n6098), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6099) );
  XNOR2_X1 U7592 ( .A(n6099), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6950) );
  AOI22_X1 U7593 ( .A1(n6305), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6664), .B2(
        n6950), .ZN(n6100) );
  XNOR2_X1 U7594 ( .A(n7420), .B(n6448), .ZN(n6110) );
  NAND2_X1 U7595 ( .A1(n6438), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6108) );
  INV_X1 U7596 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6847) );
  OR2_X1 U7597 ( .A1(n6022), .A2(n6847), .ZN(n6107) );
  OR2_X1 U7598 ( .A1(n6102), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7599 ( .A1(n6116), .A2(n6103), .ZN(n7108) );
  OR2_X1 U7600 ( .A1(n4482), .A2(n7108), .ZN(n6106) );
  INV_X1 U7601 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6104) );
  OR2_X1 U7602 ( .A1(n6361), .A2(n6104), .ZN(n6105) );
  NAND4_X1 U7603 ( .A1(n6108), .A2(n6107), .A3(n6106), .A4(n6105), .ZN(n8719)
         );
  NAND2_X1 U7604 ( .A1(n8719), .A2(n10078), .ZN(n6109) );
  XNOR2_X1 U7605 ( .A(n6110), .B(n6109), .ZN(n7010) );
  NAND2_X1 U7606 ( .A1(n6659), .A2(n6547), .ZN(n6114) );
  OR2_X1 U7607 ( .A1(n6111), .A2(n5968), .ZN(n6112) );
  XNOR2_X1 U7608 ( .A(n6112), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7019) );
  AOI22_X1 U7609 ( .A1(n6305), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6664), .B2(
        n7019), .ZN(n6113) );
  NAND2_X2 U7610 ( .A1(n6114), .A2(n6113), .ZN(n10064) );
  XNOR2_X1 U7611 ( .A(n10064), .B(n6428), .ZN(n6125) );
  NAND2_X1 U7612 ( .A1(n6438), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6122) );
  INV_X1 U7613 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6958) );
  OR2_X1 U7614 ( .A1(n6022), .A2(n6958), .ZN(n6121) );
  NAND2_X1 U7615 ( .A1(n6116), .A2(n6115), .ZN(n6117) );
  NAND2_X1 U7616 ( .A1(n6132), .A2(n6117), .ZN(n7411) );
  OR2_X1 U7617 ( .A1(n4482), .A2(n7411), .ZN(n6120) );
  INV_X1 U7618 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6118) );
  OR2_X1 U7619 ( .A1(n6361), .A2(n6118), .ZN(n6119) );
  NAND4_X1 U7620 ( .A1(n6122), .A2(n6121), .A3(n6120), .A4(n6119), .ZN(n8718)
         );
  NAND2_X1 U7621 ( .A1(n8718), .A2(n10078), .ZN(n6123) );
  XNOR2_X1 U7622 ( .A(n6125), .B(n6123), .ZN(n7075) );
  INV_X1 U7623 ( .A(n6123), .ZN(n6124) );
  NAND2_X1 U7624 ( .A1(n6125), .A2(n6124), .ZN(n6126) );
  INV_X1 U7625 ( .A(n7321), .ZN(n6144) );
  NAND2_X1 U7626 ( .A1(n6127), .A2(n6547), .ZN(n6130) );
  AND2_X1 U7627 ( .A1(n6111), .A2(n6128), .ZN(n6184) );
  XNOR2_X1 U7628 ( .A(n6147), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7211) );
  AOI22_X1 U7629 ( .A1(n6305), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6664), .B2(
        n7211), .ZN(n6129) );
  NAND2_X1 U7630 ( .A1(n6498), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6137) );
  INV_X1 U7631 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7026) );
  OR2_X1 U7632 ( .A1(n6022), .A2(n7026), .ZN(n6136) );
  AND2_X1 U7633 ( .A1(n6132), .A2(n6131), .ZN(n6133) );
  OR2_X1 U7634 ( .A1(n6133), .A2(n6154), .ZN(n7480) );
  OR2_X1 U7635 ( .A1(n4482), .A2(n7480), .ZN(n6135) );
  INV_X1 U7636 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7481) );
  OR2_X1 U7637 ( .A1(n6037), .A2(n7481), .ZN(n6134) );
  NAND4_X1 U7638 ( .A1(n6137), .A2(n6136), .A3(n6135), .A4(n6134), .ZN(n8717)
         );
  NAND2_X1 U7639 ( .A1(n8717), .A2(n10078), .ZN(n6139) );
  NAND2_X1 U7640 ( .A1(n6138), .A2(n6139), .ZN(n6145) );
  INV_X1 U7641 ( .A(n6138), .ZN(n6141) );
  INV_X1 U7642 ( .A(n6139), .ZN(n6140) );
  NAND2_X1 U7643 ( .A1(n6141), .A2(n6140), .ZN(n6142) );
  NAND2_X1 U7644 ( .A1(n6145), .A2(n6142), .ZN(n7324) );
  NAND2_X1 U7645 ( .A1(n6144), .A2(n6143), .ZN(n7322) );
  NAND2_X1 U7646 ( .A1(n7322), .A2(n6145), .ZN(n7360) );
  NAND2_X1 U7647 ( .A1(n6678), .A2(n6547), .ZN(n6153) );
  INV_X1 U7648 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7649 ( .A1(n6147), .A2(n6146), .ZN(n6148) );
  NAND2_X1 U7650 ( .A1(n6148), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6150) );
  INV_X1 U7651 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6149) );
  OR2_X1 U7652 ( .A1(n6150), .A2(n6149), .ZN(n6151) );
  NAND2_X1 U7653 ( .A1(n6150), .A2(n6149), .ZN(n6166) );
  AOI22_X1 U7654 ( .A1(n6305), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6664), .B2(
        n7589), .ZN(n6152) );
  XNOR2_X1 U7655 ( .A(n7462), .B(n6448), .ZN(n6161) );
  NAND2_X1 U7656 ( .A1(n6438), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6160) );
  INV_X1 U7657 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7218) );
  OR2_X1 U7658 ( .A1(n6022), .A2(n7218), .ZN(n6159) );
  NOR2_X1 U7659 ( .A1(n6154), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6155) );
  OR2_X1 U7660 ( .A1(n6170), .A2(n6155), .ZN(n7459) );
  OR2_X1 U7661 ( .A1(n4482), .A2(n7459), .ZN(n6158) );
  INV_X1 U7662 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n6156) );
  OR2_X1 U7663 ( .A1(n6361), .A2(n6156), .ZN(n6157) );
  NAND4_X1 U7664 ( .A1(n6160), .A2(n6159), .A3(n6158), .A4(n6157), .ZN(n8716)
         );
  NAND2_X1 U7665 ( .A1(n8716), .A2(n10078), .ZN(n6162) );
  XNOR2_X1 U7666 ( .A(n6161), .B(n6162), .ZN(n7359) );
  INV_X1 U7667 ( .A(n6161), .ZN(n6164) );
  INV_X1 U7668 ( .A(n6162), .ZN(n6163) );
  NAND2_X1 U7669 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  NAND2_X1 U7670 ( .A1(n6682), .A2(n6547), .ZN(n6169) );
  NAND2_X1 U7671 ( .A1(n6166), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6167) );
  XNOR2_X1 U7672 ( .A(n6167), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8731) );
  AOI22_X1 U7673 ( .A1(n6305), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8731), .B2(
        n6664), .ZN(n6168) );
  XNOR2_X1 U7674 ( .A(n7632), .B(n6428), .ZN(n6179) );
  NAND2_X1 U7675 ( .A1(n6438), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6176) );
  INV_X1 U7676 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7594) );
  OR2_X1 U7677 ( .A1(n6022), .A2(n7594), .ZN(n6175) );
  OR2_X1 U7678 ( .A1(n6170), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7679 ( .A1(n6189), .A2(n6171), .ZN(n7722) );
  OR2_X1 U7680 ( .A1(n4482), .A2(n7722), .ZN(n6174) );
  INV_X1 U7681 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n6172) );
  OR2_X1 U7682 ( .A1(n6361), .A2(n6172), .ZN(n6173) );
  NAND4_X1 U7683 ( .A1(n6176), .A2(n6175), .A3(n6174), .A4(n6173), .ZN(n8715)
         );
  NAND2_X1 U7684 ( .A1(n8715), .A2(n10078), .ZN(n6177) );
  INV_X1 U7685 ( .A(n6177), .ZN(n6178) );
  AND2_X1 U7686 ( .A1(n6179), .A2(n6178), .ZN(n6180) );
  INV_X1 U7687 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6181) );
  AND2_X1 U7688 ( .A1(n6182), .A2(n6181), .ZN(n6183) );
  NAND2_X1 U7689 ( .A1(n6184), .A2(n6183), .ZN(n6199) );
  NAND2_X1 U7690 ( .A1(n6199), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6185) );
  XNOR2_X1 U7691 ( .A(n6185), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7769) );
  AOI22_X1 U7692 ( .A1(n6305), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6664), .B2(
        n7769), .ZN(n6186) );
  NAND2_X1 U7693 ( .A1(n6498), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6194) );
  INV_X1 U7694 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7614) );
  OR2_X1 U7695 ( .A1(n6037), .A2(n7614), .ZN(n6193) );
  INV_X1 U7696 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7598) );
  OR2_X1 U7697 ( .A1(n6022), .A2(n7598), .ZN(n6192) );
  INV_X1 U7698 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7699 ( .A1(n6189), .A2(n6188), .ZN(n6190) );
  NAND2_X1 U7700 ( .A1(n6203), .A2(n6190), .ZN(n7613) );
  OR2_X1 U7701 ( .A1(n4482), .A2(n7613), .ZN(n6191) );
  NAND4_X1 U7702 ( .A1(n6194), .A2(n6193), .A3(n6192), .A4(n6191), .ZN(n8714)
         );
  AND2_X1 U7703 ( .A1(n8714), .A2(n10078), .ZN(n6196) );
  INV_X1 U7704 ( .A(n6195), .ZN(n6198) );
  INV_X1 U7705 ( .A(n6196), .ZN(n6197) );
  NAND2_X1 U7706 ( .A1(n6198), .A2(n6197), .ZN(n7569) );
  NAND2_X1 U7707 ( .A1(n6902), .A2(n6547), .ZN(n6201) );
  NAND2_X1 U7708 ( .A1(n6252), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6216) );
  XNOR2_X1 U7709 ( .A(n6216), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7826) );
  AOI22_X1 U7710 ( .A1(n6305), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6664), .B2(
        n7826), .ZN(n6200) );
  XNOR2_X1 U7711 ( .A(n9057), .B(n6428), .ZN(n6209) );
  NAND2_X1 U7712 ( .A1(n6498), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6208) );
  INV_X1 U7713 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7658) );
  OR2_X1 U7714 ( .A1(n6037), .A2(n7658), .ZN(n6207) );
  INV_X1 U7715 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6202) );
  OR2_X1 U7716 ( .A1(n6022), .A2(n6202), .ZN(n6206) );
  INV_X1 U7717 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7669) );
  NAND2_X1 U7718 ( .A1(n6203), .A2(n7669), .ZN(n6204) );
  NAND2_X1 U7719 ( .A1(n6223), .A2(n6204), .ZN(n7668) );
  OR2_X1 U7720 ( .A1(n4482), .A2(n7668), .ZN(n6205) );
  NAND4_X1 U7721 ( .A1(n6208), .A2(n6207), .A3(n6206), .A4(n6205), .ZN(n8713)
         );
  AND2_X1 U7722 ( .A1(n8713), .A2(n10078), .ZN(n6210) );
  NAND2_X1 U7723 ( .A1(n6209), .A2(n6210), .ZN(n6215) );
  INV_X1 U7724 ( .A(n6209), .ZN(n6212) );
  INV_X1 U7725 ( .A(n6210), .ZN(n6211) );
  NAND2_X1 U7726 ( .A1(n6212), .A2(n6211), .ZN(n6213) );
  NAND2_X1 U7727 ( .A1(n6215), .A2(n6213), .ZN(n7665) );
  INV_X1 U7728 ( .A(n7665), .ZN(n6214) );
  NAND2_X1 U7729 ( .A1(n6945), .A2(n6547), .ZN(n6221) );
  NAND2_X1 U7730 ( .A1(n6216), .A2(n6249), .ZN(n6217) );
  NAND2_X1 U7731 ( .A1(n6217), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U7732 ( .A1(n6218), .A2(n6250), .ZN(n6261) );
  OR2_X1 U7733 ( .A1(n6218), .A2(n6250), .ZN(n6219) );
  AOI22_X1 U7734 ( .A1(n6305), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8006), .B2(
        n6664), .ZN(n6220) );
  XNOR2_X1 U7735 ( .A(n7841), .B(n6448), .ZN(n6231) );
  INV_X1 U7736 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6222) );
  AND2_X1 U7737 ( .A1(n6223), .A2(n6222), .ZN(n6224) );
  NOR2_X1 U7738 ( .A1(n6265), .A2(n6224), .ZN(n7757) );
  INV_X1 U7739 ( .A(n4482), .ZN(n6225) );
  NAND2_X1 U7740 ( .A1(n7757), .A2(n6225), .ZN(n6229) );
  NAND2_X1 U7741 ( .A1(n6062), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6228) );
  NAND2_X1 U7742 ( .A1(n6498), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6227) );
  INV_X1 U7743 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7758) );
  OR2_X1 U7744 ( .A1(n6037), .A2(n7758), .ZN(n6226) );
  NAND4_X1 U7745 ( .A1(n6229), .A2(n6228), .A3(n6227), .A4(n6226), .ZN(n8712)
         );
  NAND2_X1 U7746 ( .A1(n8712), .A2(n10078), .ZN(n6230) );
  XNOR2_X1 U7747 ( .A(n6231), .B(n6230), .ZN(n7836) );
  NAND2_X1 U7748 ( .A1(n6231), .A2(n6230), .ZN(n6232) );
  NAND2_X1 U7749 ( .A1(n7059), .A2(n6547), .ZN(n6236) );
  NAND2_X1 U7750 ( .A1(n6233), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6234) );
  XNOR2_X1 U7751 ( .A(n6234), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8753) );
  AOI22_X1 U7752 ( .A1(n6305), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6664), .B2(
        n8753), .ZN(n6235) );
  XNOR2_X1 U7753 ( .A(n9051), .B(n6428), .ZN(n6243) );
  NAND2_X1 U7754 ( .A1(n6438), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6242) );
  INV_X1 U7755 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8778) );
  OR2_X1 U7756 ( .A1(n6022), .A2(n8778), .ZN(n6241) );
  OAI21_X1 U7757 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(n6237), .A(n6292), .ZN(
        n7985) );
  OR2_X1 U7758 ( .A1(n4482), .A2(n7985), .ZN(n6240) );
  INV_X1 U7759 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n6238) );
  OR2_X1 U7760 ( .A1(n6361), .A2(n6238), .ZN(n6239) );
  NAND4_X1 U7761 ( .A1(n6242), .A2(n6241), .A3(n6240), .A4(n6239), .ZN(n8967)
         );
  AND2_X1 U7762 ( .A1(n8967), .A2(n10078), .ZN(n6244) );
  NAND2_X1 U7763 ( .A1(n6243), .A2(n6244), .ZN(n6286) );
  INV_X1 U7764 ( .A(n6243), .ZN(n6246) );
  INV_X1 U7765 ( .A(n6244), .ZN(n6245) );
  NAND2_X1 U7766 ( .A1(n6246), .A2(n6245), .ZN(n6247) );
  NAND2_X1 U7767 ( .A1(n7005), .A2(n6547), .ZN(n6255) );
  NAND3_X1 U7768 ( .A1(n6250), .A2(n6249), .A3(n6248), .ZN(n6251) );
  OAI21_X1 U7769 ( .B1(n6252), .B2(n6251), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6253) );
  XNOR2_X1 U7770 ( .A(n6253), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8757) );
  AOI22_X1 U7771 ( .A1(n6305), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6664), .B2(
        n8757), .ZN(n6254) );
  XNOR2_X1 U7772 ( .A(n9632), .B(n6448), .ZN(n7981) );
  OR2_X1 U7773 ( .A1(n6267), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6257) );
  NAND2_X1 U7774 ( .A1(n6257), .A2(n6256), .ZN(n7877) );
  AOI22_X1 U7775 ( .A1(n6438), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n6062), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n6260) );
  INV_X1 U7776 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n6258) );
  OR2_X1 U7777 ( .A1(n6361), .A2(n6258), .ZN(n6259) );
  OAI211_X1 U7778 ( .C1(n7877), .C2(n4482), .A(n6260), .B(n6259), .ZN(n8710)
         );
  NAND2_X1 U7779 ( .A1(n8710), .A2(n10078), .ZN(n6278) );
  NAND2_X1 U7780 ( .A1(n7981), .A2(n6278), .ZN(n7983) );
  NAND2_X1 U7781 ( .A1(n7001), .A2(n6547), .ZN(n6264) );
  NAND2_X1 U7782 ( .A1(n6261), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6262) );
  XNOR2_X1 U7783 ( .A(n6262), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8746) );
  AOI22_X1 U7784 ( .A1(n8746), .A2(n6664), .B1(n6305), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6263) );
  XNOR2_X1 U7785 ( .A(n7815), .B(n6448), .ZN(n6276) );
  NOR2_X1 U7786 ( .A1(n6265), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6266) );
  OR2_X1 U7787 ( .A1(n6267), .A2(n6266), .ZN(n7812) );
  INV_X1 U7788 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n6268) );
  OR2_X1 U7789 ( .A1(n6361), .A2(n6268), .ZN(n6270) );
  INV_X1 U7790 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7813) );
  OR2_X1 U7791 ( .A1(n6037), .A2(n7813), .ZN(n6269) );
  AND2_X1 U7792 ( .A1(n6270), .A2(n6269), .ZN(n6273) );
  INV_X1 U7793 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6271) );
  OR2_X1 U7794 ( .A1(n6022), .A2(n6271), .ZN(n6272) );
  OAI211_X1 U7795 ( .C1(n7812), .C2(n4482), .A(n6273), .B(n6272), .ZN(n8711)
         );
  NAND2_X1 U7796 ( .A1(n8711), .A2(n10078), .ZN(n6626) );
  NAND2_X1 U7797 ( .A1(n6276), .A2(n6626), .ZN(n6274) );
  AND2_X1 U7798 ( .A1(n7983), .A2(n6274), .ZN(n6275) );
  INV_X1 U7799 ( .A(n7982), .ZN(n6284) );
  INV_X1 U7800 ( .A(n7981), .ZN(n6282) );
  INV_X1 U7801 ( .A(n6276), .ZN(n7979) );
  INV_X1 U7802 ( .A(n6626), .ZN(n6277) );
  NAND2_X1 U7803 ( .A1(n7979), .A2(n6277), .ZN(n6279) );
  NAND2_X1 U7804 ( .A1(n6279), .A2(n6278), .ZN(n6281) );
  INV_X1 U7805 ( .A(n6278), .ZN(n7980) );
  INV_X1 U7806 ( .A(n6279), .ZN(n6280) );
  AOI22_X1 U7807 ( .A1(n6282), .A2(n6281), .B1(n7980), .B2(n6280), .ZN(n6283)
         );
  AOI21_X1 U7808 ( .B1(n6625), .B2(n6285), .A(n5042), .ZN(n7984) );
  NAND2_X1 U7809 ( .A1(n7262), .A2(n6547), .ZN(n6289) );
  XNOR2_X1 U7810 ( .A(n6287), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8774) );
  AOI22_X1 U7811 ( .A1(n6305), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6664), .B2(
        n8774), .ZN(n6288) );
  XNOR2_X1 U7812 ( .A(n9045), .B(n6428), .ZN(n6299) );
  NAND2_X1 U7813 ( .A1(n6062), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6298) );
  OR2_X1 U7814 ( .A1(n6037), .A2(n8771), .ZN(n6297) );
  INV_X1 U7815 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U7816 ( .A1(n6292), .A2(n6291), .ZN(n6293) );
  NAND2_X1 U7817 ( .A1(n6310), .A2(n6293), .ZN(n7912) );
  OR2_X1 U7818 ( .A1(n4482), .A2(n7912), .ZN(n6296) );
  INV_X1 U7819 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n6294) );
  OR2_X1 U7820 ( .A1(n6361), .A2(n6294), .ZN(n6295) );
  NAND4_X1 U7821 ( .A1(n6298), .A2(n6297), .A3(n6296), .A4(n6295), .ZN(n8709)
         );
  AND2_X1 U7822 ( .A1(n8709), .A2(n10078), .ZN(n6300) );
  NAND2_X1 U7823 ( .A1(n6299), .A2(n6300), .ZN(n7993) );
  INV_X1 U7824 ( .A(n6299), .ZN(n6302) );
  INV_X1 U7825 ( .A(n6300), .ZN(n6301) );
  NAND2_X1 U7826 ( .A1(n6302), .A2(n6301), .ZN(n6303) );
  NAND2_X1 U7827 ( .A1(n7357), .A2(n6547), .ZN(n6307) );
  AOI22_X1 U7828 ( .A1(n6305), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6304), .B2(
        n6664), .ZN(n6306) );
  XNOR2_X1 U7829 ( .A(n9042), .B(n6428), .ZN(n6319) );
  INV_X1 U7830 ( .A(n6319), .ZN(n6316) );
  NAND2_X1 U7831 ( .A1(n6498), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6315) );
  INV_X1 U7832 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6308) );
  OR2_X1 U7833 ( .A1(n6037), .A2(n6308), .ZN(n6314) );
  INV_X1 U7834 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8792) );
  OR2_X1 U7835 ( .A1(n6022), .A2(n8792), .ZN(n6313) );
  INV_X1 U7836 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8001) );
  NAND2_X1 U7837 ( .A1(n6310), .A2(n8001), .ZN(n6311) );
  NAND2_X1 U7838 ( .A1(n6327), .A2(n6311), .ZN(n8000) );
  OR2_X1 U7839 ( .A1(n4482), .A2(n8000), .ZN(n6312) );
  NAND4_X1 U7840 ( .A1(n6315), .A2(n6314), .A3(n6313), .A4(n6312), .ZN(n8969)
         );
  NAND2_X1 U7841 ( .A1(n8969), .A2(n10078), .ZN(n6318) );
  NAND2_X1 U7842 ( .A1(n6316), .A2(n6318), .ZN(n6317) );
  AND2_X1 U7843 ( .A1(n7911), .A2(n6317), .ZN(n6321) );
  INV_X1 U7844 ( .A(n6317), .ZN(n6320) );
  XNOR2_X1 U7845 ( .A(n6319), .B(n6318), .ZN(n7997) );
  AND2_X1 U7846 ( .A1(n7997), .A2(n7993), .ZN(n7994) );
  NAND2_X1 U7847 ( .A1(n7514), .A2(n6547), .ZN(n6323) );
  OR2_X1 U7848 ( .A1(n8436), .A2(n7549), .ZN(n6322) );
  XNOR2_X1 U7849 ( .A(n9035), .B(n6428), .ZN(n6334) );
  NAND2_X1 U7850 ( .A1(n6438), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6333) );
  INV_X1 U7851 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n6324) );
  OR2_X1 U7852 ( .A1(n6022), .A2(n6324), .ZN(n6332) );
  INV_X1 U7853 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U7854 ( .A1(n6327), .A2(n6326), .ZN(n6328) );
  NAND2_X1 U7855 ( .A1(n6343), .A2(n6328), .ZN(n8046) );
  OR2_X1 U7856 ( .A1(n4482), .A2(n8046), .ZN(n6331) );
  INV_X1 U7857 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n6329) );
  OR2_X1 U7858 ( .A1(n6361), .A2(n6329), .ZN(n6330) );
  NAND4_X1 U7859 ( .A1(n6333), .A2(n6332), .A3(n6331), .A4(n6330), .ZN(n8939)
         );
  AND2_X1 U7860 ( .A1(n8939), .A2(n10078), .ZN(n6335) );
  NAND2_X1 U7861 ( .A1(n6334), .A2(n6335), .ZN(n6339) );
  INV_X1 U7862 ( .A(n6334), .ZN(n6337) );
  INV_X1 U7863 ( .A(n6335), .ZN(n6336) );
  NAND2_X1 U7864 ( .A1(n6337), .A2(n6336), .ZN(n6338) );
  NAND2_X1 U7865 ( .A1(n6339), .A2(n6338), .ZN(n8045) );
  NAND2_X1 U7866 ( .A1(n7586), .A2(n6547), .ZN(n6341) );
  OR2_X1 U7867 ( .A1(n8436), .A2(n7587), .ZN(n6340) );
  XNOR2_X1 U7868 ( .A(n9030), .B(n6428), .ZN(n6351) );
  NAND2_X1 U7869 ( .A1(n6438), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6348) );
  INV_X1 U7870 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n10271) );
  OR2_X1 U7871 ( .A1(n6022), .A2(n10271), .ZN(n6347) );
  INV_X1 U7872 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10390) );
  NAND2_X1 U7873 ( .A1(n6343), .A2(n10390), .ZN(n6344) );
  NAND2_X1 U7874 ( .A1(n6358), .A2(n6344), .ZN(n8932) );
  OR2_X1 U7875 ( .A1(n4482), .A2(n8932), .ZN(n6346) );
  INV_X1 U7876 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n10222) );
  OR2_X1 U7877 ( .A1(n6361), .A2(n10222), .ZN(n6345) );
  NAND4_X1 U7878 ( .A1(n6348), .A2(n6347), .A3(n6346), .A4(n6345), .ZN(n8708)
         );
  NAND2_X1 U7879 ( .A1(n8708), .A2(n10078), .ZN(n6349) );
  XNOR2_X1 U7880 ( .A(n6351), .B(n6349), .ZN(n8657) );
  NAND2_X1 U7881 ( .A1(n8658), .A2(n8657), .ZN(n8656) );
  INV_X1 U7882 ( .A(n6349), .ZN(n6350) );
  NAND2_X1 U7883 ( .A1(n6351), .A2(n6350), .ZN(n6352) );
  NAND2_X1 U7884 ( .A1(n7621), .A2(n6547), .ZN(n6354) );
  OR2_X1 U7885 ( .A1(n8436), .A2(n10341), .ZN(n6353) );
  XNOR2_X1 U7886 ( .A(n9025), .B(n6448), .ZN(n6367) );
  NAND2_X1 U7887 ( .A1(n6438), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6365) );
  INV_X1 U7888 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6355) );
  OR2_X1 U7889 ( .A1(n6022), .A2(n6355), .ZN(n6364) );
  INV_X1 U7890 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U7891 ( .A1(n6358), .A2(n6357), .ZN(n6359) );
  NAND2_X1 U7892 ( .A1(n6372), .A2(n6359), .ZN(n8918) );
  OR2_X1 U7893 ( .A1(n4482), .A2(n8918), .ZN(n6363) );
  INV_X1 U7894 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n6360) );
  OR2_X1 U7895 ( .A1(n6361), .A2(n6360), .ZN(n6362) );
  NAND4_X1 U7896 ( .A1(n6365), .A2(n6364), .A3(n6363), .A4(n6362), .ZN(n8938)
         );
  NAND2_X1 U7897 ( .A1(n8938), .A2(n10078), .ZN(n8683) );
  INV_X1 U7898 ( .A(n6366), .ZN(n6368) );
  NAND2_X1 U7899 ( .A1(n6368), .A2(n6367), .ZN(n6369) );
  NAND2_X1 U7900 ( .A1(n7782), .A2(n6547), .ZN(n6371) );
  OR2_X1 U7901 ( .A1(n8436), .A2(n10218), .ZN(n6370) );
  XNOR2_X1 U7902 ( .A(n9020), .B(n6428), .ZN(n6378) );
  XNOR2_X1 U7903 ( .A(n6380), .B(n6378), .ZN(n8648) );
  NAND2_X1 U7904 ( .A1(n6062), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6377) );
  INV_X1 U7905 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8909) );
  OR2_X1 U7906 ( .A1(n6037), .A2(n8909), .ZN(n6376) );
  INV_X1 U7907 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U7908 ( .A1(n6372), .A2(n8651), .ZN(n6373) );
  NAND2_X1 U7909 ( .A1(n6398), .A2(n6373), .ZN(n8908) );
  OR2_X1 U7910 ( .A1(n4482), .A2(n8908), .ZN(n6375) );
  INV_X1 U7911 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n10348) );
  OR2_X1 U7912 ( .A1(n6361), .A2(n10348), .ZN(n6374) );
  NAND4_X1 U7913 ( .A1(n6377), .A2(n6376), .A3(n6375), .A4(n6374), .ZN(n8883)
         );
  AND2_X1 U7914 ( .A1(n8883), .A2(n10078), .ZN(n8650) );
  NAND2_X1 U7915 ( .A1(n8648), .A2(n8650), .ZN(n8649) );
  INV_X1 U7916 ( .A(n6378), .ZN(n6379) );
  OR2_X1 U7917 ( .A1(n6380), .A2(n6379), .ZN(n6381) );
  NAND2_X1 U7918 ( .A1(n7845), .A2(n6547), .ZN(n6383) );
  OR2_X1 U7919 ( .A1(n8436), .A2(n7846), .ZN(n6382) );
  NAND2_X2 U7920 ( .A1(n6383), .A2(n6382), .ZN(n9014) );
  XNOR2_X1 U7921 ( .A(n9014), .B(n6448), .ZN(n6389) );
  XNOR2_X1 U7922 ( .A(n6391), .B(n6389), .ZN(n8676) );
  NAND2_X1 U7923 ( .A1(n6438), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6388) );
  INV_X1 U7924 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n10206) );
  OR2_X1 U7925 ( .A1(n6022), .A2(n10206), .ZN(n6387) );
  INV_X1 U7926 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8677) );
  XNOR2_X1 U7927 ( .A(n6398), .B(n8677), .ZN(n8886) );
  OR2_X1 U7928 ( .A1(n4482), .A2(n8886), .ZN(n6386) );
  INV_X1 U7929 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n6384) );
  OR2_X1 U7930 ( .A1(n6361), .A2(n6384), .ZN(n6385) );
  NAND4_X1 U7931 ( .A1(n6388), .A2(n6387), .A3(n6386), .A4(n6385), .ZN(n8900)
         );
  AND2_X1 U7932 ( .A1(n8900), .A2(n10078), .ZN(n8675) );
  NAND2_X1 U7933 ( .A1(n8676), .A2(n8675), .ZN(n8674) );
  INV_X1 U7934 ( .A(n6389), .ZN(n6390) );
  NAND2_X1 U7935 ( .A1(n6391), .A2(n6390), .ZN(n6392) );
  NAND2_X1 U7936 ( .A1(n8674), .A2(n6392), .ZN(n8668) );
  NAND2_X1 U7937 ( .A1(n6393), .A2(n6547), .ZN(n6395) );
  OR2_X1 U7938 ( .A1(n8436), .A2(n7895), .ZN(n6394) );
  XNOR2_X1 U7939 ( .A(n9011), .B(n6428), .ZN(n6405) );
  NAND2_X1 U7940 ( .A1(n6062), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6404) );
  INV_X1 U7941 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n10243) );
  OR2_X1 U7942 ( .A1(n6037), .A2(n10243), .ZN(n6403) );
  INV_X1 U7943 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6396) );
  OAI21_X1 U7944 ( .B1(n6398), .B2(n8677), .A(n6396), .ZN(n6399) );
  NAND2_X1 U7945 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_24__SCAN_IN), 
        .ZN(n6397) );
  NAND2_X1 U7946 ( .A1(n6399), .A2(n6414), .ZN(n8868) );
  OR2_X1 U7947 ( .A1(n4482), .A2(n8868), .ZN(n6402) );
  INV_X1 U7948 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n6400) );
  OR2_X1 U7949 ( .A1(n6361), .A2(n6400), .ZN(n6401) );
  NAND4_X1 U7950 ( .A1(n6404), .A2(n6403), .A3(n6402), .A4(n6401), .ZN(n8882)
         );
  AND2_X1 U7951 ( .A1(n8882), .A2(n10078), .ZN(n6406) );
  INV_X1 U7952 ( .A(n6405), .ZN(n6408) );
  INV_X1 U7953 ( .A(n6406), .ZN(n6407) );
  NAND2_X1 U7954 ( .A1(n6408), .A2(n6407), .ZN(n8665) );
  NAND2_X1 U7955 ( .A1(n7896), .A2(n6547), .ZN(n6410) );
  OR2_X1 U7956 ( .A1(n8436), .A2(n10335), .ZN(n6409) );
  XNOR2_X1 U7957 ( .A(n9005), .B(n6448), .ZN(n6421) );
  NAND2_X1 U7958 ( .A1(n6062), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6420) );
  INV_X1 U7959 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n6411) );
  OR2_X1 U7960 ( .A1(n6037), .A2(n6411), .ZN(n6419) );
  INV_X1 U7961 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U7962 ( .A1(n6414), .A2(n6413), .ZN(n6415) );
  NAND2_X1 U7963 ( .A1(n6441), .A2(n6415), .ZN(n8849) );
  INV_X1 U7964 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n6416) );
  OR2_X1 U7965 ( .A1(n6361), .A2(n6416), .ZN(n6417) );
  NAND4_X1 U7966 ( .A1(n6420), .A2(n6419), .A3(n6418), .A4(n6417), .ZN(n8707)
         );
  NAND2_X1 U7967 ( .A1(n8707), .A2(n10078), .ZN(n6422) );
  XNOR2_X1 U7968 ( .A(n6421), .B(n6422), .ZN(n8694) );
  INV_X1 U7969 ( .A(n6421), .ZN(n6424) );
  INV_X1 U7970 ( .A(n6422), .ZN(n6423) );
  NAND2_X1 U7971 ( .A1(n6424), .A2(n6423), .ZN(n6425) );
  NAND2_X1 U7972 ( .A1(n7945), .A2(n6547), .ZN(n6427) );
  OR2_X1 U7973 ( .A1(n8436), .A2(n7949), .ZN(n6426) );
  XNOR2_X1 U7974 ( .A(n8999), .B(n6428), .ZN(n6437) );
  NAND2_X1 U7975 ( .A1(n6438), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6434) );
  INV_X1 U7976 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10381) );
  OR2_X1 U7977 ( .A1(n6022), .A2(n10381), .ZN(n6433) );
  INV_X1 U7978 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10322) );
  XNOR2_X1 U7979 ( .A(n6441), .B(n10322), .ZN(n8830) );
  OR2_X1 U7980 ( .A1(n4482), .A2(n8830), .ZN(n6432) );
  INV_X1 U7981 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6430) );
  OR2_X1 U7982 ( .A1(n6361), .A2(n6430), .ZN(n6431) );
  NAND4_X1 U7983 ( .A1(n6434), .A2(n6433), .A3(n6432), .A4(n6431), .ZN(n8706)
         );
  NAND2_X1 U7984 ( .A1(n8706), .A2(n10078), .ZN(n6435) );
  XNOR2_X1 U7985 ( .A(n6437), .B(n6435), .ZN(n8642) );
  INV_X1 U7986 ( .A(n6435), .ZN(n6436) );
  NAND2_X1 U7987 ( .A1(n6438), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6447) );
  INV_X1 U7988 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6439) );
  OR2_X1 U7989 ( .A1(n6022), .A2(n6439), .ZN(n6446) );
  INV_X1 U7990 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6440) );
  OAI21_X1 U7991 ( .B1(n6441), .B2(n10322), .A(n6440), .ZN(n6442) );
  NAND2_X1 U7992 ( .A1(n6442), .A2(n6609), .ZN(n6507) );
  OR2_X1 U7993 ( .A1(n4482), .A2(n6507), .ZN(n6445) );
  INV_X1 U7994 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6443) );
  OR2_X1 U7995 ( .A1(n6361), .A2(n6443), .ZN(n6444) );
  NAND4_X1 U7996 ( .A1(n6447), .A2(n6446), .A3(n6445), .A4(n6444), .ZN(n8705)
         );
  NAND2_X1 U7997 ( .A1(n8705), .A2(n10078), .ZN(n6449) );
  XNOR2_X1 U7998 ( .A(n6449), .B(n6448), .ZN(n6450) );
  XNOR2_X1 U7999 ( .A(n6451), .B(n6450), .ZN(n6490) );
  INV_X1 U8000 ( .A(n6490), .ZN(n6489) );
  NAND2_X1 U8001 ( .A1(n6452), .A2(n6457), .ZN(n6453) );
  NAND2_X1 U8002 ( .A1(n6453), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6484) );
  INV_X1 U8003 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U8004 ( .A1(n6484), .A2(n6483), .ZN(n6486) );
  NAND2_X1 U8005 ( .A1(n6486), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6454) );
  INV_X1 U8006 ( .A(P2_B_REG_SCAN_IN), .ZN(n6455) );
  XNOR2_X1 U8007 ( .A(n7844), .B(n6455), .ZN(n6461) );
  INV_X1 U8008 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6456) );
  NAND2_X1 U8009 ( .A1(n6457), .A2(n6456), .ZN(n6458) );
  NAND2_X1 U8010 ( .A1(n6462), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6460) );
  INV_X1 U8011 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n10257) );
  XNOR2_X1 U8012 ( .A(n6460), .B(n10257), .ZN(n7894) );
  NAND2_X1 U8013 ( .A1(n6461), .A2(n7894), .ZN(n6466) );
  OAI21_X1 U8014 ( .B1(n6462), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6463) );
  MUX2_X1 U8015 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6463), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6465) );
  NAND2_X1 U8016 ( .A1(n6465), .A2(n6464), .ZN(n7899) );
  INV_X1 U8017 ( .A(n7899), .ZN(n6478) );
  NOR2_X1 U8018 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .ZN(
        n6470) );
  NOR4_X1 U8019 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6469) );
  NOR4_X1 U8020 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6468) );
  NOR4_X1 U8021 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n6467) );
  AND4_X1 U8022 ( .A1(n6470), .A2(n6469), .A3(n6468), .A4(n6467), .ZN(n6476)
         );
  NOR4_X1 U8023 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6474) );
  NOR4_X1 U8024 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6473) );
  NOR4_X1 U8025 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6472) );
  NOR4_X1 U8026 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6471) );
  AND4_X1 U8027 ( .A1(n6474), .A2(n6473), .A3(n6472), .A4(n6471), .ZN(n6475)
         );
  NAND2_X1 U8028 ( .A1(n6476), .A2(n6475), .ZN(n6477) );
  AND2_X1 U8029 ( .A1(n10018), .A2(n6477), .ZN(n6586) );
  INV_X1 U8030 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10336) );
  NAND2_X1 U8031 ( .A1(n10018), .A2(n10336), .ZN(n6480) );
  NOR2_X1 U8032 ( .A1(n7844), .A2(n6478), .ZN(n10021) );
  INV_X1 U8033 ( .A(n10021), .ZN(n6479) );
  NAND2_X1 U8034 ( .A1(n6480), .A2(n6479), .ZN(n6599) );
  INV_X1 U8035 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10023) );
  NAND2_X1 U8036 ( .A1(n10018), .A2(n10023), .ZN(n6481) );
  NAND2_X1 U8037 ( .A1(n7899), .A2(n7894), .ZN(n10022) );
  NAND2_X1 U8038 ( .A1(n6481), .A2(n10022), .ZN(n6598) );
  NOR2_X1 U8039 ( .A1(n7899), .A2(n7894), .ZN(n6482) );
  NAND2_X1 U8040 ( .A1(n7844), .A2(n6482), .ZN(n6689) );
  OR2_X1 U8041 ( .A1(n6484), .A2(n6483), .ZN(n6485) );
  NAND2_X1 U8042 ( .A1(n6486), .A2(n6485), .ZN(n6663) );
  NOR2_X1 U8043 ( .A1(n6504), .A2(n10019), .ZN(n6496) );
  AND2_X1 U8044 ( .A1(n8587), .A2(n8618), .ZN(n6495) );
  NAND2_X1 U8045 ( .A1(n8626), .A2(n10027), .ZN(n10076) );
  NAND2_X1 U8046 ( .A1(n8628), .A2(n8622), .ZN(n6666) );
  AND2_X1 U8047 ( .A1(n10076), .A2(n6666), .ZN(n6488) );
  NAND2_X1 U8048 ( .A1(n6489), .A2(n9628), .ZN(n6511) );
  INV_X1 U8049 ( .A(n6496), .ZN(n6493) );
  OR2_X1 U8050 ( .A1(n6491), .A2(n8587), .ZN(n6607) );
  AND2_X1 U8051 ( .A1(n7622), .A2(n6304), .ZN(n6492) );
  NAND2_X1 U8052 ( .A1(n10070), .A2(n8443), .ZN(n6587) );
  NAND2_X1 U8053 ( .A1(n6496), .A2(n6495), .ZN(n9635) );
  INV_X1 U8054 ( .A(n4474), .ZN(n6694) );
  INV_X1 U8055 ( .A(n8687), .ZN(n8048) );
  NAND2_X1 U8056 ( .A1(n6062), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U8057 ( .A1(n6498), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6502) );
  OR2_X1 U8058 ( .A1(n4482), .A2(n6609), .ZN(n6501) );
  INV_X1 U8059 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6499) );
  OR2_X1 U8060 ( .A1(n6037), .A2(n6499), .ZN(n6500) );
  NAND4_X1 U8061 ( .A1(n6503), .A2(n6502), .A3(n6501), .A4(n6500), .ZN(n8704)
         );
  NAND2_X1 U8062 ( .A1(n8048), .A2(n8704), .ZN(n6510) );
  INV_X1 U8063 ( .A(n8686), .ZN(n8047) );
  NAND2_X1 U8064 ( .A1(n8047), .A2(n8706), .ZN(n6509) );
  NAND2_X1 U8065 ( .A1(n6504), .A2(n6587), .ZN(n6910) );
  INV_X1 U8066 ( .A(n6666), .ZN(n6691) );
  NAND2_X1 U8067 ( .A1(n8626), .A2(n6691), .ZN(n6584) );
  AND3_X1 U8068 ( .A1(n6689), .A2(n6663), .A3(n6584), .ZN(n6505) );
  NAND2_X1 U8069 ( .A1(n6910), .A2(n6505), .ZN(n6506) );
  INV_X1 U8070 ( .A(n6507), .ZN(n8815) );
  INV_X2 U8071 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  AOI22_X1 U8072 ( .A1(n9631), .A2(n8815), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6508) );
  INV_X1 U8073 ( .A(n8967), .ZN(n8448) );
  NAND2_X1 U8074 ( .A1(n6514), .A2(n6581), .ZN(n6554) );
  NAND2_X1 U8075 ( .A1(n6554), .A2(n8471), .ZN(n7086) );
  NAND2_X1 U8076 ( .A1(n7086), .A2(n7087), .ZN(n6516) );
  INV_X1 U8077 ( .A(n4480), .ZN(n6514) );
  NAND2_X1 U8078 ( .A1(n6514), .A2(n6513), .ZN(n6515) );
  NAND2_X1 U8079 ( .A1(n6516), .A2(n6515), .ZN(n7141) );
  NAND2_X1 U8080 ( .A1(n7273), .A2(n10037), .ZN(n6518) );
  NAND2_X1 U8081 ( .A1(n8723), .A2(n6519), .ZN(n8477) );
  NAND2_X1 U8082 ( .A1(n8458), .A2(n8477), .ZN(n8590) );
  NAND2_X1 U8083 ( .A1(n6991), .A2(n6519), .ZN(n6520) );
  NOR2_X1 U8084 ( .A1(n8722), .A2(n10052), .ZN(n7063) );
  INV_X1 U8085 ( .A(n7063), .ZN(n8459) );
  NAND2_X1 U8086 ( .A1(n7137), .A2(n8591), .ZN(n6522) );
  NAND2_X1 U8087 ( .A1(n4670), .A2(n10052), .ZN(n6521) );
  NOR2_X1 U8088 ( .A1(n8721), .A2(n7069), .ZN(n6524) );
  NAND2_X1 U8089 ( .A1(n7229), .A2(n7069), .ZN(n8460) );
  NAND2_X1 U8090 ( .A1(n8460), .A2(n8479), .ZN(n8592) );
  OR2_X1 U8091 ( .A1(n8592), .A2(n7163), .ZN(n6523) );
  INV_X1 U8092 ( .A(n8720), .ZN(n6525) );
  OR2_X1 U8093 ( .A1(n6525), .A2(n7236), .ZN(n8481) );
  NAND2_X1 U8094 ( .A1(n7236), .A2(n6525), .ZN(n8485) );
  INV_X1 U8095 ( .A(n8594), .ZN(n7226) );
  OR2_X1 U8096 ( .A1(n7420), .A2(n7407), .ZN(n8487) );
  NAND2_X1 U8097 ( .A1(n7420), .A2(n7407), .ZN(n8486) );
  INV_X1 U8098 ( .A(n8595), .ZN(n6526) );
  OR2_X1 U8099 ( .A1(n7420), .A2(n8719), .ZN(n6527) );
  INV_X1 U8100 ( .A(n8718), .ZN(n7326) );
  OR2_X1 U8101 ( .A1(n10064), .A2(n7326), .ZN(n8491) );
  NAND2_X1 U8102 ( .A1(n10064), .A2(n7326), .ZN(n8490) );
  NAND2_X1 U8103 ( .A1(n8491), .A2(n8490), .ZN(n7403) );
  INV_X1 U8104 ( .A(n7403), .ZN(n8596) );
  INV_X1 U8105 ( .A(n6528), .ZN(n6529) );
  INV_X1 U8106 ( .A(n8717), .ZN(n7406) );
  NAND2_X1 U8107 ( .A1(n8497), .A2(n8500), .ZN(n8598) );
  NAND2_X1 U8108 ( .A1(n10064), .A2(n8718), .ZN(n7467) );
  NAND2_X1 U8109 ( .A1(n7462), .A2(n8716), .ZN(n6530) );
  INV_X1 U8110 ( .A(n8716), .ZN(n7517) );
  OR2_X1 U8111 ( .A1(n7462), .A2(n7517), .ZN(n8503) );
  NAND2_X1 U8112 ( .A1(n7462), .A2(n7517), .ZN(n8501) );
  NAND2_X1 U8113 ( .A1(n8503), .A2(n8501), .ZN(n8600) );
  INV_X1 U8114 ( .A(n8715), .ZN(n7611) );
  OR2_X1 U8115 ( .A1(n7632), .A2(n7611), .ZN(n8505) );
  NAND2_X1 U8116 ( .A1(n7632), .A2(n7611), .ZN(n8498) );
  NAND2_X1 U8117 ( .A1(n7632), .A2(n8715), .ZN(n6531) );
  INV_X1 U8118 ( .A(n8714), .ZN(n7670) );
  OR2_X1 U8119 ( .A1(n7616), .A2(n7670), .ZN(n8511) );
  NAND2_X1 U8120 ( .A1(n7616), .A2(n7670), .ZN(n8510) );
  INV_X1 U8121 ( .A(n8713), .ZN(n7753) );
  OR2_X1 U8122 ( .A1(n9057), .A2(n7753), .ZN(n8455) );
  NAND2_X1 U8123 ( .A1(n9057), .A2(n7753), .ZN(n8454) );
  NAND2_X1 U8124 ( .A1(n8455), .A2(n8454), .ZN(n7650) );
  NAND2_X1 U8125 ( .A1(n9057), .A2(n8713), .ZN(n6533) );
  NAND2_X1 U8126 ( .A1(n7841), .A2(n7807), .ZN(n8516) );
  NAND2_X1 U8127 ( .A1(n8515), .A2(n8516), .ZN(n8605) );
  OR2_X1 U8128 ( .A1(n7841), .A2(n8712), .ZN(n6534) );
  INV_X1 U8129 ( .A(n8711), .ZN(n7754) );
  NOR2_X1 U8130 ( .A1(n7815), .A2(n7754), .ZN(n8521) );
  INV_X1 U8131 ( .A(n8521), .ZN(n6535) );
  NAND2_X1 U8132 ( .A1(n7815), .A2(n7754), .ZN(n8520) );
  OR2_X1 U8133 ( .A1(n7815), .A2(n8711), .ZN(n6536) );
  INV_X1 U8134 ( .A(n8710), .ZN(n7987) );
  OR2_X1 U8135 ( .A1(n9632), .A2(n7987), .ZN(n8453) );
  AND2_X1 U8136 ( .A1(n9632), .A2(n7987), .ZN(n6566) );
  INV_X1 U8137 ( .A(n6566), .ZN(n8452) );
  NAND2_X1 U8138 ( .A1(n9632), .A2(n8710), .ZN(n6539) );
  XNOR2_X1 U8139 ( .A(n9051), .B(n8967), .ZN(n8607) );
  INV_X1 U8140 ( .A(n9045), .ZN(n8978) );
  INV_X1 U8141 ( .A(n8709), .ZN(n7986) );
  INV_X1 U8142 ( .A(n8969), .ZN(n8957) );
  INV_X1 U8143 ( .A(n8939), .ZN(n8659) );
  NAND2_X1 U8144 ( .A1(n9035), .A2(n8659), .ZN(n8539) );
  NAND2_X1 U8145 ( .A1(n8537), .A2(n8539), .ZN(n8955) );
  INV_X1 U8146 ( .A(n9030), .ZN(n8935) );
  NAND2_X1 U8147 ( .A1(n9025), .A2(n8660), .ZN(n8541) );
  NAND2_X1 U8148 ( .A1(n8546), .A2(n8541), .ZN(n8922) );
  INV_X1 U8149 ( .A(n9025), .ZN(n8921) );
  OR2_X1 U8150 ( .A1(n9020), .A2(n8924), .ZN(n8445) );
  NAND2_X1 U8151 ( .A1(n9020), .A2(n8924), .ZN(n8549) );
  NAND2_X1 U8152 ( .A1(n8904), .A2(n8903), .ZN(n8905) );
  OAI21_X1 U8153 ( .B1(n4655), .B2(n8924), .A(n8905), .ZN(n8891) );
  NAND2_X1 U8154 ( .A1(n9014), .A2(n8669), .ZN(n8551) );
  NAND2_X1 U8155 ( .A1(n9005), .A2(n8837), .ZN(n8561) );
  INV_X1 U8156 ( .A(n9005), .ZN(n8852) );
  INV_X1 U8157 ( .A(n8836), .ZN(n8563) );
  INV_X1 U8158 ( .A(SI_28_), .ZN(n6543) );
  NAND2_X1 U8159 ( .A1(n6544), .A2(n6543), .ZN(n6545) );
  INV_X1 U8160 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9596) );
  INV_X1 U8161 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9088) );
  MUX2_X1 U8162 ( .A(n9596), .B(n9088), .S(n4481), .Z(n8053) );
  XNOR2_X1 U8163 ( .A(n8053), .B(SI_29_), .ZN(n6546) );
  NAND2_X1 U8164 ( .A1(n9086), .A2(n6547), .ZN(n6549) );
  OR2_X1 U8165 ( .A1(n8436), .A2(n9088), .ZN(n6548) );
  INV_X1 U8166 ( .A(n8704), .ZN(n8822) );
  XNOR2_X1 U8167 ( .A(n6550), .B(n8614), .ZN(n6619) );
  INV_X1 U8168 ( .A(n10070), .ZN(n9063) );
  NAND2_X1 U8169 ( .A1(n6617), .A2(n7622), .ZN(n6552) );
  AND2_X1 U8170 ( .A1(n6666), .A2(n8618), .ZN(n6551) );
  NAND2_X1 U8171 ( .A1(n6552), .A2(n6551), .ZN(n7961) );
  INV_X1 U8172 ( .A(n7157), .ZN(n6553) );
  NAND2_X1 U8173 ( .A1(n6553), .A2(n10026), .ZN(n8635) );
  NAND2_X1 U8174 ( .A1(n7272), .A2(n8467), .ZN(n6556) );
  NAND2_X1 U8175 ( .A1(n8460), .A2(n8459), .ZN(n8456) );
  INV_X1 U8176 ( .A(n8485), .ZN(n6558) );
  INV_X1 U8177 ( .A(n8497), .ZN(n6560) );
  AND2_X1 U8178 ( .A1(n8490), .A2(n8500), .ZN(n6559) );
  OR2_X1 U8179 ( .A1(n6560), .A2(n6559), .ZN(n6561) );
  NAND2_X1 U8180 ( .A1(n6562), .A2(n6561), .ZN(n7449) );
  NAND2_X1 U8181 ( .A1(n7449), .A2(n8503), .ZN(n6563) );
  NAND2_X1 U8182 ( .A1(n6563), .A2(n8501), .ZN(n7627) );
  AND2_X1 U8183 ( .A1(n8510), .A2(n8498), .ZN(n8506) );
  OR2_X1 U8184 ( .A1(n9051), .A2(n8448), .ZN(n8451) );
  NAND2_X1 U8185 ( .A1(n9045), .A2(n7986), .ZN(n8584) );
  NAND2_X1 U8186 ( .A1(n8965), .A2(n8584), .ZN(n8029) );
  OR2_X1 U8187 ( .A1(n9042), .A2(n8957), .ZN(n8536) );
  NAND2_X1 U8188 ( .A1(n9042), .A2(n8957), .ZN(n8950) );
  NAND2_X1 U8189 ( .A1(n8536), .A2(n8950), .ZN(n8028) );
  NOR2_X1 U8190 ( .A1(n9045), .A2(n7986), .ZN(n8586) );
  NOR2_X1 U8191 ( .A1(n8028), .A2(n8586), .ZN(n6567) );
  NAND2_X1 U8192 ( .A1(n8029), .A2(n6567), .ZN(n8951) );
  INV_X1 U8193 ( .A(n8950), .ZN(n6568) );
  NOR2_X1 U8194 ( .A1(n8955), .A2(n6568), .ZN(n6569) );
  XNOR2_X1 U8195 ( .A(n9030), .B(n8959), .ZN(n8611) );
  NAND2_X1 U8196 ( .A1(n9030), .A2(n8959), .ZN(n8538) );
  INV_X1 U8197 ( .A(n8897), .ZN(n6572) );
  INV_X1 U8198 ( .A(n8882), .ZN(n8695) );
  OR2_X1 U8199 ( .A1(n9011), .A2(n8695), .ZN(n8556) );
  NOR2_X1 U8200 ( .A1(n8999), .A2(n8821), .ZN(n8564) );
  XNOR2_X1 U8201 ( .A(n8430), .B(n8571), .ZN(n6574) );
  OR2_X1 U8202 ( .A1(n8587), .A2(n8443), .ZN(n8442) );
  NAND2_X1 U8203 ( .A1(n8442), .A2(n8620), .ZN(n8971) );
  INV_X1 U8204 ( .A(n8627), .ZN(n6575) );
  AOI21_X1 U8205 ( .B1(n6575), .B2(P2_B_REG_SCAN_IN), .A(n8958), .ZN(n8800) );
  INV_X1 U8206 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6578) );
  NAND2_X1 U8207 ( .A1(n6062), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6577) );
  INV_X1 U8208 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n10269) );
  OR2_X1 U8209 ( .A1(n6361), .A2(n10269), .ZN(n6576) );
  OAI211_X1 U8210 ( .C1(n6037), .C2(n6578), .A(n6577), .B(n6576), .ZN(n8703)
         );
  INV_X1 U8211 ( .A(n9632), .ZN(n9637) );
  INV_X1 U8212 ( .A(n7815), .ZN(n7884) );
  OR2_X1 U8213 ( .A1(n6581), .A2(n10026), .ZN(n7153) );
  NAND2_X1 U8214 ( .A1(n10039), .A2(n6519), .ZN(n7269) );
  OR2_X1 U8215 ( .A1(n7269), .A2(n7136), .ZN(n7133) );
  INV_X1 U8216 ( .A(n7236), .ZN(n10057) );
  INV_X1 U8217 ( .A(n7420), .ZN(n7107) );
  NAND2_X1 U8218 ( .A1(n7232), .A2(n7107), .ZN(n7412) );
  INV_X1 U8219 ( .A(n7462), .ZN(n10071) );
  INV_X1 U8220 ( .A(n7632), .ZN(n7725) );
  NAND2_X1 U8221 ( .A1(n8039), .A2(n8973), .ZN(n8946) );
  NOR2_X2 U8222 ( .A1(n8946), .A2(n9035), .ZN(n8945) );
  NAND2_X1 U8223 ( .A1(n8852), .A2(n8866), .ZN(n8846) );
  NAND2_X1 U8224 ( .A1(n8817), .A2(n8829), .ZN(n8812) );
  AOI21_X1 U8225 ( .B1(n6606), .B2(n8812), .A(n8804), .ZN(n6614) );
  AOI22_X1 U8226 ( .A1(n6614), .A2(n10035), .B1(n9058), .B2(n6606), .ZN(n6582)
         );
  INV_X1 U8227 ( .A(n6584), .ZN(n6585) );
  OR2_X1 U8228 ( .A1(n10019), .A2(n6585), .ZN(n6908) );
  NAND2_X1 U8229 ( .A1(n6598), .A2(n6587), .ZN(n6588) );
  INV_X1 U8230 ( .A(n6599), .ZN(n6589) );
  INV_X1 U8231 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6590) );
  NAND2_X1 U8232 ( .A1(n6592), .A2(n6591), .ZN(P2_U3549) );
  NAND2_X1 U8233 ( .A1(n6594), .A2(n10086), .ZN(n6597) );
  OR2_X1 U8234 ( .A1(n10086), .A2(n6595), .ZN(n6596) );
  NAND2_X1 U8235 ( .A1(n6597), .A2(n6596), .ZN(P2_U3517) );
  INV_X1 U8236 ( .A(n6598), .ZN(n6600) );
  AND2_X1 U8237 ( .A1(n6600), .A2(n6599), .ZN(n6603) );
  INV_X1 U8238 ( .A(n6601), .ZN(n6602) );
  NAND2_X1 U8239 ( .A1(n6603), .A2(n6602), .ZN(n6605) );
  OR2_X1 U8240 ( .A1(n6605), .A2(n6304), .ZN(n7106) );
  NOR2_X2 U8241 ( .A1(n7106), .A2(n10078), .ZN(n8984) );
  INV_X1 U8242 ( .A(n6606), .ZN(n6612) );
  INV_X1 U8243 ( .A(n6607), .ZN(n6608) );
  INV_X1 U8244 ( .A(n6609), .ZN(n6610) );
  INV_X1 U8245 ( .A(n8907), .ZN(n8974) );
  AOI22_X1 U8246 ( .A1(n4476), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n6610), .B2(
        n8974), .ZN(n6611) );
  OAI21_X1 U8247 ( .B1(n6612), .B2(n8977), .A(n6611), .ZN(n6613) );
  AOI21_X1 U8248 ( .B1(n6614), .B2(n8984), .A(n6613), .ZN(n6615) );
  OR2_X1 U8249 ( .A1(n6617), .A2(n8618), .ZN(n7267) );
  NAND2_X1 U8250 ( .A1(n7961), .A2(n7267), .ZN(n6618) );
  INV_X1 U8251 ( .A(n7778), .ZN(n6620) );
  NOR2_X1 U8252 ( .A1(n6621), .A2(n6620), .ZN(n6792) );
  AND2_X2 U8253 ( .A1(n6792), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  NAND2_X1 U8254 ( .A1(n8262), .A2(n6621), .ZN(n6622) );
  NAND2_X1 U8255 ( .A1(n6622), .A2(n7778), .ZN(n9751) );
  NAND2_X1 U8256 ( .A1(n9751), .A2(n9755), .ZN(n6623) );
  NAND2_X1 U8257 ( .A1(n6623), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8258 ( .A(n10025), .ZN(n6624) );
  OR2_X2 U8259 ( .A1(n6689), .A2(n6624), .ZN(n8724) );
  INV_X1 U8260 ( .A(n8724), .ZN(P2_U3966) );
  XNOR2_X1 U8261 ( .A(n6625), .B(n7979), .ZN(n6627) );
  NOR2_X1 U8262 ( .A1(n6627), .A2(n6626), .ZN(n7978) );
  AOI211_X1 U8263 ( .C1(n6627), .C2(n6626), .A(n8701), .B(n7978), .ZN(n6631)
         );
  NOR2_X1 U8264 ( .A1(n7884), .A2(n8692), .ZN(n6630) );
  INV_X1 U8265 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8742) );
  OAI22_X1 U8266 ( .A1(n8698), .A2(n7812), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8742), .ZN(n6629) );
  OAI22_X1 U8267 ( .A1(n7807), .A2(n8686), .B1(n8687), .B2(n7987), .ZN(n6628)
         );
  OR4_X1 U8268 ( .A1(n6631), .A2(n6630), .A3(n6629), .A4(n6628), .ZN(P2_U3243)
         );
  NAND2_X1 U8269 ( .A1(n6633), .A2(P2_U3152), .ZN(n8428) );
  AND2_X1 U8270 ( .A1(n4481), .A2(P2_U3152), .ZN(n7781) );
  OAI222_X1 U8271 ( .A1(n8428), .A2(n6632), .B1(n4477), .B2(n6637), .C1(
        P2_U3152), .C2(n6701), .ZN(P2_U3357) );
  INV_X1 U8272 ( .A(n6781), .ZN(n6885) );
  INV_X1 U8273 ( .A(n6634), .ZN(n6642) );
  NAND2_X1 U8274 ( .A1(n4481), .A2(P1_U3084), .ZN(n9595) );
  OAI222_X1 U8275 ( .A1(n6885), .A2(P1_U3084), .B1(n9599), .B2(n6642), .C1(
        n6635), .C2(n9595), .ZN(P1_U3349) );
  INV_X1 U8276 ( .A(n9595), .ZN(n9592) );
  AOI22_X1 U8277 ( .A1(n9592), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n9214), .ZN(n6636) );
  OAI21_X1 U8278 ( .B1(n6637), .B2(n9599), .A(n6636), .ZN(P1_U3352) );
  AOI22_X1 U8279 ( .A1(n9592), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n6892), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6638) );
  OAI21_X1 U8280 ( .B1(n6648), .B2(n9599), .A(n6638), .ZN(P1_U3351) );
  AOI22_X1 U8281 ( .A1(n6809), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n9592), .ZN(n6639) );
  OAI21_X1 U8282 ( .B1(n6643), .B2(n9599), .A(n6639), .ZN(P1_U3350) );
  INV_X1 U8283 ( .A(n6640), .ZN(n6645) );
  INV_X1 U8284 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6641) );
  OAI222_X1 U8285 ( .A1(n9771), .A2(P1_U3084), .B1(n9599), .B2(n6645), .C1(
        n6641), .C2(n9595), .ZN(P1_U3348) );
  INV_X1 U8286 ( .A(n8428), .ZN(n7006) );
  OAI222_X1 U8287 ( .A1(n9087), .A2(n4596), .B1(n4477), .B2(n6642), .C1(
        P2_U3152), .C2(n6725), .ZN(P2_U3354) );
  OAI222_X1 U8288 ( .A1(n9087), .A2(n6644), .B1(n4477), .B2(n6643), .C1(
        P2_U3152), .C2(n6710), .ZN(P2_U3355) );
  INV_X1 U8289 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6646) );
  INV_X1 U8290 ( .A(n6747), .ZN(n6739) );
  OAI222_X1 U8291 ( .A1(n9087), .A2(n6646), .B1(n4477), .B2(n6645), .C1(
        P2_U3152), .C2(n6739), .ZN(P2_U3353) );
  OAI222_X1 U8292 ( .A1(n9087), .A2(n6649), .B1(n4477), .B2(n6648), .C1(
        P2_U3152), .C2(n6647), .ZN(P2_U3356) );
  INV_X1 U8293 ( .A(n6789), .ZN(n9786) );
  INV_X1 U8294 ( .A(n6650), .ZN(n6652) );
  INV_X1 U8295 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6651) );
  OAI222_X1 U8296 ( .A1(n9786), .A2(P1_U3084), .B1(n9599), .B2(n6652), .C1(
        n6651), .C2(n9595), .ZN(P1_U3347) );
  INV_X1 U8297 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6653) );
  INV_X1 U8298 ( .A(n6844), .ZN(n6755) );
  OAI222_X1 U8299 ( .A1(n9087), .A2(n6653), .B1(n4477), .B2(n6652), .C1(
        P2_U3152), .C2(n6755), .ZN(P2_U3352) );
  NAND2_X1 U8300 ( .A1(n8337), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6654) );
  OAI21_X1 U8301 ( .B1(n6859), .B2(n8337), .A(n6654), .ZN(P1_U3441) );
  INV_X1 U8302 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6656) );
  INV_X1 U8303 ( .A(n6655), .ZN(n6658) );
  INV_X1 U8304 ( .A(n6950), .ZN(n6957) );
  OAI222_X1 U8305 ( .A1(n9087), .A2(n6656), .B1(n4477), .B2(n6658), .C1(
        P2_U3152), .C2(n6957), .ZN(P2_U3351) );
  OAI222_X1 U8306 ( .A1(n6774), .A2(P1_U3084), .B1(n9599), .B2(n6658), .C1(
        n6657), .C2(n9595), .ZN(P1_U3346) );
  INV_X1 U8307 ( .A(n6659), .ZN(n6661) );
  OAI222_X1 U8308 ( .A1(n6827), .A2(P1_U3084), .B1(n9599), .B2(n6661), .C1(
        n6660), .C2(n9595), .ZN(P1_U3345) );
  INV_X1 U8309 ( .A(n7019), .ZN(n7025) );
  OAI222_X1 U8310 ( .A1(n8428), .A2(n6662), .B1(n4477), .B2(n6661), .C1(
        P2_U3152), .C2(n7025), .ZN(P2_U3350) );
  OR2_X1 U8311 ( .A1(n6663), .A2(P2_U3152), .ZN(n8631) );
  NAND2_X1 U8312 ( .A1(n10019), .A2(n8631), .ZN(n6665) );
  NAND2_X1 U8313 ( .A1(n6665), .A2(n6664), .ZN(n6668) );
  OR2_X1 U8314 ( .A1(n10019), .A2(n6666), .ZN(n6667) );
  AND2_X1 U8315 ( .A1(n6668), .A2(n6667), .ZN(n8799) );
  NOR2_X1 U8316 ( .A1(n10013), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8317 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6674) );
  INV_X1 U8318 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n6672) );
  NAND2_X1 U8319 ( .A1(n6062), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6671) );
  INV_X1 U8320 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6669) );
  OR2_X1 U8321 ( .A1(n6361), .A2(n6669), .ZN(n6670) );
  OAI211_X1 U8322 ( .C1(n6037), .C2(n6672), .A(n6671), .B(n6670), .ZN(n8801)
         );
  NAND2_X1 U8323 ( .A1(n8801), .A2(P2_U3966), .ZN(n6673) );
  OAI21_X1 U8324 ( .B1(P2_U3966), .B2(n6674), .A(n6673), .ZN(P2_U3583) );
  NAND2_X1 U8325 ( .A1(n7157), .A2(P2_U3966), .ZN(n6675) );
  OAI21_X1 U8326 ( .B1(P2_U3966), .B2(n5176), .A(n6675), .ZN(P2_U3552) );
  INV_X1 U8327 ( .A(n6127), .ZN(n6677) );
  AOI22_X1 U8328 ( .A1(n9816), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9592), .ZN(n6676) );
  OAI21_X1 U8329 ( .B1(n6677), .B2(n9599), .A(n6676), .ZN(P1_U3344) );
  INV_X1 U8330 ( .A(n7211), .ZN(n7217) );
  OAI222_X1 U8331 ( .A1(n8428), .A2(n10383), .B1(n4477), .B2(n6677), .C1(n7217), .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8332 ( .A(n6678), .ZN(n6681) );
  AOI22_X1 U8333 ( .A1(n7589), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n7006), .ZN(n6679) );
  OAI21_X1 U8334 ( .B1(n6681), .B2(n4477), .A(n6679), .ZN(P2_U3348) );
  AOI22_X1 U8335 ( .A1(n9823), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9592), .ZN(n6680) );
  OAI21_X1 U8336 ( .B1(n6681), .B2(n9599), .A(n6680), .ZN(P1_U3343) );
  INV_X1 U8337 ( .A(n6682), .ZN(n6685) );
  AOI22_X1 U8338 ( .A1(n8731), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n7006), .ZN(n6683) );
  OAI21_X1 U8339 ( .B1(n6685), .B2(n4477), .A(n6683), .ZN(P2_U3347) );
  OAI222_X1 U8340 ( .A1(P1_U3084), .A2(n7493), .B1(n9599), .B2(n6685), .C1(
        n6684), .C2(n9595), .ZN(P1_U3342) );
  INV_X1 U8341 ( .A(n6701), .ZN(n9605) );
  INV_X1 U8342 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6686) );
  INV_X1 U8343 ( .A(n6687), .ZN(n9602) );
  NOR3_X1 U8344 ( .A1(n10015), .A2(n10008), .A3(n9602), .ZN(n9601) );
  XNOR2_X1 U8345 ( .A(n9617), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n9614) );
  NOR2_X1 U8346 ( .A1(n9615), .A2(n9614), .ZN(n9613) );
  AOI21_X1 U8347 ( .B1(n9617), .B2(P2_REG2_REG_2__SCAN_IN), .A(n9613), .ZN(
        n6696) );
  NAND2_X1 U8348 ( .A1(n6717), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6688) );
  OAI21_X1 U8349 ( .B1(n6717), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6688), .ZN(
        n6695) );
  OR2_X1 U8350 ( .A1(n6689), .A2(P2_U3152), .ZN(n6690) );
  OAI211_X1 U8351 ( .C1(n10019), .C2(n6691), .A(n8631), .B(n6690), .ZN(n6693)
         );
  NAND2_X1 U8352 ( .A1(n6693), .A2(n6692), .ZN(n6704) );
  AND2_X1 U8353 ( .A1(n6704), .A2(n8724), .ZN(n6697) );
  NOR2_X1 U8354 ( .A1(n6697), .A2(n8627), .ZN(n10009) );
  NAND2_X1 U8355 ( .A1(n10009), .A2(n6694), .ZN(n9612) );
  AOI211_X1 U8356 ( .C1(n6696), .C2(n6695), .A(n6713), .B(n9612), .ZN(n6712)
         );
  INV_X1 U8357 ( .A(n6697), .ZN(n6698) );
  AND2_X1 U8358 ( .A1(n4474), .A2(n6698), .ZN(n9618) );
  NOR2_X1 U8359 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6039), .ZN(n6699) );
  AOI21_X1 U8360 ( .B1(n10013), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6699), .ZN(
        n6709) );
  NAND2_X1 U8361 ( .A1(n9617), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6702) );
  MUX2_X1 U8362 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6700), .S(n9617), .Z(n9620)
         );
  XNOR2_X1 U8363 ( .A(n6701), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n9608) );
  NAND3_X1 U8364 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n9608), .ZN(n9606) );
  OAI21_X1 U8365 ( .B1(n6701), .B2(n10352), .A(n9606), .ZN(n9621) );
  NAND2_X1 U8366 ( .A1(n9620), .A2(n9621), .ZN(n9619) );
  NAND2_X1 U8367 ( .A1(n6702), .A2(n9619), .ZN(n6707) );
  MUX2_X1 U8368 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6703), .S(n6717), .Z(n6706)
         );
  INV_X1 U8369 ( .A(n6704), .ZN(n6705) );
  NAND2_X1 U8370 ( .A1(n6706), .A2(n6707), .ZN(n6718) );
  OAI211_X1 U8371 ( .C1(n6707), .C2(n6706), .A(n10010), .B(n6718), .ZN(n6708)
         );
  OAI211_X1 U8372 ( .C1(n10005), .C2(n6710), .A(n6709), .B(n6708), .ZN(n6711)
         );
  OR2_X1 U8373 ( .A1(n6712), .A2(n6711), .ZN(P2_U3248) );
  NAND2_X1 U8374 ( .A1(n6732), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6714) );
  OAI21_X1 U8375 ( .B1(n6732), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6714), .ZN(
        n6715) );
  AOI211_X1 U8376 ( .C1(n6716), .C2(n6715), .A(n6728), .B(n9612), .ZN(n6727)
         );
  NOR2_X1 U8377 ( .A1(n6038), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6987) );
  AOI21_X1 U8378 ( .B1(n10013), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6987), .ZN(
        n6724) );
  NAND2_X1 U8379 ( .A1(n6717), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6719) );
  NAND2_X1 U8380 ( .A1(n6719), .A2(n6718), .ZN(n6722) );
  MUX2_X1 U8381 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6720), .S(n6732), .Z(n6721)
         );
  NAND2_X1 U8382 ( .A1(n6721), .A2(n6722), .ZN(n6733) );
  OAI211_X1 U8383 ( .C1(n6722), .C2(n6721), .A(n10010), .B(n6733), .ZN(n6723)
         );
  OAI211_X1 U8384 ( .C1(n10005), .C2(n6725), .A(n6724), .B(n6723), .ZN(n6726)
         );
  OR2_X1 U8385 ( .A1(n6727), .A2(n6726), .ZN(P2_U3249) );
  NAND2_X1 U8386 ( .A1(n6747), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6729) );
  OAI21_X1 U8387 ( .B1(n6747), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6729), .ZN(
        n6730) );
  NOR2_X1 U8388 ( .A1(n6731), .A2(n6730), .ZN(n6742) );
  AOI211_X1 U8389 ( .C1(n6731), .C2(n6730), .A(n6742), .B(n9612), .ZN(n6741)
         );
  INV_X1 U8390 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10408) );
  NOR2_X1 U8391 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10408), .ZN(n6998) );
  AOI21_X1 U8392 ( .B1(n10013), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6998), .ZN(
        n6738) );
  NAND2_X1 U8393 ( .A1(n6732), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6734) );
  NAND2_X1 U8394 ( .A1(n6734), .A2(n6733), .ZN(n6736) );
  MUX2_X1 U8395 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n7074), .S(n6747), .Z(n6735)
         );
  NAND2_X1 U8396 ( .A1(n6735), .A2(n6736), .ZN(n6748) );
  OAI211_X1 U8397 ( .C1(n6736), .C2(n6735), .A(n10010), .B(n6748), .ZN(n6737)
         );
  OAI211_X1 U8398 ( .C1(n10005), .C2(n6739), .A(n6738), .B(n6737), .ZN(n6740)
         );
  OR2_X1 U8399 ( .A1(n6741), .A2(n6740), .ZN(P2_U3250) );
  NAND2_X1 U8400 ( .A1(n6844), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6743) );
  OAI21_X1 U8401 ( .B1(n6844), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6743), .ZN(
        n6744) );
  AOI211_X1 U8402 ( .C1(n6745), .C2(n6744), .A(n6840), .B(n9612), .ZN(n6757)
         );
  NAND2_X1 U8403 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7041) );
  INV_X1 U8404 ( .A(n7041), .ZN(n6746) );
  AOI21_X1 U8405 ( .B1(n10013), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6746), .ZN(
        n6754) );
  NAND2_X1 U8406 ( .A1(n6747), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6749) );
  NAND2_X1 U8407 ( .A1(n6749), .A2(n6748), .ZN(n6752) );
  MUX2_X1 U8408 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6750), .S(n6844), .Z(n6751)
         );
  NAND2_X1 U8409 ( .A1(n6751), .A2(n6752), .ZN(n6845) );
  OAI211_X1 U8410 ( .C1(n6752), .C2(n6751), .A(n10010), .B(n6845), .ZN(n6753)
         );
  OAI211_X1 U8411 ( .C1(n10005), .C2(n6755), .A(n6754), .B(n6753), .ZN(n6756)
         );
  OR2_X1 U8412 ( .A1(n6757), .A2(n6756), .ZN(P2_U3251) );
  NOR2_X1 U8413 ( .A1(n6789), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6769) );
  NAND2_X1 U8414 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6784), .ZN(n6767) );
  INV_X1 U8415 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6758) );
  MUX2_X1 U8416 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6758), .S(n6784), .Z(n9774)
         );
  INV_X1 U8417 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6766) );
  MUX2_X1 U8418 ( .A(n6766), .B(P1_REG1_REG_4__SCAN_IN), .S(n6781), .Z(n6883)
         );
  XNOR2_X1 U8419 ( .A(n6892), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n6890) );
  INV_X1 U8420 ( .A(n6890), .ZN(n6761) );
  INV_X1 U8421 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6759) );
  MUX2_X1 U8422 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6759), .S(n9214), .Z(n9219)
         );
  AND2_X1 U8423 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9220) );
  NAND2_X1 U8424 ( .A1(n9219), .A2(n9220), .ZN(n9218) );
  NAND2_X1 U8425 ( .A1(n9214), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6760) );
  NAND2_X1 U8426 ( .A1(n9218), .A2(n6760), .ZN(n6891) );
  NAND2_X1 U8427 ( .A1(n6761), .A2(n6891), .ZN(n6763) );
  NAND2_X1 U8428 ( .A1(n6892), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6762) );
  NAND2_X1 U8429 ( .A1(n6763), .A2(n6762), .ZN(n6801) );
  INV_X1 U8430 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6764) );
  MUX2_X1 U8431 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6764), .S(n6809), .Z(n6802)
         );
  NAND2_X1 U8432 ( .A1(n6801), .A2(n6802), .ZN(n6800) );
  NAND2_X1 U8433 ( .A1(n6809), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6765) );
  NAND2_X1 U8434 ( .A1(n6800), .A2(n6765), .ZN(n6884) );
  NOR2_X1 U8435 ( .A1(n6883), .A2(n6884), .ZN(n6882) );
  AOI21_X1 U8436 ( .B1(n6885), .B2(n6766), .A(n6882), .ZN(n9775) );
  NAND2_X1 U8437 ( .A1(n9774), .A2(n9775), .ZN(n9773) );
  NAND2_X1 U8438 ( .A1(n6767), .A2(n9773), .ZN(n9790) );
  INV_X1 U8439 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6768) );
  MUX2_X1 U8440 ( .A(n6768), .B(P1_REG1_REG_6__SCAN_IN), .S(n6789), .Z(n9789)
         );
  NOR2_X1 U8441 ( .A1(n9790), .A2(n9789), .ZN(n9788) );
  NOR2_X1 U8442 ( .A1(n6769), .A2(n9788), .ZN(n6771) );
  INV_X1 U8443 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9998) );
  AOI22_X1 U8444 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6774), .B1(n6829), .B2(
        n9998), .ZN(n6770) );
  NOR2_X1 U8445 ( .A1(n6771), .A2(n6770), .ZN(n6816) );
  AOI21_X1 U8446 ( .B1(n6771), .B2(n6770), .A(n6816), .ZN(n6799) );
  NAND2_X1 U8447 ( .A1(n6876), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7951) );
  INV_X1 U8448 ( .A(n8345), .ZN(n6874) );
  NOR2_X1 U8449 ( .A1(n7951), .A2(n6874), .ZN(n6772) );
  NAND2_X1 U8450 ( .A1(n9751), .A2(n6772), .ZN(n9921) );
  NOR2_X1 U8451 ( .A1(n7951), .A2(n8345), .ZN(n6773) );
  AOI22_X1 U8452 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6829), .B1(n6774), .B2(
        n5297), .ZN(n6791) );
  INV_X1 U8453 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6775) );
  NAND2_X1 U8454 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6871) );
  INV_X1 U8455 ( .A(n6871), .ZN(n9216) );
  NAND2_X1 U8456 ( .A1(n9214), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6776) );
  NAND2_X1 U8457 ( .A1(n9215), .A2(n6776), .ZN(n6894) );
  INV_X1 U8458 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6777) );
  XNOR2_X1 U8459 ( .A(n6892), .B(n6777), .ZN(n6895) );
  NAND2_X1 U8460 ( .A1(n6894), .A2(n6895), .ZN(n6893) );
  NAND2_X1 U8461 ( .A1(n6892), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U8462 ( .A1(n6893), .A2(n6778), .ZN(n6804) );
  INV_X1 U8463 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6779) );
  XNOR2_X1 U8464 ( .A(n6809), .B(n6779), .ZN(n6805) );
  NAND2_X1 U8465 ( .A1(n6809), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6780) );
  XNOR2_X1 U8466 ( .A(n6781), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n6878) );
  NAND2_X1 U8467 ( .A1(n6885), .A2(n6782), .ZN(n6783) );
  NOR2_X1 U8468 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6784), .ZN(n6785) );
  AOI21_X1 U8469 ( .B1(n6784), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6785), .ZN(
        n9766) );
  NAND2_X1 U8470 ( .A1(n9765), .A2(n9766), .ZN(n9764) );
  INV_X1 U8471 ( .A(n6785), .ZN(n6786) );
  NAND2_X1 U8472 ( .A1(n9764), .A2(n6786), .ZN(n9781) );
  OR2_X1 U8473 ( .A1(n6789), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6788) );
  NAND2_X1 U8474 ( .A1(n6789), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6787) );
  NAND2_X1 U8475 ( .A1(n6788), .A2(n6787), .ZN(n9780) );
  NOR2_X1 U8476 ( .A1(n9781), .A2(n9780), .ZN(n9779) );
  OAI21_X1 U8477 ( .B1(n6791), .B2(n6790), .A(n6828), .ZN(n6797) );
  INV_X1 U8478 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6795) );
  NAND2_X1 U8479 ( .A1(n6874), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7947) );
  NOR2_X1 U8480 ( .A1(n6876), .A2(n7947), .ZN(n6793) );
  NAND2_X1 U8481 ( .A1(n9751), .A2(n6793), .ZN(n9914) );
  INV_X1 U8482 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10369) );
  NOR2_X1 U8483 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10369), .ZN(n7179) );
  AOI21_X1 U8484 ( .B1(n9883), .B2(n6829), .A(n7179), .ZN(n6794) );
  OAI21_X1 U8485 ( .B1(n9924), .B2(n6795), .A(n6794), .ZN(n6796) );
  AOI21_X1 U8486 ( .B1(n9911), .B2(n6797), .A(n6796), .ZN(n6798) );
  OAI21_X1 U8487 ( .B1(n6799), .B2(n9921), .A(n6798), .ZN(P1_U3248) );
  INV_X1 U8488 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10347) );
  NOR2_X1 U8489 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6925), .ZN(n6924) );
  INV_X1 U8490 ( .A(n9921), .ZN(n9900) );
  OAI211_X1 U8491 ( .C1(n6802), .C2(n6801), .A(n9900), .B(n6800), .ZN(n6807)
         );
  OAI211_X1 U8492 ( .C1(n6805), .C2(n6804), .A(n9911), .B(n6803), .ZN(n6806)
         );
  NAND2_X1 U8493 ( .A1(n6807), .A2(n6806), .ZN(n6808) );
  AOI211_X1 U8494 ( .C1(n9883), .C2(n6809), .A(n6924), .B(n6808), .ZN(n6810)
         );
  OAI21_X1 U8495 ( .B1(n10347), .B2(n9924), .A(n6810), .ZN(P1_U3244) );
  INV_X1 U8496 ( .A(n6811), .ZN(n6814) );
  INV_X1 U8497 ( .A(n7769), .ZN(n7765) );
  OAI222_X1 U8498 ( .A1(n8428), .A2(n6812), .B1(n4477), .B2(n6814), .C1(
        P2_U3152), .C2(n7765), .ZN(P2_U3346) );
  OAI222_X1 U8499 ( .A1(n7494), .A2(P1_U3084), .B1(n9599), .B2(n6814), .C1(
        n6813), .C2(n9595), .ZN(P1_U3341) );
  NOR2_X1 U8500 ( .A1(n9823), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6821) );
  NOR2_X1 U8501 ( .A1(n9816), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6819) );
  INV_X1 U8502 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10000) );
  MUX2_X1 U8503 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10000), .S(n9803), .Z(n9797)
         );
  NOR2_X1 U8504 ( .A1(n6829), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6815) );
  OR2_X1 U8505 ( .A1(n6816), .A2(n6815), .ZN(n9799) );
  INV_X1 U8506 ( .A(n9799), .ZN(n6817) );
  NAND2_X1 U8507 ( .A1(n9797), .A2(n6817), .ZN(n9800) );
  OAI21_X1 U8508 ( .B1(n6827), .B2(n10000), .A(n9800), .ZN(n9818) );
  INV_X1 U8509 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6818) );
  MUX2_X1 U8510 ( .A(n6818), .B(P1_REG1_REG_9__SCAN_IN), .S(n9816), .Z(n9819)
         );
  NOR2_X1 U8511 ( .A1(n9818), .A2(n9819), .ZN(n9817) );
  NOR2_X1 U8512 ( .A1(n6819), .A2(n9817), .ZN(n9835) );
  INV_X1 U8513 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6820) );
  MUX2_X1 U8514 ( .A(n6820), .B(P1_REG1_REG_10__SCAN_IN), .S(n9823), .Z(n9834)
         );
  NOR2_X1 U8515 ( .A1(n9835), .A2(n9834), .ZN(n9833) );
  NOR2_X1 U8516 ( .A1(n6821), .A2(n9833), .ZN(n6823) );
  INV_X1 U8517 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9743) );
  AOI22_X1 U8518 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n7493), .B1(n7487), .B2(
        n9743), .ZN(n6822) );
  NOR2_X1 U8519 ( .A1(n6823), .A2(n6822), .ZN(n7492) );
  AOI21_X1 U8520 ( .B1(n6823), .B2(n6822), .A(n7492), .ZN(n6839) );
  INV_X1 U8521 ( .A(n9924), .ZN(n9762) );
  INV_X1 U8522 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6824) );
  NOR2_X1 U8523 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6824), .ZN(n7641) );
  NOR2_X1 U8524 ( .A1(n9914), .A2(n7493), .ZN(n6825) );
  AOI211_X1 U8525 ( .C1(n9762), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n7641), .B(
        n6825), .ZN(n6838) );
  NOR2_X1 U8526 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7487), .ZN(n6826) );
  AOI21_X1 U8527 ( .B1(n7487), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6826), .ZN(
        n6835) );
  AOI22_X1 U8528 ( .A1(n9803), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7443), .B2(
        n6827), .ZN(n9795) );
  OAI21_X1 U8529 ( .B1(n9803), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6830), .ZN(
        n9813) );
  NAND2_X1 U8530 ( .A1(n9816), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6831) );
  OAI21_X1 U8531 ( .B1(n9816), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6831), .ZN(
        n9812) );
  NOR2_X1 U8532 ( .A1(n9813), .A2(n9812), .ZN(n9811) );
  OR2_X1 U8533 ( .A1(n9823), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6833) );
  NAND2_X1 U8534 ( .A1(n9823), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6832) );
  NAND2_X1 U8535 ( .A1(n6833), .A2(n6832), .ZN(n9825) );
  OAI21_X1 U8536 ( .B1(n6835), .B2(n6834), .A(n7486), .ZN(n6836) );
  NAND2_X1 U8537 ( .A1(n6836), .A2(n9911), .ZN(n6837) );
  OAI211_X1 U8538 ( .C1(n6839), .C2(n9921), .A(n6838), .B(n6837), .ZN(P1_U3252) );
  INV_X1 U8539 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6841) );
  MUX2_X1 U8540 ( .A(n6841), .B(P2_REG2_REG_7__SCAN_IN), .S(n6950), .Z(n6842)
         );
  AOI211_X1 U8541 ( .C1(n6843), .C2(n6842), .A(n6949), .B(n9612), .ZN(n6853)
         );
  AND2_X1 U8542 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7013) );
  AOI21_X1 U8543 ( .B1(n10013), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7013), .ZN(
        n6851) );
  NAND2_X1 U8544 ( .A1(n6844), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6846) );
  NAND2_X1 U8545 ( .A1(n6846), .A2(n6845), .ZN(n6849) );
  MUX2_X1 U8546 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6847), .S(n6950), .Z(n6848)
         );
  NAND2_X1 U8547 ( .A1(n6848), .A2(n6849), .ZN(n6956) );
  OAI211_X1 U8548 ( .C1(n6849), .C2(n6848), .A(n10010), .B(n6956), .ZN(n6850)
         );
  OAI211_X1 U8549 ( .C1(n10005), .C2(n6957), .A(n6851), .B(n6850), .ZN(n6852)
         );
  OR2_X1 U8550 ( .A1(n6853), .A2(n6852), .ZN(P2_U3252) );
  INV_X1 U8551 ( .A(n7052), .ZN(n6857) );
  AND2_X1 U8552 ( .A1(n6854), .A2(n7192), .ZN(n7280) );
  INV_X1 U8553 ( .A(n7280), .ZN(n6855) );
  OAI21_X1 U8554 ( .B1(n7192), .B2(n6854), .A(n6855), .ZN(n8274) );
  NAND2_X1 U8555 ( .A1(n8338), .A2(n7052), .ZN(n6856) );
  INV_X1 U8556 ( .A(n7186), .ZN(n8069) );
  OAI22_X1 U8557 ( .A1(n8274), .A2(n6856), .B1(n8069), .B2(n9670), .ZN(n7056)
         );
  AOI21_X1 U8558 ( .B1(n7192), .B2(n6857), .A(n7056), .ZN(n6982) );
  INV_X1 U8559 ( .A(n6858), .ZN(n6860) );
  AND2_X1 U8560 ( .A1(n6860), .A2(n6859), .ZN(n6862) );
  AND2_X2 U8561 ( .A1(n8259), .A2(n8139), .ZN(n8258) );
  NAND2_X1 U8562 ( .A1(n9950), .A2(n5907), .ZN(n6861) );
  INV_X1 U8563 ( .A(n9928), .ZN(n7049) );
  INV_X1 U8564 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6863) );
  OR2_X1 U8565 ( .A1(n9992), .A2(n6863), .ZN(n6864) );
  OAI21_X1 U8566 ( .B1(n6982), .B2(n9990), .A(n6864), .ZN(P1_U3454) );
  INV_X1 U8567 ( .A(n9170), .ZN(n9199) );
  INV_X1 U8568 ( .A(n7192), .ZN(n8067) );
  INV_X1 U8569 ( .A(n6865), .ZN(n6866) );
  AOI21_X1 U8570 ( .B1(n7047), .B2(n6866), .A(n9170), .ZN(n6942) );
  NAND2_X1 U8571 ( .A1(n6942), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6870) );
  OAI21_X1 U8572 ( .B1(n4568), .B2(n6868), .A(n6867), .ZN(n6873) );
  AOI22_X1 U8573 ( .A1(n9660), .A2(n6873), .B1(n9196), .B2(n7186), .ZN(n6869)
         );
  OAI211_X1 U8574 ( .C1(n9199), .C2(n8067), .A(n6870), .B(n6869), .ZN(P1_U3230) );
  NAND2_X1 U8575 ( .A1(n6874), .A2(n6871), .ZN(n6872) );
  NAND2_X1 U8576 ( .A1(n6876), .A2(n6872), .ZN(n9753) );
  AOI21_X1 U8577 ( .B1(n6873), .B2(n8345), .A(n9753), .ZN(n6877) );
  INV_X1 U8578 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10395) );
  NAND2_X1 U8579 ( .A1(n6874), .A2(n10395), .ZN(n6875) );
  AOI21_X1 U8580 ( .B1(n6876), .B2(n6875), .A(P1_IR_REG_0__SCAN_IN), .ZN(n9752) );
  NOR3_X1 U8581 ( .A1(n6877), .A2(n9752), .A3(n9211), .ZN(n6899) );
  NOR2_X1 U8582 ( .A1(n9924), .A2(n10365), .ZN(n6889) );
  XNOR2_X1 U8583 ( .A(n6879), .B(n6878), .ZN(n6880) );
  NAND2_X1 U8584 ( .A1(n9911), .A2(n6880), .ZN(n6881) );
  NAND2_X1 U8585 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n6968) );
  NAND2_X1 U8586 ( .A1(n6881), .A2(n6968), .ZN(n6888) );
  AOI21_X1 U8587 ( .B1(n6884), .B2(n6883), .A(n6882), .ZN(n6886) );
  OAI22_X1 U8588 ( .A1(n6886), .A2(n9921), .B1(n9914), .B2(n6885), .ZN(n6887)
         );
  OR4_X1 U8589 ( .A1(n6899), .A2(n6889), .A3(n6888), .A4(n6887), .ZN(P1_U3245)
         );
  XOR2_X1 U8590 ( .A(n6891), .B(n6890), .Z(n6898) );
  AOI22_X1 U8591 ( .A1(n9883), .A2(n6892), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        P1_U3084), .ZN(n6897) );
  OAI211_X1 U8592 ( .C1(n6895), .C2(n6894), .A(n9911), .B(n6893), .ZN(n6896)
         );
  OAI211_X1 U8593 ( .C1(n6898), .C2(n9921), .A(n6897), .B(n6896), .ZN(n6900)
         );
  AOI211_X1 U8594 ( .C1(n9762), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n6900), .B(
        n6899), .ZN(n6901) );
  INV_X1 U8595 ( .A(n6901), .ZN(P1_U3243) );
  INV_X1 U8596 ( .A(n9858), .ZN(n7495) );
  INV_X1 U8597 ( .A(n6902), .ZN(n6904) );
  OAI222_X1 U8598 ( .A1(P1_U3084), .A2(n7495), .B1(n9599), .B2(n6904), .C1(
        n6903), .C2(n9595), .ZN(P1_U3340) );
  INV_X1 U8599 ( .A(n7826), .ZN(n7821) );
  OAI222_X1 U8600 ( .A1(n8428), .A2(n6905), .B1(n4477), .B2(n6904), .C1(n7821), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  XNOR2_X1 U8601 ( .A(n6907), .B(n6906), .ZN(n6913) );
  AOI22_X1 U8602 ( .A1(n8047), .A2(n4480), .B1(n8048), .B2(n8723), .ZN(n6912)
         );
  INV_X1 U8603 ( .A(n6908), .ZN(n6909) );
  NAND2_X1 U8604 ( .A1(n6910), .A2(n6909), .ZN(n8638) );
  AOI22_X1 U8605 ( .A1(n6494), .A2(n7152), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n8638), .ZN(n6911) );
  OAI211_X1 U8606 ( .C1(n6913), .C2(n8701), .A(n6912), .B(n6911), .ZN(P2_U3239) );
  NAND2_X1 U8607 ( .A1(n6915), .A2(n6914), .ZN(n6916) );
  AOI21_X1 U8608 ( .B1(n6917), .B2(n6916), .A(n8701), .ZN(n6918) );
  AOI21_X1 U8609 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n8638), .A(n6918), .ZN(
        n6920) );
  AOI22_X1 U8610 ( .A1(n8047), .A2(n7157), .B1(n8048), .B2(n6517), .ZN(n6919)
         );
  OAI211_X1 U8611 ( .C1(n6513), .C2(n8692), .A(n6920), .B(n6919), .ZN(P2_U3224) );
  XOR2_X1 U8612 ( .A(n6922), .B(n6921), .Z(n6928) );
  NOR2_X1 U8613 ( .A1(n9193), .A2(n7344), .ZN(n6923) );
  AOI211_X1 U8614 ( .C1(n9196), .C2(n9212), .A(n6924), .B(n6923), .ZN(n6927)
         );
  AOI22_X1 U8615 ( .A1(n9191), .A2(n6925), .B1(n9170), .B2(n7351), .ZN(n6926)
         );
  OAI211_X1 U8616 ( .C1(n6928), .C2(n9186), .A(n6927), .B(n6926), .ZN(P1_U3216) );
  XNOR2_X1 U8617 ( .A(n6930), .B(n6929), .ZN(n6932) );
  XNOR2_X1 U8618 ( .A(n6932), .B(n6931), .ZN(n6937) );
  AOI22_X1 U8619 ( .A1(n9655), .A2(n6854), .B1(n9196), .B2(n5204), .ZN(n6934)
         );
  OAI21_X1 U8620 ( .B1(n9199), .B2(n9934), .A(n6934), .ZN(n6935) );
  AOI21_X1 U8621 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6942), .A(n6935), .ZN(
        n6936) );
  OAI21_X1 U8622 ( .B1(n9186), .B2(n6937), .A(n6936), .ZN(P1_U3220) );
  XOR2_X1 U8623 ( .A(n6938), .B(n6939), .Z(n6944) );
  INV_X1 U8624 ( .A(n7315), .ZN(n9939) );
  AOI22_X1 U8625 ( .A1(n9655), .A2(n7186), .B1(n9196), .B2(n9213), .ZN(n6940)
         );
  OAI21_X1 U8626 ( .B1(n9199), .B2(n9939), .A(n6940), .ZN(n6941) );
  AOI21_X1 U8627 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n6942), .A(n6941), .ZN(
        n6943) );
  OAI21_X1 U8628 ( .B1(n9186), .B2(n6944), .A(n6943), .ZN(P1_U3235) );
  INV_X1 U8629 ( .A(n6945), .ZN(n6947) );
  OAI222_X1 U8630 ( .A1(P1_U3084), .A2(n9238), .B1(n9599), .B2(n6947), .C1(
        n6946), .C2(n9595), .ZN(P1_U3339) );
  INV_X1 U8631 ( .A(n8006), .ZN(n8013) );
  OAI222_X1 U8632 ( .A1(n8428), .A2(n6948), .B1(n4477), .B2(n6947), .C1(n8013), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8633 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6951) );
  MUX2_X1 U8634 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6951), .S(n7019), .Z(n6952)
         );
  INV_X1 U8635 ( .A(n6952), .ZN(n6953) );
  NOR2_X1 U8636 ( .A1(n6954), .A2(n6953), .ZN(n7018) );
  AOI211_X1 U8637 ( .C1(n6954), .C2(n6953), .A(n7018), .B(n9612), .ZN(n6964)
         );
  NAND2_X1 U8638 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7078) );
  INV_X1 U8639 ( .A(n7078), .ZN(n6955) );
  AOI21_X1 U8640 ( .B1(n10013), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6955), .ZN(
        n6962) );
  OAI21_X1 U8641 ( .B1(n6957), .B2(n6847), .A(n6956), .ZN(n6960) );
  MUX2_X1 U8642 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6958), .S(n7019), .Z(n6959)
         );
  NAND2_X1 U8643 ( .A1(n6959), .A2(n6960), .ZN(n7024) );
  OAI211_X1 U8644 ( .C1(n6960), .C2(n6959), .A(n10010), .B(n7024), .ZN(n6961)
         );
  OAI211_X1 U8645 ( .C1(n10005), .C2(n7025), .A(n6962), .B(n6961), .ZN(n6963)
         );
  OR2_X1 U8646 ( .A1(n6964), .A2(n6963), .ZN(P2_U3253) );
  XNOR2_X1 U8647 ( .A(n6966), .B(n6965), .ZN(n6967) );
  INV_X1 U8648 ( .A(n9210), .ZN(n7301) );
  OAI21_X1 U8649 ( .B1(n9652), .B2(n7301), .A(n6968), .ZN(n6969) );
  AOI21_X1 U8650 ( .B1(n9655), .B2(n9213), .A(n6969), .ZN(n6971) );
  AOI22_X1 U8651 ( .A1(n9191), .A2(n7331), .B1(n9170), .B2(n7332), .ZN(n6970)
         );
  OAI211_X1 U8652 ( .C1(n6972), .C2(n9186), .A(n6971), .B(n6970), .ZN(P1_U3228) );
  XNOR2_X1 U8653 ( .A(n6973), .B(n6974), .ZN(n6979) );
  NAND2_X1 U8654 ( .A1(n9631), .A2(n6039), .ZN(n6975) );
  OAI21_X1 U8655 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6039), .A(n6975), .ZN(n6977) );
  OAI22_X1 U8656 ( .A1(n8692), .A2(n6519), .B1(n8687), .B2(n4670), .ZN(n6976)
         );
  AOI211_X1 U8657 ( .C1(n8047), .C2(n6517), .A(n6977), .B(n6976), .ZN(n6978)
         );
  OAI21_X1 U8658 ( .B1(n8701), .B2(n6979), .A(n6978), .ZN(P2_U3220) );
  NAND2_X1 U8659 ( .A1(n10002), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6981) );
  OAI21_X1 U8660 ( .B1(n6982), .B2(n10002), .A(n6981), .ZN(P1_U3523) );
  NAND2_X1 U8661 ( .A1(n6983), .A2(n6984), .ZN(n6985) );
  AOI21_X1 U8662 ( .B1(n6986), .B2(n6985), .A(n8701), .ZN(n6994) );
  OAI22_X1 U8663 ( .A1(n8692), .A2(n10052), .B1(n8687), .B2(n7229), .ZN(n6993)
         );
  INV_X1 U8664 ( .A(n6987), .ZN(n6990) );
  INV_X1 U8665 ( .A(n7131), .ZN(n6988) );
  NAND2_X1 U8666 ( .A1(n9631), .A2(n6988), .ZN(n6989) );
  OAI211_X1 U8667 ( .C1(n8686), .C2(n6991), .A(n6990), .B(n6989), .ZN(n6992)
         );
  OR3_X1 U8668 ( .A1(n6994), .A2(n6993), .A3(n6992), .ZN(P2_U3232) );
  XNOR2_X1 U8669 ( .A(n7034), .B(n7033), .ZN(n7000) );
  INV_X1 U8670 ( .A(n9635), .ZN(n8696) );
  NAND2_X1 U8671 ( .A1(n8722), .A2(n8966), .ZN(n6996) );
  NAND2_X1 U8672 ( .A1(n8720), .A2(n8968), .ZN(n6995) );
  NAND2_X1 U8673 ( .A1(n6996), .A2(n6995), .ZN(n7067) );
  OAI22_X1 U8674 ( .A1(n8692), .A2(n7163), .B1(n8698), .B2(n7164), .ZN(n6997)
         );
  AOI211_X1 U8675 ( .C1(n8696), .C2(n7067), .A(n6998), .B(n6997), .ZN(n6999)
         );
  OAI21_X1 U8676 ( .B1(n7000), .B2(n8701), .A(n6999), .ZN(P2_U3229) );
  INV_X1 U8677 ( .A(n7001), .ZN(n7004) );
  INV_X1 U8678 ( .A(n8746), .ZN(n8014) );
  OAI222_X1 U8679 ( .A1(n8428), .A2(n7002), .B1(n4477), .B2(n7004), .C1(
        P2_U3152), .C2(n8014), .ZN(P2_U3343) );
  OAI222_X1 U8680 ( .A1(n9240), .A2(P1_U3084), .B1(n9599), .B2(n7004), .C1(
        n7003), .C2(n9595), .ZN(P1_U3338) );
  INV_X1 U8681 ( .A(n7005), .ZN(n7009) );
  AOI22_X1 U8682 ( .A1(n8757), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n7006), .ZN(n7007) );
  OAI21_X1 U8683 ( .B1(n7009), .B2(n4477), .A(n7007), .ZN(P2_U3342) );
  INV_X1 U8684 ( .A(n9882), .ZN(n9242) );
  OAI222_X1 U8685 ( .A1(P1_U3084), .A2(n9242), .B1(n9599), .B2(n7009), .C1(
        n7008), .C2(n9595), .ZN(P1_U3337) );
  XNOR2_X1 U8686 ( .A(n7011), .B(n7010), .ZN(n7017) );
  INV_X1 U8687 ( .A(n7108), .ZN(n7014) );
  AOI22_X1 U8688 ( .A1(n8966), .A2(n8720), .B1(n8718), .B2(n8968), .ZN(n7102)
         );
  NOR2_X1 U8689 ( .A1(n9635), .A2(n7102), .ZN(n7012) );
  AOI211_X1 U8690 ( .C1(n9631), .C2(n7014), .A(n7013), .B(n7012), .ZN(n7016)
         );
  NAND2_X1 U8691 ( .A1(n6494), .A2(n7420), .ZN(n7015) );
  OAI211_X1 U8692 ( .C1(n7017), .C2(n8701), .A(n7016), .B(n7015), .ZN(P2_U3215) );
  AOI21_X1 U8693 ( .B1(n7019), .B2(P2_REG2_REG_8__SCAN_IN), .A(n7018), .ZN(
        n7022) );
  NAND2_X1 U8694 ( .A1(n7211), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7020) );
  OAI21_X1 U8695 ( .B1(n7211), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7020), .ZN(
        n7021) );
  NOR2_X1 U8696 ( .A1(n7022), .A2(n7021), .ZN(n7210) );
  AOI211_X1 U8697 ( .C1(n7022), .C2(n7021), .A(n7210), .B(n9612), .ZN(n7032)
         );
  NAND2_X1 U8698 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7325) );
  INV_X1 U8699 ( .A(n7325), .ZN(n7023) );
  AOI21_X1 U8700 ( .B1(n10013), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7023), .ZN(
        n7030) );
  OAI21_X1 U8701 ( .B1(n7025), .B2(n6958), .A(n7024), .ZN(n7028) );
  MUX2_X1 U8702 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7026), .S(n7211), .Z(n7027)
         );
  NAND2_X1 U8703 ( .A1(n7027), .A2(n7028), .ZN(n7216) );
  OAI211_X1 U8704 ( .C1(n7028), .C2(n7027), .A(n10010), .B(n7216), .ZN(n7029)
         );
  OAI211_X1 U8705 ( .C1(n10005), .C2(n7217), .A(n7030), .B(n7029), .ZN(n7031)
         );
  OR2_X1 U8706 ( .A1(n7032), .A2(n7031), .ZN(P2_U3254) );
  OR2_X1 U8707 ( .A1(n7034), .A2(n7033), .ZN(n7037) );
  AND2_X1 U8708 ( .A1(n7037), .A2(n7035), .ZN(n7039) );
  NAND2_X1 U8709 ( .A1(n7037), .A2(n7036), .ZN(n7038) );
  OAI21_X1 U8710 ( .B1(n7040), .B2(n7039), .A(n7038), .ZN(n7045) );
  OAI22_X1 U8711 ( .A1(n8692), .A2(n10057), .B1(n8687), .B2(n7407), .ZN(n7044)
         );
  NAND2_X1 U8712 ( .A1(n8047), .A2(n8721), .ZN(n7042) );
  OAI211_X1 U8713 ( .C1(n8698), .C2(n7233), .A(n7042), .B(n7041), .ZN(n7043)
         );
  AOI211_X1 U8714 ( .C1(n7045), .C2(n9628), .A(n7044), .B(n7043), .ZN(n7046)
         );
  INV_X1 U8715 ( .A(n7046), .ZN(P2_U3241) );
  AND2_X1 U8716 ( .A1(n7048), .A2(n7047), .ZN(n7394) );
  NAND2_X1 U8717 ( .A1(n7394), .A2(n7049), .ZN(n7051) );
  AND2_X1 U8718 ( .A1(n9931), .A2(n5907), .ZN(n7050) );
  INV_X1 U8719 ( .A(n9709), .ZN(n9478) );
  NAND2_X1 U8720 ( .A1(n4555), .A2(n9960), .ZN(n9266) );
  OAI21_X1 U8721 ( .B1(n9691), .B2(n9713), .A(n7192), .ZN(n7058) );
  INV_X1 U8722 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7054) );
  NOR2_X1 U8723 ( .A1(n9693), .A2(n7054), .ZN(n7055) );
  OAI21_X1 U8724 ( .B1(n7056), .B2(n7055), .A(n9478), .ZN(n7057) );
  OAI211_X1 U8725 ( .C1(n10395), .C2(n9478), .A(n7058), .B(n7057), .ZN(
        P1_U3291) );
  INV_X1 U8726 ( .A(n7059), .ZN(n7084) );
  AOI22_X1 U8727 ( .A1(n9234), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9592), .ZN(n7060) );
  OAI21_X1 U8728 ( .B1(n7084), .B2(n9599), .A(n7060), .ZN(P1_U3336) );
  XOR2_X1 U8729 ( .A(n7061), .B(n8592), .Z(n7169) );
  OR2_X1 U8730 ( .A1(n7062), .A2(n7063), .ZN(n7065) );
  NAND2_X1 U8731 ( .A1(n7065), .A2(n7064), .ZN(n7066) );
  XNOR2_X1 U8732 ( .A(n8592), .B(n7066), .ZN(n7068) );
  AOI21_X1 U8733 ( .B1(n7068), .B2(n8971), .A(n7067), .ZN(n7172) );
  AOI211_X1 U8734 ( .C1(n7069), .C2(n7133), .A(n10078), .B(n7230), .ZN(n7168)
         );
  AOI21_X1 U8735 ( .B1(n9058), .B2(n7069), .A(n7168), .ZN(n7070) );
  OAI211_X1 U8736 ( .C1(n7169), .C2(n9054), .A(n7172), .B(n7070), .ZN(n7072)
         );
  NAND2_X1 U8737 ( .A1(n7072), .A2(n10086), .ZN(n7071) );
  OAI21_X1 U8738 ( .B1(n10086), .B2(n6064), .A(n7071), .ZN(P2_U3466) );
  INV_X1 U8739 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7074) );
  NAND2_X1 U8740 ( .A1(n7072), .A2(n10098), .ZN(n7073) );
  OAI21_X1 U8741 ( .B1(n10098), .B2(n7074), .A(n7073), .ZN(P2_U3525) );
  XNOR2_X1 U8742 ( .A(n7076), .B(n7075), .ZN(n7083) );
  INV_X1 U8743 ( .A(n7411), .ZN(n7077) );
  NAND2_X1 U8744 ( .A1(n9631), .A2(n7077), .ZN(n7079) );
  NAND2_X1 U8745 ( .A1(n7079), .A2(n7078), .ZN(n7081) );
  OAI22_X1 U8746 ( .A1(n7407), .A2(n8686), .B1(n8687), .B2(n7406), .ZN(n7080)
         );
  AOI211_X1 U8747 ( .C1(n10064), .C2(n6494), .A(n7081), .B(n7080), .ZN(n7082)
         );
  OAI21_X1 U8748 ( .B1(n7083), .B2(n8701), .A(n7082), .ZN(P2_U3223) );
  INV_X1 U8749 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7085) );
  INV_X1 U8750 ( .A(n8753), .ZN(n8777) );
  OAI222_X1 U8751 ( .A1(n8428), .A2(n7085), .B1(n4477), .B2(n7084), .C1(n8777), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8752 ( .A(n8981), .ZN(n8906) );
  XNOR2_X1 U8753 ( .A(n7086), .B(n7087), .ZN(n10034) );
  NAND2_X1 U8754 ( .A1(n6581), .A2(n10026), .ZN(n7088) );
  NAND3_X1 U8755 ( .A1(n7153), .A2(n10035), .A3(n7088), .ZN(n10031) );
  OAI22_X1 U8756 ( .A1(n7106), .A2(n10031), .B1(n7089), .B2(n8907), .ZN(n7090)
         );
  AOI21_X1 U8757 ( .B1(n8906), .B2(n10034), .A(n7090), .ZN(n7099) );
  INV_X1 U8758 ( .A(n8471), .ZN(n7091) );
  NOR2_X1 U8759 ( .A1(n8464), .A2(n7091), .ZN(n8589) );
  INV_X1 U8760 ( .A(n8635), .ZN(n7092) );
  NAND2_X1 U8761 ( .A1(n7086), .A2(n7092), .ZN(n7093) );
  NAND2_X1 U8762 ( .A1(n7093), .A2(n8971), .ZN(n7094) );
  OR2_X1 U8763 ( .A1(n8589), .A2(n7094), .ZN(n7096) );
  AOI22_X1 U8764 ( .A1(n8966), .A2(n7157), .B1(n6517), .B2(n8968), .ZN(n7095)
         );
  NAND2_X1 U8765 ( .A1(n7096), .A2(n7095), .ZN(n10032) );
  MUX2_X1 U8766 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10032), .S(n8877), .Z(n7097)
         );
  INV_X1 U8767 ( .A(n7097), .ZN(n7098) );
  OAI211_X1 U8768 ( .C1(n6513), .C2(n8977), .A(n7099), .B(n7098), .ZN(P2_U3295) );
  XNOR2_X1 U8769 ( .A(n7100), .B(n8595), .ZN(n7422) );
  XNOR2_X1 U8770 ( .A(n7101), .B(n8595), .ZN(n7103) );
  OAI21_X1 U8771 ( .B1(n7103), .B2(n8953), .A(n7102), .ZN(n7418) );
  NAND2_X1 U8772 ( .A1(n7418), .A2(n8877), .ZN(n7113) );
  INV_X1 U8773 ( .A(n7232), .ZN(n7105) );
  INV_X1 U8774 ( .A(n7412), .ZN(n7104) );
  AOI211_X1 U8775 ( .C1(n7420), .C2(n7105), .A(n10078), .B(n7104), .ZN(n7419)
         );
  INV_X1 U8776 ( .A(n7106), .ZN(n7111) );
  NOR2_X1 U8777 ( .A1(n8977), .A2(n7107), .ZN(n7110) );
  OAI22_X1 U8778 ( .A1(n8877), .A2(n6841), .B1(n7108), .B2(n8907), .ZN(n7109)
         );
  AOI211_X1 U8779 ( .C1(n7419), .C2(n7111), .A(n7110), .B(n7109), .ZN(n7112)
         );
  OAI211_X1 U8780 ( .C1(n7422), .C2(n8981), .A(n7113), .B(n7112), .ZN(P2_U3289) );
  INV_X1 U8781 ( .A(n7114), .ZN(n7120) );
  INV_X1 U8782 ( .A(n7115), .ZN(n7116) );
  OR2_X1 U8783 ( .A1(n7117), .A2(n7116), .ZN(n7372) );
  NAND2_X1 U8784 ( .A1(n7117), .A2(n7116), .ZN(n7118) );
  NAND2_X1 U8785 ( .A1(n7372), .A2(n7118), .ZN(n7119) );
  NOR2_X1 U8786 ( .A1(n7119), .A2(n7120), .ZN(n7375) );
  AOI21_X1 U8787 ( .B1(n7120), .B2(n7119), .A(n7375), .ZN(n7126) );
  NOR2_X1 U8788 ( .A1(n7246), .A2(n9976), .ZN(n9955) );
  INV_X1 U8789 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7121) );
  NOR2_X1 U8790 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7121), .ZN(n9768) );
  AOI21_X1 U8791 ( .B1(n9196), .B2(n9209), .A(n9768), .ZN(n7123) );
  NAND2_X1 U8792 ( .A1(n9655), .A2(n9212), .ZN(n7122) );
  OAI211_X1 U8793 ( .C1(n9665), .C2(n7244), .A(n7123), .B(n7122), .ZN(n7124)
         );
  AOI21_X1 U8794 ( .B1(n9659), .B2(n9955), .A(n7124), .ZN(n7125) );
  OAI21_X1 U8795 ( .B1(n7126), .B2(n9186), .A(n7125), .ZN(P1_U3225) );
  INV_X1 U8796 ( .A(n8591), .ZN(n7127) );
  XNOR2_X1 U8797 ( .A(n7062), .B(n7127), .ZN(n7128) );
  NAND2_X1 U8798 ( .A1(n7128), .A2(n8971), .ZN(n7130) );
  AOI22_X1 U8799 ( .A1(n8966), .A2(n8723), .B1(n8721), .B2(n8968), .ZN(n7129)
         );
  NAND2_X1 U8800 ( .A1(n7130), .A2(n7129), .ZN(n10056) );
  INV_X1 U8801 ( .A(n10056), .ZN(n7140) );
  INV_X1 U8802 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10350) );
  OAI22_X1 U8803 ( .A1(n8877), .A2(n10350), .B1(n7131), .B2(n8907), .ZN(n7135)
         );
  INV_X1 U8804 ( .A(n8984), .ZN(n7880) );
  NAND2_X1 U8805 ( .A1(n7269), .A2(n7136), .ZN(n7132) );
  NAND2_X1 U8806 ( .A1(n7133), .A2(n7132), .ZN(n10053) );
  NOR2_X1 U8807 ( .A1(n7880), .A2(n10053), .ZN(n7134) );
  AOI211_X1 U8808 ( .C1(n7963), .C2(n7136), .A(n7135), .B(n7134), .ZN(n7139)
         );
  XNOR2_X1 U8809 ( .A(n8591), .B(n7137), .ZN(n10051) );
  NAND2_X1 U8810 ( .A1(n10051), .A2(n8906), .ZN(n7138) );
  OAI211_X1 U8811 ( .C1(n4476), .C2(n7140), .A(n7139), .B(n7138), .ZN(P2_U3292) );
  XNOR2_X1 U8812 ( .A(n8588), .B(n7141), .ZN(n10041) );
  INV_X1 U8813 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7142) );
  NOR2_X1 U8814 ( .A1(n8877), .A2(n7142), .ZN(n7151) );
  NAND2_X1 U8815 ( .A1(n7143), .A2(n8588), .ZN(n7144) );
  NAND2_X1 U8816 ( .A1(n7145), .A2(n7144), .ZN(n7146) );
  NAND2_X1 U8817 ( .A1(n7146), .A2(n8971), .ZN(n7148) );
  AOI22_X1 U8818 ( .A1(n8966), .A2(n4480), .B1(n8723), .B2(n8968), .ZN(n7147)
         );
  AND2_X1 U8819 ( .A1(n7148), .A2(n7147), .ZN(n10044) );
  OAI22_X1 U8820 ( .A1(n10044), .A2(n4476), .B1(n7149), .B2(n8907), .ZN(n7150)
         );
  AOI211_X1 U8821 ( .C1(n8906), .C2(n10041), .A(n7151), .B(n7150), .ZN(n7156)
         );
  INV_X1 U8822 ( .A(n10039), .ZN(n7154) );
  NAND2_X1 U8823 ( .A1(n7153), .A2(n7152), .ZN(n10036) );
  NAND3_X1 U8824 ( .A1(n8984), .A2(n7154), .A3(n10036), .ZN(n7155) );
  OAI211_X1 U8825 ( .C1(n10037), .C2(n8977), .A(n7156), .B(n7155), .ZN(
        P2_U3294) );
  INV_X1 U8826 ( .A(n10026), .ZN(n8632) );
  NAND2_X1 U8827 ( .A1(n7157), .A2(n8632), .ZN(n8633) );
  NAND2_X1 U8828 ( .A1(n8635), .A2(n8633), .ZN(n10028) );
  INV_X1 U8829 ( .A(n10028), .ZN(n7162) );
  AOI22_X1 U8830 ( .A1(n10028), .A2(n8971), .B1(n8968), .B2(n4480), .ZN(n10030) );
  OAI22_X1 U8831 ( .A1(n4476), .A2(n10030), .B1(n7158), .B2(n8907), .ZN(n7159)
         );
  AOI21_X1 U8832 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n4476), .A(n7159), .ZN(
        n7161) );
  OAI21_X1 U8833 ( .B1(n8984), .B2(n7963), .A(n10026), .ZN(n7160) );
  OAI211_X1 U8834 ( .C1(n7162), .C2(n8981), .A(n7161), .B(n7160), .ZN(P2_U3296) );
  NOR2_X1 U8835 ( .A1(n4476), .A2(n6304), .ZN(n8871) );
  NOR2_X1 U8836 ( .A1(n8977), .A2(n7163), .ZN(n7167) );
  INV_X1 U8837 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7165) );
  OAI22_X1 U8838 ( .A1(n8877), .A2(n7165), .B1(n7164), .B2(n8907), .ZN(n7166)
         );
  AOI211_X1 U8839 ( .C1(n7168), .C2(n8871), .A(n7167), .B(n7166), .ZN(n7171)
         );
  OR2_X1 U8840 ( .A1(n7169), .A2(n8981), .ZN(n7170) );
  OAI211_X1 U8841 ( .C1(n7172), .C2(n4476), .A(n7171), .B(n7170), .ZN(P2_U3291) );
  INV_X1 U8842 ( .A(n7173), .ZN(n7177) );
  OAI21_X1 U8843 ( .B1(n7177), .B2(n7175), .A(n7174), .ZN(n7176) );
  OAI211_X1 U8844 ( .C1(n7178), .C2(n7177), .A(n9660), .B(n7176), .ZN(n7185)
         );
  INV_X1 U8845 ( .A(n7427), .ZN(n7398) );
  NOR2_X1 U8846 ( .A1(n7398), .A2(n9976), .ZN(n9974) );
  INV_X1 U8847 ( .A(n7395), .ZN(n7182) );
  AOI21_X1 U8848 ( .B1(n9196), .B2(n9654), .A(n7179), .ZN(n7181) );
  NAND2_X1 U8849 ( .A1(n9655), .A2(n9209), .ZN(n7180) );
  OAI211_X1 U8850 ( .C1(n9665), .C2(n7182), .A(n7181), .B(n7180), .ZN(n7183)
         );
  AOI21_X1 U8851 ( .B1(n9659), .B2(n9974), .A(n7183), .ZN(n7184) );
  NAND2_X1 U8852 ( .A1(n7185), .A2(n7184), .ZN(P1_U3211) );
  INV_X1 U8853 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7207) );
  NAND2_X1 U8854 ( .A1(n7186), .A2(n6933), .ZN(n7187) );
  NAND2_X1 U8855 ( .A1(n7279), .A2(n7187), .ZN(n7308) );
  NAND2_X1 U8856 ( .A1(n7344), .A2(n7315), .ZN(n7195) );
  NAND2_X1 U8857 ( .A1(n5204), .A2(n9939), .ZN(n8071) );
  NAND2_X1 U8858 ( .A1(n7344), .A2(n9939), .ZN(n7340) );
  INV_X1 U8859 ( .A(n9213), .ZN(n7310) );
  NAND2_X1 U8860 ( .A1(n7310), .A2(n9945), .ZN(n7191) );
  AND2_X1 U8861 ( .A1(n7340), .A2(n7191), .ZN(n7190) );
  NAND2_X1 U8862 ( .A1(n9213), .A2(n9945), .ZN(n8074) );
  INV_X1 U8863 ( .A(n9212), .ZN(n7343) );
  NAND2_X1 U8864 ( .A1(n7343), .A2(n7332), .ZN(n7386) );
  NAND2_X1 U8865 ( .A1(n9212), .A2(n7250), .ZN(n8304) );
  NAND2_X1 U8866 ( .A1(n7386), .A2(n8304), .ZN(n7249) );
  XNOR2_X1 U8867 ( .A(n4563), .B(n7249), .ZN(n7337) );
  AND2_X1 U8868 ( .A1(n7349), .A2(n7332), .ZN(n7193) );
  OR2_X1 U8869 ( .A1(n7193), .A2(n7241), .ZN(n7335) );
  OAI22_X1 U8870 ( .A1(n7335), .A2(n9986), .B1(n7250), .B2(n9976), .ZN(n7205)
         );
  NAND2_X1 U8871 ( .A1(n8069), .A2(n6933), .ZN(n7194) );
  NAND2_X1 U8872 ( .A1(n7196), .A2(n8074), .ZN(n7388) );
  XOR2_X1 U8873 ( .A(n7249), .B(n7388), .Z(n7204) );
  OR2_X1 U8874 ( .A1(n8259), .A2(n9430), .ZN(n7198) );
  OR2_X1 U8875 ( .A1(n5907), .A2(n5153), .ZN(n7197) );
  OR2_X1 U8876 ( .A1(n8262), .A2(n5919), .ZN(n9668) );
  AOI22_X1 U8877 ( .A1(n9705), .A2(n9213), .B1(n9210), .B2(n9702), .ZN(n7203)
         );
  NAND2_X1 U8878 ( .A1(n8259), .A2(n9430), .ZN(n7201) );
  MUX2_X1 U8879 ( .A(n7201), .B(n7200), .S(n7199), .Z(n9674) );
  INV_X1 U8880 ( .A(n9674), .ZN(n9968) );
  NAND2_X1 U8881 ( .A1(n7337), .A2(n9968), .ZN(n7202) );
  OAI211_X1 U8882 ( .C1(n7204), .C2(n9426), .A(n7203), .B(n7202), .ZN(n7330)
         );
  AOI211_X1 U8883 ( .C1(n9950), .C2(n7337), .A(n7205), .B(n7330), .ZN(n7208)
         );
  OR2_X1 U8884 ( .A1(n7208), .A2(n9990), .ZN(n7206) );
  OAI21_X1 U8885 ( .B1(n9992), .B2(n7207), .A(n7206), .ZN(P1_U3466) );
  OR2_X1 U8886 ( .A1(n7208), .A2(n10002), .ZN(n7209) );
  OAI21_X1 U8887 ( .B1(n10004), .B2(n6766), .A(n7209), .ZN(P1_U3527) );
  NAND2_X1 U8888 ( .A1(n7589), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7212) );
  OAI21_X1 U8889 ( .B1(n7589), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7212), .ZN(
        n7213) );
  AOI211_X1 U8890 ( .C1(n7214), .C2(n7213), .A(n7588), .B(n9612), .ZN(n7224)
         );
  INV_X1 U8891 ( .A(n7589), .ZN(n7596) );
  NAND2_X1 U8892 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7362) );
  INV_X1 U8893 ( .A(n7362), .ZN(n7215) );
  AOI21_X1 U8894 ( .B1(n10013), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7215), .ZN(
        n7222) );
  OAI21_X1 U8895 ( .B1(n7217), .B2(n7026), .A(n7216), .ZN(n7220) );
  MUX2_X1 U8896 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7218), .S(n7589), .Z(n7219)
         );
  NAND2_X1 U8897 ( .A1(n7219), .A2(n7220), .ZN(n7595) );
  OAI211_X1 U8898 ( .C1(n7220), .C2(n7219), .A(n10010), .B(n7595), .ZN(n7221)
         );
  OAI211_X1 U8899 ( .C1(n10005), .C2(n7596), .A(n7222), .B(n7221), .ZN(n7223)
         );
  OR2_X1 U8900 ( .A1(n7224), .A2(n7223), .ZN(P2_U3255) );
  XNOR2_X1 U8901 ( .A(n7225), .B(n8594), .ZN(n10061) );
  INV_X1 U8902 ( .A(n10061), .ZN(n7240) );
  XNOR2_X1 U8903 ( .A(n7227), .B(n7226), .ZN(n7228) );
  OAI222_X1 U8904 ( .A1(n8958), .A2(n7407), .B1(n8956), .B2(n7229), .C1(n7228), 
        .C2(n8953), .ZN(n10059) );
  NOR2_X1 U8905 ( .A1(n7230), .A2(n10057), .ZN(n7231) );
  OR2_X1 U8906 ( .A1(n7232), .A2(n7231), .ZN(n10058) );
  OAI22_X1 U8907 ( .A1(n8877), .A2(n7234), .B1(n7233), .B2(n8907), .ZN(n7235)
         );
  AOI21_X1 U8908 ( .B1(n7963), .B2(n7236), .A(n7235), .ZN(n7237) );
  OAI21_X1 U8909 ( .B1(n7880), .B2(n10058), .A(n7237), .ZN(n7238) );
  AOI21_X1 U8910 ( .B1(n10059), .B2(n8877), .A(n7238), .ZN(n7239) );
  OAI21_X1 U8911 ( .B1(n8981), .B2(n7240), .A(n7239), .ZN(P2_U3290) );
  INV_X1 U8912 ( .A(n7241), .ZN(n7243) );
  INV_X1 U8913 ( .A(n7303), .ZN(n7242) );
  AOI211_X1 U8914 ( .C1(n7294), .C2(n7243), .A(n9986), .B(n7242), .ZN(n9954)
         );
  NOR2_X1 U8915 ( .A1(n9693), .A2(n7244), .ZN(n7248) );
  INV_X1 U8916 ( .A(n9209), .ZN(n7382) );
  NAND2_X1 U8917 ( .A1(n7388), .A2(n7386), .ZN(n7245) );
  NAND2_X1 U8918 ( .A1(n7301), .A2(n7294), .ZN(n8307) );
  AND2_X1 U8919 ( .A1(n8307), .A2(n8305), .ZN(n7256) );
  XNOR2_X1 U8920 ( .A(n7299), .B(n7256), .ZN(n7247) );
  OAI222_X1 U8921 ( .A1(n9670), .A2(n7382), .B1(n9668), .B2(n7343), .C1(n9426), 
        .C2(n7247), .ZN(n9956) );
  AOI211_X1 U8922 ( .C1(n9954), .C2(n9430), .A(n7248), .B(n9956), .ZN(n7261)
         );
  AOI22_X1 U8923 ( .A1(n9713), .A2(n7294), .B1(n9709), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n7260) );
  NAND2_X1 U8924 ( .A1(n7343), .A2(n7250), .ZN(n7251) );
  NAND2_X1 U8925 ( .A1(n7252), .A2(n7251), .ZN(n7255) );
  INV_X1 U8926 ( .A(n7255), .ZN(n7254) );
  NAND2_X1 U8927 ( .A1(n7254), .A2(n7253), .ZN(n7296) );
  NAND2_X1 U8928 ( .A1(n7255), .A2(n7256), .ZN(n9952) );
  NAND2_X1 U8929 ( .A1(n8338), .A2(n7257), .ZN(n7258) );
  NAND3_X1 U8930 ( .A1(n7296), .A2(n9952), .A3(n9469), .ZN(n7259) );
  OAI211_X1 U8931 ( .C1(n7261), .C2(n9678), .A(n7260), .B(n7259), .ZN(P1_U3286) );
  INV_X1 U8932 ( .A(n9233), .ZN(n9915) );
  INV_X1 U8933 ( .A(n7262), .ZN(n7264) );
  INV_X1 U8934 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7263) );
  OAI222_X1 U8935 ( .A1(n9915), .A2(P1_U3084), .B1(n9599), .B2(n7264), .C1(
        n7263), .C2(n9595), .ZN(P1_U3335) );
  INV_X1 U8936 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7265) );
  INV_X1 U8937 ( .A(n8774), .ZN(n8788) );
  OAI222_X1 U8938 ( .A1(n8428), .A2(n7265), .B1(n4477), .B2(n7264), .C1(
        P2_U3152), .C2(n8788), .ZN(P2_U3340) );
  XNOR2_X1 U8939 ( .A(n7266), .B(n8467), .ZN(n10045) );
  INV_X1 U8940 ( .A(n7267), .ZN(n7268) );
  NAND2_X1 U8941 ( .A1(n8877), .A2(n7268), .ZN(n7966) );
  OAI21_X1 U8942 ( .B1(n10039), .B2(n6519), .A(n7269), .ZN(n10046) );
  AOI22_X1 U8943 ( .A1(n4476), .A2(P2_REG2_REG_3__SCAN_IN), .B1(n8974), .B2(
        n6039), .ZN(n7270) );
  OAI21_X1 U8944 ( .B1(n7880), .B2(n10046), .A(n7270), .ZN(n7271) );
  XNOR2_X1 U8945 ( .A(n7272), .B(n8467), .ZN(n7275) );
  OAI22_X1 U8946 ( .A1(n7273), .A2(n8956), .B1(n4670), .B2(n8958), .ZN(n7274)
         );
  AOI21_X1 U8947 ( .B1(n7275), .B2(n8971), .A(n7274), .ZN(n7276) );
  OAI21_X1 U8948 ( .B1(n10045), .B2(n7961), .A(n7276), .ZN(n10047) );
  NAND2_X1 U8949 ( .A1(n10047), .A2(n8877), .ZN(n7277) );
  OAI211_X1 U8950 ( .C1(n10045), .C2(n7966), .A(n7278), .B(n7277), .ZN(
        P2_U3293) );
  NAND2_X1 U8951 ( .A1(n7281), .A2(n8139), .ZN(n7282) );
  NOR2_X1 U8952 ( .A1(n9678), .A2(n7282), .ZN(n9692) );
  INV_X1 U8953 ( .A(n9692), .ZN(n7721) );
  AOI22_X1 U8954 ( .A1(n9705), .A2(n6854), .B1(n5204), .B2(n9702), .ZN(n7288)
         );
  OAI21_X1 U8955 ( .B1(n7283), .B2(n7285), .A(n7284), .ZN(n7286) );
  NAND2_X1 U8956 ( .A1(n7286), .A2(n9700), .ZN(n7287) );
  OAI211_X1 U8957 ( .C1(n9932), .C2(n9674), .A(n7288), .B(n7287), .ZN(n9935)
         );
  INV_X1 U8958 ( .A(n7314), .ZN(n7289) );
  OAI211_X1 U8959 ( .C1(n9934), .C2(n8067), .A(n7289), .B(n9960), .ZN(n9933)
         );
  INV_X1 U8960 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7290) );
  OAI22_X1 U8961 ( .A1(n9933), .A2(n8139), .B1(n9693), .B2(n7290), .ZN(n7291)
         );
  OAI21_X1 U8962 ( .B1(n9935), .B2(n7291), .A(n9478), .ZN(n7293) );
  AOI22_X1 U8963 ( .A1(n9713), .A2(n6933), .B1(n9709), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7292) );
  OAI211_X1 U8964 ( .C1(n9932), .C2(n7721), .A(n7293), .B(n7292), .ZN(P1_U3290) );
  NAND2_X1 U8965 ( .A1(n9210), .A2(n7294), .ZN(n7295) );
  NAND2_X1 U8966 ( .A1(n7382), .A2(n9958), .ZN(n8308) );
  INV_X1 U8967 ( .A(n9958), .ZN(n7381) );
  NAND2_X1 U8968 ( .A1(n7381), .A2(n9209), .ZN(n8153) );
  NAND2_X1 U8969 ( .A1(n8308), .A2(n8153), .ZN(n8143) );
  OAI21_X1 U8970 ( .B1(n7297), .B2(n8143), .A(n7384), .ZN(n9967) );
  INV_X1 U8971 ( .A(n9967), .ZN(n9964) );
  INV_X1 U8972 ( .A(n9208), .ZN(n7438) );
  INV_X1 U8973 ( .A(n8305), .ZN(n7298) );
  XNOR2_X1 U8974 ( .A(n8146), .B(n8143), .ZN(n7300) );
  OAI222_X1 U8975 ( .A1(n9670), .A2(n7438), .B1(n9668), .B2(n7301), .C1(n7300), 
        .C2(n9426), .ZN(n9966) );
  NAND2_X1 U8976 ( .A1(n9966), .A2(n9478), .ZN(n7307) );
  OR2_X1 U8977 ( .A1(n7303), .A2(n9958), .ZN(n7392) );
  INV_X1 U8978 ( .A(n7392), .ZN(n7302) );
  AOI21_X1 U8979 ( .B1(n9958), .B2(n7303), .A(n7302), .ZN(n9961) );
  INV_X1 U8980 ( .A(n9693), .ZN(n9679) );
  AOI22_X1 U8981 ( .A1(n9678), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7368), .B2(
        n9679), .ZN(n7304) );
  OAI21_X1 U8982 ( .B1(n9475), .B2(n7381), .A(n7304), .ZN(n7305) );
  AOI21_X1 U8983 ( .B1(n9961), .B2(n9691), .A(n7305), .ZN(n7306) );
  OAI211_X1 U8984 ( .C1(n9415), .C2(n9964), .A(n7307), .B(n7306), .ZN(P1_U3285) );
  XOR2_X1 U8985 ( .A(n8273), .B(n8073), .Z(n7313) );
  NAND2_X1 U8986 ( .A1(n7308), .A2(n8273), .ZN(n7309) );
  NAND2_X1 U8987 ( .A1(n7341), .A2(n7309), .ZN(n9943) );
  OAI22_X1 U8988 ( .A1(n8069), .A2(n9668), .B1(n7310), .B2(n9670), .ZN(n7311)
         );
  AOI21_X1 U8989 ( .B1(n9943), .B2(n9968), .A(n7311), .ZN(n7312) );
  OAI21_X1 U8990 ( .B1(n7313), .B2(n9426), .A(n7312), .ZN(n9941) );
  INV_X1 U8991 ( .A(n9941), .ZN(n7320) );
  OAI21_X1 U8992 ( .B1(n9939), .B2(n7314), .A(n4776), .ZN(n9940) );
  AOI22_X1 U8993 ( .A1(n9709), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9679), .ZN(n7317) );
  NAND2_X1 U8994 ( .A1(n9713), .A2(n7315), .ZN(n7316) );
  OAI211_X1 U8995 ( .C1(n9266), .C2(n9940), .A(n7317), .B(n7316), .ZN(n7318)
         );
  AOI21_X1 U8996 ( .B1(n9692), .B2(n9943), .A(n7318), .ZN(n7319) );
  OAI21_X1 U8997 ( .B1(n9709), .B2(n7320), .A(n7319), .ZN(P1_U3289) );
  INV_X1 U8998 ( .A(n7322), .ZN(n7323) );
  AOI21_X1 U8999 ( .B1(n7321), .B2(n7324), .A(n7323), .ZN(n7329) );
  OAI21_X1 U9000 ( .B1(n8698), .B2(n7480), .A(n7325), .ZN(n7328) );
  OAI22_X1 U9001 ( .A1(n7326), .A2(n8686), .B1(n8687), .B2(n7517), .ZN(n7327)
         );
  OAI21_X1 U9002 ( .B1(n7329), .B2(n8701), .A(n4497), .ZN(P2_U3233) );
  INV_X1 U9003 ( .A(n7330), .ZN(n7339) );
  AOI22_X1 U9004 ( .A1(n9709), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7331), .B2(
        n9679), .ZN(n7334) );
  NAND2_X1 U9005 ( .A1(n9713), .A2(n7332), .ZN(n7333) );
  OAI211_X1 U9006 ( .C1(n9266), .C2(n7335), .A(n7334), .B(n7333), .ZN(n7336)
         );
  AOI21_X1 U9007 ( .B1(n7337), .B2(n9692), .A(n7336), .ZN(n7338) );
  OAI21_X1 U9008 ( .B1(n7339), .B2(n9678), .A(n7338), .ZN(P1_U3287) );
  NAND2_X1 U9009 ( .A1(n7341), .A2(n7340), .ZN(n7342) );
  XNOR2_X1 U9010 ( .A(n7342), .B(n4486), .ZN(n7348) );
  XNOR2_X1 U9011 ( .A(n8301), .B(n4486), .ZN(n7346) );
  OAI22_X1 U9012 ( .A1(n7344), .A2(n9668), .B1(n7343), .B2(n9670), .ZN(n7345)
         );
  AOI21_X1 U9013 ( .B1(n7346), .B2(n9700), .A(n7345), .ZN(n7347) );
  OAI21_X1 U9014 ( .B1(n7348), .B2(n9674), .A(n7347), .ZN(n9947) );
  INV_X1 U9015 ( .A(n9947), .ZN(n7356) );
  INV_X1 U9016 ( .A(n7348), .ZN(n9949) );
  OAI21_X1 U9017 ( .B1(n7350), .B2(n9945), .A(n7349), .ZN(n9946) );
  AOI22_X1 U9018 ( .A1(n9709), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9679), .B2(
        n6925), .ZN(n7353) );
  NAND2_X1 U9019 ( .A1(n9713), .A2(n7351), .ZN(n7352) );
  OAI211_X1 U9020 ( .C1(n9266), .C2(n9946), .A(n7353), .B(n7352), .ZN(n7354)
         );
  AOI21_X1 U9021 ( .B1(n9949), .B2(n9692), .A(n7354), .ZN(n7355) );
  OAI21_X1 U9022 ( .B1(n7356), .B2(n9678), .A(n7355), .ZN(P1_U3288) );
  INV_X1 U9023 ( .A(n7357), .ZN(n8426) );
  OAI222_X1 U9024 ( .A1(P1_U3084), .A2(n9430), .B1(n9599), .B2(n8426), .C1(
        n7358), .C2(n9595), .ZN(P1_U3334) );
  XNOR2_X1 U9025 ( .A(n7360), .B(n7359), .ZN(n7367) );
  INV_X1 U9026 ( .A(n7459), .ZN(n7361) );
  NAND2_X1 U9027 ( .A1(n9631), .A2(n7361), .ZN(n7363) );
  NAND2_X1 U9028 ( .A1(n7363), .A2(n7362), .ZN(n7365) );
  OAI22_X1 U9029 ( .A1(n7406), .A2(n8686), .B1(n8687), .B2(n7611), .ZN(n7364)
         );
  AOI211_X1 U9030 ( .C1(n7462), .C2(n6494), .A(n7365), .B(n7364), .ZN(n7366)
         );
  OAI21_X1 U9031 ( .B1(n7367), .B2(n8701), .A(n7366), .ZN(P2_U3219) );
  INV_X1 U9032 ( .A(n7368), .ZN(n7371) );
  AND2_X1 U9033 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9783) );
  AOI21_X1 U9034 ( .B1(n9655), .B2(n9210), .A(n9783), .ZN(n7370) );
  NAND2_X1 U9035 ( .A1(n9196), .A2(n9208), .ZN(n7369) );
  OAI211_X1 U9036 ( .C1(n9665), .C2(n7371), .A(n7370), .B(n7369), .ZN(n7379)
         );
  INV_X1 U9037 ( .A(n7372), .ZN(n7373) );
  OR3_X1 U9038 ( .A1(n7375), .A2(n7374), .A3(n7373), .ZN(n7377) );
  AOI21_X1 U9039 ( .B1(n7377), .B2(n7376), .A(n9186), .ZN(n7378) );
  AOI211_X1 U9040 ( .C1(n9170), .C2(n9958), .A(n7379), .B(n7378), .ZN(n7380)
         );
  INV_X1 U9041 ( .A(n7380), .ZN(P1_U3237) );
  NAND2_X1 U9042 ( .A1(n7382), .A2(n7381), .ZN(n7383) );
  OR2_X1 U9043 ( .A1(n7438), .A2(n7427), .ZN(n8154) );
  NAND2_X1 U9044 ( .A1(n7427), .A2(n7438), .ZN(n8147) );
  NAND2_X1 U9045 ( .A1(n8154), .A2(n8147), .ZN(n8277) );
  INV_X1 U9046 ( .A(n8277), .ZN(n7433) );
  XNOR2_X1 U9047 ( .A(n7426), .B(n7433), .ZN(n9971) );
  NAND2_X1 U9048 ( .A1(n8153), .A2(n8305), .ZN(n7385) );
  NAND2_X1 U9049 ( .A1(n7385), .A2(n8308), .ZN(n7387) );
  NAND2_X1 U9050 ( .A1(n7387), .A2(n8304), .ZN(n8275) );
  NAND3_X1 U9051 ( .A1(n8308), .A2(n8307), .A3(n7386), .ZN(n8312) );
  NAND2_X1 U9052 ( .A1(n8312), .A2(n7387), .ZN(n8066) );
  XNOR2_X1 U9053 ( .A(n7434), .B(n7433), .ZN(n7389) );
  NAND2_X1 U9054 ( .A1(n7389), .A2(n9700), .ZN(n7391) );
  AOI22_X1 U9055 ( .A1(n9705), .A2(n9209), .B1(n9654), .B2(n9702), .ZN(n7390)
         );
  NAND2_X1 U9056 ( .A1(n7391), .A2(n7390), .ZN(n9972) );
  INV_X1 U9057 ( .A(n7439), .ZN(n7441) );
  AOI211_X1 U9058 ( .C1(n7427), .C2(n7392), .A(n9986), .B(n7441), .ZN(n9973)
         );
  NOR2_X1 U9059 ( .A1(n9928), .A2(n8139), .ZN(n7393) );
  AND2_X1 U9060 ( .A1(n7394), .A2(n7393), .ZN(n7941) );
  NAND2_X1 U9061 ( .A1(n9973), .A2(n7941), .ZN(n7397) );
  AOI22_X1 U9062 ( .A1(n9678), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7395), .B2(
        n9679), .ZN(n7396) );
  OAI211_X1 U9063 ( .C1(n7398), .C2(n9475), .A(n7397), .B(n7396), .ZN(n7399)
         );
  AOI21_X1 U9064 ( .B1(n9478), .B2(n9972), .A(n7399), .ZN(n7400) );
  OAI21_X1 U9065 ( .B1(n9971), .B2(n9415), .A(n7400), .ZN(P1_U3284) );
  OR2_X1 U9066 ( .A1(n7401), .A2(n8596), .ZN(n7469) );
  NAND2_X1 U9067 ( .A1(n7401), .A2(n8596), .ZN(n7402) );
  NAND2_X1 U9068 ( .A1(n7469), .A2(n7402), .ZN(n10063) );
  OR2_X1 U9069 ( .A1(n7404), .A2(n7403), .ZN(n7472) );
  OAI21_X1 U9070 ( .B1(n7405), .B2(n8596), .A(n7472), .ZN(n7409) );
  OAI22_X1 U9071 ( .A1(n7407), .A2(n8956), .B1(n7406), .B2(n8958), .ZN(n7408)
         );
  AOI21_X1 U9072 ( .B1(n7409), .B2(n8971), .A(n7408), .ZN(n7410) );
  OAI21_X1 U9073 ( .B1(n10063), .B2(n7961), .A(n7410), .ZN(n10067) );
  NAND2_X1 U9074 ( .A1(n10067), .A2(n8877), .ZN(n7417) );
  OAI22_X1 U9075 ( .A1(n8877), .A2(n6951), .B1(n7411), .B2(n8907), .ZN(n7415)
         );
  NAND2_X1 U9076 ( .A1(n7412), .A2(n10064), .ZN(n7413) );
  NAND2_X1 U9077 ( .A1(n7478), .A2(n7413), .ZN(n10066) );
  NOR2_X1 U9078 ( .A1(n10066), .A2(n7880), .ZN(n7414) );
  AOI211_X1 U9079 ( .C1(n7963), .C2(n10064), .A(n7415), .B(n7414), .ZN(n7416)
         );
  OAI211_X1 U9080 ( .C1(n10063), .C2(n7966), .A(n7417), .B(n7416), .ZN(
        P2_U3288) );
  AOI211_X1 U9081 ( .C1(n9058), .C2(n7420), .A(n7419), .B(n7418), .ZN(n7421)
         );
  OAI21_X1 U9082 ( .B1(n9054), .B2(n7422), .A(n7421), .ZN(n7424) );
  NAND2_X1 U9083 ( .A1(n7424), .A2(n10098), .ZN(n7423) );
  OAI21_X1 U9084 ( .B1(n10098), .B2(n6847), .A(n7423), .ZN(P2_U3527) );
  NAND2_X1 U9085 ( .A1(n7424), .A2(n10086), .ZN(n7425) );
  OAI21_X1 U9086 ( .B1(n10086), .B2(n6104), .A(n7425), .ZN(P2_U3472) );
  INV_X1 U9087 ( .A(n9654), .ZN(n8160) );
  OR2_X1 U9088 ( .A1(n8165), .A2(n8160), .ZN(n8149) );
  NAND2_X1 U9089 ( .A1(n8165), .A2(n8160), .ZN(n8086) );
  AND2_X1 U9090 ( .A1(n8149), .A2(n8086), .ZN(n7436) );
  OR2_X1 U9091 ( .A1(n9208), .A2(n7427), .ZN(n7428) );
  NAND2_X1 U9092 ( .A1(n7429), .A2(n7428), .ZN(n7430) );
  INV_X1 U9093 ( .A(n7523), .ZN(n7432) );
  AOI21_X1 U9094 ( .B1(n7436), .B2(n7430), .A(n7432), .ZN(n9981) );
  INV_X1 U9095 ( .A(n9981), .ZN(n7448) );
  INV_X1 U9096 ( .A(n9207), .ZN(n8159) );
  XNOR2_X1 U9097 ( .A(n7526), .B(n7431), .ZN(n7437) );
  OAI222_X1 U9098 ( .A1(n9670), .A2(n8159), .B1(n9668), .B2(n7438), .C1(n7437), 
        .C2(n9426), .ZN(n9980) );
  INV_X1 U9099 ( .A(n8165), .ZN(n9977) );
  INV_X1 U9100 ( .A(n7555), .ZN(n7440) );
  OAI21_X1 U9101 ( .B1(n9977), .B2(n7441), .A(n7440), .ZN(n9978) );
  INV_X1 U9102 ( .A(n7442), .ZN(n7510) );
  OAI22_X1 U9103 ( .A1(n9478), .A2(n7443), .B1(n7510), .B2(n9693), .ZN(n7444)
         );
  AOI21_X1 U9104 ( .B1(n9713), .B2(n8165), .A(n7444), .ZN(n7445) );
  OAI21_X1 U9105 ( .B1(n9978), .B2(n9266), .A(n7445), .ZN(n7446) );
  AOI21_X1 U9106 ( .B1(n9980), .B2(n9478), .A(n7446), .ZN(n7447) );
  OAI21_X1 U9107 ( .B1(n7448), .B2(n9415), .A(n7447), .ZN(P1_U3283) );
  XNOR2_X1 U9108 ( .A(n7449), .B(n7457), .ZN(n7450) );
  NAND2_X1 U9109 ( .A1(n7450), .A2(n8971), .ZN(n7452) );
  AOI22_X1 U9110 ( .A1(n8966), .A2(n8717), .B1(n8715), .B2(n8968), .ZN(n7451)
         );
  NAND2_X1 U9111 ( .A1(n7452), .A2(n7451), .ZN(n10074) );
  INV_X1 U9112 ( .A(n10074), .ZN(n7466) );
  AND2_X1 U9113 ( .A1(n7454), .A2(n7453), .ZN(n7456) );
  NOR2_X1 U9114 ( .A1(n7456), .A2(n7457), .ZN(n7455) );
  AOI21_X1 U9115 ( .B1(n7457), .B2(n7456), .A(n7455), .ZN(n10075) );
  NOR2_X1 U9116 ( .A1(n7477), .A2(n10071), .ZN(n7458) );
  OR2_X1 U9117 ( .A1(n7630), .A2(n7458), .ZN(n10072) );
  INV_X1 U9118 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7460) );
  OAI22_X1 U9119 ( .A1(n8877), .A2(n7460), .B1(n7459), .B2(n8907), .ZN(n7461)
         );
  AOI21_X1 U9120 ( .B1(n7462), .B2(n7963), .A(n7461), .ZN(n7463) );
  OAI21_X1 U9121 ( .B1(n10072), .B2(n7880), .A(n7463), .ZN(n7464) );
  AOI21_X1 U9122 ( .B1(n10075), .B2(n8906), .A(n7464), .ZN(n7465) );
  OAI21_X1 U9123 ( .B1(n4476), .B2(n7466), .A(n7465), .ZN(P2_U3286) );
  AND2_X1 U9124 ( .A1(n7469), .A2(n7467), .ZN(n7471) );
  NAND2_X1 U9125 ( .A1(n7469), .A2(n7468), .ZN(n7470) );
  OAI21_X1 U9126 ( .B1(n7471), .B2(n8598), .A(n7470), .ZN(n7560) );
  INV_X1 U9127 ( .A(n7961), .ZN(n7655) );
  NAND2_X1 U9128 ( .A1(n7472), .A2(n8490), .ZN(n7473) );
  XNOR2_X1 U9129 ( .A(n8598), .B(n7473), .ZN(n7475) );
  AOI22_X1 U9130 ( .A1(n8966), .A2(n8718), .B1(n8716), .B2(n8968), .ZN(n7474)
         );
  OAI21_X1 U9131 ( .B1(n7475), .B2(n8953), .A(n7474), .ZN(n7476) );
  AOI21_X1 U9132 ( .B1(n7560), .B2(n7655), .A(n7476), .ZN(n7563) );
  NOR2_X1 U9133 ( .A1(n7479), .A2(n8977), .ZN(n7483) );
  OAI22_X1 U9134 ( .A1(n8877), .A2(n7481), .B1(n7480), .B2(n8907), .ZN(n7482)
         );
  AOI211_X1 U9135 ( .C1(n7561), .C2(n8984), .A(n7483), .B(n7482), .ZN(n7485)
         );
  INV_X1 U9136 ( .A(n7966), .ZN(n7661) );
  NAND2_X1 U9137 ( .A1(n7560), .A2(n7661), .ZN(n7484) );
  OAI211_X1 U9138 ( .C1(n7563), .C2(n4476), .A(n7485), .B(n7484), .ZN(P2_U3287) );
  INV_X1 U9139 ( .A(n7494), .ZN(n9845) );
  OAI21_X1 U9140 ( .B1(n7487), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7486), .ZN(
        n9841) );
  XOR2_X1 U9141 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n7494), .Z(n9842) );
  NOR2_X1 U9142 ( .A1(n9841), .A2(n9842), .ZN(n9840) );
  INV_X1 U9143 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9695) );
  MUX2_X1 U9144 ( .A(n9695), .B(P1_REG2_REG_13__SCAN_IN), .S(n9858), .Z(n9854)
         );
  INV_X1 U9145 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7488) );
  NAND2_X1 U9146 ( .A1(n7489), .A2(n7488), .ZN(n9226) );
  OAI21_X1 U9147 ( .B1(n7489), .B2(n7488), .A(n9226), .ZN(n7502) );
  INV_X1 U9148 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7491) );
  INV_X1 U9149 ( .A(n9238), .ZN(n7496) );
  AND2_X1 U9150 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7903) );
  AOI21_X1 U9151 ( .B1(n9883), .B2(n7496), .A(n7903), .ZN(n7490) );
  OAI21_X1 U9152 ( .B1(n9924), .B2(n7491), .A(n7490), .ZN(n7501) );
  INV_X1 U9153 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10205) );
  INV_X1 U9154 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9735) );
  AOI21_X1 U9155 ( .B1(n9743), .B2(n7493), .A(n7492), .ZN(n9848) );
  MUX2_X1 U9156 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9735), .S(n7494), .Z(n9847)
         );
  NOR2_X1 U9157 ( .A1(n9848), .A2(n9847), .ZN(n9846) );
  AOI21_X1 U9158 ( .B1(n9735), .B2(n7494), .A(n9846), .ZN(n9861) );
  MUX2_X1 U9159 ( .A(n10205), .B(P1_REG1_REG_13__SCAN_IN), .S(n9858), .Z(n9860) );
  NOR2_X1 U9160 ( .A1(n9861), .A2(n9860), .ZN(n9859) );
  AOI21_X1 U9161 ( .B1(n10205), .B2(n7495), .A(n9859), .ZN(n7498) );
  INV_X1 U9162 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U9163 ( .A1(n7496), .A2(n10283), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n9238), .ZN(n7497) );
  NOR2_X1 U9164 ( .A1(n7498), .A2(n7497), .ZN(n9237) );
  AOI21_X1 U9165 ( .B1(n7498), .B2(n7497), .A(n9237), .ZN(n7499) );
  NOR2_X1 U9166 ( .A1(n7499), .A2(n9921), .ZN(n7500) );
  AOI211_X1 U9167 ( .C1(n7502), .C2(n9911), .A(n7501), .B(n7500), .ZN(n7503)
         );
  INV_X1 U9168 ( .A(n7503), .ZN(P1_U3255) );
  AOI21_X1 U9169 ( .B1(n7507), .B2(n7505), .A(n7504), .ZN(n7506) );
  AOI21_X1 U9170 ( .B1(n4559), .B2(n7507), .A(n7506), .ZN(n7513) );
  AND2_X1 U9171 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9802) );
  AOI21_X1 U9172 ( .B1(n9196), .B2(n9207), .A(n9802), .ZN(n7509) );
  NAND2_X1 U9173 ( .A1(n9655), .A2(n9208), .ZN(n7508) );
  OAI211_X1 U9174 ( .C1(n9665), .C2(n7510), .A(n7509), .B(n7508), .ZN(n7511)
         );
  AOI21_X1 U9175 ( .B1(n9170), .B2(n8165), .A(n7511), .ZN(n7512) );
  OAI21_X1 U9176 ( .B1(n7513), .B2(n9186), .A(n7512), .ZN(P1_U3219) );
  INV_X1 U9177 ( .A(n7514), .ZN(n7548) );
  OAI222_X1 U9178 ( .A1(n5153), .A2(P1_U3084), .B1(n9599), .B2(n7548), .C1(
        n7515), .C2(n9595), .ZN(P1_U3333) );
  XNOR2_X1 U9179 ( .A(n4558), .B(n7516), .ZN(n7521) );
  INV_X1 U9180 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8729) );
  OAI22_X1 U9181 ( .A1(n8698), .A2(n7722), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8729), .ZN(n7519) );
  OAI22_X1 U9182 ( .A1(n7517), .A2(n8686), .B1(n8687), .B2(n7670), .ZN(n7518)
         );
  AOI211_X1 U9183 ( .C1(n7632), .C2(n6494), .A(n7519), .B(n7518), .ZN(n7520)
         );
  OAI21_X1 U9184 ( .B1(n7521), .B2(n8701), .A(n7520), .ZN(P2_U3238) );
  NAND2_X1 U9185 ( .A1(n8165), .A2(n9654), .ZN(n7522) );
  OR2_X1 U9186 ( .A1(n8166), .A2(n9207), .ZN(n7524) );
  INV_X1 U9187 ( .A(n9206), .ZN(n9651) );
  NAND2_X1 U9188 ( .A1(n7706), .A2(n9651), .ZN(n8178) );
  NAND2_X1 U9189 ( .A1(n8173), .A2(n8178), .ZN(n8279) );
  NAND2_X1 U9190 ( .A1(n7525), .A2(n8279), .ZN(n7708) );
  OAI21_X1 U9191 ( .B1(n7525), .B2(n8279), .A(n7708), .ZN(n7578) );
  INV_X1 U9192 ( .A(n7578), .ZN(n7537) );
  OR2_X1 U9193 ( .A1(n8166), .A2(n8159), .ZN(n8150) );
  AND2_X1 U9194 ( .A1(n8150), .A2(n8149), .ZN(n8094) );
  NAND2_X1 U9195 ( .A1(n8166), .A2(n8159), .ZN(n8156) );
  INV_X1 U9196 ( .A(n8279), .ZN(n7527) );
  OAI211_X1 U9197 ( .C1(n5040), .C2(n7527), .A(n7709), .B(n9700), .ZN(n7529)
         );
  AOI22_X1 U9198 ( .A1(n9702), .A2(n9205), .B1(n9207), .B2(n9705), .ZN(n7528)
         );
  NAND2_X1 U9199 ( .A1(n7529), .A2(n7528), .ZN(n7576) );
  INV_X1 U9200 ( .A(n7706), .ZN(n7534) );
  INV_X1 U9201 ( .A(n8166), .ZN(n9658) );
  NAND2_X1 U9202 ( .A1(n7555), .A2(n9658), .ZN(n7554) );
  INV_X1 U9203 ( .A(n7715), .ZN(n7530) );
  AOI211_X1 U9204 ( .C1(n7706), .C2(n7554), .A(n9986), .B(n7530), .ZN(n7577)
         );
  NAND2_X1 U9205 ( .A1(n7577), .A2(n7941), .ZN(n7533) );
  AOI22_X1 U9206 ( .A1(n9678), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7531), .B2(
        n9679), .ZN(n7532) );
  OAI211_X1 U9207 ( .C1(n7534), .C2(n9475), .A(n7533), .B(n7532), .ZN(n7535)
         );
  AOI21_X1 U9208 ( .B1(n9478), .B2(n7576), .A(n7535), .ZN(n7536) );
  OAI21_X1 U9209 ( .B1(n7537), .B2(n9415), .A(n7536), .ZN(P1_U3281) );
  XNOR2_X1 U9210 ( .A(n7539), .B(n7538), .ZN(n7540) );
  XNOR2_X1 U9211 ( .A(n7541), .B(n7540), .ZN(n7547) );
  AND2_X1 U9212 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9828) );
  AOI21_X1 U9213 ( .B1(n9655), .B2(n9207), .A(n9828), .ZN(n7543) );
  NAND2_X1 U9214 ( .A1(n9196), .A2(n9205), .ZN(n7542) );
  OAI211_X1 U9215 ( .C1(n9665), .C2(n7544), .A(n7543), .B(n7542), .ZN(n7545)
         );
  AOI21_X1 U9216 ( .B1(n9170), .B2(n7706), .A(n7545), .ZN(n7546) );
  OAI21_X1 U9217 ( .B1(n7547), .B2(n9186), .A(n7546), .ZN(P1_U3215) );
  OAI222_X1 U9218 ( .A1(n9087), .A2(n7549), .B1(P2_U3152), .B2(n8587), .C1(
        n4477), .C2(n7548), .ZN(P2_U3338) );
  NAND2_X1 U9219 ( .A1(n7550), .A2(n8149), .ZN(n7551) );
  NAND2_X1 U9220 ( .A1(n8150), .A2(n8156), .ZN(n8278) );
  XNOR2_X1 U9221 ( .A(n7551), .B(n8278), .ZN(n7552) );
  AOI222_X1 U9222 ( .A1(n9700), .A2(n7552), .B1(n9206), .B2(n9702), .C1(n9654), 
        .C2(n9705), .ZN(n9984) );
  XOR2_X1 U9223 ( .A(n8278), .B(n7553), .Z(n9989) );
  NAND2_X1 U9224 ( .A1(n9989), .A2(n9469), .ZN(n7559) );
  OAI22_X1 U9225 ( .A1(n9478), .A2(n4757), .B1(n9664), .B2(n9693), .ZN(n7557)
         );
  OAI21_X1 U9226 ( .B1(n7555), .B2(n9658), .A(n7554), .ZN(n9985) );
  NOR2_X1 U9227 ( .A1(n9985), .A2(n9266), .ZN(n7556) );
  AOI211_X1 U9228 ( .C1(n9713), .C2(n8166), .A(n7557), .B(n7556), .ZN(n7558)
         );
  OAI211_X1 U9229 ( .C1(n9709), .C2(n9984), .A(n7559), .B(n7558), .ZN(P1_U3282) );
  INV_X1 U9230 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10318) );
  INV_X1 U9231 ( .A(n7560), .ZN(n7564) );
  OAI211_X1 U9232 ( .C1(n7564), .C2(n9063), .A(n7563), .B(n7562), .ZN(n7566)
         );
  NAND2_X1 U9233 ( .A1(n7566), .A2(n10086), .ZN(n7565) );
  OAI21_X1 U9234 ( .B1(n10086), .B2(n10318), .A(n7565), .ZN(P2_U3478) );
  NAND2_X1 U9235 ( .A1(n7566), .A2(n10098), .ZN(n7567) );
  OAI21_X1 U9236 ( .B1(n10098), .B2(n7026), .A(n7567), .ZN(P2_U3529) );
  NAND2_X1 U9237 ( .A1(n7569), .A2(n7568), .ZN(n7570) );
  XNOR2_X1 U9238 ( .A(n7571), .B(n7570), .ZN(n7575) );
  AOI22_X1 U9239 ( .A1(n8047), .A2(n8715), .B1(n8048), .B2(n8713), .ZN(n7572)
         );
  NAND2_X1 U9240 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7601) );
  OAI211_X1 U9241 ( .C1(n7613), .C2(n8698), .A(n7572), .B(n7601), .ZN(n7573)
         );
  AOI21_X1 U9242 ( .B1(n7616), .B2(n6494), .A(n7573), .ZN(n7574) );
  OAI21_X1 U9243 ( .B1(n7575), .B2(n8701), .A(n7574), .ZN(P2_U3226) );
  INV_X1 U9244 ( .A(n9950), .ZN(n9963) );
  AOI211_X1 U9245 ( .C1(n7578), .C2(n9988), .A(n7577), .B(n7576), .ZN(n7585)
         );
  NAND2_X1 U9246 ( .A1(n9992), .A2(n9959), .ZN(n9588) );
  INV_X1 U9247 ( .A(n9588), .ZN(n7581) );
  INV_X1 U9248 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7579) );
  NOR2_X1 U9249 ( .A1(n9992), .A2(n7579), .ZN(n7580) );
  AOI21_X1 U9250 ( .B1(n7706), .B2(n7581), .A(n7580), .ZN(n7582) );
  OAI21_X1 U9251 ( .B1(n7585), .B2(n9990), .A(n7582), .ZN(P1_U3484) );
  NAND2_X1 U9252 ( .A1(n10004), .A2(n9959), .ZN(n9551) );
  INV_X1 U9253 ( .A(n9551), .ZN(n7583) );
  AOI22_X1 U9254 ( .A1(n7706), .A2(n7583), .B1(n10002), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7584) );
  OAI21_X1 U9255 ( .B1(n7585), .B2(n10002), .A(n7584), .ZN(P1_U3533) );
  INV_X1 U9256 ( .A(n7586), .ZN(n8061) );
  OAI222_X1 U9257 ( .A1(n9087), .A2(n7587), .B1(P2_U3152), .B2(n8443), .C1(
        n4477), .C2(n8061), .ZN(P2_U3337) );
  NOR2_X1 U9258 ( .A1(n8731), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7590) );
  AOI21_X1 U9259 ( .B1(n8731), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7590), .ZN(
        n8727) );
  NAND2_X1 U9260 ( .A1(n7769), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7591) );
  OAI21_X1 U9261 ( .B1(n7769), .B2(P2_REG2_REG_12__SCAN_IN), .A(n7591), .ZN(
        n7592) );
  NOR2_X1 U9262 ( .A1(n7592), .A2(n7593), .ZN(n7768) );
  AOI211_X1 U9263 ( .C1(n7593), .C2(n7592), .A(n7768), .B(n9612), .ZN(n7607)
         );
  INV_X1 U9264 ( .A(n10010), .ZN(n8023) );
  NAND2_X1 U9265 ( .A1(n8731), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7597) );
  MUX2_X1 U9266 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7594), .S(n8731), .Z(n8733)
         );
  OAI21_X1 U9267 ( .B1(n7596), .B2(n7218), .A(n7595), .ZN(n8734) );
  NAND2_X1 U9268 ( .A1(n8733), .A2(n8734), .ZN(n8732) );
  NAND2_X1 U9269 ( .A1(n7597), .A2(n8732), .ZN(n7600) );
  MUX2_X1 U9270 ( .A(n7598), .B(P2_REG1_REG_12__SCAN_IN), .S(n7769), .Z(n7599)
         );
  NOR2_X1 U9271 ( .A1(n7600), .A2(n7599), .ZN(n7764) );
  AOI21_X1 U9272 ( .B1(n7600), .B2(n7599), .A(n7764), .ZN(n7605) );
  INV_X1 U9273 ( .A(n7601), .ZN(n7602) );
  AOI21_X1 U9274 ( .B1(n10013), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7602), .ZN(
        n7604) );
  NAND2_X1 U9275 ( .A1(n9618), .A2(n7769), .ZN(n7603) );
  OAI211_X1 U9276 ( .C1(n8023), .C2(n7605), .A(n7604), .B(n7603), .ZN(n7606)
         );
  OR2_X1 U9277 ( .A1(n7607), .A2(n7606), .ZN(P2_U3257) );
  XNOR2_X1 U9278 ( .A(n7608), .B(n8603), .ZN(n10083) );
  INV_X1 U9279 ( .A(n10083), .ZN(n7620) );
  NAND2_X1 U9280 ( .A1(n7626), .A2(n8498), .ZN(n7609) );
  XOR2_X1 U9281 ( .A(n8603), .B(n7609), .Z(n7610) );
  OAI222_X1 U9282 ( .A1(n8958), .A2(n7753), .B1(n8956), .B2(n7611), .C1(n7610), 
        .C2(n8953), .ZN(n10080) );
  INV_X1 U9283 ( .A(n7616), .ZN(n10077) );
  INV_X1 U9284 ( .A(n7612), .ZN(n7657) );
  OAI21_X1 U9285 ( .B1(n4556), .B2(n10077), .A(n7657), .ZN(n10079) );
  OAI22_X1 U9286 ( .A1(n8877), .A2(n7614), .B1(n7613), .B2(n8907), .ZN(n7615)
         );
  AOI21_X1 U9287 ( .B1(n7616), .B2(n7963), .A(n7615), .ZN(n7617) );
  OAI21_X1 U9288 ( .B1(n10079), .B2(n7880), .A(n7617), .ZN(n7618) );
  AOI21_X1 U9289 ( .B1(n10080), .B2(n8877), .A(n7618), .ZN(n7619) );
  OAI21_X1 U9290 ( .B1(n8981), .B2(n7620), .A(n7619), .ZN(P2_U3284) );
  INV_X1 U9291 ( .A(n7621), .ZN(n7624) );
  OAI222_X1 U9292 ( .A1(n9087), .A2(n10341), .B1(n4477), .B2(n7624), .C1(n7622), .C2(P2_U3152), .ZN(P2_U3336) );
  OAI222_X1 U9293 ( .A1(P1_U3084), .A2(n8259), .B1(n9599), .B2(n7624), .C1(
        n7623), .C2(n9595), .ZN(P1_U3331) );
  XNOR2_X1 U9294 ( .A(n7625), .B(n8601), .ZN(n7731) );
  OAI21_X1 U9295 ( .B1(n7628), .B2(n7627), .A(n7626), .ZN(n7629) );
  AOI222_X1 U9296 ( .A1(n8971), .A2(n7629), .B1(n8714), .B2(n8968), .C1(n8716), 
        .C2(n8966), .ZN(n7726) );
  INV_X1 U9297 ( .A(n7630), .ZN(n7631) );
  AOI21_X1 U9298 ( .B1(n7632), .B2(n7631), .A(n4556), .ZN(n7729) );
  AOI22_X1 U9299 ( .A1(n7729), .A2(n10035), .B1(n9058), .B2(n7632), .ZN(n7633)
         );
  OAI211_X1 U9300 ( .C1(n9054), .C2(n7731), .A(n7726), .B(n7633), .ZN(n7635)
         );
  NAND2_X1 U9301 ( .A1(n7635), .A2(n10098), .ZN(n7634) );
  OAI21_X1 U9302 ( .B1(n10098), .B2(n7594), .A(n7634), .ZN(P2_U3531) );
  NAND2_X1 U9303 ( .A1(n7635), .A2(n10086), .ZN(n7636) );
  OAI21_X1 U9304 ( .B1(n10086), .B2(n6172), .A(n7636), .ZN(P2_U3484) );
  XNOR2_X1 U9305 ( .A(n7637), .B(n7638), .ZN(n7645) );
  INV_X1 U9306 ( .A(n7639), .ZN(n7713) );
  INV_X1 U9307 ( .A(n9704), .ZN(n7799) );
  NOR2_X1 U9308 ( .A1(n9652), .A2(n7799), .ZN(n7640) );
  AOI211_X1 U9309 ( .C1(n9655), .C2(n9206), .A(n7641), .B(n7640), .ZN(n7642)
         );
  OAI21_X1 U9310 ( .B1(n9665), .B2(n7713), .A(n7642), .ZN(n7643) );
  AOI21_X1 U9311 ( .B1(n9170), .B2(n9737), .A(n7643), .ZN(n7644) );
  OAI21_X1 U9312 ( .B1(n7645), .B2(n9186), .A(n7644), .ZN(P1_U3234) );
  NAND2_X1 U9313 ( .A1(n7646), .A2(n6564), .ZN(n7647) );
  NAND2_X1 U9314 ( .A1(n7649), .A2(n7650), .ZN(n7651) );
  AOI21_X1 U9315 ( .B1(n7652), .B2(n7651), .A(n8953), .ZN(n7654) );
  OAI22_X1 U9316 ( .A1(n7807), .A2(n8958), .B1(n7670), .B2(n8956), .ZN(n7653)
         );
  AOI211_X1 U9317 ( .C1(n9056), .C2(n7655), .A(n7654), .B(n7653), .ZN(n9061)
         );
  INV_X1 U9318 ( .A(n7656), .ZN(n7756) );
  AOI21_X1 U9319 ( .B1(n9057), .B2(n7657), .A(n7756), .ZN(n9059) );
  INV_X1 U9320 ( .A(n9057), .ZN(n7675) );
  NOR2_X1 U9321 ( .A1(n7675), .A2(n8977), .ZN(n7660) );
  OAI22_X1 U9322 ( .A1(n8877), .A2(n7658), .B1(n7668), .B2(n8907), .ZN(n7659)
         );
  AOI211_X1 U9323 ( .C1(n9059), .C2(n8984), .A(n7660), .B(n7659), .ZN(n7663)
         );
  NAND2_X1 U9324 ( .A1(n9056), .A2(n7661), .ZN(n7662) );
  OAI211_X1 U9325 ( .C1(n9061), .C2(n4476), .A(n7663), .B(n7662), .ZN(P2_U3283) );
  AOI21_X1 U9326 ( .B1(n7664), .B2(n7665), .A(n8701), .ZN(n7667) );
  NAND2_X1 U9327 ( .A1(n7667), .A2(n7666), .ZN(n7674) );
  INV_X1 U9328 ( .A(n7668), .ZN(n7672) );
  NOR2_X1 U9329 ( .A1(n7669), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7774) );
  OAI22_X1 U9330 ( .A1(n7670), .A2(n8686), .B1(n8687), .B2(n7807), .ZN(n7671)
         );
  AOI211_X1 U9331 ( .C1(n9631), .C2(n7672), .A(n7774), .B(n7671), .ZN(n7673)
         );
  OAI211_X1 U9332 ( .C1(n7675), .C2(n8692), .A(n7674), .B(n7673), .ZN(P2_U3236) );
  INV_X1 U9333 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10510) );
  NOR2_X1 U9334 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7676) );
  AOI21_X1 U9335 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7676), .ZN(n10106) );
  NOR2_X1 U9336 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7677) );
  AOI21_X1 U9337 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7677), .ZN(n10109) );
  NOR2_X1 U9338 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7678) );
  AOI21_X1 U9339 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7678), .ZN(n10112) );
  NOR2_X1 U9340 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7679) );
  AOI21_X1 U9341 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7679), .ZN(n10115) );
  NOR2_X1 U9342 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7680) );
  AOI21_X1 U9343 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7680), .ZN(n10118) );
  NOR2_X1 U9344 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7686) );
  XOR2_X1 U9345 ( .A(n10365), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10521) );
  NAND2_X1 U9346 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7684) );
  XNOR2_X1 U9347 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n10347), .ZN(n10519) );
  NAND2_X1 U9348 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7682) );
  XOR2_X1 U9349 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10504) );
  AOI21_X1 U9350 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10099) );
  INV_X1 U9351 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10103) );
  NAND3_X1 U9352 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10101) );
  OAI21_X1 U9353 ( .B1(n10099), .B2(n10103), .A(n10101), .ZN(n10503) );
  NAND2_X1 U9354 ( .A1(n10504), .A2(n10503), .ZN(n7681) );
  NAND2_X1 U9355 ( .A1(n7682), .A2(n7681), .ZN(n10518) );
  NAND2_X1 U9356 ( .A1(n10519), .A2(n10518), .ZN(n7683) );
  NAND2_X1 U9357 ( .A1(n7684), .A2(n7683), .ZN(n10520) );
  NOR2_X1 U9358 ( .A1(n10521), .A2(n10520), .ZN(n7685) );
  NOR2_X1 U9359 ( .A1(n7686), .A2(n7685), .ZN(n7687) );
  NOR2_X1 U9360 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7687), .ZN(n10505) );
  AND2_X1 U9361 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7687), .ZN(n10506) );
  NOR2_X1 U9362 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10506), .ZN(n7688) );
  NOR2_X1 U9363 ( .A1(n10505), .A2(n7688), .ZN(n7689) );
  NAND2_X1 U9364 ( .A1(n7689), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7691) );
  INV_X1 U9365 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9794) );
  XNOR2_X1 U9366 ( .A(n7689), .B(n9794), .ZN(n10502) );
  NAND2_X1 U9367 ( .A1(n10502), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7690) );
  NAND2_X1 U9368 ( .A1(n7691), .A2(n7690), .ZN(n7692) );
  NAND2_X1 U9369 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7692), .ZN(n7694) );
  XNOR2_X1 U9370 ( .A(n6795), .B(n7692), .ZN(n10516) );
  NAND2_X1 U9371 ( .A1(n10516), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7693) );
  NAND2_X1 U9372 ( .A1(n7694), .A2(n7693), .ZN(n7695) );
  NAND2_X1 U9373 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7695), .ZN(n7697) );
  INV_X1 U9374 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9809) );
  XNOR2_X1 U9375 ( .A(n9809), .B(n7695), .ZN(n10517) );
  NAND2_X1 U9376 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10517), .ZN(n7696) );
  NAND2_X1 U9377 ( .A1(n7697), .A2(n7696), .ZN(n7698) );
  AND2_X1 U9378 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7698), .ZN(n7699) );
  INV_X1 U9379 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10515) );
  XNOR2_X1 U9380 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7698), .ZN(n10514) );
  NOR2_X1 U9381 ( .A1(n10515), .A2(n10514), .ZN(n10513) );
  NOR2_X1 U9382 ( .A1(n7699), .A2(n10513), .ZN(n10127) );
  NAND2_X1 U9383 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7700) );
  OAI21_X1 U9384 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7700), .ZN(n10126) );
  NOR2_X1 U9385 ( .A1(n10127), .A2(n10126), .ZN(n10125) );
  AOI21_X1 U9386 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10125), .ZN(n10124) );
  NAND2_X1 U9387 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7701) );
  OAI21_X1 U9388 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7701), .ZN(n10123) );
  NOR2_X1 U9389 ( .A1(n10124), .A2(n10123), .ZN(n10122) );
  AOI21_X1 U9390 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10122), .ZN(n10121) );
  NOR2_X1 U9391 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7702) );
  AOI21_X1 U9392 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7702), .ZN(n10120) );
  NAND2_X1 U9393 ( .A1(n10121), .A2(n10120), .ZN(n10119) );
  OAI21_X1 U9394 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10119), .ZN(n10117) );
  NAND2_X1 U9395 ( .A1(n10118), .A2(n10117), .ZN(n10116) );
  OAI21_X1 U9396 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10116), .ZN(n10114) );
  NAND2_X1 U9397 ( .A1(n10115), .A2(n10114), .ZN(n10113) );
  OAI21_X1 U9398 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10113), .ZN(n10111) );
  NAND2_X1 U9399 ( .A1(n10112), .A2(n10111), .ZN(n10110) );
  OAI21_X1 U9400 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10110), .ZN(n10108) );
  NAND2_X1 U9401 ( .A1(n10109), .A2(n10108), .ZN(n10107) );
  OAI21_X1 U9402 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10107), .ZN(n10105) );
  NAND2_X1 U9403 ( .A1(n10106), .A2(n10105), .ZN(n10104) );
  OAI21_X1 U9404 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10104), .ZN(n10509) );
  NOR2_X1 U9405 ( .A1(n10510), .A2(n10509), .ZN(n7703) );
  NAND2_X1 U9406 ( .A1(n10510), .A2(n10509), .ZN(n10508) );
  OAI21_X1 U9407 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7703), .A(n10508), .ZN(
        n7705) );
  XNOR2_X1 U9408 ( .A(n4597), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7704) );
  XNOR2_X1 U9409 ( .A(n7705), .B(n7704), .ZN(ADD_1071_U4) );
  OR2_X1 U9410 ( .A1(n7706), .A2(n9206), .ZN(n7707) );
  NAND2_X1 U9411 ( .A1(n7708), .A2(n7707), .ZN(n7735) );
  INV_X1 U9412 ( .A(n9205), .ZN(n7789) );
  OR2_X1 U9413 ( .A1(n9737), .A2(n7789), .ZN(n7856) );
  NAND2_X1 U9414 ( .A1(n9737), .A2(n7789), .ZN(n8083) );
  XNOR2_X1 U9415 ( .A(n7735), .B(n8283), .ZN(n9736) );
  AOI22_X1 U9416 ( .A1(n9702), .A2(n9704), .B1(n9206), .B2(n9705), .ZN(n7712)
         );
  NAND2_X1 U9417 ( .A1(n7710), .A2(n8283), .ZN(n7732) );
  OAI211_X1 U9418 ( .C1(n7710), .C2(n8283), .A(n7732), .B(n9700), .ZN(n7711)
         );
  OAI211_X1 U9419 ( .C1(n9736), .C2(n9674), .A(n7712), .B(n7711), .ZN(n9740)
         );
  NAND2_X1 U9420 ( .A1(n9740), .A2(n9478), .ZN(n7720) );
  OAI22_X1 U9421 ( .A1(n9478), .A2(n7714), .B1(n7713), .B2(n9693), .ZN(n7718)
         );
  AND2_X1 U9422 ( .A1(n7715), .A2(n9737), .ZN(n7716) );
  OR2_X1 U9423 ( .A1(n7716), .A2(n7743), .ZN(n9739) );
  NOR2_X1 U9424 ( .A1(n9739), .A2(n9266), .ZN(n7717) );
  AOI211_X1 U9425 ( .C1(n9713), .C2(n9737), .A(n7718), .B(n7717), .ZN(n7719)
         );
  OAI211_X1 U9426 ( .C1(n9736), .C2(n7721), .A(n7720), .B(n7719), .ZN(P1_U3280) );
  INV_X1 U9427 ( .A(n7722), .ZN(n7723) );
  AOI22_X1 U9428 ( .A1(n4476), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7723), .B2(
        n8974), .ZN(n7724) );
  OAI21_X1 U9429 ( .B1(n7725), .B2(n8977), .A(n7724), .ZN(n7728) );
  NOR2_X1 U9430 ( .A1(n7726), .A2(n4476), .ZN(n7727) );
  AOI211_X1 U9431 ( .C1(n7729), .C2(n8984), .A(n7728), .B(n7727), .ZN(n7730)
         );
  OAI21_X1 U9432 ( .B1(n8981), .B2(n7731), .A(n7730), .ZN(P2_U3285) );
  NAND2_X1 U9433 ( .A1(n7851), .A2(n7799), .ZN(n8179) );
  XOR2_X1 U9434 ( .A(n7855), .B(n8282), .Z(n7733) );
  AOI222_X1 U9435 ( .A1(n9700), .A2(n7733), .B1(n9205), .B2(n9705), .C1(n9204), 
        .C2(n9702), .ZN(n9731) );
  NAND2_X1 U9436 ( .A1(n9737), .A2(n9205), .ZN(n7734) );
  NAND2_X1 U9437 ( .A1(n7735), .A2(n7734), .ZN(n7737) );
  OR2_X1 U9438 ( .A1(n9737), .A2(n9205), .ZN(n7736) );
  NAND2_X1 U9439 ( .A1(n7737), .A2(n7736), .ZN(n7738) );
  AND2_X1 U9440 ( .A1(n7738), .A2(n8282), .ZN(n9729) );
  INV_X1 U9441 ( .A(n9729), .ZN(n7741) );
  INV_X1 U9442 ( .A(n7738), .ZN(n7740) );
  INV_X1 U9443 ( .A(n8282), .ZN(n7739) );
  NAND3_X1 U9444 ( .A1(n7741), .A2(n9469), .A3(n7853), .ZN(n7749) );
  INV_X1 U9445 ( .A(n7851), .ZN(n9732) );
  INV_X1 U9446 ( .A(n9687), .ZN(n7742) );
  OAI211_X1 U9447 ( .C1(n9732), .C2(n7743), .A(n7742), .B(n9960), .ZN(n9730)
         );
  INV_X1 U9448 ( .A(n7941), .ZN(n7746) );
  AOI22_X1 U9449 ( .A1(n9678), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7791), .B2(
        n9679), .ZN(n7745) );
  NAND2_X1 U9450 ( .A1(n7851), .A2(n9713), .ZN(n7744) );
  OAI211_X1 U9451 ( .C1(n9730), .C2(n7746), .A(n7745), .B(n7744), .ZN(n7747)
         );
  INV_X1 U9452 ( .A(n7747), .ZN(n7748) );
  OAI211_X1 U9453 ( .C1(n9731), .C2(n9678), .A(n7749), .B(n7748), .ZN(P1_U3279) );
  XNOR2_X1 U9454 ( .A(n7750), .B(n5018), .ZN(n9646) );
  INV_X1 U9455 ( .A(n9646), .ZN(n7763) );
  XNOR2_X1 U9456 ( .A(n7751), .B(n8605), .ZN(n7752) );
  OAI222_X1 U9457 ( .A1(n8958), .A2(n7754), .B1(n8956), .B2(n7753), .C1(n7752), 
        .C2(n8953), .ZN(n9644) );
  INV_X1 U9458 ( .A(n7841), .ZN(n9642) );
  INV_X1 U9459 ( .A(n7810), .ZN(n7755) );
  OAI21_X1 U9460 ( .B1(n9642), .B2(n7756), .A(n7755), .ZN(n9643) );
  INV_X1 U9461 ( .A(n7757), .ZN(n7839) );
  OAI22_X1 U9462 ( .A1(n8877), .A2(n7758), .B1(n7839), .B2(n8907), .ZN(n7759)
         );
  AOI21_X1 U9463 ( .B1(n7841), .B2(n7963), .A(n7759), .ZN(n7760) );
  OAI21_X1 U9464 ( .B1(n9643), .B2(n7880), .A(n7760), .ZN(n7761) );
  AOI21_X1 U9465 ( .B1(n9644), .B2(n8877), .A(n7761), .ZN(n7762) );
  OAI21_X1 U9466 ( .B1(n8981), .B2(n7763), .A(n7762), .ZN(P2_U3282) );
  AOI21_X1 U9467 ( .B1(n7765), .B2(n7598), .A(n7764), .ZN(n7767) );
  AOI22_X1 U9468 ( .A1(n7826), .A2(n6202), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7821), .ZN(n7766) );
  NOR2_X1 U9469 ( .A1(n7767), .A2(n7766), .ZN(n7820) );
  AOI21_X1 U9470 ( .B1(n7767), .B2(n7766), .A(n7820), .ZN(n7777) );
  AOI22_X1 U9471 ( .A1(n7826), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7658), .B2(
        n7821), .ZN(n7770) );
  OAI21_X1 U9472 ( .B1(n7771), .B2(n7770), .A(n7825), .ZN(n7772) );
  INV_X1 U9473 ( .A(n9612), .ZN(n10011) );
  NAND2_X1 U9474 ( .A1(n7772), .A2(n10011), .ZN(n7776) );
  NOR2_X1 U9475 ( .A1(n10005), .A2(n7821), .ZN(n7773) );
  AOI211_X1 U9476 ( .C1(P2_ADDR_REG_13__SCAN_IN), .C2(n10013), .A(n7774), .B(
        n7773), .ZN(n7775) );
  OAI211_X1 U9477 ( .C1(n7777), .C2(n8023), .A(n7776), .B(n7775), .ZN(P2_U3258) );
  INV_X1 U9478 ( .A(n7782), .ZN(n7780) );
  NAND2_X1 U9479 ( .A1(n9592), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7779) );
  OR2_X1 U9480 ( .A1(n7778), .A2(P1_U3084), .ZN(n8342) );
  OAI211_X1 U9481 ( .C1(n7780), .C2(n9599), .A(n7779), .B(n8342), .ZN(P1_U3330) );
  NAND2_X1 U9482 ( .A1(n7782), .A2(n7781), .ZN(n7783) );
  OAI211_X1 U9483 ( .C1(n10218), .C2(n9087), .A(n7783), .B(n8631), .ZN(
        P2_U3335) );
  OAI21_X1 U9484 ( .B1(n7786), .B2(n7785), .A(n7784), .ZN(n7787) );
  NAND2_X1 U9485 ( .A1(n7787), .A2(n9660), .ZN(n7793) );
  AND2_X1 U9486 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9844) );
  AOI21_X1 U9487 ( .B1(n9196), .B2(n9204), .A(n9844), .ZN(n7788) );
  OAI21_X1 U9488 ( .B1(n7789), .B2(n9193), .A(n7788), .ZN(n7790) );
  AOI21_X1 U9489 ( .B1(n7791), .B2(n9191), .A(n7790), .ZN(n7792) );
  OAI211_X1 U9490 ( .C1(n9732), .C2(n9199), .A(n7793), .B(n7792), .ZN(P1_U3222) );
  NAND2_X1 U9491 ( .A1(n5480), .A2(n7795), .ZN(n7796) );
  XNOR2_X1 U9492 ( .A(n7797), .B(n7796), .ZN(n7804) );
  NOR2_X1 U9493 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7798), .ZN(n9857) );
  NOR2_X1 U9494 ( .A1(n9193), .A2(n7799), .ZN(n7800) );
  AOI211_X1 U9495 ( .C1(n9196), .C2(n9703), .A(n9857), .B(n7800), .ZN(n7801)
         );
  OAI21_X1 U9496 ( .B1(n9665), .B2(n9694), .A(n7801), .ZN(n7802) );
  AOI21_X1 U9497 ( .B1(n9712), .B2(n9170), .A(n7802), .ZN(n7803) );
  OAI21_X1 U9498 ( .B1(n7804), .B2(n9186), .A(n7803), .ZN(P1_U3232) );
  XNOR2_X1 U9499 ( .A(n7805), .B(n8519), .ZN(n7806) );
  OAI222_X1 U9500 ( .A1(n8958), .A2(n7987), .B1(n8956), .B2(n7807), .C1(n8953), 
        .C2(n7806), .ZN(n7886) );
  INV_X1 U9501 ( .A(n7886), .ZN(n7819) );
  OAI21_X1 U9502 ( .B1(n7809), .B2(n8606), .A(n7808), .ZN(n7888) );
  NOR2_X1 U9503 ( .A1(n7884), .A2(n7810), .ZN(n7811) );
  OR2_X1 U9504 ( .A1(n7876), .A2(n7811), .ZN(n7885) );
  OAI22_X1 U9505 ( .A1(n8877), .A2(n7813), .B1(n7812), .B2(n8907), .ZN(n7814)
         );
  AOI21_X1 U9506 ( .B1(n7815), .B2(n7963), .A(n7814), .ZN(n7816) );
  OAI21_X1 U9507 ( .B1(n7885), .B2(n7880), .A(n7816), .ZN(n7817) );
  AOI21_X1 U9508 ( .B1(n7888), .B2(n8906), .A(n7817), .ZN(n7818) );
  OAI21_X1 U9509 ( .B1(n7819), .B2(n4476), .A(n7818), .ZN(P2_U3281) );
  AOI21_X1 U9510 ( .B1(n7821), .B2(n6202), .A(n7820), .ZN(n7823) );
  INV_X1 U9511 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9647) );
  AOI22_X1 U9512 ( .A1(n8006), .A2(n9647), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n8013), .ZN(n7822) );
  NOR2_X1 U9513 ( .A1(n7823), .A2(n7822), .ZN(n8012) );
  AOI21_X1 U9514 ( .B1(n7823), .B2(n7822), .A(n8012), .ZN(n7834) );
  NOR2_X1 U9515 ( .A1(n8006), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7824) );
  AOI21_X1 U9516 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8006), .A(n7824), .ZN(
        n7828) );
  OAI21_X1 U9517 ( .B1(n7828), .B2(n7827), .A(n8005), .ZN(n7829) );
  NAND2_X1 U9518 ( .A1(n7829), .A2(n10011), .ZN(n7833) );
  INV_X1 U9519 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7830) );
  NAND2_X1 U9520 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7837) );
  OAI21_X1 U9521 ( .B1(n8799), .B2(n7830), .A(n7837), .ZN(n7831) );
  AOI21_X1 U9522 ( .B1(n9618), .B2(n8006), .A(n7831), .ZN(n7832) );
  OAI211_X1 U9523 ( .C1(n7834), .C2(n8023), .A(n7833), .B(n7832), .ZN(P2_U3259) );
  AOI21_X1 U9524 ( .B1(n7836), .B2(n7835), .A(n4560), .ZN(n7843) );
  AOI22_X1 U9525 ( .A1(n8047), .A2(n8713), .B1(n8048), .B2(n8711), .ZN(n7838)
         );
  OAI211_X1 U9526 ( .C1(n7839), .C2(n8698), .A(n7838), .B(n7837), .ZN(n7840)
         );
  AOI21_X1 U9527 ( .B1(n7841), .B2(n6494), .A(n7840), .ZN(n7842) );
  OAI21_X1 U9528 ( .B1(n7843), .B2(n8701), .A(n7842), .ZN(P2_U3217) );
  INV_X1 U9529 ( .A(n7844), .ZN(n7847) );
  INV_X1 U9530 ( .A(n7845), .ZN(n7849) );
  OAI222_X1 U9531 ( .A1(P2_U3152), .A2(n7847), .B1(n4477), .B2(n7849), .C1(
        n7846), .C2(n9087), .ZN(P2_U3334) );
  OAI222_X1 U9532 ( .A1(n7850), .A2(P1_U3084), .B1(n9599), .B2(n7849), .C1(
        n7848), .C2(n9595), .ZN(P1_U3329) );
  INV_X1 U9533 ( .A(n9703), .ZN(n9669) );
  XNOR2_X1 U9534 ( .A(n8082), .B(n9669), .ZN(n8285) );
  NAND2_X1 U9535 ( .A1(n7851), .A2(n9704), .ZN(n7852) );
  OR2_X1 U9536 ( .A1(n9712), .A2(n9204), .ZN(n7854) );
  XOR2_X1 U9537 ( .A(n8285), .B(n7934), .Z(n9549) );
  INV_X1 U9538 ( .A(n9549), .ZN(n7868) );
  INV_X1 U9539 ( .A(n7856), .ZN(n7857) );
  NAND2_X1 U9540 ( .A1(n8179), .A2(n7857), .ZN(n7858) );
  AND2_X1 U9541 ( .A1(n7858), .A2(n8184), .ZN(n8097) );
  INV_X1 U9542 ( .A(n9204), .ZN(n7906) );
  OR2_X1 U9543 ( .A1(n9712), .A2(n7906), .ZN(n8187) );
  NAND2_X1 U9544 ( .A1(n9712), .A2(n7906), .ZN(n8191) );
  NAND2_X1 U9545 ( .A1(n8187), .A2(n8191), .ZN(n9696) );
  INV_X1 U9546 ( .A(n8285), .ZN(n7860) );
  XNOR2_X1 U9547 ( .A(n7928), .B(n7860), .ZN(n7861) );
  NAND2_X1 U9548 ( .A1(n7861), .A2(n9700), .ZN(n7863) );
  AOI22_X1 U9549 ( .A1(n9705), .A2(n9204), .B1(n9203), .B2(n9702), .ZN(n7862)
         );
  NAND2_X1 U9550 ( .A1(n7863), .A2(n7862), .ZN(n9547) );
  INV_X1 U9551 ( .A(n8082), .ZN(n9589) );
  INV_X1 U9552 ( .A(n9712), .ZN(n9723) );
  AOI211_X1 U9553 ( .C1(n8082), .C2(n9689), .A(n9986), .B(n4542), .ZN(n9548)
         );
  NAND2_X1 U9554 ( .A1(n9548), .A2(n7941), .ZN(n7865) );
  AOI22_X1 U9555 ( .A1(n9678), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7902), .B2(
        n9679), .ZN(n7864) );
  OAI211_X1 U9556 ( .C1(n9589), .C2(n9475), .A(n7865), .B(n7864), .ZN(n7866)
         );
  AOI21_X1 U9557 ( .B1(n9478), .B2(n9547), .A(n7866), .ZN(n7867) );
  OAI21_X1 U9558 ( .B1(n7868), .B2(n9415), .A(n7867), .ZN(P1_U3277) );
  XNOR2_X1 U9559 ( .A(n7869), .B(n6537), .ZN(n7872) );
  NAND2_X1 U9560 ( .A1(n8711), .A2(n8966), .ZN(n7871) );
  NAND2_X1 U9561 ( .A1(n8967), .A2(n8968), .ZN(n7870) );
  AND2_X1 U9562 ( .A1(n7871), .A2(n7870), .ZN(n9636) );
  OAI21_X1 U9563 ( .B1(n7872), .B2(n8953), .A(n9636), .ZN(n9640) );
  INV_X1 U9564 ( .A(n9640), .ZN(n7883) );
  INV_X1 U9565 ( .A(n7873), .ZN(n7874) );
  AOI21_X1 U9566 ( .B1(n8522), .B2(n7875), .A(n7874), .ZN(n9641) );
  OAI21_X1 U9567 ( .B1(n9637), .B2(n7876), .A(n4561), .ZN(n9638) );
  INV_X1 U9568 ( .A(n7877), .ZN(n9630) );
  AOI22_X1 U9569 ( .A1(n4476), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n9630), .B2(
        n8974), .ZN(n7879) );
  NAND2_X1 U9570 ( .A1(n9632), .A2(n7963), .ZN(n7878) );
  OAI211_X1 U9571 ( .C1(n9638), .C2(n7880), .A(n7879), .B(n7878), .ZN(n7881)
         );
  AOI21_X1 U9572 ( .B1(n9641), .B2(n8906), .A(n7881), .ZN(n7882) );
  OAI21_X1 U9573 ( .B1(n4476), .B2(n7883), .A(n7882), .ZN(P2_U3280) );
  OAI22_X1 U9574 ( .A1(n7885), .A2(n10078), .B1(n7884), .B2(n10076), .ZN(n7887) );
  AOI211_X1 U9575 ( .C1(n10082), .C2(n7888), .A(n7887), .B(n7886), .ZN(n7890)
         );
  MUX2_X1 U9576 ( .A(n6268), .B(n7890), .S(n10086), .Z(n7889) );
  INV_X1 U9577 ( .A(n7889), .ZN(P2_U3496) );
  MUX2_X1 U9578 ( .A(n6271), .B(n7890), .S(n10098), .Z(n7891) );
  INV_X1 U9579 ( .A(n7891), .ZN(P2_U3535) );
  INV_X1 U9580 ( .A(n6393), .ZN(n7893) );
  OAI222_X1 U9581 ( .A1(P1_U3084), .A2(n7892), .B1(n9599), .B2(n7893), .C1(
        n10217), .C2(n9595), .ZN(P1_U3328) );
  OAI222_X1 U9582 ( .A1(n7895), .A2(n9087), .B1(P2_U3152), .B2(n7894), .C1(
        n4477), .C2(n7893), .ZN(P2_U3333) );
  INV_X1 U9583 ( .A(n5886), .ZN(n7897) );
  INV_X1 U9584 ( .A(n7896), .ZN(n7898) );
  OAI222_X1 U9585 ( .A1(n7897), .A2(P1_U3084), .B1(n9599), .B2(n7898), .C1(
        n10321), .C2(n9595), .ZN(P1_U3327) );
  OAI222_X1 U9586 ( .A1(P2_U3152), .A2(n7899), .B1(n4477), .B2(n7898), .C1(
        n10335), .C2(n9087), .ZN(P2_U3332) );
  XOR2_X1 U9587 ( .A(n7901), .B(n7900), .Z(n7909) );
  NAND2_X1 U9588 ( .A1(n9191), .A2(n7902), .ZN(n7905) );
  AOI21_X1 U9589 ( .B1(n9196), .B2(n9203), .A(n7903), .ZN(n7904) );
  OAI211_X1 U9590 ( .C1(n7906), .C2(n9193), .A(n7905), .B(n7904), .ZN(n7907)
         );
  AOI21_X1 U9591 ( .B1(n8082), .B2(n9170), .A(n7907), .ZN(n7908) );
  OAI21_X1 U9592 ( .B1(n7909), .B2(n9186), .A(n7908), .ZN(P1_U3213) );
  NAND2_X1 U9593 ( .A1(n7910), .A2(n7911), .ZN(n7995) );
  OAI211_X1 U9594 ( .C1(n7910), .C2(n7911), .A(n7995), .B(n9628), .ZN(n7915)
         );
  INV_X1 U9595 ( .A(n7912), .ZN(n8975) );
  AND2_X1 U9596 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8782) );
  OAI22_X1 U9597 ( .A1(n8448), .A2(n8686), .B1(n8687), .B2(n8957), .ZN(n7913)
         );
  AOI211_X1 U9598 ( .C1(n9631), .C2(n8975), .A(n8782), .B(n7913), .ZN(n7914)
         );
  OAI211_X1 U9599 ( .C1(n8978), .C2(n8692), .A(n7915), .B(n7914), .ZN(P2_U3240) );
  INV_X1 U9600 ( .A(n7920), .ZN(n7917) );
  OAI21_X1 U9601 ( .B1(n7917), .B2(n7916), .A(n9660), .ZN(n7927) );
  AOI21_X1 U9602 ( .B1(n7920), .B2(n7919), .A(n7918), .ZN(n7926) );
  INV_X1 U9603 ( .A(n9463), .ZN(n9671) );
  NOR2_X1 U9604 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7921), .ZN(n9869) );
  AOI21_X1 U9605 ( .B1(n9655), .B2(n9703), .A(n9869), .ZN(n7922) );
  OAI21_X1 U9606 ( .B1(n9671), .B2(n9652), .A(n7922), .ZN(n7924) );
  NAND2_X1 U9607 ( .A1(n9682), .A2(n9959), .ZN(n9716) );
  INV_X1 U9608 ( .A(n9659), .ZN(n9151) );
  NOR2_X1 U9609 ( .A1(n9716), .A2(n9151), .ZN(n7923) );
  AOI211_X1 U9610 ( .C1(n9680), .C2(n9191), .A(n7924), .B(n7923), .ZN(n7925)
         );
  OAI21_X1 U9611 ( .B1(n7927), .B2(n7926), .A(n7925), .ZN(P1_U3239) );
  OR2_X1 U9612 ( .A1(n8082), .A2(n9669), .ZN(n8194) );
  INV_X1 U9613 ( .A(n9203), .ZN(n7971) );
  NAND2_X1 U9614 ( .A1(n9682), .A2(n7971), .ZN(n8198) );
  NAND2_X1 U9615 ( .A1(n9667), .A2(n8198), .ZN(n8397) );
  OR2_X1 U9616 ( .A1(n9682), .A2(n7971), .ZN(n8199) );
  NAND2_X1 U9617 ( .A1(n8397), .A2(n8199), .ZN(n7929) );
  OR2_X1 U9618 ( .A1(n8372), .A2(n9671), .ZN(n8203) );
  NAND2_X1 U9619 ( .A1(n8372), .A2(n9671), .ZN(n8204) );
  NAND2_X1 U9620 ( .A1(n8203), .A2(n8204), .ZN(n8370) );
  XNOR2_X1 U9621 ( .A(n7929), .B(n8370), .ZN(n7930) );
  NAND2_X1 U9622 ( .A1(n7930), .A2(n9700), .ZN(n7932) );
  AOI22_X1 U9623 ( .A1(n9443), .A2(n9702), .B1(n9705), .B2(n9203), .ZN(n7931)
         );
  NAND2_X1 U9624 ( .A1(n7932), .A2(n7931), .ZN(n9543) );
  INV_X1 U9625 ( .A(n9543), .ZN(n7944) );
  AND2_X1 U9626 ( .A1(n8082), .A2(n9703), .ZN(n7933) );
  OAI22_X1 U9627 ( .A1(n7934), .A2(n7933), .B1(n9703), .B2(n8082), .ZN(n9673)
         );
  NOR2_X1 U9628 ( .A1(n9682), .A2(n9203), .ZN(n7935) );
  OR2_X1 U9629 ( .A1(n9673), .A2(n7935), .ZN(n7937) );
  NAND2_X1 U9630 ( .A1(n9682), .A2(n9203), .ZN(n7936) );
  NAND2_X1 U9631 ( .A1(n7937), .A2(n7936), .ZN(n8371) );
  INV_X1 U9632 ( .A(n8370), .ZN(n8201) );
  XNOR2_X1 U9633 ( .A(n8371), .B(n8201), .ZN(n9545) );
  NAND2_X1 U9634 ( .A1(n9545), .A2(n9469), .ZN(n7943) );
  INV_X1 U9635 ( .A(n8372), .ZN(n9584) );
  AOI211_X1 U9636 ( .C1(n8372), .C2(n4495), .A(n9986), .B(n9470), .ZN(n9544)
         );
  NOR2_X1 U9637 ( .A1(n9584), .A2(n9475), .ZN(n7940) );
  INV_X1 U9638 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7938) );
  OAI22_X1 U9639 ( .A1(n9478), .A2(n7938), .B1(n7974), .B2(n9693), .ZN(n7939)
         );
  AOI211_X1 U9640 ( .C1(n9544), .C2(n7941), .A(n7940), .B(n7939), .ZN(n7942)
         );
  OAI211_X1 U9641 ( .C1(n9709), .C2(n7944), .A(n7943), .B(n7942), .ZN(P1_U3275) );
  INV_X1 U9642 ( .A(n7945), .ZN(n7948) );
  NAND2_X1 U9643 ( .A1(n9592), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7946) );
  OAI211_X1 U9644 ( .C1(n7948), .C2(n9599), .A(n7947), .B(n7946), .ZN(P1_U3326) );
  OAI222_X1 U9645 ( .A1(n9087), .A2(n7949), .B1(n4477), .B2(n7948), .C1(n8627), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U9646 ( .A(n7950), .ZN(n8059) );
  NAND2_X1 U9647 ( .A1(n9592), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n7952) );
  OAI211_X1 U9648 ( .C1(n8059), .C2(n9599), .A(n7952), .B(n7951), .ZN(P1_U3325) );
  AND2_X1 U9649 ( .A1(n7953), .A2(n8607), .ZN(n7954) );
  NOR2_X1 U9650 ( .A1(n7955), .A2(n7954), .ZN(n9055) );
  XOR2_X1 U9651 ( .A(n7956), .B(n8607), .Z(n7957) );
  AOI222_X1 U9652 ( .A1(n8971), .A2(n7957), .B1(n8709), .B2(n8968), .C1(n8710), 
        .C2(n8966), .ZN(n9053) );
  AOI21_X1 U9653 ( .B1(n4561), .B2(n9051), .A(n10078), .ZN(n7958) );
  AND2_X1 U9654 ( .A1(n7958), .A2(n4483), .ZN(n9050) );
  NOR2_X1 U9655 ( .A1(n8907), .A2(n7985), .ZN(n7959) );
  AOI21_X1 U9656 ( .B1(n9050), .B2(n8618), .A(n7959), .ZN(n7960) );
  OAI211_X1 U9657 ( .C1(n9055), .C2(n7961), .A(n9053), .B(n7960), .ZN(n7962)
         );
  NAND2_X1 U9658 ( .A1(n7962), .A2(n8877), .ZN(n7965) );
  AOI22_X1 U9659 ( .A1(n9051), .A2(n7963), .B1(n4476), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n7964) );
  OAI211_X1 U9660 ( .C1(n9055), .C2(n7966), .A(n7965), .B(n7964), .ZN(P2_U3279) );
  XOR2_X1 U9661 ( .A(n7968), .B(n7967), .Z(n7969) );
  XNOR2_X1 U9662 ( .A(n7970), .B(n7969), .ZN(n7977) );
  AND2_X1 U9663 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9881) );
  NOR2_X1 U9664 ( .A1(n9193), .A2(n7971), .ZN(n7972) );
  AOI211_X1 U9665 ( .C1(n9196), .C2(n9443), .A(n9881), .B(n7972), .ZN(n7973)
         );
  OAI21_X1 U9666 ( .B1(n7974), .B2(n9665), .A(n7973), .ZN(n7975) );
  AOI21_X1 U9667 ( .B1(n8372), .B2(n9170), .A(n7975), .ZN(n7976) );
  OAI21_X1 U9668 ( .B1(n7977), .B2(n9186), .A(n7976), .ZN(P1_U3224) );
  AOI21_X1 U9669 ( .B1(n6625), .B2(n7979), .A(n7978), .ZN(n9627) );
  XNOR2_X1 U9670 ( .A(n7981), .B(n7980), .ZN(n9626) );
  NAND2_X1 U9671 ( .A1(n9627), .A2(n9626), .ZN(n9625) );
  AOI21_X1 U9672 ( .B1(n9625), .B2(n7983), .A(n7982), .ZN(n7992) );
  NAND2_X1 U9673 ( .A1(n7984), .A2(n9628), .ZN(n7991) );
  INV_X1 U9674 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10279) );
  OAI22_X1 U9675 ( .A1(n8698), .A2(n7985), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10279), .ZN(n7989) );
  OAI22_X1 U9676 ( .A1(n7987), .A2(n8686), .B1(n8687), .B2(n7986), .ZN(n7988)
         );
  AOI211_X1 U9677 ( .C1(n9051), .C2(n6494), .A(n7989), .B(n7988), .ZN(n7990)
         );
  OAI21_X1 U9678 ( .B1(n7992), .B2(n7991), .A(n7990), .ZN(P2_U3230) );
  AND2_X1 U9679 ( .A1(n7995), .A2(n7993), .ZN(n7998) );
  NAND2_X1 U9680 ( .A1(n7995), .A2(n7994), .ZN(n7996) );
  OAI21_X1 U9681 ( .B1(n7998), .B2(n7997), .A(n7996), .ZN(n7999) );
  NAND2_X1 U9682 ( .A1(n7999), .A2(n9628), .ZN(n8004) );
  INV_X1 U9683 ( .A(n8000), .ZN(n8036) );
  AOI22_X1 U9684 ( .A1(n8966), .A2(n8709), .B1(n8939), .B2(n8968), .ZN(n8032)
         );
  OAI22_X1 U9685 ( .A1(n9635), .A2(n8032), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8001), .ZN(n8002) );
  AOI21_X1 U9686 ( .B1(n8036), .B2(n9631), .A(n8002), .ZN(n8003) );
  OAI211_X1 U9687 ( .C1(n8039), .C2(n8692), .A(n8004), .B(n8003), .ZN(P2_U3221) );
  OAI21_X1 U9688 ( .B1(n8006), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8005), .ZN(
        n8007) );
  NAND2_X1 U9689 ( .A1(n8014), .A2(n8007), .ZN(n8008) );
  XNOR2_X1 U9690 ( .A(n8007), .B(n8746), .ZN(n8740) );
  NAND2_X1 U9691 ( .A1(n8740), .A2(n7813), .ZN(n8739) );
  NAND2_X1 U9692 ( .A1(n8008), .A2(n8739), .ZN(n8011) );
  NAND2_X1 U9693 ( .A1(n8757), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8009) );
  OAI21_X1 U9694 ( .B1(n8757), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8009), .ZN(
        n8010) );
  NOR2_X1 U9695 ( .A1(n8010), .A2(n8011), .ZN(n8752) );
  AOI211_X1 U9696 ( .C1(n8011), .C2(n8010), .A(n8752), .B(n9612), .ZN(n8026)
         );
  AOI21_X1 U9697 ( .B1(n8013), .B2(n9647), .A(n8012), .ZN(n8015) );
  NAND2_X1 U9698 ( .A1(n8746), .A2(n8015), .ZN(n8016) );
  XNOR2_X1 U9699 ( .A(n8015), .B(n8014), .ZN(n8745) );
  NAND2_X1 U9700 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8745), .ZN(n8744) );
  NAND2_X1 U9701 ( .A1(n8016), .A2(n8744), .ZN(n8019) );
  INV_X1 U9702 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8017) );
  MUX2_X1 U9703 ( .A(n8017), .B(P2_REG1_REG_16__SCAN_IN), .S(n8757), .Z(n8018)
         );
  NOR2_X1 U9704 ( .A1(n8018), .A2(n8019), .ZN(n8758) );
  AOI21_X1 U9705 ( .B1(n8019), .B2(n8018), .A(n8758), .ZN(n8024) );
  NAND2_X1 U9706 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n9633) );
  INV_X1 U9707 ( .A(n9633), .ZN(n8020) );
  AOI21_X1 U9708 ( .B1(n10013), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8020), .ZN(
        n8022) );
  NAND2_X1 U9709 ( .A1(n9618), .A2(n8757), .ZN(n8021) );
  OAI211_X1 U9710 ( .C1(n8024), .C2(n8023), .A(n8022), .B(n8021), .ZN(n8025)
         );
  OR2_X1 U9711 ( .A1(n8026), .A2(n8025), .ZN(P2_U3261) );
  XNOR2_X1 U9712 ( .A(n8027), .B(n8028), .ZN(n9044) );
  INV_X1 U9713 ( .A(n8951), .ZN(n8031) );
  INV_X1 U9714 ( .A(n8586), .ZN(n8533) );
  INV_X1 U9715 ( .A(n8028), .ZN(n8609) );
  AOI21_X1 U9716 ( .B1(n8029), .B2(n8533), .A(n8609), .ZN(n8030) );
  OAI21_X1 U9717 ( .B1(n8031), .B2(n8030), .A(n8971), .ZN(n8033) );
  NAND2_X1 U9718 ( .A1(n8033), .A2(n8032), .ZN(n9040) );
  INV_X1 U9719 ( .A(n8973), .ZN(n8035) );
  INV_X1 U9720 ( .A(n8946), .ZN(n8034) );
  AOI211_X1 U9721 ( .C1(n9042), .C2(n8035), .A(n10078), .B(n8034), .ZN(n9041)
         );
  NAND2_X1 U9722 ( .A1(n9041), .A2(n8871), .ZN(n8038) );
  AOI22_X1 U9723 ( .A1(n4476), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8036), .B2(
        n8974), .ZN(n8037) );
  OAI211_X1 U9724 ( .C1(n8039), .C2(n8977), .A(n8038), .B(n8037), .ZN(n8040)
         );
  AOI21_X1 U9725 ( .B1(n9040), .B2(n8877), .A(n8040), .ZN(n8041) );
  OAI21_X1 U9726 ( .B1(n9044), .B2(n8981), .A(n8041), .ZN(P2_U3277) );
  INV_X1 U9727 ( .A(n8042), .ZN(n8043) );
  AOI211_X1 U9728 ( .C1(n8045), .C2(n8044), .A(n8701), .B(n8043), .ZN(n8052)
         );
  INV_X1 U9729 ( .A(n9035), .ZN(n8949) );
  INV_X1 U9730 ( .A(n8046), .ZN(n8947) );
  AOI22_X1 U9731 ( .A1(n9631), .A2(n8947), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8050) );
  AOI22_X1 U9732 ( .A1(n8048), .A2(n8708), .B1(n8047), .B2(n8969), .ZN(n8049)
         );
  OAI211_X1 U9733 ( .C1(n8949), .C2(n8692), .A(n8050), .B(n8049), .ZN(n8051)
         );
  OR2_X1 U9734 ( .A1(n8052), .A2(n8051), .ZN(P2_U3235) );
  INV_X1 U9735 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8058) );
  INV_X1 U9736 ( .A(n8053), .ZN(n8054) );
  NAND2_X1 U9737 ( .A1(n8054), .A2(SI_29_), .ZN(n8055) );
  MUX2_X1 U9738 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n4481), .Z(n8125) );
  INV_X1 U9739 ( .A(n8432), .ZN(n8641) );
  OAI222_X1 U9740 ( .A1(n9595), .A2(n8058), .B1(n9599), .B2(n8641), .C1(
        P1_U3084), .C2(n8057), .ZN(P1_U3323) );
  OAI222_X1 U9741 ( .A1(n4477), .A2(n8059), .B1(P2_U3152), .B2(n4474), .C1(
        n10290), .C2(n9087), .ZN(P2_U3330) );
  OAI222_X1 U9742 ( .A1(n5907), .A2(P1_U3084), .B1(n9599), .B2(n8061), .C1(
        n8060), .C2(n9595), .ZN(P1_U3332) );
  NAND2_X1 U9743 ( .A1(n5210), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8064) );
  NAND2_X1 U9744 ( .A1(n8133), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8063) );
  NAND2_X1 U9745 ( .A1(n5382), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8062) );
  NAND3_X1 U9746 ( .A1(n8064), .A2(n8063), .A3(n8062), .ZN(n9257) );
  NAND2_X1 U9747 ( .A1(n8356), .A2(n9257), .ZN(n8263) );
  NAND2_X1 U9748 ( .A1(n9489), .A2(n8065), .ZN(n8245) );
  INV_X1 U9749 ( .A(n8066), .ZN(n8093) );
  NAND2_X1 U9750 ( .A1(n6854), .A2(n8067), .ZN(n8068) );
  OAI211_X1 U9751 ( .C1(n8069), .C2(n6933), .A(n8297), .B(n8068), .ZN(n8070)
         );
  NAND2_X1 U9752 ( .A1(n8070), .A2(n7195), .ZN(n8072) );
  OAI21_X1 U9753 ( .B1(n8073), .B2(n8072), .A(n8071), .ZN(n8077) );
  NAND2_X1 U9754 ( .A1(n8154), .A2(n8074), .ZN(n8075) );
  NOR2_X1 U9755 ( .A1(n8275), .A2(n8075), .ZN(n8302) );
  INV_X1 U9756 ( .A(n8302), .ZN(n8076) );
  AOI21_X1 U9757 ( .B1(n8077), .B2(n8303), .A(n8076), .ZN(n8092) );
  INV_X1 U9758 ( .A(n9327), .ZN(n9194) );
  INV_X1 U9759 ( .A(n9352), .ZN(n9322) );
  NAND2_X1 U9760 ( .A1(n9331), .A2(n9322), .ZN(n8407) );
  NAND2_X1 U9761 ( .A1(n8265), .A2(n8407), .ZN(n8228) );
  INV_X1 U9762 ( .A(n9351), .ZN(n9380) );
  NAND2_X1 U9763 ( .A1(n9514), .A2(n9380), .ZN(n8288) );
  INV_X1 U9764 ( .A(n9402), .ZN(n8078) );
  INV_X1 U9765 ( .A(n9202), .ZN(n9428) );
  NAND2_X1 U9766 ( .A1(n9408), .A2(n9428), .ZN(n8209) );
  INV_X1 U9767 ( .A(n8209), .ZN(n8270) );
  NAND2_X1 U9768 ( .A1(n8269), .A2(n8270), .ZN(n8079) );
  AND2_X1 U9769 ( .A1(n8079), .A2(n9364), .ZN(n8080) );
  NAND2_X1 U9770 ( .A1(n8288), .A2(n8080), .ZN(n8111) );
  INV_X1 U9771 ( .A(n8111), .ZN(n8081) );
  INV_X1 U9772 ( .A(n9444), .ZN(n9180) );
  NAND2_X1 U9773 ( .A1(n9431), .A2(n9180), .ZN(n9396) );
  INV_X1 U9774 ( .A(n9367), .ZN(n9147) );
  NAND2_X1 U9775 ( .A1(n9509), .A2(n9147), .ZN(n8268) );
  AND3_X1 U9776 ( .A1(n8081), .A2(n9396), .A3(n8268), .ZN(n8105) );
  INV_X1 U9777 ( .A(n8105), .ZN(n8091) );
  INV_X1 U9778 ( .A(n9464), .ZN(n9427) );
  NAND2_X1 U9779 ( .A1(n9452), .A2(n9427), .ZN(n8399) );
  INV_X1 U9780 ( .A(n9443), .ZN(n8106) );
  NAND2_X1 U9781 ( .A1(n9474), .A2(n8106), .ZN(n8202) );
  NAND2_X1 U9782 ( .A1(n8399), .A2(n8202), .ZN(n8141) );
  INV_X1 U9783 ( .A(n8204), .ZN(n8395) );
  NAND2_X1 U9784 ( .A1(n8082), .A2(n9669), .ZN(n8192) );
  NAND2_X1 U9785 ( .A1(n8179), .A2(n8083), .ZN(n8185) );
  NAND2_X1 U9786 ( .A1(n8178), .A2(n8156), .ZN(n8084) );
  AND2_X1 U9787 ( .A1(n8084), .A2(n8173), .ZN(n8085) );
  OR2_X1 U9788 ( .A1(n8185), .A2(n8085), .ZN(n8096) );
  INV_X1 U9789 ( .A(n8096), .ZN(n8087) );
  AND2_X1 U9790 ( .A1(n8086), .A2(n8147), .ZN(n8157) );
  AND4_X1 U9791 ( .A1(n8192), .A2(n8087), .A3(n8157), .A4(n8191), .ZN(n8088)
         );
  NAND2_X1 U9792 ( .A1(n8198), .A2(n8088), .ZN(n8089) );
  OR3_X1 U9793 ( .A1(n8141), .A2(n8395), .A3(n8089), .ZN(n8090) );
  OR3_X1 U9794 ( .A1(n8228), .A2(n8091), .A3(n8090), .ZN(n8316) );
  AOI211_X1 U9795 ( .C1(n8093), .C2(n8154), .A(n8092), .B(n8316), .ZN(n8116)
         );
  INV_X1 U9796 ( .A(n8141), .ZN(n8104) );
  AND2_X1 U9797 ( .A1(n8203), .A2(n8199), .ZN(n8396) );
  AND2_X1 U9798 ( .A1(n8173), .A2(n8094), .ZN(n8095) );
  NOR2_X1 U9799 ( .A1(n8096), .A2(n8095), .ZN(n8099) );
  AND2_X1 U9800 ( .A1(n8097), .A2(n8187), .ZN(n8189) );
  INV_X1 U9801 ( .A(n8189), .ZN(n8098) );
  OAI21_X1 U9802 ( .B1(n8099), .B2(n8098), .A(n8191), .ZN(n8100) );
  NAND2_X1 U9803 ( .A1(n8100), .A2(n8194), .ZN(n8101) );
  NAND3_X1 U9804 ( .A1(n8101), .A2(n8198), .A3(n8192), .ZN(n8102) );
  AOI21_X1 U9805 ( .B1(n8396), .B2(n8102), .A(n8395), .ZN(n8103) );
  NAND3_X1 U9806 ( .A1(n8105), .A2(n8104), .A3(n8103), .ZN(n8114) );
  OR2_X1 U9807 ( .A1(n9331), .A2(n9322), .ZN(n8267) );
  NAND2_X1 U9808 ( .A1(n8404), .A2(n8269), .ZN(n8220) );
  NAND2_X1 U9809 ( .A1(n9396), .A2(n8399), .ZN(n8211) );
  OR2_X1 U9810 ( .A1(n9452), .A2(n9427), .ZN(n8272) );
  NAND2_X1 U9811 ( .A1(n8272), .A2(n8398), .ZN(n8142) );
  INV_X1 U9812 ( .A(n8142), .ZN(n8107) );
  NOR2_X1 U9813 ( .A1(n8211), .A2(n8107), .ZN(n8110) );
  NOR2_X1 U9814 ( .A1(n9408), .A2(n9428), .ZN(n9401) );
  OR2_X1 U9815 ( .A1(n9431), .A2(n9180), .ZN(n8271) );
  INV_X1 U9816 ( .A(n8271), .ZN(n8108) );
  NOR2_X1 U9817 ( .A1(n9401), .A2(n8108), .ZN(n8210) );
  INV_X1 U9818 ( .A(n8210), .ZN(n8109) );
  OR3_X1 U9819 ( .A1(n8220), .A2(n8110), .A3(n8109), .ZN(n8112) );
  NAND2_X1 U9820 ( .A1(n8111), .A2(n8404), .ZN(n8217) );
  NAND3_X1 U9821 ( .A1(n8112), .A2(n8217), .A3(n8268), .ZN(n8113) );
  AND4_X1 U9822 ( .A1(n8114), .A2(n8267), .A3(n8113), .A4(n8405), .ZN(n8115)
         );
  INV_X1 U9823 ( .A(n9287), .ZN(n9321) );
  OR2_X1 U9824 ( .A1(n9494), .A2(n9321), .ZN(n8266) );
  OAI211_X1 U9825 ( .C1(n8115), .C2(n8228), .A(n8266), .B(n8409), .ZN(n8318)
         );
  NOR2_X1 U9826 ( .A1(n8116), .A2(n8318), .ZN(n8117) );
  INV_X1 U9827 ( .A(n8413), .ZN(n8234) );
  NAND2_X1 U9828 ( .A1(n9494), .A2(n9321), .ZN(n8412) );
  NAND2_X1 U9829 ( .A1(n8420), .A2(n9253), .ZN(n9254) );
  OAI211_X1 U9830 ( .C1(n8234), .C2(n8412), .A(n9254), .B(n8245), .ZN(n8319)
         );
  AOI21_X1 U9831 ( .B1(n9285), .B2(n8117), .A(n8319), .ZN(n8121) );
  NAND2_X1 U9832 ( .A1(n9086), .A2(n8132), .ZN(n8119) );
  NAND2_X1 U9833 ( .A1(n8131), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8118) );
  INV_X1 U9834 ( .A(n9201), .ZN(n8120) );
  NAND2_X1 U9835 ( .A1(n8264), .A2(n8249), .ZN(n8324) );
  NAND2_X1 U9836 ( .A1(n9485), .A2(n8120), .ZN(n8322) );
  OAI21_X1 U9837 ( .B1(n8121), .B2(n8324), .A(n8322), .ZN(n8122) );
  NOR2_X1 U9838 ( .A1(n8356), .A2(n9257), .ZN(n8294) );
  AOI21_X1 U9839 ( .B1(n8263), .B2(n8122), .A(n8294), .ZN(n8138) );
  INV_X1 U9840 ( .A(n8123), .ZN(n8124) );
  NAND2_X1 U9841 ( .A1(n8124), .A2(SI_30_), .ZN(n8128) );
  NAND2_X1 U9842 ( .A1(n8126), .A2(n8125), .ZN(n8127) );
  MUX2_X1 U9843 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n4481), .Z(n8129) );
  XNOR2_X1 U9844 ( .A(n8129), .B(SI_31_), .ZN(n8130) );
  NAND2_X1 U9845 ( .A1(n5210), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8136) );
  NAND2_X1 U9846 ( .A1(n8133), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8135) );
  NAND2_X1 U9847 ( .A1(n5382), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8134) );
  NAND3_X1 U9848 ( .A1(n8136), .A2(n8135), .A3(n8134), .ZN(n9200) );
  NOR2_X1 U9849 ( .A1(n8369), .A2(n9200), .ZN(n8296) );
  INV_X1 U9850 ( .A(n8369), .ZN(n8357) );
  INV_X1 U9851 ( .A(n9200), .ZN(n8137) );
  INV_X1 U9852 ( .A(n8326), .ZN(n8298) );
  OAI21_X1 U9853 ( .B1(n8138), .B2(n8296), .A(n8298), .ZN(n8140) );
  XNOR2_X1 U9854 ( .A(n8140), .B(n8139), .ZN(n8336) );
  MUX2_X1 U9855 ( .A(n8142), .B(n8141), .S(n8258), .Z(n8208) );
  INV_X1 U9856 ( .A(n8192), .ZN(n8197) );
  INV_X1 U9857 ( .A(n8143), .ZN(n8144) );
  INV_X1 U9858 ( .A(n8146), .ZN(n8148) );
  AND4_X1 U9859 ( .A1(n8150), .A2(n8154), .A3(n8149), .A4(n8213), .ZN(n8151)
         );
  NAND3_X1 U9860 ( .A1(n8152), .A2(n8151), .A3(n8173), .ZN(n8183) );
  AND2_X1 U9861 ( .A1(n8154), .A2(n8153), .ZN(n8310) );
  NAND2_X1 U9862 ( .A1(n8155), .A2(n8310), .ZN(n8177) );
  AND4_X1 U9863 ( .A1(n8178), .A2(n8157), .A3(n8258), .A4(n8156), .ZN(n8176)
         );
  OAI21_X1 U9864 ( .B1(n9207), .B2(n9654), .A(n8258), .ZN(n8158) );
  AOI21_X1 U9865 ( .B1(n8165), .B2(n8159), .A(n8158), .ZN(n8163) );
  OR3_X1 U9866 ( .A1(n8160), .A2(n8159), .A3(n8165), .ZN(n8161) );
  NAND2_X1 U9867 ( .A1(n8166), .A2(n8161), .ZN(n8162) );
  NAND3_X1 U9868 ( .A1(n8178), .A2(n8163), .A3(n8162), .ZN(n8172) );
  NOR2_X1 U9869 ( .A1(n9654), .A2(n8258), .ZN(n8164) );
  NAND2_X1 U9870 ( .A1(n8165), .A2(n8164), .ZN(n8169) );
  OAI21_X1 U9871 ( .B1(n8258), .B2(n9207), .A(n8169), .ZN(n8167) );
  NAND2_X1 U9872 ( .A1(n8167), .A2(n8166), .ZN(n8168) );
  OAI21_X1 U9873 ( .B1(n8169), .B2(n9207), .A(n8168), .ZN(n8170) );
  NAND2_X1 U9874 ( .A1(n8173), .A2(n8170), .ZN(n8171) );
  OAI211_X1 U9875 ( .C1(n8173), .C2(n8213), .A(n8172), .B(n8171), .ZN(n8175)
         );
  INV_X1 U9876 ( .A(n8184), .ZN(n8174) );
  NAND2_X1 U9877 ( .A1(n8179), .A2(n8178), .ZN(n8180) );
  NAND2_X1 U9878 ( .A1(n8180), .A2(n8213), .ZN(n8181) );
  NAND4_X1 U9879 ( .A1(n8183), .A2(n8283), .A3(n8182), .A4(n8181), .ZN(n8190)
         );
  NAND2_X1 U9880 ( .A1(n8185), .A2(n8184), .ZN(n8186) );
  NAND4_X1 U9881 ( .A1(n8190), .A2(n8258), .A3(n8191), .A4(n8186), .ZN(n8196)
         );
  NAND2_X1 U9882 ( .A1(n8194), .A2(n8187), .ZN(n8188) );
  NAND2_X1 U9883 ( .A1(n8188), .A2(n8192), .ZN(n8195) );
  NAND2_X1 U9884 ( .A1(n8190), .A2(n8189), .ZN(n8193) );
  MUX2_X1 U9885 ( .A(n8199), .B(n8198), .S(n8258), .Z(n8200) );
  MUX2_X1 U9886 ( .A(n8204), .B(n8203), .S(n8258), .Z(n8205) );
  AND2_X1 U9887 ( .A1(n8209), .A2(n9396), .ZN(n8400) );
  OAI21_X1 U9888 ( .B1(n8212), .B2(n8211), .A(n8210), .ZN(n8214) );
  AND2_X1 U9889 ( .A1(n8217), .A2(n8268), .ZN(n8218) );
  OAI211_X1 U9890 ( .C1(n8220), .C2(n8219), .A(n8407), .B(n8218), .ZN(n8224)
         );
  INV_X1 U9891 ( .A(n9401), .ZN(n9375) );
  INV_X1 U9892 ( .A(n9364), .ZN(n8402) );
  NAND2_X1 U9893 ( .A1(n8222), .A2(n8267), .ZN(n8223) );
  INV_X1 U9894 ( .A(n8405), .ZN(n8225) );
  INV_X1 U9895 ( .A(n8268), .ZN(n8226) );
  AND2_X1 U9896 ( .A1(n8267), .A2(n8226), .ZN(n8227) );
  OR2_X1 U9897 ( .A1(n8228), .A2(n8227), .ZN(n8229) );
  INV_X1 U9898 ( .A(n8407), .ZN(n8230) );
  OAI211_X1 U9899 ( .C1(n8230), .C2(n8405), .A(n8409), .B(n8267), .ZN(n8231)
         );
  AOI21_X1 U9900 ( .B1(n8265), .B2(n9287), .A(n8234), .ZN(n8237) );
  INV_X1 U9901 ( .A(n8245), .ZN(n8235) );
  AOI21_X1 U9902 ( .B1(n8409), .B2(n9494), .A(n8235), .ZN(n8236) );
  MUX2_X1 U9903 ( .A(n8237), .B(n8236), .S(n8258), .Z(n8238) );
  AOI21_X1 U9904 ( .B1(n8239), .B2(n9285), .A(n8238), .ZN(n8248) );
  AOI21_X1 U9905 ( .B1(n8241), .B2(n8265), .A(n9287), .ZN(n8240) );
  NOR2_X1 U9906 ( .A1(n8240), .A2(n9494), .ZN(n8244) );
  AOI21_X1 U9907 ( .B1(n8241), .B2(n8409), .A(n9494), .ZN(n8242) );
  NOR2_X1 U9908 ( .A1(n8242), .A2(n9287), .ZN(n8243) );
  MUX2_X1 U9909 ( .A(n8245), .B(n8413), .S(n8258), .Z(n8246) );
  OR2_X1 U9910 ( .A1(n8249), .A2(n8258), .ZN(n8255) );
  INV_X1 U9911 ( .A(n9485), .ZN(n8252) );
  OAI21_X1 U9912 ( .B1(n9201), .B2(n9254), .A(n8252), .ZN(n8250) );
  MUX2_X1 U9913 ( .A(n9201), .B(n8250), .S(n8258), .Z(n8251) );
  NOR2_X1 U9914 ( .A1(n8296), .A2(n8258), .ZN(n8253) );
  AOI21_X1 U9915 ( .B1(n9200), .B2(n9257), .A(n8356), .ZN(n8321) );
  MUX2_X1 U9916 ( .A(n9201), .B(n9485), .S(n8213), .Z(n8256) );
  OAI211_X1 U9917 ( .C1(n8213), .C2(n9254), .A(n8256), .B(n8255), .ZN(n8257)
         );
  OAI21_X1 U9918 ( .B1(n9430), .B2(n8262), .A(n8261), .ZN(n8332) );
  INV_X1 U9919 ( .A(n8263), .ZN(n8295) );
  INV_X1 U9920 ( .A(n9255), .ZN(n8292) );
  NAND2_X1 U9921 ( .A1(n8266), .A2(n8412), .ZN(n9301) );
  NAND2_X1 U9922 ( .A1(n8267), .A2(n8407), .ZN(n9329) );
  NAND2_X1 U9923 ( .A1(n8405), .A2(n8268), .ZN(n9342) );
  OR2_X1 U9924 ( .A1(n9401), .A2(n8270), .ZN(n9397) );
  INV_X1 U9925 ( .A(n9672), .ZN(n9666) );
  NAND4_X1 U9926 ( .A1(n8274), .A2(n4486), .A3(n8273), .A4(n7283), .ZN(n8276)
         );
  OR4_X1 U9927 ( .A1(n8277), .A2(n8276), .A3(n8312), .A4(n8275), .ZN(n8280) );
  NOR4_X1 U9928 ( .A1(n8280), .A2(n8279), .A3(n8278), .A4(n7431), .ZN(n8281)
         );
  NAND4_X1 U9929 ( .A1(n7859), .A2(n8283), .A3(n8282), .A4(n8281), .ZN(n8284)
         );
  NOR4_X1 U9930 ( .A1(n8370), .A2(n8285), .A3(n9666), .A4(n8284), .ZN(n8286)
         );
  NAND4_X1 U9931 ( .A1(n9433), .A2(n9467), .A3(n9449), .A4(n8286), .ZN(n8287)
         );
  NOR4_X1 U9932 ( .A1(n9342), .A2(n9387), .A3(n9397), .A4(n8287), .ZN(n8289)
         );
  NAND2_X1 U9933 ( .A1(n8404), .A2(n8288), .ZN(n9358) );
  INV_X1 U9934 ( .A(n9358), .ZN(n9365) );
  NAND2_X1 U9935 ( .A1(n8289), .A2(n9365), .ZN(n8290) );
  NOR4_X1 U9936 ( .A1(n9318), .A2(n9301), .A3(n9329), .A4(n8290), .ZN(n8291)
         );
  NAND4_X1 U9937 ( .A1(n8292), .A2(n9285), .A3(n8414), .A4(n8291), .ZN(n8293)
         );
  NOR4_X1 U9938 ( .A1(n8296), .A2(n8295), .A3(n8294), .A4(n8293), .ZN(n8299)
         );
  AOI21_X1 U9939 ( .B1(n8299), .B2(n8298), .A(n8297), .ZN(n8330) );
  NAND2_X1 U9940 ( .A1(n8302), .A2(n8301), .ZN(n8314) );
  INV_X1 U9941 ( .A(n8303), .ZN(n8311) );
  NAND2_X1 U9942 ( .A1(n8305), .A2(n8304), .ZN(n8306) );
  NAND3_X1 U9943 ( .A1(n8308), .A2(n8307), .A3(n8306), .ZN(n8309) );
  OAI211_X1 U9944 ( .C1(n8312), .C2(n8311), .A(n8310), .B(n8309), .ZN(n8313)
         );
  NAND2_X1 U9945 ( .A1(n8314), .A2(n8313), .ZN(n8315) );
  NOR2_X1 U9946 ( .A1(n8316), .A2(n8315), .ZN(n8317) );
  NOR2_X1 U9947 ( .A1(n8318), .A2(n8317), .ZN(n8320) );
  AOI21_X1 U9948 ( .B1(n8320), .B2(n8413), .A(n8319), .ZN(n8325) );
  INV_X1 U9949 ( .A(n8321), .ZN(n8323) );
  OAI211_X1 U9950 ( .C1(n8325), .C2(n8324), .A(n8323), .B(n8322), .ZN(n8327)
         );
  AOI211_X1 U9951 ( .C1(n4806), .C2(n8327), .A(n5907), .B(n8326), .ZN(n8328)
         );
  NOR2_X1 U9952 ( .A1(n8330), .A2(n8328), .ZN(n8329) );
  MUX2_X1 U9953 ( .A(n8330), .B(n8329), .S(n9430), .Z(n8331) );
  AOI21_X1 U9954 ( .B1(n8333), .B2(n8332), .A(n8331), .ZN(n8335) );
  NOR4_X1 U9955 ( .A1(n8338), .A2(n8337), .A3(n5919), .A4(n8345), .ZN(n8341)
         );
  OAI21_X1 U9956 ( .B1(n8339), .B2(n8342), .A(P1_B_REG_SCAN_IN), .ZN(n8340) );
  OAI22_X1 U9957 ( .A1(n8343), .A2(n8342), .B1(n8341), .B2(n8340), .ZN(
        P1_U3240) );
  INV_X1 U9958 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n8347) );
  INV_X1 U9959 ( .A(n9494), .ZN(n9300) );
  INV_X1 U9960 ( .A(n9509), .ZN(n9347) );
  INV_X1 U9961 ( .A(n9474), .ZN(n9580) );
  NAND2_X1 U9962 ( .A1(n9470), .A2(n9580), .ZN(n9471) );
  NAND2_X1 U9963 ( .A1(n9300), .A2(n9312), .ZN(n9295) );
  XNOR2_X1 U9964 ( .A(n8356), .B(n4502), .ZN(n8352) );
  INV_X1 U9965 ( .A(P1_B_REG_SCAN_IN), .ZN(n8344) );
  NOR2_X1 U9966 ( .A1(n8345), .A2(n8344), .ZN(n8346) );
  NOR2_X1 U9967 ( .A1(n9670), .A2(n8346), .ZN(n9258) );
  AND2_X1 U9968 ( .A1(n9258), .A2(n9200), .ZN(n8359) );
  AOI21_X1 U9969 ( .B1(n8352), .B2(n9960), .A(n8359), .ZN(n8349) );
  MUX2_X1 U9970 ( .A(n8347), .B(n8349), .S(n9992), .Z(n8348) );
  OAI21_X1 U9971 ( .B1(n8356), .B2(n9588), .A(n8348), .ZN(P1_U3521) );
  INV_X1 U9972 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8350) );
  MUX2_X1 U9973 ( .A(n8350), .B(n8349), .S(n10004), .Z(n8351) );
  OAI21_X1 U9974 ( .B1(n8356), .B2(n9551), .A(n8351), .ZN(P1_U3553) );
  NAND2_X1 U9975 ( .A1(n8352), .A2(n9691), .ZN(n8355) );
  INV_X1 U9976 ( .A(n8359), .ZN(n8353) );
  NOR2_X1 U9977 ( .A1(n9678), .A2(n8353), .ZN(n8366) );
  AOI21_X1 U9978 ( .B1(n9709), .B2(P1_REG2_REG_30__SCAN_IN), .A(n8366), .ZN(
        n8354) );
  OAI211_X1 U9979 ( .C1(n8356), .C2(n9475), .A(n8355), .B(n8354), .ZN(P1_U3262) );
  INV_X1 U9980 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8360) );
  XNOR2_X1 U9981 ( .A(n8358), .B(n8357), .ZN(n8365) );
  AOI21_X1 U9982 ( .B1(n8365), .B2(n9960), .A(n8359), .ZN(n8362) );
  MUX2_X1 U9983 ( .A(n8360), .B(n8362), .S(n9992), .Z(n8361) );
  OAI21_X1 U9984 ( .B1(n8369), .B2(n9588), .A(n8361), .ZN(P1_U3522) );
  INV_X1 U9985 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8363) );
  MUX2_X1 U9986 ( .A(n8363), .B(n8362), .S(n10004), .Z(n8364) );
  OAI21_X1 U9987 ( .B1(n8369), .B2(n9551), .A(n8364), .ZN(P1_U3554) );
  NAND2_X1 U9988 ( .A1(n8365), .A2(n9691), .ZN(n8368) );
  AOI21_X1 U9989 ( .B1(n9709), .B2(P1_REG2_REG_31__SCAN_IN), .A(n8366), .ZN(
        n8367) );
  OAI211_X1 U9990 ( .C1(n8369), .C2(n9475), .A(n8368), .B(n8367), .ZN(P1_U3261) );
  NAND2_X1 U9991 ( .A1(n8371), .A2(n8370), .ZN(n8374) );
  NAND2_X1 U9992 ( .A1(n8372), .A2(n9463), .ZN(n8373) );
  NAND2_X1 U9993 ( .A1(n8374), .A2(n8373), .ZN(n9468) );
  OR2_X1 U9994 ( .A1(n9474), .A2(n9443), .ZN(n8375) );
  NAND2_X1 U9995 ( .A1(n9408), .A2(n9202), .ZN(n8380) );
  INV_X1 U9996 ( .A(n8380), .ZN(n8378) );
  OR2_X1 U9997 ( .A1(n9408), .A2(n9202), .ZN(n8376) );
  OR2_X1 U9998 ( .A1(n9431), .A2(n9444), .ZN(n9392) );
  AND2_X1 U9999 ( .A1(n8376), .A2(n9392), .ZN(n8377) );
  NOR2_X1 U10000 ( .A1(n8378), .A2(n8377), .ZN(n8382) );
  OR2_X1 U10001 ( .A1(n9449), .A2(n8382), .ZN(n9383) );
  NAND2_X1 U10002 ( .A1(n9452), .A2(n9464), .ZN(n9432) );
  NAND2_X1 U10003 ( .A1(n9431), .A2(n9444), .ZN(n8379) );
  AND2_X1 U10004 ( .A1(n9432), .A2(n8379), .ZN(n9391) );
  AND2_X1 U10005 ( .A1(n9391), .A2(n8380), .ZN(n8381) );
  OR2_X1 U10006 ( .A1(n8382), .A2(n8381), .ZN(n9384) );
  OR2_X1 U10007 ( .A1(n9514), .A2(n9351), .ZN(n8386) );
  AND2_X1 U10008 ( .A1(n9509), .A2(n9367), .ZN(n8387) );
  NOR2_X1 U10009 ( .A1(n9331), .A2(n9352), .ZN(n8388) );
  NAND2_X1 U10010 ( .A1(n9331), .A2(n9352), .ZN(n8389) );
  OR2_X1 U10011 ( .A1(n9313), .A2(n9327), .ZN(n8390) );
  NAND2_X1 U10012 ( .A1(n9494), .A2(n9287), .ZN(n8391) );
  OAI22_X1 U10013 ( .A1(n9280), .A2(n9285), .B1(n9304), .B2(n9489), .ZN(n8393)
         );
  INV_X1 U10014 ( .A(n8393), .ZN(n8392) );
  NAND2_X1 U10015 ( .A1(n8392), .A2(n8415), .ZN(n9252) );
  NAND2_X1 U10016 ( .A1(n8393), .A2(n8414), .ZN(n8394) );
  NAND2_X1 U10017 ( .A1(n9252), .A2(n8394), .ZN(n9279) );
  AOI21_X2 U10018 ( .B1(n8397), .B2(n8396), .A(n8395), .ZN(n9461) );
  INV_X1 U10019 ( .A(n9449), .ZN(n9438) );
  NOR2_X1 U10020 ( .A1(n9387), .A2(n9401), .ZN(n8401) );
  NOR2_X1 U10021 ( .A1(n9358), .A2(n8402), .ZN(n8403) );
  INV_X1 U10022 ( .A(n9342), .ZN(n9349) );
  INV_X1 U10023 ( .A(n8410), .ZN(n9303) );
  INV_X1 U10024 ( .A(n8414), .ZN(n8415) );
  OAI21_X1 U10025 ( .B1(n4509), .B2(n8416), .A(n9700), .ZN(n8418) );
  AOI22_X1 U10026 ( .A1(n9201), .A2(n9702), .B1(n9304), .B2(n9705), .ZN(n8417)
         );
  AOI21_X1 U10027 ( .B1(n8420), .B2(n9281), .A(n9986), .ZN(n8421) );
  AND2_X1 U10028 ( .A1(n8421), .A2(n9263), .ZN(n9271) );
  OAI21_X1 U10029 ( .B1(n9275), .B2(n9588), .A(n4511), .ZN(P1_U3519) );
  INV_X1 U10030 ( .A(n8424), .ZN(n8425) );
  OAI222_X1 U10031 ( .A1(n8428), .A2(n8427), .B1(n4477), .B2(n8426), .C1(n8618), .C2(P2_U3152), .ZN(P2_U3339) );
  INV_X1 U10032 ( .A(n8433), .ZN(n8435) );
  INV_X1 U10033 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n10340) );
  NOR2_X1 U10034 ( .A1(n8436), .A2(n10340), .ZN(n8431) );
  INV_X1 U10035 ( .A(n8992), .ZN(n8806) );
  AND2_X1 U10036 ( .A1(n8992), .A2(n8703), .ZN(n8444) );
  OAI21_X1 U10037 ( .B1(n8435), .B2(n8806), .A(n8434), .ZN(n8439) );
  INV_X1 U10038 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9082) );
  INV_X1 U10039 ( .A(n8581), .ZN(n8438) );
  INV_X1 U10040 ( .A(n8703), .ZN(n8437) );
  NAND2_X1 U10041 ( .A1(n8806), .A2(n8437), .ZN(n8577) );
  NOR2_X1 U10042 ( .A1(n8987), .A2(n8801), .ZN(n8582) );
  AOI21_X1 U10043 ( .B1(n8439), .B2(n8616), .A(n8582), .ZN(n8440) );
  XNOR2_X1 U10044 ( .A(n8440), .B(n6304), .ZN(n8441) );
  NOR2_X1 U10045 ( .A1(n8582), .A2(n8444), .ZN(n8617) );
  OR3_X1 U10046 ( .A1(n8618), .A2(n8628), .A3(n8443), .ZN(n8580) );
  INV_X1 U10047 ( .A(n8444), .ZN(n8578) );
  INV_X1 U10048 ( .A(n8580), .ZN(n8572) );
  OR3_X1 U10049 ( .A1(n8993), .A2(n8838), .A3(n8572), .ZN(n8570) );
  INV_X1 U10050 ( .A(n8892), .ZN(n8447) );
  INV_X1 U10051 ( .A(n8445), .ZN(n8446) );
  OAI21_X1 U10052 ( .B1(n8447), .B2(n8446), .A(n8572), .ZN(n8548) );
  NAND2_X1 U10053 ( .A1(n9051), .A2(n8448), .ZN(n8449) );
  AND2_X1 U10054 ( .A1(n8584), .A2(n8449), .ZN(n8450) );
  MUX2_X1 U10055 ( .A(n8451), .B(n8450), .S(n8572), .Z(n8528) );
  MUX2_X1 U10056 ( .A(n8453), .B(n8452), .S(n8580), .Z(n8526) );
  MUX2_X1 U10057 ( .A(n8455), .B(n8454), .S(n8580), .Z(n8514) );
  MUX2_X1 U10058 ( .A(n8457), .B(n8456), .S(n8572), .Z(n8480) );
  AND2_X1 U10059 ( .A1(n8459), .A2(n8458), .ZN(n8461) );
  OAI211_X1 U10060 ( .C1(n8480), .C2(n8461), .A(n8485), .B(n8460), .ZN(n8462)
         );
  NAND2_X1 U10061 ( .A1(n8462), .A2(n8580), .ZN(n8470) );
  INV_X1 U10062 ( .A(n8480), .ZN(n8468) );
  AND2_X1 U10063 ( .A1(n8633), .A2(n8622), .ZN(n8463) );
  OAI211_X1 U10064 ( .C1(n8464), .C2(n8463), .A(n8474), .B(n8471), .ZN(n8465)
         );
  NAND3_X1 U10065 ( .A1(n8465), .A2(n8473), .A3(n8580), .ZN(n8466) );
  NAND3_X1 U10066 ( .A1(n8468), .A2(n8467), .A3(n8466), .ZN(n8469) );
  NAND2_X1 U10067 ( .A1(n8471), .A2(n8633), .ZN(n8472) );
  NAND3_X1 U10068 ( .A1(n6554), .A2(n8473), .A3(n8472), .ZN(n8475) );
  NAND3_X1 U10069 ( .A1(n8475), .A2(n8572), .A3(n8474), .ZN(n8476) );
  AOI22_X1 U10070 ( .A1(n8480), .A2(n8479), .B1(n8478), .B2(n8477), .ZN(n8483)
         );
  INV_X1 U10071 ( .A(n8481), .ZN(n8482) );
  OAI21_X1 U10072 ( .B1(n8483), .B2(n8482), .A(n8572), .ZN(n8484) );
  MUX2_X1 U10073 ( .A(n8487), .B(n8486), .S(n8580), .Z(n8488) );
  NAND3_X1 U10074 ( .A1(n8489), .A2(n8596), .A3(n8488), .ZN(n8496) );
  INV_X1 U10075 ( .A(n8490), .ZN(n8493) );
  NAND2_X1 U10076 ( .A1(n8497), .A2(n8491), .ZN(n8492) );
  MUX2_X1 U10077 ( .A(n8493), .B(n8492), .S(n8580), .Z(n8494) );
  INV_X1 U10078 ( .A(n8494), .ZN(n8495) );
  NAND3_X1 U10079 ( .A1(n8496), .A2(n8500), .A3(n8495), .ZN(n8502) );
  NAND3_X1 U10080 ( .A1(n8502), .A2(n8503), .A3(n8497), .ZN(n8499) );
  NAND3_X1 U10081 ( .A1(n8502), .A2(n8501), .A3(n8500), .ZN(n8504) );
  NAND2_X1 U10082 ( .A1(n8511), .A2(n8505), .ZN(n8507) );
  MUX2_X1 U10083 ( .A(n8507), .B(n4577), .S(n8580), .Z(n8508) );
  INV_X1 U10084 ( .A(n8508), .ZN(n8509) );
  MUX2_X1 U10085 ( .A(n8511), .B(n8510), .S(n8572), .Z(n8512) );
  NAND3_X1 U10086 ( .A1(n8514), .A2(n8513), .A3(n5018), .ZN(n8518) );
  MUX2_X1 U10087 ( .A(n8516), .B(n8515), .S(n8580), .Z(n8517) );
  AND3_X1 U10088 ( .A1(n8519), .A2(n8518), .A3(n8517), .ZN(n8524) );
  MUX2_X1 U10089 ( .A(n5008), .B(n8521), .S(n8572), .Z(n8523) );
  OAI21_X1 U10090 ( .B1(n8524), .B2(n8523), .A(n8522), .ZN(n8525) );
  NAND3_X1 U10091 ( .A1(n8607), .A2(n8526), .A3(n8525), .ZN(n8527) );
  NAND2_X1 U10092 ( .A1(n8528), .A2(n8527), .ZN(n8534) );
  NAND2_X1 U10093 ( .A1(n8534), .A2(n8584), .ZN(n8529) );
  NAND3_X1 U10094 ( .A1(n8529), .A2(n8536), .A3(n8533), .ZN(n8530) );
  NAND3_X1 U10095 ( .A1(n8530), .A2(n8539), .A3(n8950), .ZN(n8531) );
  OR2_X1 U10096 ( .A1(n9030), .A2(n8959), .ZN(n8540) );
  NAND3_X1 U10097 ( .A1(n8531), .A2(n8537), .A3(n8540), .ZN(n8532) );
  NAND3_X1 U10098 ( .A1(n8541), .A2(n8532), .A3(n8538), .ZN(n8544) );
  NAND2_X1 U10099 ( .A1(n8534), .A2(n8533), .ZN(n8535) );
  AND2_X1 U10100 ( .A1(n8542), .A2(n8541), .ZN(n8543) );
  MUX2_X1 U10101 ( .A(n8544), .B(n8543), .S(n8572), .Z(n8545) );
  OAI211_X1 U10102 ( .C1(n8572), .C2(n8546), .A(n8545), .B(n6571), .ZN(n8547)
         );
  NAND2_X1 U10103 ( .A1(n8548), .A2(n8547), .ZN(n8552) );
  AOI21_X1 U10104 ( .B1(n8551), .B2(n8549), .A(n8572), .ZN(n8550) );
  OAI21_X1 U10105 ( .B1(n8572), .B2(n8553), .A(n8872), .ZN(n8559) );
  AND2_X1 U10106 ( .A1(n9011), .A2(n8695), .ZN(n8555) );
  NAND2_X1 U10107 ( .A1(n8560), .A2(n8572), .ZN(n8554) );
  OAI21_X1 U10108 ( .B1(n8854), .B2(n8555), .A(n8554), .ZN(n8558) );
  INV_X1 U10109 ( .A(n8556), .ZN(n8855) );
  NAND2_X1 U10110 ( .A1(n8855), .A2(n8572), .ZN(n8557) );
  MUX2_X1 U10111 ( .A(n8561), .B(n8560), .S(n8580), .Z(n8562) );
  NAND2_X1 U10112 ( .A1(n8999), .A2(n8821), .ZN(n8566) );
  INV_X1 U10113 ( .A(n8564), .ZN(n8565) );
  MUX2_X1 U10114 ( .A(n8566), .B(n8565), .S(n8572), .Z(n8567) );
  NAND3_X1 U10115 ( .A1(n8993), .A2(n8838), .A3(n8572), .ZN(n8568) );
  NAND4_X1 U10116 ( .A1(n8571), .A2(n8570), .A3(n8569), .A4(n8568), .ZN(n8576)
         );
  MUX2_X1 U10117 ( .A(n8574), .B(n8573), .S(n8572), .Z(n8575) );
  NAND4_X1 U10118 ( .A1(n8578), .A2(n8577), .A3(n8576), .A4(n8575), .ZN(n8579)
         );
  MUX2_X1 U10119 ( .A(n8582), .B(n8581), .S(n8580), .Z(n8583) );
  INV_X1 U10120 ( .A(n8872), .ZN(n8864) );
  INV_X1 U10121 ( .A(n8584), .ZN(n8585) );
  NOR2_X1 U10122 ( .A1(n8586), .A2(n8585), .ZN(n8980) );
  INV_X1 U10123 ( .A(n8587), .ZN(n8621) );
  NAND4_X1 U10124 ( .A1(n8589), .A2(n8621), .A3(n6555), .A4(n8633), .ZN(n8593)
         );
  NOR4_X1 U10125 ( .A1(n8593), .A2(n8592), .A3(n8591), .A4(n8590), .ZN(n8597)
         );
  NAND4_X1 U10126 ( .A1(n8597), .A2(n8596), .A3(n8595), .A4(n8594), .ZN(n8599)
         );
  NOR4_X1 U10127 ( .A1(n8601), .A2(n8600), .A3(n8599), .A4(n8598), .ZN(n8602)
         );
  NAND3_X1 U10128 ( .A1(n6564), .A2(n8603), .A3(n8602), .ZN(n8604) );
  NOR4_X1 U10129 ( .A1(n6537), .A2(n8606), .A3(n8605), .A4(n8604), .ZN(n8608)
         );
  NAND4_X1 U10130 ( .A1(n8609), .A2(n8980), .A3(n8608), .A4(n8607), .ZN(n8610)
         );
  NOR4_X1 U10131 ( .A1(n8903), .A2(n8922), .A3(n8955), .A4(n8610), .ZN(n8612)
         );
  NAND4_X1 U10132 ( .A1(n8844), .A2(n8892), .A3(n8612), .A4(n6570), .ZN(n8613)
         );
  NOR4_X1 U10133 ( .A1(n8614), .A2(n8864), .A3(n8836), .A4(n8613), .ZN(n8615)
         );
  NAND4_X1 U10134 ( .A1(n8617), .A2(n8616), .A3(n8615), .A4(n8810), .ZN(n8619)
         );
  XNOR2_X1 U10135 ( .A(n8619), .B(n8618), .ZN(n8623) );
  OAI22_X1 U10136 ( .A1(n8623), .A2(n8622), .B1(n8621), .B2(n8620), .ZN(n8624)
         );
  NOR4_X1 U10137 ( .A1(n10019), .A2(n8627), .A3(n8626), .A4(n8956), .ZN(n8630)
         );
  OAI21_X1 U10138 ( .B1(n8631), .B2(n8628), .A(P2_B_REG_SCAN_IN), .ZN(n8629)
         );
  OAI22_X1 U10139 ( .A1(n4536), .A2(n8631), .B1(n8630), .B2(n8629), .ZN(
        P2_U3244) );
  NOR2_X1 U10140 ( .A1(n8692), .A2(n8632), .ZN(n8637) );
  MUX2_X1 U10141 ( .A(n8633), .B(n8632), .S(n10035), .Z(n8634) );
  AOI21_X1 U10142 ( .B1(n8635), .B2(n8634), .A(n8701), .ZN(n8636) );
  AOI211_X1 U10143 ( .C1(P2_REG3_REG_0__SCAN_IN), .C2(n8638), .A(n8637), .B(
        n8636), .ZN(n8639) );
  OAI21_X1 U10144 ( .B1(n6514), .B2(n8687), .A(n8639), .ZN(P2_U3234) );
  OAI222_X1 U10145 ( .A1(n9087), .A2(n10340), .B1(n4477), .B2(n8641), .C1(
        n8640), .C2(P2_U3152), .ZN(P2_U3328) );
  XNOR2_X1 U10146 ( .A(n8643), .B(n8642), .ZN(n8647) );
  OAI22_X1 U10147 ( .A1(n8698), .A2(n8830), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10322), .ZN(n8645) );
  OAI22_X1 U10148 ( .A1(n8838), .A2(n8687), .B1(n8686), .B2(n8837), .ZN(n8644)
         );
  AOI211_X1 U10149 ( .C1(n8999), .C2(n6494), .A(n8645), .B(n8644), .ZN(n8646)
         );
  OAI21_X1 U10150 ( .B1(n8647), .B2(n8701), .A(n8646), .ZN(P2_U3216) );
  OAI211_X1 U10151 ( .C1(n8648), .C2(n8650), .A(n8649), .B(n9628), .ZN(n8655)
         );
  OAI22_X1 U10152 ( .A1(n8698), .A2(n8908), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8651), .ZN(n8653) );
  OAI22_X1 U10153 ( .A1(n8669), .A2(n8687), .B1(n8686), .B2(n8660), .ZN(n8652)
         );
  AOI211_X1 U10154 ( .C1(n9020), .C2(n6494), .A(n8653), .B(n8652), .ZN(n8654)
         );
  NAND2_X1 U10155 ( .A1(n8655), .A2(n8654), .ZN(P2_U3218) );
  OAI211_X1 U10156 ( .C1(n8658), .C2(n8657), .A(n8656), .B(n9628), .ZN(n8664)
         );
  OAI22_X1 U10157 ( .A1(n8698), .A2(n8932), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10390), .ZN(n8662) );
  OAI22_X1 U10158 ( .A1(n8660), .A2(n8687), .B1(n8686), .B2(n8659), .ZN(n8661)
         );
  AOI211_X1 U10159 ( .C1(n9030), .C2(n6494), .A(n8662), .B(n8661), .ZN(n8663)
         );
  NAND2_X1 U10160 ( .A1(n8664), .A2(n8663), .ZN(P2_U3225) );
  NOR2_X1 U10161 ( .A1(n4720), .A2(n8666), .ZN(n8667) );
  XNOR2_X1 U10162 ( .A(n8668), .B(n8667), .ZN(n8673) );
  OAI22_X1 U10163 ( .A1(n8669), .A2(n8956), .B1(n8837), .B2(n8958), .ZN(n8874)
         );
  AOI22_X1 U10164 ( .A1(n8696), .A2(n8874), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8670) );
  OAI21_X1 U10165 ( .B1(n8868), .B2(n8698), .A(n8670), .ZN(n8671) );
  AOI21_X1 U10166 ( .B1(n9011), .B2(n6494), .A(n8671), .ZN(n8672) );
  OAI21_X1 U10167 ( .B1(n8673), .B2(n8701), .A(n8672), .ZN(P2_U3227) );
  OAI211_X1 U10168 ( .C1(n8676), .C2(n8675), .A(n8674), .B(n9628), .ZN(n8681)
         );
  OAI22_X1 U10169 ( .A1(n8698), .A2(n8886), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8677), .ZN(n8679) );
  OAI22_X1 U10170 ( .A1(n8924), .A2(n8686), .B1(n8687), .B2(n8695), .ZN(n8678)
         );
  AOI211_X1 U10171 ( .C1(n9014), .C2(n6494), .A(n8679), .B(n8678), .ZN(n8680)
         );
  NAND2_X1 U10172 ( .A1(n8681), .A2(n8680), .ZN(P2_U3231) );
  OAI21_X1 U10173 ( .B1(n8684), .B2(n8683), .A(n8682), .ZN(n8685) );
  NAND2_X1 U10174 ( .A1(n8685), .A2(n9628), .ZN(n8691) );
  NOR2_X1 U10175 ( .A1(n8698), .A2(n8918), .ZN(n8689) );
  OAI22_X1 U10176 ( .A1(n8924), .A2(n8687), .B1(n8686), .B2(n8959), .ZN(n8688)
         );
  AOI211_X1 U10177 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3152), .A(n8689), 
        .B(n8688), .ZN(n8690) );
  OAI211_X1 U10178 ( .C1(n8921), .C2(n8692), .A(n8691), .B(n8690), .ZN(
        P2_U3237) );
  XNOR2_X1 U10179 ( .A(n8693), .B(n8694), .ZN(n8702) );
  OAI22_X1 U10180 ( .A1(n8695), .A2(n8956), .B1(n8821), .B2(n8958), .ZN(n8859)
         );
  AOI22_X1 U10181 ( .A1(n8696), .A2(n8859), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8697) );
  OAI21_X1 U10182 ( .B1(n8849), .B2(n8698), .A(n8697), .ZN(n8699) );
  AOI21_X1 U10183 ( .B1(n9005), .B2(n6494), .A(n8699), .ZN(n8700) );
  OAI21_X1 U10184 ( .B1(n8702), .B2(n8701), .A(n8700), .ZN(P2_U3242) );
  MUX2_X1 U10185 ( .A(n8703), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8724), .Z(
        P2_U3582) );
  MUX2_X1 U10186 ( .A(n8704), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8724), .Z(
        P2_U3581) );
  MUX2_X1 U10187 ( .A(n8705), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8724), .Z(
        P2_U3580) );
  MUX2_X1 U10188 ( .A(n8706), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8724), .Z(
        P2_U3579) );
  MUX2_X1 U10189 ( .A(n8707), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8724), .Z(
        P2_U3578) );
  MUX2_X1 U10190 ( .A(n8882), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8724), .Z(
        P2_U3577) );
  MUX2_X1 U10191 ( .A(n8900), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8724), .Z(
        P2_U3576) );
  MUX2_X1 U10192 ( .A(n8883), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8724), .Z(
        P2_U3575) );
  MUX2_X1 U10193 ( .A(n8938), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8724), .Z(
        P2_U3574) );
  MUX2_X1 U10194 ( .A(n8708), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8724), .Z(
        P2_U3573) );
  MUX2_X1 U10195 ( .A(n8939), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8724), .Z(
        P2_U3572) );
  MUX2_X1 U10196 ( .A(n8969), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8724), .Z(
        P2_U3571) );
  MUX2_X1 U10197 ( .A(n8709), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8724), .Z(
        P2_U3570) );
  MUX2_X1 U10198 ( .A(n8967), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8724), .Z(
        P2_U3569) );
  MUX2_X1 U10199 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8710), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10200 ( .A(n8711), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8724), .Z(
        P2_U3567) );
  MUX2_X1 U10201 ( .A(n8712), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8724), .Z(
        P2_U3566) );
  MUX2_X1 U10202 ( .A(n8713), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8724), .Z(
        P2_U3565) );
  MUX2_X1 U10203 ( .A(n8714), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8724), .Z(
        P2_U3564) );
  MUX2_X1 U10204 ( .A(n8715), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8724), .Z(
        P2_U3563) );
  MUX2_X1 U10205 ( .A(n8716), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8724), .Z(
        P2_U3562) );
  MUX2_X1 U10206 ( .A(n8717), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8724), .Z(
        P2_U3561) );
  MUX2_X1 U10207 ( .A(n8718), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8724), .Z(
        P2_U3560) );
  MUX2_X1 U10208 ( .A(n8719), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8724), .Z(
        P2_U3559) );
  MUX2_X1 U10209 ( .A(n8720), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8724), .Z(
        P2_U3558) );
  MUX2_X1 U10210 ( .A(n8721), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8724), .Z(
        P2_U3557) );
  MUX2_X1 U10211 ( .A(n8722), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8724), .Z(
        P2_U3556) );
  MUX2_X1 U10212 ( .A(n8723), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8724), .Z(
        P2_U3555) );
  MUX2_X1 U10213 ( .A(n6517), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8724), .Z(
        P2_U3554) );
  MUX2_X1 U10214 ( .A(n4480), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8724), .Z(
        P2_U3553) );
  OAI21_X1 U10215 ( .B1(n8727), .B2(n8726), .A(n8725), .ZN(n8728) );
  NAND2_X1 U10216 ( .A1(n10011), .A2(n8728), .ZN(n8738) );
  NOR2_X1 U10217 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8729), .ZN(n8730) );
  AOI21_X1 U10218 ( .B1(n10013), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8730), .ZN(
        n8737) );
  NAND2_X1 U10219 ( .A1(n9618), .A2(n8731), .ZN(n8736) );
  OAI211_X1 U10220 ( .C1(n8734), .C2(n8733), .A(n10010), .B(n8732), .ZN(n8735)
         );
  NAND4_X1 U10221 ( .A1(n8738), .A2(n8737), .A3(n8736), .A4(n8735), .ZN(
        P2_U3256) );
  OAI21_X1 U10222 ( .B1(n8740), .B2(n7813), .A(n8739), .ZN(n8741) );
  NAND2_X1 U10223 ( .A1(n8741), .A2(n10011), .ZN(n8750) );
  NOR2_X1 U10224 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8742), .ZN(n8743) );
  AOI21_X1 U10225 ( .B1(n10013), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8743), .ZN(
        n8749) );
  OAI211_X1 U10226 ( .C1(n8745), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10010), .B(
        n8744), .ZN(n8748) );
  NAND2_X1 U10227 ( .A1(n9618), .A2(n8746), .ZN(n8747) );
  NAND4_X1 U10228 ( .A1(n8750), .A2(n8749), .A3(n8748), .A4(n8747), .ZN(
        P2_U3260) );
  NAND2_X1 U10229 ( .A1(n8753), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8768) );
  OAI21_X1 U10230 ( .B1(n8753), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8768), .ZN(
        n8754) );
  AOI211_X1 U10231 ( .C1(n8755), .C2(n8754), .A(n8766), .B(n9612), .ZN(n8765)
         );
  NOR2_X1 U10232 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10279), .ZN(n8756) );
  AOI21_X1 U10233 ( .B1(n10013), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8756), .ZN(
        n8763) );
  INV_X1 U10234 ( .A(n8757), .ZN(n8759) );
  AOI21_X1 U10235 ( .B1(n8759), .B2(n8017), .A(n8758), .ZN(n8761) );
  XNOR2_X1 U10236 ( .A(n8777), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8760) );
  NAND2_X1 U10237 ( .A1(n8760), .A2(n8761), .ZN(n8776) );
  OAI211_X1 U10238 ( .C1(n8761), .C2(n8760), .A(n10010), .B(n8776), .ZN(n8762)
         );
  OAI211_X1 U10239 ( .C1(n10005), .C2(n8777), .A(n8763), .B(n8762), .ZN(n8764)
         );
  OR2_X1 U10240 ( .A1(n8765), .A2(n8764), .ZN(P2_U3262) );
  INV_X1 U10241 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8771) );
  INV_X1 U10242 ( .A(n8766), .ZN(n8767) );
  NAND2_X1 U10243 ( .A1(n8768), .A2(n8767), .ZN(n8769) );
  AOI211_X1 U10244 ( .C1(n8771), .C2(n8770), .A(n4518), .B(n9612), .ZN(n8772)
         );
  INV_X1 U10245 ( .A(n8772), .ZN(n8787) );
  INV_X1 U10246 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8773) );
  NAND2_X1 U10247 ( .A1(n8788), .A2(n8773), .ZN(n8790) );
  NAND2_X1 U10248 ( .A1(n8774), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8775) );
  NAND2_X1 U10249 ( .A1(n8790), .A2(n8775), .ZN(n8780) );
  OAI21_X1 U10250 ( .B1(n8778), .B2(n8777), .A(n8776), .ZN(n8779) );
  OR2_X1 U10251 ( .A1(n8780), .A2(n8779), .ZN(n8791) );
  NAND2_X1 U10252 ( .A1(n8780), .A2(n8779), .ZN(n8781) );
  NAND2_X1 U10253 ( .A1(n8791), .A2(n8781), .ZN(n8785) );
  INV_X1 U10254 ( .A(n8782), .ZN(n8783) );
  OAI21_X1 U10255 ( .B1(n8799), .B2(n10510), .A(n8783), .ZN(n8784) );
  AOI21_X1 U10256 ( .B1(n10010), .B2(n8785), .A(n8784), .ZN(n8786) );
  OAI211_X1 U10257 ( .C1(n10005), .C2(n8788), .A(n8787), .B(n8786), .ZN(
        P2_U3263) );
  XNOR2_X1 U10258 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8789), .ZN(n8795) );
  NAND2_X1 U10259 ( .A1(n8791), .A2(n8790), .ZN(n8793) );
  XNOR2_X1 U10260 ( .A(n8793), .B(n8792), .ZN(n8796) );
  INV_X1 U10261 ( .A(n8796), .ZN(n8794) );
  AOI22_X1 U10262 ( .A1(n8795), .A2(n10011), .B1(n8794), .B2(n10010), .ZN(
        n8797) );
  NAND2_X1 U10263 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8798) );
  NAND2_X1 U10264 ( .A1(n8992), .A2(n8804), .ZN(n8988) );
  NAND2_X1 U10265 ( .A1(n8986), .A2(n8984), .ZN(n8803) );
  NAND2_X1 U10266 ( .A1(n8801), .A2(n8800), .ZN(n8990) );
  NOR2_X1 U10267 ( .A1(n4476), .A2(n8990), .ZN(n8807) );
  AOI21_X1 U10268 ( .B1(n4476), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8807), .ZN(
        n8802) );
  OAI211_X1 U10269 ( .C1(n8987), .C2(n8977), .A(n8803), .B(n8802), .ZN(
        P2_U3265) );
  INV_X1 U10270 ( .A(n8804), .ZN(n8805) );
  NAND2_X1 U10271 ( .A1(n8806), .A2(n8805), .ZN(n8989) );
  NAND3_X1 U10272 ( .A1(n8989), .A2(n8984), .A3(n8988), .ZN(n8809) );
  AOI21_X1 U10273 ( .B1(n4476), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8807), .ZN(
        n8808) );
  OAI211_X1 U10274 ( .C1(n8992), .C2(n8977), .A(n8809), .B(n8808), .ZN(
        P2_U3266) );
  XNOR2_X1 U10275 ( .A(n8811), .B(n8810), .ZN(n8998) );
  INV_X1 U10276 ( .A(n8829), .ZN(n8814) );
  INV_X1 U10277 ( .A(n8812), .ZN(n8813) );
  AOI21_X1 U10278 ( .B1(n8993), .B2(n8814), .A(n8813), .ZN(n8994) );
  AOI22_X1 U10279 ( .A1(n4476), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8815), .B2(
        n8974), .ZN(n8816) );
  OAI21_X1 U10280 ( .B1(n8817), .B2(n8977), .A(n8816), .ZN(n8826) );
  AOI211_X1 U10281 ( .C1(n8820), .C2(n8819), .A(n8953), .B(n8818), .ZN(n8824)
         );
  OAI22_X1 U10282 ( .A1(n8822), .A2(n8958), .B1(n8821), .B2(n8956), .ZN(n8823)
         );
  NOR2_X1 U10283 ( .A1(n8824), .A2(n8823), .ZN(n8996) );
  NOR2_X1 U10284 ( .A1(n8996), .A2(n4476), .ZN(n8825) );
  AOI211_X1 U10285 ( .C1(n8994), .C2(n8984), .A(n8826), .B(n8825), .ZN(n8827)
         );
  OAI21_X1 U10286 ( .B1(n8998), .B2(n8981), .A(n8827), .ZN(P2_U3268) );
  XNOR2_X1 U10287 ( .A(n8828), .B(n8836), .ZN(n9003) );
  AOI21_X1 U10288 ( .B1(n8999), .B2(n8846), .A(n8829), .ZN(n9000) );
  INV_X1 U10289 ( .A(n8999), .ZN(n8833) );
  INV_X1 U10290 ( .A(n8830), .ZN(n8831) );
  AOI22_X1 U10291 ( .A1(n4476), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8831), .B2(
        n8974), .ZN(n8832) );
  OAI21_X1 U10292 ( .B1(n8833), .B2(n8977), .A(n8832), .ZN(n8842) );
  AOI211_X1 U10293 ( .C1(n8836), .C2(n8835), .A(n8953), .B(n8834), .ZN(n8840)
         );
  OAI22_X1 U10294 ( .A1(n8838), .A2(n8958), .B1(n8837), .B2(n8956), .ZN(n8839)
         );
  NOR2_X1 U10295 ( .A1(n8840), .A2(n8839), .ZN(n9002) );
  NOR2_X1 U10296 ( .A1(n9002), .A2(n4476), .ZN(n8841) );
  AOI211_X1 U10297 ( .C1(n9000), .C2(n8984), .A(n8842), .B(n8841), .ZN(n8843)
         );
  OAI21_X1 U10298 ( .B1(n9003), .B2(n8981), .A(n8843), .ZN(P2_U3269) );
  XNOR2_X1 U10299 ( .A(n8845), .B(n8844), .ZN(n9008) );
  INV_X1 U10300 ( .A(n8866), .ZN(n8848) );
  INV_X1 U10301 ( .A(n8846), .ZN(n8847) );
  AOI211_X1 U10302 ( .C1(n9005), .C2(n8848), .A(n10078), .B(n8847), .ZN(n9004)
         );
  INV_X1 U10303 ( .A(n8849), .ZN(n8850) );
  AOI22_X1 U10304 ( .A1(n4476), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8850), .B2(
        n8974), .ZN(n8851) );
  OAI21_X1 U10305 ( .B1(n8852), .B2(n8977), .A(n8851), .ZN(n8862) );
  INV_X1 U10306 ( .A(n8853), .ZN(n8856) );
  OAI21_X1 U10307 ( .B1(n8856), .B2(n8855), .A(n8854), .ZN(n8858) );
  AOI21_X1 U10308 ( .B1(n8858), .B2(n8857), .A(n8953), .ZN(n8860) );
  NOR2_X1 U10309 ( .A1(n8860), .A2(n8859), .ZN(n9007) );
  NOR2_X1 U10310 ( .A1(n9007), .A2(n4476), .ZN(n8861) );
  AOI211_X1 U10311 ( .C1(n9004), .C2(n8871), .A(n8862), .B(n8861), .ZN(n8863)
         );
  OAI21_X1 U10312 ( .B1(n9008), .B2(n8981), .A(n8863), .ZN(P2_U3270) );
  XNOR2_X1 U10313 ( .A(n8865), .B(n8864), .ZN(n9013) );
  AOI211_X1 U10314 ( .C1(n9011), .C2(n8867), .A(n10078), .B(n8866), .ZN(n9010)
         );
  NOR2_X1 U10315 ( .A1(n4923), .A2(n8977), .ZN(n8870) );
  OAI22_X1 U10316 ( .A1(n8877), .A2(n10243), .B1(n8868), .B2(n8907), .ZN(n8869) );
  AOI211_X1 U10317 ( .C1(n9010), .C2(n8871), .A(n8870), .B(n8869), .ZN(n8879)
         );
  OAI211_X1 U10318 ( .C1(n8873), .C2(n8872), .A(n8853), .B(n8971), .ZN(n8876)
         );
  INV_X1 U10319 ( .A(n8874), .ZN(n8875) );
  NAND2_X1 U10320 ( .A1(n8876), .A2(n8875), .ZN(n9009) );
  NAND2_X1 U10321 ( .A1(n9009), .A2(n8877), .ZN(n8878) );
  OAI211_X1 U10322 ( .C1(n9013), .C2(n8981), .A(n8879), .B(n8878), .ZN(
        P2_U3271) );
  OAI211_X1 U10323 ( .C1(n8892), .C2(n8881), .A(n8880), .B(n8971), .ZN(n8885)
         );
  AOI22_X1 U10324 ( .A1(n8966), .A2(n8883), .B1(n8882), .B2(n8968), .ZN(n8884)
         );
  XNOR2_X1 U10325 ( .A(n4541), .B(n9014), .ZN(n9015) );
  INV_X1 U10326 ( .A(n8886), .ZN(n8887) );
  AOI22_X1 U10327 ( .A1(n4476), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8887), .B2(
        n8974), .ZN(n8888) );
  OAI21_X1 U10328 ( .B1(n8889), .B2(n8977), .A(n8888), .ZN(n8894) );
  AOI21_X1 U10329 ( .B1(n8892), .B2(n8891), .A(n8890), .ZN(n9018) );
  NOR2_X1 U10330 ( .A1(n9018), .A2(n8981), .ZN(n8893) );
  AOI211_X1 U10331 ( .C1(n9015), .C2(n8984), .A(n8894), .B(n8893), .ZN(n8895)
         );
  OAI21_X1 U10332 ( .B1(n4476), .B2(n9017), .A(n8895), .ZN(P2_U3272) );
  NAND2_X1 U10333 ( .A1(n8897), .A2(n8903), .ZN(n8898) );
  NAND2_X1 U10334 ( .A1(n8896), .A2(n8898), .ZN(n8899) );
  NAND2_X1 U10335 ( .A1(n8899), .A2(n8971), .ZN(n8902) );
  AOI22_X1 U10336 ( .A1(n8968), .A2(n8900), .B1(n8938), .B2(n8966), .ZN(n8901)
         );
  OR2_X1 U10337 ( .A1(n8904), .A2(n8903), .ZN(n9019) );
  NAND3_X1 U10338 ( .A1(n9019), .A2(n8905), .A3(n8906), .ZN(n8913) );
  AOI21_X1 U10339 ( .B1(n9020), .B2(n8915), .A(n4541), .ZN(n9021) );
  NOR2_X1 U10340 ( .A1(n4655), .A2(n8977), .ZN(n8911) );
  OAI22_X1 U10341 ( .A1(n8877), .A2(n8909), .B1(n8908), .B2(n8907), .ZN(n8910)
         );
  AOI211_X1 U10342 ( .C1(n9021), .C2(n8984), .A(n8911), .B(n8910), .ZN(n8912)
         );
  OAI211_X1 U10343 ( .C1(n4476), .C2(n9023), .A(n8913), .B(n8912), .ZN(
        P2_U3273) );
  XOR2_X1 U10344 ( .A(n8914), .B(n8922), .Z(n9029) );
  INV_X1 U10345 ( .A(n8915), .ZN(n8916) );
  AOI21_X1 U10346 ( .B1(n9025), .B2(n8917), .A(n8916), .ZN(n9026) );
  INV_X1 U10347 ( .A(n8918), .ZN(n8919) );
  AOI22_X1 U10348 ( .A1(n4476), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8919), .B2(
        n8974), .ZN(n8920) );
  OAI21_X1 U10349 ( .B1(n8921), .B2(n8977), .A(n8920), .ZN(n8929) );
  AOI21_X1 U10350 ( .B1(n8923), .B2(n8922), .A(n8953), .ZN(n8927) );
  OAI22_X1 U10351 ( .A1(n8924), .A2(n8958), .B1(n8959), .B2(n8956), .ZN(n8925)
         );
  AOI21_X1 U10352 ( .B1(n8927), .B2(n8926), .A(n8925), .ZN(n9028) );
  NOR2_X1 U10353 ( .A1(n9028), .A2(n4476), .ZN(n8928) );
  AOI211_X1 U10354 ( .C1(n9026), .C2(n8984), .A(n8929), .B(n8928), .ZN(n8930)
         );
  OAI21_X1 U10355 ( .B1(n9029), .B2(n8981), .A(n8930), .ZN(P2_U3274) );
  XNOR2_X1 U10356 ( .A(n8931), .B(n6570), .ZN(n9034) );
  XNOR2_X1 U10357 ( .A(n8945), .B(n9030), .ZN(n9031) );
  INV_X1 U10358 ( .A(n8932), .ZN(n8933) );
  AOI22_X1 U10359 ( .A1(n4476), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8933), .B2(
        n8974), .ZN(n8934) );
  OAI21_X1 U10360 ( .B1(n8935), .B2(n8977), .A(n8934), .ZN(n8942) );
  OAI21_X1 U10361 ( .B1(n8937), .B2(n6570), .A(n8936), .ZN(n8940) );
  AOI222_X1 U10362 ( .A1(n8971), .A2(n8940), .B1(n8939), .B2(n8966), .C1(n8938), .C2(n8968), .ZN(n9033) );
  NOR2_X1 U10363 ( .A1(n9033), .A2(n4476), .ZN(n8941) );
  AOI211_X1 U10364 ( .C1(n9031), .C2(n8984), .A(n8942), .B(n8941), .ZN(n8943)
         );
  OAI21_X1 U10365 ( .B1(n9034), .B2(n8981), .A(n8943), .ZN(P2_U3275) );
  XNOR2_X1 U10366 ( .A(n8944), .B(n8955), .ZN(n9039) );
  AOI21_X1 U10367 ( .B1(n9035), .B2(n8946), .A(n8945), .ZN(n9036) );
  AOI22_X1 U10368 ( .A1(n4476), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8947), .B2(
        n8974), .ZN(n8948) );
  OAI21_X1 U10369 ( .B1(n8949), .B2(n8977), .A(n8948), .ZN(n8963) );
  NAND2_X1 U10370 ( .A1(n8951), .A2(n8950), .ZN(n8954) );
  AOI211_X1 U10371 ( .C1(n8955), .C2(n8954), .A(n8953), .B(n5026), .ZN(n8961)
         );
  OAI22_X1 U10372 ( .A1(n8959), .A2(n8958), .B1(n8957), .B2(n8956), .ZN(n8960)
         );
  NOR2_X1 U10373 ( .A1(n8961), .A2(n8960), .ZN(n9038) );
  NOR2_X1 U10374 ( .A1(n9038), .A2(n4476), .ZN(n8962) );
  AOI211_X1 U10375 ( .C1(n9036), .C2(n8984), .A(n8963), .B(n8962), .ZN(n8964)
         );
  OAI21_X1 U10376 ( .B1(n9039), .B2(n8981), .A(n8964), .ZN(P2_U3276) );
  XOR2_X1 U10377 ( .A(n8980), .B(n8965), .Z(n8970) );
  AOI222_X1 U10378 ( .A1(n8971), .A2(n8970), .B1(n8969), .B2(n8968), .C1(n8967), .C2(n8966), .ZN(n9048) );
  AND2_X1 U10379 ( .A1(n9045), .A2(n4483), .ZN(n8972) );
  NOR2_X1 U10380 ( .A1(n8973), .A2(n8972), .ZN(n9046) );
  AOI22_X1 U10381 ( .A1(n4476), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8975), .B2(
        n8974), .ZN(n8976) );
  OAI21_X1 U10382 ( .B1(n8978), .B2(n8977), .A(n8976), .ZN(n8983) );
  XOR2_X1 U10383 ( .A(n8980), .B(n8979), .Z(n9049) );
  NOR2_X1 U10384 ( .A1(n9049), .A2(n8981), .ZN(n8982) );
  AOI211_X1 U10385 ( .C1(n9046), .C2(n8984), .A(n8983), .B(n8982), .ZN(n8985)
         );
  OAI21_X1 U10386 ( .B1(n4476), .B2(n9048), .A(n8985), .ZN(P2_U3278) );
  MUX2_X1 U10387 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9064), .S(n10098), .Z(
        P2_U3551) );
  NAND3_X1 U10388 ( .A1(n8989), .A2(n10035), .A3(n8988), .ZN(n8991) );
  OAI211_X1 U10389 ( .C1(n8992), .C2(n10076), .A(n8991), .B(n8990), .ZN(n9065)
         );
  MUX2_X1 U10390 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9065), .S(n10098), .Z(
        P2_U3550) );
  AOI22_X1 U10391 ( .A1(n8994), .A2(n10035), .B1(n9058), .B2(n8993), .ZN(n8995) );
  OAI21_X1 U10392 ( .B1(n8998), .B2(n9054), .A(n8997), .ZN(n9066) );
  MUX2_X1 U10393 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9066), .S(n10098), .Z(
        P2_U3548) );
  AOI22_X1 U10394 ( .A1(n9000), .A2(n10035), .B1(n9058), .B2(n8999), .ZN(n9001) );
  OAI211_X1 U10395 ( .C1(n9003), .C2(n9054), .A(n9002), .B(n9001), .ZN(n9067)
         );
  MUX2_X1 U10396 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9067), .S(n10098), .Z(
        P2_U3547) );
  AOI21_X1 U10397 ( .B1(n9058), .B2(n9005), .A(n9004), .ZN(n9006) );
  OAI211_X1 U10398 ( .C1(n9008), .C2(n9054), .A(n9007), .B(n9006), .ZN(n9068)
         );
  MUX2_X1 U10399 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9068), .S(n10098), .Z(
        P2_U3546) );
  AOI211_X1 U10400 ( .C1(n9058), .C2(n9011), .A(n9010), .B(n9009), .ZN(n9012)
         );
  OAI21_X1 U10401 ( .B1(n9013), .B2(n9054), .A(n9012), .ZN(n9069) );
  MUX2_X1 U10402 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9069), .S(n10098), .Z(
        P2_U3545) );
  AOI22_X1 U10403 ( .A1(n9015), .A2(n10035), .B1(n9058), .B2(n9014), .ZN(n9016) );
  OAI211_X1 U10404 ( .C1(n9018), .C2(n9054), .A(n9017), .B(n9016), .ZN(n9070)
         );
  MUX2_X1 U10405 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9070), .S(n10098), .Z(
        P2_U3544) );
  NAND3_X1 U10406 ( .A1(n9019), .A2(n8905), .A3(n10082), .ZN(n9024) );
  AOI22_X1 U10407 ( .A1(n9021), .A2(n10035), .B1(n9058), .B2(n9020), .ZN(n9022) );
  NAND3_X1 U10408 ( .A1(n9024), .A2(n9023), .A3(n9022), .ZN(n9071) );
  MUX2_X1 U10409 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9071), .S(n10098), .Z(
        P2_U3543) );
  AOI22_X1 U10410 ( .A1(n9026), .A2(n10035), .B1(n9058), .B2(n9025), .ZN(n9027) );
  OAI211_X1 U10411 ( .C1(n9029), .C2(n9054), .A(n9028), .B(n9027), .ZN(n9072)
         );
  MUX2_X1 U10412 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9072), .S(n10098), .Z(
        P2_U3542) );
  AOI22_X1 U10413 ( .A1(n9031), .A2(n10035), .B1(n9058), .B2(n9030), .ZN(n9032) );
  OAI211_X1 U10414 ( .C1(n9034), .C2(n9054), .A(n9033), .B(n9032), .ZN(n9073)
         );
  MUX2_X1 U10415 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9073), .S(n10098), .Z(
        P2_U3541) );
  AOI22_X1 U10416 ( .A1(n9036), .A2(n10035), .B1(n9058), .B2(n9035), .ZN(n9037) );
  OAI211_X1 U10417 ( .C1(n9039), .C2(n9054), .A(n9038), .B(n9037), .ZN(n9074)
         );
  MUX2_X1 U10418 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9074), .S(n10098), .Z(
        P2_U3540) );
  AOI211_X1 U10419 ( .C1(n9058), .C2(n9042), .A(n9041), .B(n9040), .ZN(n9043)
         );
  OAI21_X1 U10420 ( .B1(n9044), .B2(n9054), .A(n9043), .ZN(n9075) );
  MUX2_X1 U10421 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9075), .S(n10098), .Z(
        P2_U3539) );
  AOI22_X1 U10422 ( .A1(n9046), .A2(n10035), .B1(n9058), .B2(n9045), .ZN(n9047) );
  OAI211_X1 U10423 ( .C1(n9049), .C2(n9054), .A(n9048), .B(n9047), .ZN(n9076)
         );
  MUX2_X1 U10424 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9076), .S(n10098), .Z(
        P2_U3538) );
  AOI21_X1 U10425 ( .B1(n9058), .B2(n9051), .A(n9050), .ZN(n9052) );
  OAI211_X1 U10426 ( .C1(n9055), .C2(n9054), .A(n9053), .B(n9052), .ZN(n9077)
         );
  MUX2_X1 U10427 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9077), .S(n10098), .Z(
        P2_U3537) );
  INV_X1 U10428 ( .A(n9056), .ZN(n9062) );
  AOI22_X1 U10429 ( .A1(n9059), .A2(n10035), .B1(n9058), .B2(n9057), .ZN(n9060) );
  OAI211_X1 U10430 ( .C1(n9063), .C2(n9062), .A(n9061), .B(n9060), .ZN(n9078)
         );
  MUX2_X1 U10431 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9078), .S(n10098), .Z(
        P2_U3533) );
  MUX2_X1 U10432 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9065), .S(n10086), .Z(
        P2_U3518) );
  MUX2_X1 U10433 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9066), .S(n10086), .Z(
        P2_U3516) );
  MUX2_X1 U10434 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9067), .S(n10086), .Z(
        P2_U3515) );
  MUX2_X1 U10435 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9068), .S(n10086), .Z(
        P2_U3514) );
  MUX2_X1 U10436 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9069), .S(n10086), .Z(
        P2_U3513) );
  MUX2_X1 U10437 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9070), .S(n10086), .Z(
        P2_U3512) );
  MUX2_X1 U10438 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9071), .S(n10086), .Z(
        P2_U3511) );
  MUX2_X1 U10439 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9072), .S(n10086), .Z(
        P2_U3510) );
  MUX2_X1 U10440 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9073), .S(n10086), .Z(
        P2_U3509) );
  MUX2_X1 U10441 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9074), .S(n10086), .Z(
        P2_U3508) );
  MUX2_X1 U10442 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9075), .S(n10086), .Z(
        P2_U3507) );
  MUX2_X1 U10443 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9076), .S(n10086), .Z(
        P2_U3505) );
  MUX2_X1 U10444 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9077), .S(n10086), .Z(
        P2_U3502) );
  MUX2_X1 U10445 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9078), .S(n10086), .Z(
        P2_U3490) );
  INV_X1 U10446 ( .A(n9079), .ZN(n9594) );
  NAND3_X1 U10447 ( .A1(n9081), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n9083) );
  OAI22_X1 U10448 ( .A1(n9080), .A2(n9083), .B1(n9082), .B2(n9087), .ZN(n9084)
         );
  INV_X1 U10449 ( .A(n9084), .ZN(n9085) );
  OAI21_X1 U10450 ( .B1(n9594), .B2(n4477), .A(n9085), .ZN(P2_U3327) );
  INV_X1 U10451 ( .A(n9086), .ZN(n9598) );
  OAI222_X1 U10452 ( .A1(n4477), .A2(n9598), .B1(P2_U3152), .B2(n9089), .C1(
        n9088), .C2(n9087), .ZN(P2_U3329) );
  MUX2_X1 U10453 ( .A(n9090), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10454 ( .A(n9092), .B(n9091), .ZN(n9093) );
  XNOR2_X1 U10455 ( .A(n9094), .B(n9093), .ZN(n9099) );
  NAND2_X1 U10456 ( .A1(n9288), .A2(n9196), .ZN(n9096) );
  AOI22_X1 U10457 ( .A1(n9282), .A2(n9191), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n9095) );
  OAI211_X1 U10458 ( .C1(n9321), .C2(n9193), .A(n9096), .B(n9095), .ZN(n9097)
         );
  AOI21_X1 U10459 ( .B1(n9489), .B2(n9170), .A(n9097), .ZN(n9098) );
  OAI21_X1 U10460 ( .B1(n9099), .B2(n9186), .A(n9098), .ZN(P1_U3212) );
  NOR2_X1 U10461 ( .A1(n5749), .A2(n9100), .ZN(n9105) );
  AOI21_X1 U10462 ( .B1(n9103), .B2(n9102), .A(n9101), .ZN(n9104) );
  OAI21_X1 U10463 ( .B1(n9105), .B2(n9104), .A(n9660), .ZN(n9110) );
  OAI22_X1 U10464 ( .A1(n9344), .A2(n9665), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9106), .ZN(n9108) );
  NOR2_X1 U10465 ( .A1(n9380), .A2(n9193), .ZN(n9107) );
  AOI211_X1 U10466 ( .C1(n9196), .C2(n9352), .A(n9108), .B(n9107), .ZN(n9109)
         );
  OAI211_X1 U10467 ( .C1(n9347), .C2(n9199), .A(n9110), .B(n9109), .ZN(
        P1_U3214) );
  INV_X1 U10468 ( .A(n9431), .ZN(n9572) );
  OAI21_X1 U10469 ( .B1(n9113), .B2(n9112), .A(n9111), .ZN(n9114) );
  NAND2_X1 U10470 ( .A1(n9114), .A2(n9660), .ZN(n9118) );
  NAND2_X1 U10471 ( .A1(n9202), .A2(n9196), .ZN(n9115) );
  NAND2_X1 U10472 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9250) );
  OAI211_X1 U10473 ( .C1(n9427), .C2(n9193), .A(n9115), .B(n9250), .ZN(n9116)
         );
  AOI21_X1 U10474 ( .B1(n9420), .B2(n9191), .A(n9116), .ZN(n9117) );
  OAI211_X1 U10475 ( .C1(n9572), .C2(n9199), .A(n9118), .B(n9117), .ZN(
        P1_U3217) );
  NAND2_X1 U10476 ( .A1(n9153), .A2(n9154), .ZN(n9152) );
  NAND2_X1 U10477 ( .A1(n9152), .A2(n9156), .ZN(n9119) );
  XOR2_X1 U10478 ( .A(n9120), .B(n9119), .Z(n9125) );
  AOI22_X1 U10479 ( .A1(n9202), .A2(n9655), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9122) );
  NAND2_X1 U10480 ( .A1(n9191), .A2(n9374), .ZN(n9121) );
  OAI211_X1 U10481 ( .C1(n9380), .C2(n9652), .A(n9122), .B(n9121), .ZN(n9123)
         );
  AOI21_X1 U10482 ( .B1(n9519), .B2(n9170), .A(n9123), .ZN(n9124) );
  OAI21_X1 U10483 ( .B1(n9125), .B2(n9186), .A(n9124), .ZN(P1_U3221) );
  NAND2_X1 U10484 ( .A1(n9126), .A2(n9144), .ZN(n9143) );
  NAND2_X1 U10485 ( .A1(n9143), .A2(n9127), .ZN(n9128) );
  XOR2_X1 U10486 ( .A(n9129), .B(n9128), .Z(n9134) );
  OAI22_X1 U10487 ( .A1(n9315), .A2(n9665), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10310), .ZN(n9131) );
  NOR2_X1 U10488 ( .A1(n9322), .A2(n9193), .ZN(n9130) );
  AOI211_X1 U10489 ( .C1(n9196), .C2(n9287), .A(n9131), .B(n9130), .ZN(n9133)
         );
  NAND2_X1 U10490 ( .A1(n9313), .A2(n9170), .ZN(n9132) );
  OAI211_X1 U10491 ( .C1(n9134), .C2(n9186), .A(n9133), .B(n9132), .ZN(
        P1_U3223) );
  XOR2_X1 U10492 ( .A(n9136), .B(n9135), .Z(n9142) );
  NOR2_X1 U10493 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9137), .ZN(n9894) );
  NOR2_X1 U10494 ( .A1(n9193), .A2(n9671), .ZN(n9138) );
  AOI211_X1 U10495 ( .C1(n9196), .C2(n9464), .A(n9894), .B(n9138), .ZN(n9139)
         );
  OAI21_X1 U10496 ( .B1(n9665), .B2(n9476), .A(n9139), .ZN(n9140) );
  AOI21_X1 U10497 ( .B1(n9474), .B2(n9170), .A(n9140), .ZN(n9141) );
  OAI21_X1 U10498 ( .B1(n9142), .B2(n9186), .A(n9141), .ZN(P1_U3226) );
  NAND2_X1 U10499 ( .A1(n9331), .A2(n9959), .ZN(n9506) );
  OAI21_X1 U10500 ( .B1(n9144), .B2(n9126), .A(n9143), .ZN(n9145) );
  NAND2_X1 U10501 ( .A1(n9145), .A2(n9660), .ZN(n9150) );
  AOI22_X1 U10502 ( .A1(n9334), .A2(n9191), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9146) );
  OAI21_X1 U10503 ( .B1(n9147), .B2(n9193), .A(n9146), .ZN(n9148) );
  AOI21_X1 U10504 ( .B1(n9196), .B2(n9327), .A(n9148), .ZN(n9149) );
  OAI211_X1 U10505 ( .C1(n9151), .C2(n9506), .A(n9150), .B(n9149), .ZN(
        P1_U3227) );
  INV_X1 U10506 ( .A(n9152), .ZN(n9157) );
  AOI21_X1 U10507 ( .B1(n9154), .B2(n9156), .A(n9153), .ZN(n9155) );
  AOI21_X1 U10508 ( .B1(n9157), .B2(n9156), .A(n9155), .ZN(n9162) );
  NAND2_X1 U10509 ( .A1(n9402), .A2(n9196), .ZN(n9159) );
  AOI22_X1 U10510 ( .A1(n9655), .A2(n9444), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9158) );
  OAI211_X1 U10511 ( .C1(n9665), .C2(n9409), .A(n9159), .B(n9158), .ZN(n9160)
         );
  AOI21_X1 U10512 ( .B1(n9408), .B2(n9170), .A(n9160), .ZN(n9161) );
  OAI21_X1 U10513 ( .B1(n9162), .B2(n9186), .A(n9161), .ZN(P1_U3231) );
  NAND2_X1 U10514 ( .A1(n9164), .A2(n9163), .ZN(n9165) );
  XOR2_X1 U10515 ( .A(n9166), .B(n9165), .Z(n9172) );
  NAND2_X1 U10516 ( .A1(n9367), .A2(n9196), .ZN(n9168) );
  AOI22_X1 U10517 ( .A1(n9402), .A2(n9655), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9167) );
  OAI211_X1 U10518 ( .C1(n9665), .C2(n9361), .A(n9168), .B(n9167), .ZN(n9169)
         );
  AOI21_X1 U10519 ( .B1(n9514), .B2(n9170), .A(n9169), .ZN(n9171) );
  OAI21_X1 U10520 ( .B1(n9172), .B2(n9186), .A(n9171), .ZN(P1_U3233) );
  INV_X1 U10521 ( .A(n9452), .ZN(n9576) );
  INV_X1 U10522 ( .A(n9176), .ZN(n9173) );
  NOR2_X1 U10523 ( .A1(n9174), .A2(n9173), .ZN(n9179) );
  AOI21_X1 U10524 ( .B1(n9177), .B2(n9176), .A(n9175), .ZN(n9178) );
  OAI21_X1 U10525 ( .B1(n9179), .B2(n9178), .A(n9660), .ZN(n9184) );
  NAND2_X1 U10526 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9912) );
  OAI21_X1 U10527 ( .B1(n9180), .B2(n9652), .A(n9912), .ZN(n9182) );
  NOR2_X1 U10528 ( .A1(n9665), .A2(n9453), .ZN(n9181) );
  AOI211_X1 U10529 ( .C1(n9655), .C2(n9443), .A(n9182), .B(n9181), .ZN(n9183)
         );
  OAI211_X1 U10530 ( .C1(n9576), .C2(n9199), .A(n9184), .B(n9183), .ZN(
        P1_U3236) );
  AOI21_X1 U10531 ( .B1(n9185), .B2(n9187), .A(n9186), .ZN(n9189) );
  NAND2_X1 U10532 ( .A1(n9189), .A2(n9188), .ZN(n9198) );
  INV_X1 U10533 ( .A(n9190), .ZN(n9298) );
  AOI22_X1 U10534 ( .A1(n9298), .A2(n9191), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9192) );
  OAI21_X1 U10535 ( .B1(n9194), .B2(n9193), .A(n9192), .ZN(n9195) );
  AOI21_X1 U10536 ( .B1(n9196), .B2(n9304), .A(n9195), .ZN(n9197) );
  OAI211_X1 U10537 ( .C1(n9300), .C2(n9199), .A(n9198), .B(n9197), .ZN(
        P1_U3238) );
  MUX2_X1 U10538 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9200), .S(P1_U4006), .Z(
        P1_U3586) );
  MUX2_X1 U10539 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9257), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10540 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9201), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10541 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9288), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10542 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9304), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10543 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9287), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10544 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9327), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10545 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9352), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10546 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9367), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10547 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9351), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10548 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9402), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10549 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9202), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10550 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9444), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10551 ( .A(n9464), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9211), .Z(
        P1_U3573) );
  MUX2_X1 U10552 ( .A(n9443), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9211), .Z(
        P1_U3572) );
  MUX2_X1 U10553 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9463), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10554 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9203), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10555 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9703), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10556 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9204), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10557 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9704), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10558 ( .A(n9205), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9211), .Z(
        P1_U3566) );
  MUX2_X1 U10559 ( .A(n9206), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9211), .Z(
        P1_U3565) );
  MUX2_X1 U10560 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9207), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10561 ( .A(n9654), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9211), .Z(
        P1_U3563) );
  MUX2_X1 U10562 ( .A(n9208), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9211), .Z(
        P1_U3562) );
  MUX2_X1 U10563 ( .A(n9209), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9211), .Z(
        P1_U3561) );
  MUX2_X1 U10564 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9210), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10565 ( .A(n9212), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9211), .Z(
        P1_U3559) );
  MUX2_X1 U10566 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9213), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10567 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n5204), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10568 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n7186), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10569 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6854), .S(P1_U4006), .Z(
        P1_U3555) );
  NAND2_X1 U10570 ( .A1(n9762), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n9224) );
  AOI22_X1 U10571 ( .A1(n9883), .A2(n9214), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        P1_U3084), .ZN(n9223) );
  OAI211_X1 U10572 ( .C1(n9217), .C2(n9216), .A(n9911), .B(n9215), .ZN(n9222)
         );
  OAI211_X1 U10573 ( .C1(n9220), .C2(n9219), .A(n9900), .B(n9218), .ZN(n9221)
         );
  NAND4_X1 U10574 ( .A1(n9224), .A2(n9223), .A3(n9222), .A4(n9221), .ZN(
        P1_U3242) );
  NAND2_X1 U10575 ( .A1(n9225), .A2(n9238), .ZN(n9227) );
  NAND2_X1 U10576 ( .A1(n9227), .A2(n9226), .ZN(n9228) );
  NOR2_X1 U10577 ( .A1(n9240), .A2(n9228), .ZN(n9229) );
  INV_X1 U10578 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9866) );
  XNOR2_X1 U10579 ( .A(n9228), .B(n9240), .ZN(n9867) );
  NOR2_X1 U10580 ( .A1(n9866), .A2(n9867), .ZN(n9865) );
  NOR2_X1 U10581 ( .A1(n9229), .A2(n9865), .ZN(n9879) );
  NAND2_X1 U10582 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9882), .ZN(n9230) );
  OAI21_X1 U10583 ( .B1(n9882), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9230), .ZN(
        n9878) );
  NOR2_X1 U10584 ( .A1(n9879), .A2(n9878), .ZN(n9877) );
  AOI21_X1 U10585 ( .B1(n9882), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9877), .ZN(
        n9891) );
  NAND2_X1 U10586 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9234), .ZN(n9231) );
  OAI21_X1 U10587 ( .B1(n9234), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9231), .ZN(
        n9892) );
  NOR2_X1 U10588 ( .A1(n9891), .A2(n9892), .ZN(n9890) );
  XNOR2_X1 U10589 ( .A(n9233), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n9907) );
  INV_X1 U10590 ( .A(n9247), .ZN(n9245) );
  INV_X1 U10591 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9537) );
  XNOR2_X1 U10592 ( .A(n9233), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9919) );
  INV_X1 U10593 ( .A(n9234), .ZN(n9897) );
  XNOR2_X1 U10594 ( .A(n9234), .B(n10394), .ZN(n9902) );
  NOR2_X1 U10595 ( .A1(n9242), .A2(n9235), .ZN(n9236) );
  AOI21_X1 U10596 ( .B1(n9235), .B2(n9242), .A(n9236), .ZN(n9885) );
  AOI21_X1 U10597 ( .B1(n9238), .B2(n10283), .A(n9237), .ZN(n9239) );
  NAND2_X1 U10598 ( .A1(n9870), .A2(n9239), .ZN(n9241) );
  XNOR2_X1 U10599 ( .A(n9240), .B(n9239), .ZN(n9872) );
  NAND2_X1 U10600 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9872), .ZN(n9871) );
  NAND2_X1 U10601 ( .A1(n9241), .A2(n9871), .ZN(n9886) );
  NAND2_X1 U10602 ( .A1(n9885), .A2(n9886), .ZN(n9884) );
  OAI21_X1 U10603 ( .B1(n9242), .B2(n9235), .A(n9884), .ZN(n9901) );
  NAND2_X1 U10604 ( .A1(n9902), .A2(n9901), .ZN(n9899) );
  OAI21_X1 U10605 ( .B1(n9897), .B2(n10394), .A(n9899), .ZN(n9918) );
  NOR2_X1 U10606 ( .A1(n9919), .A2(n9918), .ZN(n9917) );
  AOI21_X1 U10607 ( .B1(n9915), .B2(n9537), .A(n9917), .ZN(n9243) );
  XOR2_X1 U10608 ( .A(n9243), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9246) );
  OAI21_X1 U10609 ( .B1(n9246), .B2(n9921), .A(n9914), .ZN(n9244) );
  AOI21_X1 U10610 ( .B1(n9245), .B2(n9911), .A(n9244), .ZN(n9249) );
  AOI22_X1 U10611 ( .A1(n9247), .A2(n9911), .B1(n9900), .B2(n9246), .ZN(n9248)
         );
  MUX2_X1 U10612 ( .A(n9249), .B(n9248), .S(n9430), .Z(n9251) );
  OAI211_X1 U10613 ( .C1(n5119), .C2(n9924), .A(n9251), .B(n9250), .ZN(
        P1_U3260) );
  INV_X1 U10614 ( .A(n9257), .ZN(n9260) );
  INV_X1 U10615 ( .A(n9258), .ZN(n9259) );
  OAI222_X1 U10616 ( .A1(n9426), .A2(n5058), .B1(n9260), .B2(n9259), .C1(n9253), .C2(n9668), .ZN(n9261) );
  INV_X1 U10617 ( .A(n9261), .ZN(n9488) );
  NAND2_X1 U10618 ( .A1(n9488), .A2(n5041), .ZN(n9269) );
  NAND2_X1 U10619 ( .A1(n9485), .A2(n9263), .ZN(n9264) );
  INV_X1 U10620 ( .A(n9486), .ZN(n9267) );
  AOI22_X1 U10621 ( .A1(n9485), .A2(n9713), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9678), .ZN(n9265) );
  OAI21_X1 U10622 ( .B1(n9267), .B2(n9266), .A(n9265), .ZN(n9268) );
  AOI21_X1 U10623 ( .B1(n9269), .B2(n9478), .A(n9268), .ZN(n9270) );
  OAI21_X1 U10624 ( .B1(n9484), .B2(n9415), .A(n9270), .ZN(P1_U3355) );
  NAND2_X1 U10625 ( .A1(n9271), .A2(n4555), .ZN(n9274) );
  AOI22_X1 U10626 ( .A1(n9272), .A2(n9679), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9709), .ZN(n9273) );
  OAI211_X1 U10627 ( .C1(n9275), .C2(n9475), .A(n9274), .B(n9273), .ZN(n9276)
         );
  AOI21_X1 U10628 ( .B1(n9277), .B2(n9478), .A(n9276), .ZN(n9278) );
  OAI21_X1 U10629 ( .B1(n9279), .B2(n9415), .A(n9278), .ZN(P1_U3263) );
  XOR2_X1 U10630 ( .A(n9280), .B(n9285), .Z(n9493) );
  AOI21_X1 U10631 ( .B1(n9489), .B2(n9295), .A(n8419), .ZN(n9490) );
  AOI22_X1 U10632 ( .A1(n9282), .A2(n9679), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9709), .ZN(n9283) );
  OAI21_X1 U10633 ( .B1(n4791), .B2(n9475), .A(n9283), .ZN(n9292) );
  OAI211_X1 U10634 ( .C1(n9286), .C2(n9285), .A(n9284), .B(n9700), .ZN(n9290)
         );
  AOI22_X1 U10635 ( .A1(n9288), .A2(n9702), .B1(n9705), .B2(n9287), .ZN(n9289)
         );
  AND2_X1 U10636 ( .A1(n9290), .A2(n9289), .ZN(n9492) );
  NOR2_X1 U10637 ( .A1(n9492), .A2(n9678), .ZN(n9291) );
  AOI211_X1 U10638 ( .C1(n9691), .C2(n9490), .A(n9292), .B(n9291), .ZN(n9293)
         );
  OAI21_X1 U10639 ( .B1(n9493), .B2(n9415), .A(n9293), .ZN(P1_U3264) );
  XOR2_X1 U10640 ( .A(n9301), .B(n9294), .Z(n9498) );
  INV_X1 U10641 ( .A(n9312), .ZN(n9297) );
  INV_X1 U10642 ( .A(n9295), .ZN(n9296) );
  AOI21_X1 U10643 ( .B1(n9494), .B2(n9297), .A(n9296), .ZN(n9495) );
  AOI22_X1 U10644 ( .A1(n9298), .A2(n9679), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9709), .ZN(n9299) );
  OAI21_X1 U10645 ( .B1(n9300), .B2(n9475), .A(n9299), .ZN(n9307) );
  OAI21_X1 U10646 ( .B1(n9303), .B2(n8411), .A(n9302), .ZN(n9305) );
  AOI222_X1 U10647 ( .A1(n9700), .A2(n9305), .B1(n9304), .B2(n9702), .C1(n9327), .C2(n9705), .ZN(n9497) );
  NOR2_X1 U10648 ( .A1(n9497), .A2(n9678), .ZN(n9306) );
  AOI211_X1 U10649 ( .C1(n9495), .C2(n9691), .A(n9307), .B(n9306), .ZN(n9308)
         );
  OAI21_X1 U10650 ( .B1(n9498), .B2(n9415), .A(n9308), .ZN(P1_U3265) );
  INV_X1 U10651 ( .A(n9309), .ZN(n9311) );
  OAI21_X1 U10652 ( .B1(n9311), .B2(n9318), .A(n9310), .ZN(n9501) );
  INV_X1 U10653 ( .A(n9501), .ZN(n9325) );
  AOI211_X1 U10654 ( .C1(n9313), .C2(n9333), .A(n9986), .B(n9312), .ZN(n9500)
         );
  INV_X1 U10655 ( .A(n9313), .ZN(n9558) );
  NOR2_X1 U10656 ( .A1(n9558), .A2(n9475), .ZN(n9317) );
  OAI22_X1 U10657 ( .A1(n9315), .A2(n9693), .B1(n9314), .B2(n9478), .ZN(n9316)
         );
  AOI211_X1 U10658 ( .C1(n9500), .C2(n4555), .A(n9317), .B(n9316), .ZN(n9324)
         );
  XNOR2_X1 U10659 ( .A(n9319), .B(n9318), .ZN(n9320) );
  OAI222_X1 U10660 ( .A1(n9668), .A2(n9322), .B1(n9670), .B2(n9321), .C1(n9320), .C2(n9426), .ZN(n9499) );
  NAND2_X1 U10661 ( .A1(n9499), .A2(n9478), .ZN(n9323) );
  OAI211_X1 U10662 ( .C1(n9325), .C2(n9415), .A(n9324), .B(n9323), .ZN(
        P1_U3266) );
  OAI21_X1 U10663 ( .B1(n4533), .B2(n8406), .A(n9326), .ZN(n9328) );
  AOI222_X1 U10664 ( .A1(n9700), .A2(n9328), .B1(n9327), .B2(n9702), .C1(n9367), .C2(n9705), .ZN(n9507) );
  XNOR2_X1 U10665 ( .A(n9330), .B(n9329), .ZN(n9504) );
  NAND2_X1 U10666 ( .A1(n9504), .A2(n9469), .ZN(n9340) );
  INV_X1 U10667 ( .A(n9331), .ZN(n9336) );
  INV_X1 U10668 ( .A(n9332), .ZN(n9343) );
  OAI211_X1 U10669 ( .C1(n9336), .C2(n9343), .A(n9960), .B(n9333), .ZN(n9505)
         );
  INV_X1 U10670 ( .A(n9505), .ZN(n9338) );
  AOI22_X1 U10671 ( .A1(n9334), .A2(n9679), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9678), .ZN(n9335) );
  OAI21_X1 U10672 ( .B1(n9336), .B2(n9475), .A(n9335), .ZN(n9337) );
  AOI21_X1 U10673 ( .B1(n9338), .B2(n4555), .A(n9337), .ZN(n9339) );
  OAI211_X1 U10674 ( .C1(n9709), .C2(n9507), .A(n9340), .B(n9339), .ZN(
        P1_U3267) );
  XNOR2_X1 U10675 ( .A(n9341), .B(n9342), .ZN(n9513) );
  AOI21_X1 U10676 ( .B1(n9509), .B2(n4787), .A(n9343), .ZN(n9510) );
  INV_X1 U10677 ( .A(n9344), .ZN(n9345) );
  AOI22_X1 U10678 ( .A1(n9345), .A2(n9679), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9709), .ZN(n9346) );
  OAI21_X1 U10679 ( .B1(n9347), .B2(n9475), .A(n9346), .ZN(n9356) );
  OAI211_X1 U10680 ( .C1(n9350), .C2(n9349), .A(n9348), .B(n9700), .ZN(n9354)
         );
  AOI22_X1 U10681 ( .A1(n9352), .A2(n9702), .B1(n9705), .B2(n9351), .ZN(n9353)
         );
  NOR2_X1 U10682 ( .A1(n9512), .A2(n9678), .ZN(n9355) );
  AOI211_X1 U10683 ( .C1(n9510), .C2(n9691), .A(n9356), .B(n9355), .ZN(n9357)
         );
  OAI21_X1 U10684 ( .B1(n9513), .B2(n9415), .A(n9357), .ZN(P1_U3268) );
  XNOR2_X1 U10685 ( .A(n9359), .B(n9358), .ZN(n9518) );
  AOI21_X1 U10686 ( .B1(n9514), .B2(n9372), .A(n9360), .ZN(n9515) );
  INV_X1 U10687 ( .A(n9361), .ZN(n9362) );
  AOI22_X1 U10688 ( .A1(n9362), .A2(n9679), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9709), .ZN(n9363) );
  OAI21_X1 U10689 ( .B1(n4785), .B2(n9475), .A(n9363), .ZN(n9370) );
  NAND2_X1 U10690 ( .A1(n9376), .A2(n9364), .ZN(n9366) );
  XNOR2_X1 U10691 ( .A(n9366), .B(n9365), .ZN(n9368) );
  AOI222_X1 U10692 ( .A1(n9700), .A2(n9368), .B1(n9402), .B2(n9705), .C1(n9367), .C2(n9702), .ZN(n9517) );
  NOR2_X1 U10693 ( .A1(n9517), .A2(n9678), .ZN(n9369) );
  AOI211_X1 U10694 ( .C1(n9515), .C2(n9691), .A(n9370), .B(n9369), .ZN(n9371)
         );
  OAI21_X1 U10695 ( .B1(n9415), .B2(n9518), .A(n9371), .ZN(P1_U3269) );
  AOI21_X1 U10696 ( .B1(n9405), .B2(n9519), .A(n9986), .ZN(n9373) );
  AND2_X1 U10697 ( .A1(n9373), .A2(n9372), .ZN(n9521) );
  AND2_X1 U10698 ( .A1(n9374), .A2(n9679), .ZN(n9381) );
  NAND2_X1 U10699 ( .A1(n9400), .A2(n9375), .ZN(n9378) );
  INV_X1 U10700 ( .A(n9376), .ZN(n9377) );
  AOI21_X1 U10701 ( .B1(n9387), .B2(n9378), .A(n9377), .ZN(n9379) );
  OAI222_X1 U10702 ( .A1(n9670), .A2(n9380), .B1(n9668), .B2(n9428), .C1(n9426), .C2(n9379), .ZN(n9520) );
  AOI211_X1 U10703 ( .C1(n9521), .C2(n9430), .A(n9381), .B(n9520), .ZN(n9390)
         );
  AOI22_X1 U10704 ( .A1(n9519), .A2(n9713), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9678), .ZN(n9389) );
  OR2_X1 U10705 ( .A1(n9382), .A2(n9383), .ZN(n9385) );
  NAND2_X1 U10706 ( .A1(n9385), .A2(n9384), .ZN(n9386) );
  XOR2_X1 U10707 ( .A(n9387), .B(n9386), .Z(n9522) );
  NAND2_X1 U10708 ( .A1(n9522), .A2(n9469), .ZN(n9388) );
  OAI211_X1 U10709 ( .C1(n9390), .C2(n9678), .A(n9389), .B(n9388), .ZN(
        P1_U3270) );
  NAND2_X1 U10710 ( .A1(n9447), .A2(n9391), .ZN(n9393) );
  AND2_X1 U10711 ( .A1(n9393), .A2(n9392), .ZN(n9394) );
  XOR2_X1 U10712 ( .A(n9397), .B(n9394), .Z(n9526) );
  INV_X1 U10713 ( .A(n9526), .ZN(n9416) );
  INV_X1 U10714 ( .A(n9395), .ZN(n9422) );
  INV_X1 U10715 ( .A(n9396), .ZN(n9398) );
  OAI21_X1 U10716 ( .B1(n9422), .B2(n9398), .A(n9397), .ZN(n9399) );
  OAI211_X1 U10717 ( .C1(n9401), .C2(n9400), .A(n9399), .B(n9700), .ZN(n9404)
         );
  AOI22_X1 U10718 ( .A1(n9402), .A2(n9702), .B1(n9705), .B2(n9444), .ZN(n9403)
         );
  NAND2_X1 U10719 ( .A1(n9404), .A2(n9403), .ZN(n9524) );
  INV_X1 U10720 ( .A(n9419), .ZN(n9407) );
  INV_X1 U10721 ( .A(n9405), .ZN(n9406) );
  AOI211_X1 U10722 ( .C1(n9408), .C2(n9407), .A(n9986), .B(n9406), .ZN(n9525)
         );
  NAND2_X1 U10723 ( .A1(n9525), .A2(n4555), .ZN(n9412) );
  INV_X1 U10724 ( .A(n9409), .ZN(n9410) );
  AOI22_X1 U10725 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(n9678), .B1(n9410), .B2(
        n9679), .ZN(n9411) );
  OAI211_X1 U10726 ( .C1(n9568), .C2(n9475), .A(n9412), .B(n9411), .ZN(n9413)
         );
  AOI21_X1 U10727 ( .B1(n9524), .B2(n9478), .A(n9413), .ZN(n9414) );
  OAI21_X1 U10728 ( .B1(n9416), .B2(n9415), .A(n9414), .ZN(P1_U3271) );
  NAND2_X1 U10729 ( .A1(n9450), .A2(n9431), .ZN(n9417) );
  NAND2_X1 U10730 ( .A1(n9417), .A2(n9960), .ZN(n9418) );
  NOR2_X1 U10731 ( .A1(n9419), .A2(n9418), .ZN(n9530) );
  AND2_X1 U10732 ( .A1(n9420), .A2(n9679), .ZN(n9429) );
  INV_X1 U10733 ( .A(n9421), .ZN(n9424) );
  INV_X1 U10734 ( .A(n9433), .ZN(n9423) );
  AOI21_X1 U10735 ( .B1(n9424), .B2(n9423), .A(n9422), .ZN(n9425) );
  OAI222_X1 U10736 ( .A1(n9670), .A2(n9428), .B1(n9668), .B2(n9427), .C1(n9426), .C2(n9425), .ZN(n9529) );
  AOI211_X1 U10737 ( .C1(n9530), .C2(n9430), .A(n9429), .B(n9529), .ZN(n9437)
         );
  AOI22_X1 U10738 ( .A1(n9431), .A2(n9713), .B1(n9709), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n9436) );
  NAND2_X1 U10739 ( .A1(n9447), .A2(n9432), .ZN(n9434) );
  XNOR2_X1 U10740 ( .A(n9434), .B(n9433), .ZN(n9531) );
  NAND2_X1 U10741 ( .A1(n9531), .A2(n9469), .ZN(n9435) );
  OAI211_X1 U10742 ( .C1(n9437), .C2(n9678), .A(n9436), .B(n9435), .ZN(
        P1_U3272) );
  NAND2_X1 U10743 ( .A1(n9439), .A2(n9438), .ZN(n9440) );
  NAND2_X1 U10744 ( .A1(n9441), .A2(n9440), .ZN(n9442) );
  NAND2_X1 U10745 ( .A1(n9442), .A2(n9700), .ZN(n9446) );
  AOI22_X1 U10746 ( .A1(n9444), .A2(n9702), .B1(n9705), .B2(n9443), .ZN(n9445)
         );
  NAND2_X1 U10747 ( .A1(n9446), .A2(n9445), .ZN(n9534) );
  INV_X1 U10748 ( .A(n9534), .ZN(n9459) );
  INV_X1 U10749 ( .A(n9447), .ZN(n9448) );
  AOI21_X1 U10750 ( .B1(n9449), .B2(n9382), .A(n9448), .ZN(n9536) );
  NAND2_X1 U10751 ( .A1(n9536), .A2(n9469), .ZN(n9458) );
  INV_X1 U10752 ( .A(n9450), .ZN(n9451) );
  AOI211_X1 U10753 ( .C1(n9452), .C2(n9471), .A(n9986), .B(n9451), .ZN(n9535)
         );
  NOR2_X1 U10754 ( .A1(n9576), .A2(n9475), .ZN(n9456) );
  OAI22_X1 U10755 ( .A1(n9478), .A2(n9454), .B1(n9453), .B2(n9693), .ZN(n9455)
         );
  AOI211_X1 U10756 ( .C1(n9535), .C2(n4555), .A(n9456), .B(n9455), .ZN(n9457)
         );
  OAI211_X1 U10757 ( .C1(n9709), .C2(n9459), .A(n9458), .B(n9457), .ZN(
        P1_U3273) );
  INV_X1 U10758 ( .A(n9467), .ZN(n9460) );
  XNOR2_X1 U10759 ( .A(n9461), .B(n9460), .ZN(n9462) );
  NAND2_X1 U10760 ( .A1(n9462), .A2(n9700), .ZN(n9466) );
  AOI22_X1 U10761 ( .A1(n9464), .A2(n9702), .B1(n9705), .B2(n9463), .ZN(n9465)
         );
  NAND2_X1 U10762 ( .A1(n9466), .A2(n9465), .ZN(n9539) );
  INV_X1 U10763 ( .A(n9539), .ZN(n9483) );
  XNOR2_X1 U10764 ( .A(n9468), .B(n9467), .ZN(n9541) );
  NAND2_X1 U10765 ( .A1(n9541), .A2(n9469), .ZN(n9482) );
  INV_X1 U10766 ( .A(n9470), .ZN(n9473) );
  INV_X1 U10767 ( .A(n9471), .ZN(n9472) );
  AOI211_X1 U10768 ( .C1(n9474), .C2(n9473), .A(n9986), .B(n9472), .ZN(n9540)
         );
  NOR2_X1 U10769 ( .A1(n9580), .A2(n9475), .ZN(n9480) );
  INV_X1 U10770 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9477) );
  OAI22_X1 U10771 ( .A1(n9478), .A2(n9477), .B1(n9476), .B2(n9693), .ZN(n9479)
         );
  AOI211_X1 U10772 ( .C1(n9540), .C2(n4555), .A(n9480), .B(n9479), .ZN(n9481)
         );
  OAI211_X1 U10773 ( .C1(n9709), .C2(n9483), .A(n9482), .B(n9481), .ZN(
        P1_U3274) );
  AOI22_X1 U10774 ( .A1(n9486), .A2(n9960), .B1(n9959), .B2(n9485), .ZN(n9487)
         );
  MUX2_X1 U10775 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9552), .S(n10004), .Z(
        P1_U3552) );
  AOI22_X1 U10776 ( .A1(n9490), .A2(n9960), .B1(n9959), .B2(n9489), .ZN(n9491)
         );
  OAI211_X1 U10777 ( .C1(n9493), .C2(n9970), .A(n9492), .B(n9491), .ZN(n9553)
         );
  MUX2_X1 U10778 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9553), .S(n10004), .Z(
        P1_U3550) );
  AOI22_X1 U10779 ( .A1(n9495), .A2(n9960), .B1(n9959), .B2(n9494), .ZN(n9496)
         );
  OAI211_X1 U10780 ( .C1(n9498), .C2(n9970), .A(n9497), .B(n9496), .ZN(n9554)
         );
  MUX2_X1 U10781 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9554), .S(n10004), .Z(
        P1_U3549) );
  INV_X1 U10782 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9502) );
  AOI211_X1 U10783 ( .C1(n9501), .C2(n9988), .A(n9500), .B(n9499), .ZN(n9555)
         );
  MUX2_X1 U10784 ( .A(n9502), .B(n9555), .S(n10004), .Z(n9503) );
  OAI21_X1 U10785 ( .B1(n9558), .B2(n9551), .A(n9503), .ZN(P1_U3548) );
  NAND2_X1 U10786 ( .A1(n9504), .A2(n9988), .ZN(n9508) );
  NAND4_X1 U10787 ( .A1(n9508), .A2(n9507), .A3(n9506), .A4(n9505), .ZN(n9559)
         );
  MUX2_X1 U10788 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9559), .S(n10004), .Z(
        P1_U3547) );
  AOI22_X1 U10789 ( .A1(n9510), .A2(n9960), .B1(n9959), .B2(n9509), .ZN(n9511)
         );
  OAI211_X1 U10790 ( .C1(n9513), .C2(n9970), .A(n9512), .B(n9511), .ZN(n9560)
         );
  MUX2_X1 U10791 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9560), .S(n10004), .Z(
        P1_U3546) );
  AOI22_X1 U10792 ( .A1(n9515), .A2(n9960), .B1(n9959), .B2(n9514), .ZN(n9516)
         );
  OAI211_X1 U10793 ( .C1(n9518), .C2(n9970), .A(n9517), .B(n9516), .ZN(n9561)
         );
  MUX2_X1 U10794 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9561), .S(n10004), .Z(
        P1_U3545) );
  INV_X1 U10795 ( .A(n9519), .ZN(n9564) );
  INV_X1 U10796 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10370) );
  AOI211_X1 U10797 ( .C1(n9522), .C2(n9988), .A(n9521), .B(n9520), .ZN(n9562)
         );
  MUX2_X1 U10798 ( .A(n10370), .B(n9562), .S(n10004), .Z(n9523) );
  OAI21_X1 U10799 ( .B1(n9564), .B2(n9551), .A(n9523), .ZN(P1_U3544) );
  AOI211_X1 U10800 ( .C1(n9526), .C2(n9988), .A(n9525), .B(n9524), .ZN(n9565)
         );
  MUX2_X1 U10801 ( .A(n9527), .B(n9565), .S(n10004), .Z(n9528) );
  OAI21_X1 U10802 ( .B1(n9568), .B2(n9551), .A(n9528), .ZN(P1_U3543) );
  INV_X1 U10803 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9532) );
  AOI211_X1 U10804 ( .C1(n9531), .C2(n9988), .A(n9530), .B(n9529), .ZN(n9569)
         );
  MUX2_X1 U10805 ( .A(n9532), .B(n9569), .S(n10004), .Z(n9533) );
  OAI21_X1 U10806 ( .B1(n9572), .B2(n9551), .A(n9533), .ZN(P1_U3542) );
  AOI211_X1 U10807 ( .C1(n9536), .C2(n9988), .A(n9535), .B(n9534), .ZN(n9573)
         );
  MUX2_X1 U10808 ( .A(n9537), .B(n9573), .S(n10004), .Z(n9538) );
  OAI21_X1 U10809 ( .B1(n9576), .B2(n9551), .A(n9538), .ZN(P1_U3541) );
  AOI211_X1 U10810 ( .C1(n9541), .C2(n9988), .A(n9540), .B(n9539), .ZN(n9577)
         );
  MUX2_X1 U10811 ( .A(n10394), .B(n9577), .S(n10004), .Z(n9542) );
  OAI21_X1 U10812 ( .B1(n9580), .B2(n9551), .A(n9542), .ZN(P1_U3540) );
  AOI211_X1 U10813 ( .C1(n9545), .C2(n9988), .A(n9544), .B(n9543), .ZN(n9581)
         );
  MUX2_X1 U10814 ( .A(n9235), .B(n9581), .S(n10004), .Z(n9546) );
  OAI21_X1 U10815 ( .B1(n9584), .B2(n9551), .A(n9546), .ZN(P1_U3539) );
  AOI211_X1 U10816 ( .C1(n9549), .C2(n9988), .A(n9548), .B(n9547), .ZN(n9585)
         );
  MUX2_X1 U10817 ( .A(n10283), .B(n9585), .S(n10004), .Z(n9550) );
  OAI21_X1 U10818 ( .B1(n9589), .B2(n9551), .A(n9550), .ZN(P1_U3537) );
  MUX2_X1 U10819 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9552), .S(n9992), .Z(
        P1_U3520) );
  MUX2_X1 U10820 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9553), .S(n9992), .Z(
        P1_U3518) );
  MUX2_X1 U10821 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9554), .S(n9992), .Z(
        P1_U3517) );
  INV_X1 U10822 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9556) );
  MUX2_X1 U10823 ( .A(n9556), .B(n9555), .S(n9992), .Z(n9557) );
  OAI21_X1 U10824 ( .B1(n9558), .B2(n9588), .A(n9557), .ZN(P1_U3516) );
  MUX2_X1 U10825 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9559), .S(n9992), .Z(
        P1_U3515) );
  MUX2_X1 U10826 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9560), .S(n9992), .Z(
        P1_U3514) );
  MUX2_X1 U10827 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9561), .S(n9992), .Z(
        P1_U3513) );
  MUX2_X1 U10828 ( .A(n10404), .B(n9562), .S(n9992), .Z(n9563) );
  OAI21_X1 U10829 ( .B1(n9564), .B2(n9588), .A(n9563), .ZN(P1_U3512) );
  INV_X1 U10830 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9566) );
  MUX2_X1 U10831 ( .A(n9566), .B(n9565), .S(n9992), .Z(n9567) );
  OAI21_X1 U10832 ( .B1(n9568), .B2(n9588), .A(n9567), .ZN(P1_U3511) );
  INV_X1 U10833 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9570) );
  MUX2_X1 U10834 ( .A(n9570), .B(n9569), .S(n9992), .Z(n9571) );
  OAI21_X1 U10835 ( .B1(n9572), .B2(n9588), .A(n9571), .ZN(P1_U3510) );
  INV_X1 U10836 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9574) );
  MUX2_X1 U10837 ( .A(n9574), .B(n9573), .S(n9992), .Z(n9575) );
  OAI21_X1 U10838 ( .B1(n9576), .B2(n9588), .A(n9575), .ZN(P1_U3508) );
  INV_X1 U10839 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9578) );
  MUX2_X1 U10840 ( .A(n9578), .B(n9577), .S(n9992), .Z(n9579) );
  OAI21_X1 U10841 ( .B1(n9580), .B2(n9588), .A(n9579), .ZN(P1_U3505) );
  INV_X1 U10842 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9582) );
  MUX2_X1 U10843 ( .A(n9582), .B(n9581), .S(n9992), .Z(n9583) );
  OAI21_X1 U10844 ( .B1(n9584), .B2(n9588), .A(n9583), .ZN(P1_U3502) );
  INV_X1 U10845 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9586) );
  MUX2_X1 U10846 ( .A(n9586), .B(n9585), .S(n9992), .Z(n9587) );
  OAI21_X1 U10847 ( .B1(n9589), .B2(n9588), .A(n9587), .ZN(P1_U3496) );
  NOR4_X1 U10848 ( .A1(n5080), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9590), .ZN(n9591) );
  AOI21_X1 U10849 ( .B1(n9592), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9591), .ZN(
        n9593) );
  OAI21_X1 U10850 ( .B1(n9594), .B2(n9599), .A(n9593), .ZN(P1_U3322) );
  OAI222_X1 U10851 ( .A1(n9599), .A2(n9598), .B1(n5082), .B2(P1_U3084), .C1(
        n9596), .C2(n9595), .ZN(P1_U3324) );
  MUX2_X1 U10852 ( .A(n9600), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10853 ( .A1(n10013), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9611) );
  NAND2_X1 U10854 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9603) );
  AOI211_X1 U10855 ( .C1(n9603), .C2(n9602), .A(n9601), .B(n9612), .ZN(n9604)
         );
  AOI21_X1 U10856 ( .B1(n9618), .B2(n9605), .A(n9604), .ZN(n9610) );
  INV_X1 U10857 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10087) );
  NOR2_X1 U10858 ( .A1(n10015), .A2(n10087), .ZN(n9607) );
  OAI211_X1 U10859 ( .C1(n9608), .C2(n9607), .A(n10010), .B(n9606), .ZN(n9609)
         );
  NAND3_X1 U10860 ( .A1(n9611), .A2(n9610), .A3(n9609), .ZN(P2_U3246) );
  AOI22_X1 U10861 ( .A1(n10013), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9624) );
  AOI211_X1 U10862 ( .C1(n9615), .C2(n9614), .A(n9613), .B(n9612), .ZN(n9616)
         );
  AOI21_X1 U10863 ( .B1(n9618), .B2(n9617), .A(n9616), .ZN(n9623) );
  OAI211_X1 U10864 ( .C1(n9621), .C2(n9620), .A(n10010), .B(n9619), .ZN(n9622)
         );
  NAND3_X1 U10865 ( .A1(n9624), .A2(n9623), .A3(n9622), .ZN(P2_U3247) );
  OAI21_X1 U10866 ( .B1(n9627), .B2(n9626), .A(n9625), .ZN(n9629) );
  AOI222_X1 U10867 ( .A1(n6494), .A2(n9632), .B1(n9631), .B2(n9630), .C1(n9629), .C2(n9628), .ZN(n9634) );
  OAI211_X1 U10868 ( .C1(n9636), .C2(n9635), .A(n9634), .B(n9633), .ZN(
        P2_U3228) );
  OAI22_X1 U10869 ( .A1(n9638), .A2(n10078), .B1(n9637), .B2(n10076), .ZN(
        n9639) );
  AOI211_X1 U10870 ( .C1(n9641), .C2(n10082), .A(n9640), .B(n9639), .ZN(n9648)
         );
  AOI22_X1 U10871 ( .A1(n10098), .A2(n9648), .B1(n8017), .B2(n10096), .ZN(
        P2_U3536) );
  OAI22_X1 U10872 ( .A1(n9643), .A2(n10078), .B1(n9642), .B2(n10076), .ZN(
        n9645) );
  AOI211_X1 U10873 ( .C1(n9646), .C2(n10082), .A(n9645), .B(n9644), .ZN(n9650)
         );
  AOI22_X1 U10874 ( .A1(n10098), .A2(n9650), .B1(n9647), .B2(n10096), .ZN(
        P2_U3534) );
  AOI22_X1 U10875 ( .A1(n10086), .A2(n9648), .B1(n6258), .B2(n10084), .ZN(
        P2_U3499) );
  INV_X1 U10876 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9649) );
  AOI22_X1 U10877 ( .A1(n10086), .A2(n9650), .B1(n9649), .B2(n10084), .ZN(
        P2_U3493) );
  OAI22_X1 U10878 ( .A1(n9652), .A2(n9651), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9810), .ZN(n9653) );
  AOI21_X1 U10879 ( .B1(n9655), .B2(n9654), .A(n9653), .ZN(n9663) );
  XNOR2_X1 U10880 ( .A(n9656), .B(n9657), .ZN(n9661) );
  NOR2_X1 U10881 ( .A1(n9658), .A2(n9976), .ZN(n9982) );
  AOI22_X1 U10882 ( .A1(n9661), .A2(n9660), .B1(n9659), .B2(n9982), .ZN(n9662)
         );
  OAI211_X1 U10883 ( .C1(n9665), .C2(n9664), .A(n9663), .B(n9662), .ZN(
        P1_U3229) );
  XNOR2_X1 U10884 ( .A(n9667), .B(n9666), .ZN(n9677) );
  OAI22_X1 U10885 ( .A1(n9671), .A2(n9670), .B1(n9669), .B2(n9668), .ZN(n9676)
         );
  XNOR2_X1 U10886 ( .A(n9673), .B(n9672), .ZN(n9681) );
  NOR2_X1 U10887 ( .A1(n9681), .A2(n9674), .ZN(n9675) );
  AOI211_X1 U10888 ( .C1(n9700), .C2(n9677), .A(n9676), .B(n9675), .ZN(n9718)
         );
  AOI222_X1 U10889 ( .A1(n9682), .A2(n9713), .B1(n9680), .B2(n9679), .C1(
        P1_REG2_REG_15__SCAN_IN), .C2(n9678), .ZN(n9685) );
  INV_X1 U10890 ( .A(n9681), .ZN(n9721) );
  OAI21_X1 U10891 ( .B1(n4778), .B2(n4542), .A(n4495), .ZN(n9717) );
  INV_X1 U10892 ( .A(n9717), .ZN(n9683) );
  AOI22_X1 U10893 ( .A1(n9721), .A2(n9692), .B1(n9691), .B2(n9683), .ZN(n9684)
         );
  OAI211_X1 U10894 ( .C1(n9709), .C2(n9718), .A(n9685), .B(n9684), .ZN(
        P1_U3276) );
  XNOR2_X1 U10895 ( .A(n9686), .B(n7859), .ZN(n9726) );
  OR2_X1 U10896 ( .A1(n9687), .A2(n9723), .ZN(n9688) );
  NAND2_X1 U10897 ( .A1(n9689), .A2(n9688), .ZN(n9724) );
  INV_X1 U10898 ( .A(n9724), .ZN(n9690) );
  AOI22_X1 U10899 ( .A1(n9726), .A2(n9692), .B1(n9691), .B2(n9690), .ZN(n9715)
         );
  OAI22_X1 U10900 ( .A1(n9478), .A2(n9695), .B1(n9694), .B2(n9693), .ZN(n9711)
         );
  NAND2_X1 U10901 ( .A1(n9697), .A2(n9696), .ZN(n9698) );
  NAND2_X1 U10902 ( .A1(n9699), .A2(n9698), .ZN(n9701) );
  NAND2_X1 U10903 ( .A1(n9701), .A2(n9700), .ZN(n9707) );
  AOI22_X1 U10904 ( .A1(n9705), .A2(n9704), .B1(n9703), .B2(n9702), .ZN(n9706)
         );
  NAND2_X1 U10905 ( .A1(n9707), .A2(n9706), .ZN(n9708) );
  AOI21_X1 U10906 ( .B1(n9726), .B2(n9968), .A(n9708), .ZN(n9728) );
  NOR2_X1 U10907 ( .A1(n9728), .A2(n9709), .ZN(n9710) );
  AOI211_X1 U10908 ( .C1(n9713), .C2(n9712), .A(n9711), .B(n9710), .ZN(n9714)
         );
  NAND2_X1 U10909 ( .A1(n9715), .A2(n9714), .ZN(P1_U3278) );
  OAI21_X1 U10910 ( .B1(n9717), .B2(n9986), .A(n9716), .ZN(n9720) );
  INV_X1 U10911 ( .A(n9718), .ZN(n9719) );
  AOI211_X1 U10912 ( .C1(n9950), .C2(n9721), .A(n9720), .B(n9719), .ZN(n9745)
         );
  INV_X1 U10913 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9722) );
  AOI22_X1 U10914 ( .A1(n10004), .A2(n9745), .B1(n9722), .B2(n10002), .ZN(
        P1_U3538) );
  OAI22_X1 U10915 ( .A1(n9724), .A2(n9986), .B1(n9723), .B2(n9976), .ZN(n9725)
         );
  AOI21_X1 U10916 ( .B1(n9726), .B2(n9950), .A(n9725), .ZN(n9727) );
  AND2_X1 U10917 ( .A1(n9728), .A2(n9727), .ZN(n9747) );
  AOI22_X1 U10918 ( .A1(n10004), .A2(n9747), .B1(n10205), .B2(n10002), .ZN(
        P1_U3536) );
  NOR2_X1 U10919 ( .A1(n9729), .A2(n9970), .ZN(n9734) );
  OAI211_X1 U10920 ( .C1(n9732), .C2(n9976), .A(n9731), .B(n9730), .ZN(n9733)
         );
  AOI21_X1 U10921 ( .B1(n9734), .B2(n7853), .A(n9733), .ZN(n9749) );
  AOI22_X1 U10922 ( .A1(n10004), .A2(n9749), .B1(n9735), .B2(n10002), .ZN(
        P1_U3535) );
  INV_X1 U10923 ( .A(n9736), .ZN(n9742) );
  INV_X1 U10924 ( .A(n9737), .ZN(n9738) );
  OAI22_X1 U10925 ( .A1(n9739), .A2(n9986), .B1(n9738), .B2(n9976), .ZN(n9741)
         );
  AOI211_X1 U10926 ( .C1(n9950), .C2(n9742), .A(n9741), .B(n9740), .ZN(n9750)
         );
  AOI22_X1 U10927 ( .A1(n10004), .A2(n9750), .B1(n9743), .B2(n10002), .ZN(
        P1_U3534) );
  INV_X1 U10928 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9744) );
  AOI22_X1 U10929 ( .A1(n9992), .A2(n9745), .B1(n9744), .B2(n9990), .ZN(
        P1_U3499) );
  INV_X1 U10930 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9746) );
  AOI22_X1 U10931 ( .A1(n9992), .A2(n9747), .B1(n9746), .B2(n9990), .ZN(
        P1_U3493) );
  INV_X1 U10932 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9748) );
  AOI22_X1 U10933 ( .A1(n9992), .A2(n9749), .B1(n9748), .B2(n9990), .ZN(
        P1_U3490) );
  AOI22_X1 U10934 ( .A1(n9992), .A2(n9750), .B1(n5411), .B2(n9990), .ZN(
        P1_U3487) );
  XNOR2_X1 U10935 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10936 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  NOR3_X1 U10937 ( .A1(n9921), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n5179), .ZN(
        n9761) );
  INV_X1 U10938 ( .A(n9751), .ZN(n9759) );
  INV_X1 U10939 ( .A(n9752), .ZN(n9757) );
  INV_X1 U10940 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10407) );
  INV_X1 U10941 ( .A(n9753), .ZN(n9754) );
  OAI21_X1 U10942 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n10407), .A(n9754), .ZN(
        n9756) );
  NAND4_X1 U10943 ( .A1(n9757), .A2(n9756), .A3(P1_STATE_REG_SCAN_IN), .A4(
        n9755), .ZN(n9758) );
  NOR2_X1 U10944 ( .A1(n9759), .A2(n9758), .ZN(n9760) );
  AOI211_X1 U10945 ( .C1(P1_ADDR_REG_0__SCAN_IN), .C2(n9762), .A(n9761), .B(
        n9760), .ZN(n9763) );
  OAI21_X1 U10946 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7054), .A(n9763), .ZN(
        P1_U3241) );
  INV_X1 U10947 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9778) );
  OAI21_X1 U10948 ( .B1(n9766), .B2(n9765), .A(n9764), .ZN(n9767) );
  NAND2_X1 U10949 ( .A1(n9911), .A2(n9767), .ZN(n9770) );
  INV_X1 U10950 ( .A(n9768), .ZN(n9769) );
  OAI211_X1 U10951 ( .C1(n9914), .C2(n9771), .A(n9770), .B(n9769), .ZN(n9772)
         );
  INV_X1 U10952 ( .A(n9772), .ZN(n9777) );
  OAI211_X1 U10953 ( .C1(n9775), .C2(n9774), .A(n9900), .B(n9773), .ZN(n9776)
         );
  OAI211_X1 U10954 ( .C1(n9778), .C2(n9924), .A(n9777), .B(n9776), .ZN(
        P1_U3246) );
  AOI21_X1 U10955 ( .B1(n9781), .B2(n9780), .A(n9779), .ZN(n9782) );
  NAND2_X1 U10956 ( .A1(n9911), .A2(n9782), .ZN(n9785) );
  INV_X1 U10957 ( .A(n9783), .ZN(n9784) );
  OAI211_X1 U10958 ( .C1(n9914), .C2(n9786), .A(n9785), .B(n9784), .ZN(n9787)
         );
  INV_X1 U10959 ( .A(n9787), .ZN(n9793) );
  AOI21_X1 U10960 ( .B1(n9790), .B2(n9789), .A(n9788), .ZN(n9791) );
  OR2_X1 U10961 ( .A1(n9791), .A2(n9921), .ZN(n9792) );
  OAI211_X1 U10962 ( .C1(n9794), .C2(n9924), .A(n9793), .B(n9792), .ZN(
        P1_U3247) );
  XOR2_X1 U10963 ( .A(n9796), .B(n9795), .Z(n9806) );
  INV_X1 U10964 ( .A(n9911), .ZN(n9876) );
  INV_X1 U10965 ( .A(n9797), .ZN(n9798) );
  NAND2_X1 U10966 ( .A1(n9799), .A2(n9798), .ZN(n9801) );
  NAND3_X1 U10967 ( .A1(n9801), .A2(n9900), .A3(n9800), .ZN(n9805) );
  AOI21_X1 U10968 ( .B1(n9883), .B2(n9803), .A(n9802), .ZN(n9804) );
  OAI211_X1 U10969 ( .C1(n9806), .C2(n9876), .A(n9805), .B(n9804), .ZN(n9807)
         );
  INV_X1 U10970 ( .A(n9807), .ZN(n9808) );
  OAI21_X1 U10971 ( .B1(n9924), .B2(n9809), .A(n9808), .ZN(P1_U3249) );
  NOR2_X1 U10972 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9810), .ZN(n9815) );
  AOI211_X1 U10973 ( .C1(n9813), .C2(n9812), .A(n9811), .B(n9876), .ZN(n9814)
         );
  AOI211_X1 U10974 ( .C1(n9883), .C2(n9816), .A(n9815), .B(n9814), .ZN(n9822)
         );
  AOI21_X1 U10975 ( .B1(n9819), .B2(n9818), .A(n9817), .ZN(n9820) );
  OR2_X1 U10976 ( .A1(n9921), .A2(n9820), .ZN(n9821) );
  OAI211_X1 U10977 ( .C1(n10515), .C2(n9924), .A(n9822), .B(n9821), .ZN(
        P1_U3250) );
  INV_X1 U10978 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9839) );
  INV_X1 U10979 ( .A(n9823), .ZN(n9831) );
  AOI21_X1 U10980 ( .B1(n9826), .B2(n9825), .A(n9824), .ZN(n9827) );
  NAND2_X1 U10981 ( .A1(n9911), .A2(n9827), .ZN(n9830) );
  INV_X1 U10982 ( .A(n9828), .ZN(n9829) );
  OAI211_X1 U10983 ( .C1(n9914), .C2(n9831), .A(n9830), .B(n9829), .ZN(n9832)
         );
  INV_X1 U10984 ( .A(n9832), .ZN(n9838) );
  AOI21_X1 U10985 ( .B1(n9835), .B2(n9834), .A(n9833), .ZN(n9836) );
  OR2_X1 U10986 ( .A1(n9836), .A2(n9921), .ZN(n9837) );
  OAI211_X1 U10987 ( .C1(n9839), .C2(n9924), .A(n9838), .B(n9837), .ZN(
        P1_U3251) );
  INV_X1 U10988 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9852) );
  AOI211_X1 U10989 ( .C1(n9842), .C2(n9841), .A(n9876), .B(n9840), .ZN(n9843)
         );
  AOI211_X1 U10990 ( .C1(n9883), .C2(n9845), .A(n9844), .B(n9843), .ZN(n9851)
         );
  AOI21_X1 U10991 ( .B1(n9848), .B2(n9847), .A(n9846), .ZN(n9849) );
  OR2_X1 U10992 ( .A1(n9849), .A2(n9921), .ZN(n9850) );
  OAI211_X1 U10993 ( .C1(n9852), .C2(n9924), .A(n9851), .B(n9850), .ZN(
        P1_U3253) );
  INV_X1 U10994 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10412) );
  AOI211_X1 U10995 ( .C1(n9855), .C2(n9854), .A(n9876), .B(n9853), .ZN(n9856)
         );
  AOI211_X1 U10996 ( .C1(n9883), .C2(n9858), .A(n9857), .B(n9856), .ZN(n9864)
         );
  AOI21_X1 U10997 ( .B1(n9861), .B2(n9860), .A(n9859), .ZN(n9862) );
  OR2_X1 U10998 ( .A1(n9862), .A2(n9921), .ZN(n9863) );
  OAI211_X1 U10999 ( .C1(n10412), .C2(n9924), .A(n9864), .B(n9863), .ZN(
        P1_U3254) );
  INV_X1 U11000 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9875) );
  AOI211_X1 U11001 ( .C1(n9867), .C2(n9866), .A(n9865), .B(n9876), .ZN(n9868)
         );
  AOI211_X1 U11002 ( .C1(n9883), .C2(n9870), .A(n9869), .B(n9868), .ZN(n9874)
         );
  OAI211_X1 U11003 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9872), .A(n9900), .B(
        n9871), .ZN(n9873) );
  OAI211_X1 U11004 ( .C1(n9875), .C2(n9924), .A(n9874), .B(n9873), .ZN(
        P1_U3256) );
  INV_X1 U11005 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9889) );
  AOI211_X1 U11006 ( .C1(n9879), .C2(n9878), .A(n9877), .B(n9876), .ZN(n9880)
         );
  AOI211_X1 U11007 ( .C1(n9883), .C2(n9882), .A(n9881), .B(n9880), .ZN(n9888)
         );
  OAI211_X1 U11008 ( .C1(n9886), .C2(n9885), .A(n9900), .B(n9884), .ZN(n9887)
         );
  OAI211_X1 U11009 ( .C1(n9889), .C2(n9924), .A(n9888), .B(n9887), .ZN(
        P1_U3257) );
  INV_X1 U11010 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9905) );
  AOI21_X1 U11011 ( .B1(n9892), .B2(n9891), .A(n9890), .ZN(n9893) );
  NAND2_X1 U11012 ( .A1(n9911), .A2(n9893), .ZN(n9896) );
  INV_X1 U11013 ( .A(n9894), .ZN(n9895) );
  OAI211_X1 U11014 ( .C1(n9897), .C2(n9914), .A(n9896), .B(n9895), .ZN(n9898)
         );
  INV_X1 U11015 ( .A(n9898), .ZN(n9904) );
  OAI211_X1 U11016 ( .C1(n9902), .C2(n9901), .A(n9900), .B(n9899), .ZN(n9903)
         );
  OAI211_X1 U11017 ( .C1(n9905), .C2(n9924), .A(n9904), .B(n9903), .ZN(
        P1_U3258) );
  INV_X1 U11018 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10511) );
  NAND2_X1 U11019 ( .A1(n9907), .A2(n9906), .ZN(n9910) );
  INV_X1 U11020 ( .A(n9908), .ZN(n9909) );
  NAND3_X1 U11021 ( .A1(n9911), .A2(n9910), .A3(n9909), .ZN(n9913) );
  OAI211_X1 U11022 ( .C1(n9915), .C2(n9914), .A(n9913), .B(n9912), .ZN(n9916)
         );
  INV_X1 U11023 ( .A(n9916), .ZN(n9923) );
  AOI21_X1 U11024 ( .B1(n9919), .B2(n9918), .A(n9917), .ZN(n9920) );
  OR2_X1 U11025 ( .A1(n9921), .A2(n9920), .ZN(n9922) );
  OAI211_X1 U11026 ( .C1(n10511), .C2(n9924), .A(n9923), .B(n9922), .ZN(
        P1_U3259) );
  AND2_X1 U11027 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9927), .ZN(P1_U3292) );
  INV_X1 U11028 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10277) );
  NOR2_X1 U11029 ( .A1(n9926), .A2(n10277), .ZN(P1_U3293) );
  AND2_X1 U11030 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9927), .ZN(P1_U3294) );
  AND2_X1 U11031 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9927), .ZN(P1_U3295) );
  AND2_X1 U11032 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9927), .ZN(P1_U3296) );
  AND2_X1 U11033 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9927), .ZN(P1_U3297) );
  AND2_X1 U11034 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9927), .ZN(P1_U3298) );
  AND2_X1 U11035 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9927), .ZN(P1_U3299) );
  AND2_X1 U11036 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9927), .ZN(P1_U3300) );
  AND2_X1 U11037 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9927), .ZN(P1_U3301) );
  AND2_X1 U11038 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9927), .ZN(P1_U3302) );
  AND2_X1 U11039 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9927), .ZN(P1_U3303) );
  AND2_X1 U11040 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9927), .ZN(P1_U3304) );
  AND2_X1 U11041 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9927), .ZN(P1_U3305) );
  INV_X1 U11042 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10413) );
  NOR2_X1 U11043 ( .A1(n9926), .A2(n10413), .ZN(P1_U3306) );
  AND2_X1 U11044 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9927), .ZN(P1_U3307) );
  AND2_X1 U11045 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9927), .ZN(P1_U3308) );
  AND2_X1 U11046 ( .A1(n9927), .A2(P1_D_REG_14__SCAN_IN), .ZN(P1_U3309) );
  AND2_X1 U11047 ( .A1(n9927), .A2(P1_D_REG_13__SCAN_IN), .ZN(P1_U3310) );
  INV_X1 U11048 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10282) );
  NOR2_X1 U11049 ( .A1(n9926), .A2(n10282), .ZN(P1_U3311) );
  AND2_X1 U11050 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9927), .ZN(P1_U3312) );
  AND2_X1 U11051 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9927), .ZN(P1_U3313) );
  AND2_X1 U11052 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9927), .ZN(P1_U3314) );
  AND2_X1 U11053 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9927), .ZN(P1_U3315) );
  AND2_X1 U11054 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9927), .ZN(P1_U3316) );
  AND2_X1 U11055 ( .A1(n9927), .A2(P1_D_REG_6__SCAN_IN), .ZN(P1_U3317) );
  AND2_X1 U11056 ( .A1(n9927), .A2(P1_D_REG_5__SCAN_IN), .ZN(P1_U3318) );
  AND2_X1 U11057 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9927), .ZN(P1_U3319) );
  AND2_X1 U11058 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9927), .ZN(P1_U3320) );
  AND2_X1 U11059 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9927), .ZN(P1_U3321) );
  NAND2_X1 U11060 ( .A1(n9928), .A2(n9931), .ZN(n9929) );
  OAI21_X1 U11061 ( .B1(n9931), .B2(n9930), .A(n9929), .ZN(P1_U3440) );
  INV_X1 U11062 ( .A(n9932), .ZN(n9937) );
  OAI21_X1 U11063 ( .B1(n9934), .B2(n9976), .A(n9933), .ZN(n9936) );
  AOI211_X1 U11064 ( .C1(n9950), .C2(n9937), .A(n9936), .B(n9935), .ZN(n9993)
         );
  INV_X1 U11065 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9938) );
  AOI22_X1 U11066 ( .A1(n9992), .A2(n9993), .B1(n9938), .B2(n9990), .ZN(
        P1_U3457) );
  OAI22_X1 U11067 ( .A1(n9940), .A2(n9986), .B1(n9939), .B2(n9976), .ZN(n9942)
         );
  AOI211_X1 U11068 ( .C1(n9950), .C2(n9943), .A(n9942), .B(n9941), .ZN(n9994)
         );
  INV_X1 U11069 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9944) );
  AOI22_X1 U11070 ( .A1(n9992), .A2(n9994), .B1(n9944), .B2(n9990), .ZN(
        P1_U3460) );
  OAI22_X1 U11071 ( .A1(n9946), .A2(n9986), .B1(n9945), .B2(n9976), .ZN(n9948)
         );
  AOI211_X1 U11072 ( .C1(n9950), .C2(n9949), .A(n9948), .B(n9947), .ZN(n9995)
         );
  INV_X1 U11073 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9951) );
  AOI22_X1 U11074 ( .A1(n9992), .A2(n9995), .B1(n9951), .B2(n9990), .ZN(
        P1_U3463) );
  AND3_X1 U11075 ( .A1(n7296), .A2(n9988), .A3(n9952), .ZN(n9953) );
  NOR4_X1 U11076 ( .A1(n9956), .A2(n9955), .A3(n9954), .A4(n9953), .ZN(n9996)
         );
  INV_X1 U11077 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9957) );
  AOI22_X1 U11078 ( .A1(n9992), .A2(n9996), .B1(n9957), .B2(n9990), .ZN(
        P1_U3469) );
  AOI22_X1 U11079 ( .A1(n9961), .A2(n9960), .B1(n9959), .B2(n9958), .ZN(n9962)
         );
  OAI21_X1 U11080 ( .B1(n9964), .B2(n9963), .A(n9962), .ZN(n9965) );
  AOI211_X1 U11081 ( .C1(n9968), .C2(n9967), .A(n9966), .B(n9965), .ZN(n9997)
         );
  INV_X1 U11082 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9969) );
  AOI22_X1 U11083 ( .A1(n9992), .A2(n9997), .B1(n9969), .B2(n9990), .ZN(
        P1_U3472) );
  NOR2_X1 U11084 ( .A1(n9971), .A2(n9970), .ZN(n9975) );
  NOR4_X1 U11085 ( .A1(n9975), .A2(n9974), .A3(n9973), .A4(n9972), .ZN(n9999)
         );
  AOI22_X1 U11086 ( .A1(n9992), .A2(n9999), .B1(n5298), .B2(n9990), .ZN(
        P1_U3475) );
  OAI22_X1 U11087 ( .A1(n9978), .A2(n9986), .B1(n9977), .B2(n9976), .ZN(n9979)
         );
  AOI211_X1 U11088 ( .C1(n9981), .C2(n9988), .A(n9980), .B(n9979), .ZN(n10001)
         );
  AOI22_X1 U11089 ( .A1(n9992), .A2(n10001), .B1(n5323), .B2(n9990), .ZN(
        P1_U3478) );
  INV_X1 U11090 ( .A(n9982), .ZN(n9983) );
  OAI211_X1 U11091 ( .C1(n9986), .C2(n9985), .A(n9984), .B(n9983), .ZN(n9987)
         );
  AOI21_X1 U11092 ( .B1(n9989), .B2(n9988), .A(n9987), .ZN(n10003) );
  INV_X1 U11093 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9991) );
  AOI22_X1 U11094 ( .A1(n9992), .A2(n10003), .B1(n9991), .B2(n9990), .ZN(
        P1_U3481) );
  AOI22_X1 U11095 ( .A1(n10004), .A2(n9993), .B1(n6759), .B2(n10002), .ZN(
        P1_U3524) );
  INV_X1 U11096 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10256) );
  AOI22_X1 U11097 ( .A1(n10004), .A2(n9994), .B1(n10256), .B2(n10002), .ZN(
        P1_U3525) );
  AOI22_X1 U11098 ( .A1(n10004), .A2(n9995), .B1(n6764), .B2(n10002), .ZN(
        P1_U3526) );
  AOI22_X1 U11099 ( .A1(n10004), .A2(n9996), .B1(n6758), .B2(n10002), .ZN(
        P1_U3528) );
  AOI22_X1 U11100 ( .A1(n10004), .A2(n9997), .B1(n6768), .B2(n10002), .ZN(
        P1_U3529) );
  AOI22_X1 U11101 ( .A1(n10004), .A2(n9999), .B1(n9998), .B2(n10002), .ZN(
        P1_U3530) );
  AOI22_X1 U11102 ( .A1(n10004), .A2(n10001), .B1(n10000), .B2(n10002), .ZN(
        P1_U3531) );
  AOI22_X1 U11103 ( .A1(n10004), .A2(n10003), .B1(n6818), .B2(n10002), .ZN(
        P1_U3532) );
  AOI21_X1 U11104 ( .B1(n10010), .B2(n10087), .A(n10015), .ZN(n10006) );
  NAND2_X1 U11105 ( .A1(n10006), .A2(n10005), .ZN(n10007) );
  AOI21_X1 U11106 ( .B1(n10009), .B2(n10008), .A(n10007), .ZN(n10017) );
  AOI22_X1 U11107 ( .A1(n10011), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10010), .ZN(n10016) );
  AOI22_X1 U11108 ( .A1(n10013), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10014) );
  OAI221_X1 U11109 ( .B1(n10017), .B2(n10016), .C1(n10017), .C2(n10015), .A(
        n10014), .ZN(P2_U3245) );
  AND2_X1 U11110 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10128), .ZN(P2_U3297) );
  AND2_X1 U11111 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10128), .ZN(P2_U3298) );
  INV_X1 U11112 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10378) );
  NOR2_X1 U11113 ( .A1(n10020), .A2(n10378), .ZN(P2_U3299) );
  INV_X1 U11114 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10323) );
  NOR2_X1 U11115 ( .A1(n10020), .A2(n10323), .ZN(P2_U3300) );
  AND2_X1 U11116 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10128), .ZN(P2_U3301) );
  AND2_X1 U11117 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10128), .ZN(P2_U3302) );
  INV_X1 U11118 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10391) );
  NOR2_X1 U11119 ( .A1(n10020), .A2(n10391), .ZN(P2_U3303) );
  AND2_X1 U11120 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10128), .ZN(P2_U3304) );
  INV_X1 U11121 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10208) );
  NOR2_X1 U11122 ( .A1(n10020), .A2(n10208), .ZN(P2_U3305) );
  AND2_X1 U11123 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10128), .ZN(P2_U3306) );
  AND2_X1 U11124 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10128), .ZN(P2_U3308) );
  AND2_X1 U11125 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10128), .ZN(P2_U3309) );
  AND2_X1 U11126 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10128), .ZN(P2_U3310) );
  AND2_X1 U11127 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10128), .ZN(P2_U3311) );
  AND2_X1 U11128 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10128), .ZN(P2_U3312) );
  AND2_X1 U11129 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10128), .ZN(P2_U3313) );
  AND2_X1 U11130 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10128), .ZN(P2_U3314) );
  INV_X1 U11131 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10265) );
  NOR2_X1 U11132 ( .A1(n10020), .A2(n10265), .ZN(P2_U3315) );
  AND2_X1 U11133 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10128), .ZN(P2_U3316) );
  INV_X1 U11134 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10353) );
  NOR2_X1 U11135 ( .A1(n10020), .A2(n10353), .ZN(P2_U3317) );
  INV_X1 U11136 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10190) );
  NOR2_X1 U11137 ( .A1(n10020), .A2(n10190), .ZN(P2_U3318) );
  INV_X1 U11138 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10294) );
  NOR2_X1 U11139 ( .A1(n10020), .A2(n10294), .ZN(P2_U3319) );
  AND2_X1 U11140 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10128), .ZN(P2_U3320) );
  INV_X1 U11141 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10264) );
  NOR2_X1 U11142 ( .A1(n10020), .A2(n10264), .ZN(P2_U3321) );
  AND2_X1 U11143 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10128), .ZN(P2_U3322) );
  INV_X1 U11144 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10410) );
  NOR2_X1 U11145 ( .A1(n10020), .A2(n10410), .ZN(P2_U3323) );
  AND2_X1 U11146 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10128), .ZN(P2_U3324) );
  AND2_X1 U11147 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10128), .ZN(P2_U3325) );
  AND2_X1 U11148 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10128), .ZN(P2_U3326) );
  AOI22_X1 U11149 ( .A1(n10025), .A2(n10021), .B1(n10336), .B2(n10128), .ZN(
        P2_U3437) );
  INV_X1 U11150 ( .A(n10022), .ZN(n10024) );
  AOI22_X1 U11151 ( .A1(n10025), .A2(n10024), .B1(n10023), .B2(n10128), .ZN(
        P2_U3438) );
  AOI22_X1 U11152 ( .A1(n10028), .A2(n10082), .B1(n10027), .B2(n10026), .ZN(
        n10029) );
  AND2_X1 U11153 ( .A1(n10030), .A2(n10029), .ZN(n10088) );
  AOI22_X1 U11154 ( .A1(n10086), .A2(n10088), .B1(n6002), .B2(n10084), .ZN(
        P2_U3451) );
  OAI21_X1 U11155 ( .B1(n6513), .B2(n10076), .A(n10031), .ZN(n10033) );
  AOI211_X1 U11156 ( .C1(n10082), .C2(n10034), .A(n10033), .B(n10032), .ZN(
        n10089) );
  AOI22_X1 U11157 ( .A1(n10086), .A2(n10089), .B1(n5971), .B2(n10084), .ZN(
        P2_U3454) );
  NAND2_X1 U11158 ( .A1(n10036), .A2(n10035), .ZN(n10038) );
  OAI22_X1 U11159 ( .A1(n10039), .A2(n10038), .B1(n10037), .B2(n10076), .ZN(
        n10040) );
  INV_X1 U11160 ( .A(n10040), .ZN(n10043) );
  NAND2_X1 U11161 ( .A1(n10041), .A2(n10082), .ZN(n10042) );
  AND3_X1 U11162 ( .A1(n10044), .A2(n10043), .A3(n10042), .ZN(n10090) );
  AOI22_X1 U11163 ( .A1(n10086), .A2(n10090), .B1(n6013), .B2(n10084), .ZN(
        P2_U3457) );
  INV_X1 U11164 ( .A(n10045), .ZN(n10049) );
  OAI22_X1 U11165 ( .A1(n10046), .A2(n10078), .B1(n6519), .B2(n10076), .ZN(
        n10048) );
  AOI211_X1 U11166 ( .C1(n10070), .C2(n10049), .A(n10048), .B(n10047), .ZN(
        n10091) );
  INV_X1 U11167 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10050) );
  AOI22_X1 U11168 ( .A1(n10086), .A2(n10091), .B1(n10050), .B2(n10084), .ZN(
        P2_U3460) );
  AND2_X1 U11169 ( .A1(n10051), .A2(n10082), .ZN(n10055) );
  OAI22_X1 U11170 ( .A1(n10053), .A2(n10078), .B1(n10052), .B2(n10076), .ZN(
        n10054) );
  NOR3_X1 U11171 ( .A1(n10056), .A2(n10055), .A3(n10054), .ZN(n10092) );
  AOI22_X1 U11172 ( .A1(n10086), .A2(n10092), .B1(n6042), .B2(n10084), .ZN(
        P2_U3463) );
  OAI22_X1 U11173 ( .A1(n10058), .A2(n10078), .B1(n10057), .B2(n10076), .ZN(
        n10060) );
  AOI211_X1 U11174 ( .C1(n10061), .C2(n10082), .A(n10060), .B(n10059), .ZN(
        n10093) );
  INV_X1 U11175 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10062) );
  AOI22_X1 U11176 ( .A1(n10086), .A2(n10093), .B1(n10062), .B2(n10084), .ZN(
        P2_U3469) );
  INV_X1 U11177 ( .A(n10063), .ZN(n10069) );
  INV_X1 U11178 ( .A(n10064), .ZN(n10065) );
  OAI22_X1 U11179 ( .A1(n10066), .A2(n10078), .B1(n10065), .B2(n10076), .ZN(
        n10068) );
  AOI211_X1 U11180 ( .C1(n10070), .C2(n10069), .A(n10068), .B(n10067), .ZN(
        n10094) );
  AOI22_X1 U11181 ( .A1(n10086), .A2(n10094), .B1(n6118), .B2(n10084), .ZN(
        P2_U3475) );
  OAI22_X1 U11182 ( .A1(n10072), .A2(n10078), .B1(n10071), .B2(n10076), .ZN(
        n10073) );
  AOI211_X1 U11183 ( .C1(n10075), .C2(n10082), .A(n10074), .B(n10073), .ZN(
        n10095) );
  AOI22_X1 U11184 ( .A1(n10086), .A2(n10095), .B1(n6156), .B2(n10084), .ZN(
        P2_U3481) );
  OAI22_X1 U11185 ( .A1(n10079), .A2(n10078), .B1(n10077), .B2(n10076), .ZN(
        n10081) );
  AOI211_X1 U11186 ( .C1(n10083), .C2(n10082), .A(n10081), .B(n10080), .ZN(
        n10097) );
  INV_X1 U11187 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10085) );
  AOI22_X1 U11188 ( .A1(n10086), .A2(n10097), .B1(n10085), .B2(n10084), .ZN(
        P2_U3487) );
  AOI22_X1 U11189 ( .A1(n10098), .A2(n10088), .B1(n10087), .B2(n10096), .ZN(
        P2_U3520) );
  AOI22_X1 U11190 ( .A1(n10098), .A2(n10089), .B1(n10352), .B2(n10096), .ZN(
        P2_U3521) );
  AOI22_X1 U11191 ( .A1(n10098), .A2(n10090), .B1(n6700), .B2(n10096), .ZN(
        P2_U3522) );
  AOI22_X1 U11192 ( .A1(n10098), .A2(n10091), .B1(n6703), .B2(n10096), .ZN(
        P2_U3523) );
  AOI22_X1 U11193 ( .A1(n10098), .A2(n10092), .B1(n6720), .B2(n10096), .ZN(
        P2_U3524) );
  AOI22_X1 U11194 ( .A1(n10098), .A2(n10093), .B1(n6750), .B2(n10096), .ZN(
        P2_U3526) );
  AOI22_X1 U11195 ( .A1(n10098), .A2(n10094), .B1(n6958), .B2(n10096), .ZN(
        P2_U3528) );
  AOI22_X1 U11196 ( .A1(n10098), .A2(n10095), .B1(n7218), .B2(n10096), .ZN(
        P2_U3530) );
  AOI22_X1 U11197 ( .A1(n10098), .A2(n10097), .B1(n7598), .B2(n10096), .ZN(
        P2_U3532) );
  INV_X1 U11198 ( .A(n10099), .ZN(n10100) );
  NAND2_X1 U11199 ( .A1(n10101), .A2(n10100), .ZN(n10102) );
  XOR2_X1 U11200 ( .A(n10103), .B(n10102), .Z(ADD_1071_U5) );
  XOR2_X1 U11201 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11202 ( .B1(n10106), .B2(n10105), .A(n10104), .ZN(ADD_1071_U56) );
  OAI21_X1 U11203 ( .B1(n10109), .B2(n10108), .A(n10107), .ZN(ADD_1071_U57) );
  OAI21_X1 U11204 ( .B1(n10112), .B2(n10111), .A(n10110), .ZN(ADD_1071_U58) );
  OAI21_X1 U11205 ( .B1(n10115), .B2(n10114), .A(n10113), .ZN(ADD_1071_U59) );
  OAI21_X1 U11206 ( .B1(n10118), .B2(n10117), .A(n10116), .ZN(ADD_1071_U60) );
  OAI21_X1 U11207 ( .B1(n10121), .B2(n10120), .A(n10119), .ZN(ADD_1071_U61) );
  AOI21_X1 U11208 ( .B1(n10124), .B2(n10123), .A(n10122), .ZN(ADD_1071_U62) );
  AOI21_X1 U11209 ( .B1(n10127), .B2(n10126), .A(n10125), .ZN(ADD_1071_U63) );
  NAND2_X1 U11210 ( .A1(n10128), .A2(P2_D_REG_21__SCAN_IN), .ZN(n10501) );
  AOI22_X1 U11211 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(keyinput192), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(keyinput131), .ZN(n10129) );
  OAI221_X1 U11212 ( .B1(P1_DATAO_REG_17__SCAN_IN), .B2(keyinput192), .C1(
        P1_DATAO_REG_19__SCAN_IN), .C2(keyinput131), .A(n10129), .ZN(n10136)
         );
  AOI22_X1 U11213 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput209), .B1(
        P1_IR_REG_4__SCAN_IN), .B2(keyinput241), .ZN(n10130) );
  OAI221_X1 U11214 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput209), .C1(
        P1_IR_REG_4__SCAN_IN), .C2(keyinput241), .A(n10130), .ZN(n10135) );
  AOI22_X1 U11215 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(keyinput139), .B1(
        P1_REG0_REG_8__SCAN_IN), .B2(keyinput236), .ZN(n10131) );
  OAI221_X1 U11216 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(keyinput139), .C1(
        P1_REG0_REG_8__SCAN_IN), .C2(keyinput236), .A(n10131), .ZN(n10134) );
  AOI22_X1 U11217 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput246), .B1(
        P2_IR_REG_21__SCAN_IN), .B2(keyinput138), .ZN(n10132) );
  OAI221_X1 U11218 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput246), .C1(
        P2_IR_REG_21__SCAN_IN), .C2(keyinput138), .A(n10132), .ZN(n10133) );
  NOR4_X1 U11219 ( .A1(n10136), .A2(n10135), .A3(n10134), .A4(n10133), .ZN(
        n10164) );
  AOI22_X1 U11220 ( .A1(P2_D_REG_29__SCAN_IN), .A2(keyinput206), .B1(
        P1_IR_REG_31__SCAN_IN), .B2(keyinput212), .ZN(n10137) );
  OAI221_X1 U11221 ( .B1(P2_D_REG_29__SCAN_IN), .B2(keyinput206), .C1(
        P1_IR_REG_31__SCAN_IN), .C2(keyinput212), .A(n10137), .ZN(n10144) );
  AOI22_X1 U11222 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput173), .B1(
        P1_REG1_REG_3__SCAN_IN), .B2(keyinput150), .ZN(n10138) );
  OAI221_X1 U11223 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput173), .C1(
        P1_REG1_REG_3__SCAN_IN), .C2(keyinput150), .A(n10138), .ZN(n10143) );
  AOI22_X1 U11224 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(keyinput160), .B1(
        P1_D_REG_13__SCAN_IN), .B2(keyinput222), .ZN(n10139) );
  OAI221_X1 U11225 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(keyinput160), .C1(
        P1_D_REG_13__SCAN_IN), .C2(keyinput222), .A(n10139), .ZN(n10142) );
  AOI22_X1 U11226 ( .A1(P2_REG1_REG_27__SCAN_IN), .A2(keyinput140), .B1(
        P1_REG3_REG_15__SCAN_IN), .B2(keyinput198), .ZN(n10140) );
  OAI221_X1 U11227 ( .B1(P2_REG1_REG_27__SCAN_IN), .B2(keyinput140), .C1(
        P1_REG3_REG_15__SCAN_IN), .C2(keyinput198), .A(n10140), .ZN(n10141) );
  NOR4_X1 U11228 ( .A1(n10144), .A2(n10143), .A3(n10142), .A4(n10141), .ZN(
        n10163) );
  AOI22_X1 U11229 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput243), .B1(
        P1_D_REG_6__SCAN_IN), .B2(keyinput229), .ZN(n10145) );
  OAI221_X1 U11230 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput243), .C1(
        P1_D_REG_6__SCAN_IN), .C2(keyinput229), .A(n10145), .ZN(n10152) );
  AOI22_X1 U11231 ( .A1(P2_REG2_REG_4__SCAN_IN), .A2(keyinput193), .B1(
        P1_D_REG_14__SCAN_IN), .B2(keyinput133), .ZN(n10146) );
  OAI221_X1 U11232 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(keyinput193), .C1(
        P1_D_REG_14__SCAN_IN), .C2(keyinput133), .A(n10146), .ZN(n10151) );
  AOI22_X1 U11233 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(keyinput154), .B1(
        P1_REG0_REG_21__SCAN_IN), .B2(keyinput216), .ZN(n10147) );
  OAI221_X1 U11234 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(keyinput154), .C1(
        P1_REG0_REG_21__SCAN_IN), .C2(keyinput216), .A(n10147), .ZN(n10150) );
  AOI22_X1 U11235 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(keyinput168), .B1(
        P1_D_REG_17__SCAN_IN), .B2(keyinput128), .ZN(n10148) );
  OAI221_X1 U11236 ( .B1(P1_DATAO_REG_30__SCAN_IN), .B2(keyinput168), .C1(
        P1_D_REG_17__SCAN_IN), .C2(keyinput128), .A(n10148), .ZN(n10149) );
  NOR4_X1 U11237 ( .A1(n10152), .A2(n10151), .A3(n10150), .A4(n10149), .ZN(
        n10162) );
  AOI22_X1 U11238 ( .A1(P2_D_REG_25__SCAN_IN), .A2(keyinput214), .B1(SI_17_), 
        .B2(keyinput251), .ZN(n10153) );
  OAI221_X1 U11239 ( .B1(P2_D_REG_25__SCAN_IN), .B2(keyinput214), .C1(SI_17_), 
        .C2(keyinput251), .A(n10153), .ZN(n10160) );
  AOI22_X1 U11240 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(keyinput245), .B1(
        P1_IR_REG_12__SCAN_IN), .B2(keyinput226), .ZN(n10154) );
  OAI221_X1 U11241 ( .B1(P2_IR_REG_12__SCAN_IN), .B2(keyinput245), .C1(
        P1_IR_REG_12__SCAN_IN), .C2(keyinput226), .A(n10154), .ZN(n10159) );
  AOI22_X1 U11242 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(keyinput182), .B1(
        P1_IR_REG_7__SCAN_IN), .B2(keyinput225), .ZN(n10155) );
  OAI221_X1 U11243 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(keyinput182), .C1(
        P1_IR_REG_7__SCAN_IN), .C2(keyinput225), .A(n10155), .ZN(n10158) );
  AOI22_X1 U11244 ( .A1(P2_D_REG_11__SCAN_IN), .A2(keyinput234), .B1(
        P1_REG1_REG_0__SCAN_IN), .B2(keyinput249), .ZN(n10156) );
  OAI221_X1 U11245 ( .B1(P2_D_REG_11__SCAN_IN), .B2(keyinput234), .C1(
        P1_REG1_REG_0__SCAN_IN), .C2(keyinput249), .A(n10156), .ZN(n10157) );
  NOR4_X1 U11246 ( .A1(n10160), .A2(n10159), .A3(n10158), .A4(n10157), .ZN(
        n10161) );
  NAND4_X1 U11247 ( .A1(n10164), .A2(n10163), .A3(n10162), .A4(n10161), .ZN(
        n10306) );
  AOI22_X1 U11248 ( .A1(P2_REG1_REG_2__SCAN_IN), .A2(keyinput233), .B1(
        P1_REG2_REG_16__SCAN_IN), .B2(keyinput129), .ZN(n10165) );
  OAI221_X1 U11249 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(keyinput233), .C1(
        P1_REG2_REG_16__SCAN_IN), .C2(keyinput129), .A(n10165), .ZN(n10172) );
  AOI22_X1 U11250 ( .A1(SI_15_), .A2(keyinput248), .B1(P1_IR_REG_25__SCAN_IN), 
        .B2(keyinput171), .ZN(n10166) );
  OAI221_X1 U11251 ( .B1(SI_15_), .B2(keyinput248), .C1(P1_IR_REG_25__SCAN_IN), 
        .C2(keyinput171), .A(n10166), .ZN(n10171) );
  AOI22_X1 U11252 ( .A1(P2_REG0_REG_1__SCAN_IN), .A2(keyinput148), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(keyinput224), .ZN(n10167) );
  OAI221_X1 U11253 ( .B1(P2_REG0_REG_1__SCAN_IN), .B2(keyinput148), .C1(
        P1_DATAO_REG_13__SCAN_IN), .C2(keyinput224), .A(n10167), .ZN(n10170)
         );
  AOI22_X1 U11254 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(keyinput215), .B1(
        P1_REG0_REG_7__SCAN_IN), .B2(keyinput165), .ZN(n10168) );
  OAI221_X1 U11255 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(keyinput215), .C1(
        P1_REG0_REG_7__SCAN_IN), .C2(keyinput165), .A(n10168), .ZN(n10169) );
  NOR4_X1 U11256 ( .A1(n10172), .A2(n10171), .A3(n10170), .A4(n10169), .ZN(
        n10202) );
  AOI22_X1 U11257 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(keyinput202), .B1(SI_16_), 
        .B2(keyinput157), .ZN(n10173) );
  OAI221_X1 U11258 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(keyinput202), .C1(SI_16_), .C2(keyinput157), .A(n10173), .ZN(n10180) );
  AOI22_X1 U11259 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(keyinput174), .B1(
        P1_REG2_REG_23__SCAN_IN), .B2(keyinput207), .ZN(n10174) );
  OAI221_X1 U11260 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(keyinput174), .C1(
        P1_REG2_REG_23__SCAN_IN), .C2(keyinput207), .A(n10174), .ZN(n10179) );
  AOI22_X1 U11261 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput163), .B1(
        P1_D_REG_5__SCAN_IN), .B2(keyinput149), .ZN(n10175) );
  OAI221_X1 U11262 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput163), .C1(
        P1_D_REG_5__SCAN_IN), .C2(keyinput149), .A(n10175), .ZN(n10178) );
  AOI22_X1 U11263 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(keyinput217), .B1(
        P2_D_REG_0__SCAN_IN), .B2(keyinput205), .ZN(n10176) );
  OAI221_X1 U11264 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(keyinput217), .C1(
        P2_D_REG_0__SCAN_IN), .C2(keyinput205), .A(n10176), .ZN(n10177) );
  NOR4_X1 U11265 ( .A1(n10180), .A2(n10179), .A3(n10178), .A4(n10177), .ZN(
        n10201) );
  AOI22_X1 U11266 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(keyinput135), .B1(
        P1_REG1_REG_18__SCAN_IN), .B2(keyinput177), .ZN(n10181) );
  OAI221_X1 U11267 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(keyinput135), .C1(
        P1_REG1_REG_18__SCAN_IN), .C2(keyinput177), .A(n10181), .ZN(n10188) );
  AOI22_X1 U11268 ( .A1(P2_REG2_REG_23__SCAN_IN), .A2(keyinput136), .B1(
        P1_REG0_REG_4__SCAN_IN), .B2(keyinput203), .ZN(n10182) );
  OAI221_X1 U11269 ( .B1(P2_REG2_REG_23__SCAN_IN), .B2(keyinput136), .C1(
        P1_REG0_REG_4__SCAN_IN), .C2(keyinput203), .A(n10182), .ZN(n10187) );
  AOI22_X1 U11270 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(keyinput159), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(keyinput190), .ZN(n10183) );
  OAI221_X1 U11271 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(keyinput159), .C1(
        P1_ADDR_REG_13__SCAN_IN), .C2(keyinput190), .A(n10183), .ZN(n10186) );
  AOI22_X1 U11272 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(keyinput235), .B1(
        P1_REG1_REG_28__SCAN_IN), .B2(keyinput180), .ZN(n10184) );
  OAI221_X1 U11273 ( .B1(P2_IR_REG_22__SCAN_IN), .B2(keyinput235), .C1(
        P1_REG1_REG_28__SCAN_IN), .C2(keyinput180), .A(n10184), .ZN(n10185) );
  NOR4_X1 U11274 ( .A1(n10188), .A2(n10187), .A3(n10186), .A4(n10185), .ZN(
        n10200) );
  AOI22_X1 U11275 ( .A1(n10369), .A2(keyinput253), .B1(keyinput175), .B2(
        n10190), .ZN(n10189) );
  OAI221_X1 U11276 ( .B1(n10369), .B2(keyinput253), .C1(n10190), .C2(
        keyinput175), .A(n10189), .ZN(n10198) );
  AOI22_X1 U11277 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(keyinput184), .B1(
        P1_REG3_REG_17__SCAN_IN), .B2(keyinput186), .ZN(n10191) );
  OAI221_X1 U11278 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(keyinput184), .C1(
        P1_REG3_REG_17__SCAN_IN), .C2(keyinput186), .A(n10191), .ZN(n10197) );
  AOI22_X1 U11279 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(keyinput254), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(keyinput130), .ZN(n10192) );
  OAI221_X1 U11280 ( .B1(P1_REG3_REG_13__SCAN_IN), .B2(keyinput254), .C1(
        P1_DATAO_REG_22__SCAN_IN), .C2(keyinput130), .A(n10192), .ZN(n10196)
         );
  XNOR2_X1 U11281 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput213), .ZN(n10194)
         );
  XNOR2_X1 U11282 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput137), .ZN(n10193)
         );
  NAND2_X1 U11283 ( .A1(n10194), .A2(n10193), .ZN(n10195) );
  NOR4_X1 U11284 ( .A1(n10198), .A2(n10197), .A3(n10196), .A4(n10195), .ZN(
        n10199) );
  NAND4_X1 U11285 ( .A1(n10202), .A2(n10201), .A3(n10200), .A4(n10199), .ZN(
        n10305) );
  AOI22_X1 U11286 ( .A1(n6782), .A2(keyinput181), .B1(keyinput134), .B2(n10365), .ZN(n10203) );
  OAI221_X1 U11287 ( .B1(n6782), .B2(keyinput181), .C1(n10365), .C2(
        keyinput134), .A(n10203), .ZN(n10215) );
  AOI22_X1 U11288 ( .A1(n10206), .A2(keyinput194), .B1(n10205), .B2(
        keyinput166), .ZN(n10204) );
  OAI221_X1 U11289 ( .B1(n10206), .B2(keyinput194), .C1(n10205), .C2(
        keyinput166), .A(n10204), .ZN(n10214) );
  INV_X1 U11290 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10209) );
  AOI22_X1 U11291 ( .A1(n10209), .A2(keyinput162), .B1(keyinput232), .B2(
        n10208), .ZN(n10207) );
  OAI221_X1 U11292 ( .B1(n10209), .B2(keyinput162), .C1(n10208), .C2(
        keyinput232), .A(n10207), .ZN(n10213) );
  XNOR2_X1 U11293 ( .A(P1_REG0_REG_27__SCAN_IN), .B(keyinput221), .ZN(n10211)
         );
  XNOR2_X1 U11294 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput155), .ZN(n10210) );
  NAND2_X1 U11295 ( .A1(n10211), .A2(n10210), .ZN(n10212) );
  NOR4_X1 U11296 ( .A1(n10215), .A2(n10214), .A3(n10213), .A4(n10212), .ZN(
        n10251) );
  AOI22_X1 U11297 ( .A1(n10218), .A2(keyinput204), .B1(n10217), .B2(
        keyinput153), .ZN(n10216) );
  OAI221_X1 U11298 ( .B1(n10218), .B2(keyinput204), .C1(n10217), .C2(
        keyinput153), .A(n10216), .ZN(n10226) );
  AOI22_X1 U11299 ( .A1(n10395), .A2(keyinput208), .B1(keyinput156), .B2(
        n10408), .ZN(n10219) );
  OAI221_X1 U11300 ( .B1(n10395), .B2(keyinput208), .C1(n10408), .C2(
        keyinput156), .A(n10219), .ZN(n10225) );
  AOI22_X1 U11301 ( .A1(n8344), .A2(keyinput219), .B1(keyinput151), .B2(n7813), 
        .ZN(n10220) );
  OAI221_X1 U11302 ( .B1(n8344), .B2(keyinput219), .C1(n7813), .C2(keyinput151), .A(n10220), .ZN(n10224) );
  AOI22_X1 U11303 ( .A1(n5652), .A2(keyinput170), .B1(keyinput250), .B2(n10222), .ZN(n10221) );
  OAI221_X1 U11304 ( .B1(n5652), .B2(keyinput170), .C1(n10222), .C2(
        keyinput250), .A(n10221), .ZN(n10223) );
  NOR4_X1 U11305 ( .A1(n10226), .A2(n10225), .A3(n10224), .A4(n10223), .ZN(
        n10250) );
  AOI22_X1 U11306 ( .A1(n9314), .A2(keyinput179), .B1(keyinput167), .B2(n6038), 
        .ZN(n10227) );
  OAI221_X1 U11307 ( .B1(n9314), .B2(keyinput179), .C1(n6038), .C2(keyinput167), .A(n10227), .ZN(n10236) );
  AOI22_X1 U11308 ( .A1(n10318), .A2(keyinput161), .B1(n10370), .B2(
        keyinput172), .ZN(n10228) );
  OAI221_X1 U11309 ( .B1(n10318), .B2(keyinput161), .C1(n10370), .C2(
        keyinput172), .A(n10228), .ZN(n10235) );
  AOI22_X1 U11310 ( .A1(n10383), .A2(keyinput199), .B1(n10230), .B2(
        keyinput242), .ZN(n10229) );
  OAI221_X1 U11311 ( .B1(n10383), .B2(keyinput199), .C1(n10230), .C2(
        keyinput242), .A(n10229), .ZN(n10234) );
  XOR2_X1 U11312 ( .A(n5260), .B(keyinput196), .Z(n10232) );
  XNOR2_X1 U11313 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput132), .ZN(n10231)
         );
  NAND2_X1 U11314 ( .A1(n10232), .A2(n10231), .ZN(n10233) );
  NOR4_X1 U11315 ( .A1(n10236), .A2(n10235), .A3(n10234), .A4(n10233), .ZN(
        n10249) );
  AOI22_X1 U11316 ( .A1(n10238), .A2(keyinput255), .B1(keyinput201), .B2(
        n10322), .ZN(n10237) );
  OAI221_X1 U11317 ( .B1(n10238), .B2(keyinput255), .C1(n10322), .C2(
        keyinput201), .A(n10237), .ZN(n10247) );
  INV_X1 U11318 ( .A(SI_29_), .ZN(n10332) );
  INV_X1 U11319 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10240) );
  AOI22_X1 U11320 ( .A1(n10332), .A2(keyinput143), .B1(n10240), .B2(
        keyinput189), .ZN(n10239) );
  OAI221_X1 U11321 ( .B1(n10332), .B2(keyinput143), .C1(n10240), .C2(
        keyinput189), .A(n10239), .ZN(n10246) );
  AOI22_X1 U11322 ( .A1(n6013), .A2(keyinput158), .B1(n10410), .B2(keyinput142), .ZN(n10241) );
  OAI221_X1 U11323 ( .B1(n6013), .B2(keyinput158), .C1(n10410), .C2(
        keyinput142), .A(n10241), .ZN(n10245) );
  AOI22_X1 U11324 ( .A1(n10243), .A2(keyinput191), .B1(n6768), .B2(keyinput231), .ZN(n10242) );
  OAI221_X1 U11325 ( .B1(n10243), .B2(keyinput191), .C1(n6768), .C2(
        keyinput231), .A(n10242), .ZN(n10244) );
  NOR4_X1 U11326 ( .A1(n10247), .A2(n10246), .A3(n10245), .A4(n10244), .ZN(
        n10248) );
  NAND4_X1 U11327 ( .A1(n10251), .A2(n10250), .A3(n10249), .A4(n10248), .ZN(
        n10304) );
  INV_X1 U11328 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n10312) );
  AOI22_X1 U11329 ( .A1(n6411), .A2(keyinput188), .B1(keyinput147), .B2(n10312), .ZN(n10252) );
  OAI221_X1 U11330 ( .B1(n6411), .B2(keyinput188), .C1(n10312), .C2(
        keyinput147), .A(n10252), .ZN(n10262) );
  INV_X1 U11331 ( .A(SI_18_), .ZN(n10254) );
  AOI22_X1 U11332 ( .A1(n10323), .A2(keyinput240), .B1(n10254), .B2(
        keyinput230), .ZN(n10253) );
  OAI221_X1 U11333 ( .B1(n10323), .B2(keyinput240), .C1(n10254), .C2(
        keyinput230), .A(n10253), .ZN(n10261) );
  AOI22_X1 U11334 ( .A1(n10257), .A2(keyinput176), .B1(n10256), .B2(
        keyinput146), .ZN(n10255) );
  OAI221_X1 U11335 ( .B1(n10257), .B2(keyinput176), .C1(n10256), .C2(
        keyinput146), .A(n10255), .ZN(n10260) );
  AOI22_X1 U11336 ( .A1(n6258), .A2(keyinput210), .B1(n10333), .B2(keyinput152), .ZN(n10258) );
  OAI221_X1 U11337 ( .B1(n6258), .B2(keyinput210), .C1(n10333), .C2(
        keyinput152), .A(n10258), .ZN(n10259) );
  NOR4_X1 U11338 ( .A1(n10262), .A2(n10261), .A3(n10260), .A4(n10259), .ZN(
        n10302) );
  AOI22_X1 U11339 ( .A1(n10265), .A2(keyinput200), .B1(keyinput211), .B2(
        n10264), .ZN(n10263) );
  OAI221_X1 U11340 ( .B1(n10265), .B2(keyinput200), .C1(n10264), .C2(
        keyinput211), .A(n10263), .ZN(n10275) );
  AOI22_X1 U11341 ( .A1(n10267), .A2(keyinput247), .B1(keyinput218), .B2(
        n10310), .ZN(n10266) );
  OAI221_X1 U11342 ( .B1(n10267), .B2(keyinput247), .C1(n10310), .C2(
        keyinput218), .A(n10266), .ZN(n10274) );
  AOI22_X1 U11343 ( .A1(n10269), .A2(keyinput164), .B1(keyinput220), .B2(
        n10347), .ZN(n10268) );
  OAI221_X1 U11344 ( .B1(n10269), .B2(keyinput164), .C1(n10347), .C2(
        keyinput220), .A(n10268), .ZN(n10273) );
  AOI22_X1 U11345 ( .A1(n10271), .A2(keyinput228), .B1(keyinput227), .B2(n6703), .ZN(n10270) );
  OAI221_X1 U11346 ( .B1(n10271), .B2(keyinput228), .C1(n6703), .C2(
        keyinput227), .A(n10270), .ZN(n10272) );
  NOR4_X1 U11347 ( .A1(n10275), .A2(n10274), .A3(n10273), .A4(n10272), .ZN(
        n10301) );
  AOI22_X1 U11348 ( .A1(n10277), .A2(keyinput252), .B1(keyinput169), .B2(n7460), .ZN(n10276) );
  OAI221_X1 U11349 ( .B1(n10277), .B2(keyinput252), .C1(n7460), .C2(
        keyinput169), .A(n10276), .ZN(n10287) );
  AOI22_X1 U11350 ( .A1(n10279), .A2(keyinput178), .B1(n9695), .B2(keyinput239), .ZN(n10278) );
  OAI221_X1 U11351 ( .B1(n10279), .B2(keyinput178), .C1(n9695), .C2(
        keyinput239), .A(n10278), .ZN(n10286) );
  AOI22_X1 U11352 ( .A1(n10352), .A2(keyinput197), .B1(n10321), .B2(
        keyinput141), .ZN(n10280) );
  OAI221_X1 U11353 ( .B1(n10352), .B2(keyinput197), .C1(n10321), .C2(
        keyinput141), .A(n10280), .ZN(n10285) );
  AOI22_X1 U11354 ( .A1(n10283), .A2(keyinput238), .B1(n10282), .B2(
        keyinput223), .ZN(n10281) );
  OAI221_X1 U11355 ( .B1(n10283), .B2(keyinput238), .C1(n10282), .C2(
        keyinput223), .A(n10281), .ZN(n10284) );
  NOR4_X1 U11356 ( .A1(n10287), .A2(n10286), .A3(n10285), .A4(n10284), .ZN(
        n10300) );
  INV_X1 U11357 ( .A(SI_6_), .ZN(n10380) );
  AOI22_X1 U11358 ( .A1(n10380), .A2(keyinput195), .B1(keyinput144), .B2(
        n10348), .ZN(n10288) );
  OAI221_X1 U11359 ( .B1(n10380), .B2(keyinput195), .C1(n10348), .C2(
        keyinput144), .A(n10288), .ZN(n10298) );
  AOI22_X1 U11360 ( .A1(n10290), .A2(keyinput237), .B1(keyinput187), .B2(
        n10394), .ZN(n10289) );
  OAI221_X1 U11361 ( .B1(n10290), .B2(keyinput237), .C1(n10394), .C2(
        keyinput187), .A(n10289), .ZN(n10297) );
  INV_X1 U11362 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n10292) );
  AOI22_X1 U11363 ( .A1(n10292), .A2(keyinput185), .B1(n5411), .B2(keyinput145), .ZN(n10291) );
  OAI221_X1 U11364 ( .B1(n10292), .B2(keyinput185), .C1(n5411), .C2(
        keyinput145), .A(n10291), .ZN(n10296) );
  AOI22_X1 U11365 ( .A1(n10335), .A2(keyinput183), .B1(keyinput244), .B2(
        n10294), .ZN(n10293) );
  OAI221_X1 U11366 ( .B1(n10335), .B2(keyinput183), .C1(n10294), .C2(
        keyinput244), .A(n10293), .ZN(n10295) );
  NOR4_X1 U11367 ( .A1(n10298), .A2(n10297), .A3(n10296), .A4(n10295), .ZN(
        n10299) );
  NAND4_X1 U11368 ( .A1(n10302), .A2(n10301), .A3(n10300), .A4(n10299), .ZN(
        n10303) );
  NOR4_X1 U11369 ( .A1(n10306), .A2(n10305), .A3(n10304), .A4(n10303), .ZN(
        n10499) );
  AOI22_X1 U11370 ( .A1(P1_REG0_REG_4__SCAN_IN), .A2(keyinput75), .B1(
        P1_IR_REG_13__SCAN_IN), .B2(keyinput27), .ZN(n10307) );
  OAI221_X1 U11371 ( .B1(P1_REG0_REG_4__SCAN_IN), .B2(keyinput75), .C1(
        P1_IR_REG_13__SCAN_IN), .C2(keyinput27), .A(n10307), .ZN(n10316) );
  AOI22_X1 U11372 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(keyinput26), .B1(
        P1_REG3_REG_20__SCAN_IN), .B2(keyinput42), .ZN(n10308) );
  OAI221_X1 U11373 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(keyinput26), .C1(
        P1_REG3_REG_20__SCAN_IN), .C2(keyinput42), .A(n10308), .ZN(n10315) );
  AOI22_X1 U11374 ( .A1(P2_REG0_REG_16__SCAN_IN), .A2(keyinput82), .B1(n10310), 
        .B2(keyinput90), .ZN(n10309) );
  OAI221_X1 U11375 ( .B1(P2_REG0_REG_16__SCAN_IN), .B2(keyinput82), .C1(n10310), .C2(keyinput90), .A(n10309), .ZN(n10314) );
  AOI22_X1 U11376 ( .A1(n10312), .A2(keyinput19), .B1(keyinput32), .B2(n10510), 
        .ZN(n10311) );
  OAI221_X1 U11377 ( .B1(n10312), .B2(keyinput19), .C1(n10510), .C2(keyinput32), .A(n10311), .ZN(n10313) );
  NOR4_X1 U11378 ( .A1(n10316), .A2(n10315), .A3(n10314), .A4(n10313), .ZN(
        n10363) );
  INV_X1 U11379 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U11380 ( .A1(n10319), .A2(keyinput46), .B1(n10318), .B2(keyinput33), 
        .ZN(n10317) );
  OAI221_X1 U11381 ( .B1(n10319), .B2(keyinput46), .C1(n10318), .C2(keyinput33), .A(n10317), .ZN(n10330) );
  AOI22_X1 U11382 ( .A1(n10322), .A2(keyinput73), .B1(n10321), .B2(keyinput13), 
        .ZN(n10320) );
  OAI221_X1 U11383 ( .B1(n10322), .B2(keyinput73), .C1(n10321), .C2(keyinput13), .A(n10320), .ZN(n10329) );
  XNOR2_X1 U11384 ( .A(n10323), .B(keyinput112), .ZN(n10328) );
  XNOR2_X1 U11385 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput85), .ZN(n10326)
         );
  XNOR2_X1 U11386 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput98), .ZN(n10325) );
  XNOR2_X1 U11387 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(keyinput109), .ZN(n10324)
         );
  NAND3_X1 U11388 ( .A1(n10326), .A2(n10325), .A3(n10324), .ZN(n10327) );
  NOR4_X1 U11389 ( .A1(n10330), .A2(n10329), .A3(n10328), .A4(n10327), .ZN(
        n10362) );
  AOI22_X1 U11390 ( .A1(n10333), .A2(keyinput24), .B1(keyinput15), .B2(n10332), 
        .ZN(n10331) );
  OAI221_X1 U11391 ( .B1(n10333), .B2(keyinput24), .C1(n10332), .C2(keyinput15), .A(n10331), .ZN(n10345) );
  AOI22_X1 U11392 ( .A1(n10336), .A2(keyinput77), .B1(n10335), .B2(keyinput55), 
        .ZN(n10334) );
  OAI221_X1 U11393 ( .B1(n10336), .B2(keyinput77), .C1(n10335), .C2(keyinput55), .A(n10334), .ZN(n10344) );
  AOI22_X1 U11394 ( .A1(n6795), .A2(keyinput89), .B1(n10338), .B2(keyinput29), 
        .ZN(n10337) );
  OAI221_X1 U11395 ( .B1(n6795), .B2(keyinput89), .C1(n10338), .C2(keyinput29), 
        .A(n10337), .ZN(n10343) );
  AOI22_X1 U11396 ( .A1(n10341), .A2(keyinput2), .B1(keyinput40), .B2(n10340), 
        .ZN(n10339) );
  OAI221_X1 U11397 ( .B1(n10341), .B2(keyinput2), .C1(n10340), .C2(keyinput40), 
        .A(n10339), .ZN(n10342) );
  NOR4_X1 U11398 ( .A1(n10345), .A2(n10344), .A3(n10343), .A4(n10342), .ZN(
        n10361) );
  AOI22_X1 U11399 ( .A1(n10348), .A2(keyinput16), .B1(keyinput92), .B2(n10347), 
        .ZN(n10346) );
  OAI221_X1 U11400 ( .B1(n10348), .B2(keyinput16), .C1(n10347), .C2(keyinput92), .A(n10346), .ZN(n10359) );
  AOI22_X1 U11401 ( .A1(n10350), .A2(keyinput65), .B1(n9314), .B2(keyinput51), 
        .ZN(n10349) );
  OAI221_X1 U11402 ( .B1(n10350), .B2(keyinput65), .C1(n9314), .C2(keyinput51), 
        .A(n10349), .ZN(n10358) );
  AOI22_X1 U11403 ( .A1(n10353), .A2(keyinput106), .B1(keyinput69), .B2(n10352), .ZN(n10351) );
  OAI221_X1 U11404 ( .B1(n10353), .B2(keyinput106), .C1(n10352), .C2(
        keyinput69), .A(n10351), .ZN(n10357) );
  XOR2_X1 U11405 ( .A(n5260), .B(keyinput68), .Z(n10355) );
  XNOR2_X1 U11406 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput84), .ZN(n10354) );
  NAND2_X1 U11407 ( .A1(n10355), .A2(n10354), .ZN(n10356) );
  NOR4_X1 U11408 ( .A1(n10359), .A2(n10358), .A3(n10357), .A4(n10356), .ZN(
        n10360) );
  NAND4_X1 U11409 ( .A1(n10363), .A2(n10362), .A3(n10361), .A4(n10360), .ZN(
        n10498) );
  AOI22_X1 U11410 ( .A1(n7460), .A2(keyinput41), .B1(keyinput6), .B2(n10365), 
        .ZN(n10364) );
  OAI221_X1 U11411 ( .B1(n7460), .B2(keyinput41), .C1(n10365), .C2(keyinput6), 
        .A(n10364), .ZN(n10376) );
  INV_X1 U11412 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10367) );
  AOI22_X1 U11413 ( .A1(n10367), .A2(keyinput11), .B1(n6764), .B2(keyinput22), 
        .ZN(n10366) );
  OAI221_X1 U11414 ( .B1(n10367), .B2(keyinput11), .C1(n6764), .C2(keyinput22), 
        .A(n10366), .ZN(n10375) );
  AOI22_X1 U11415 ( .A1(n10370), .A2(keyinput44), .B1(n10369), .B2(keyinput125), .ZN(n10368) );
  OAI221_X1 U11416 ( .B1(n10370), .B2(keyinput44), .C1(n10369), .C2(
        keyinput125), .A(n10368), .ZN(n10374) );
  XNOR2_X1 U11417 ( .A(P2_REG0_REG_21__SCAN_IN), .B(keyinput122), .ZN(n10372)
         );
  XNOR2_X1 U11418 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput43), .ZN(n10371) );
  NAND2_X1 U11419 ( .A1(n10372), .A2(n10371), .ZN(n10373) );
  NOR4_X1 U11420 ( .A1(n10376), .A2(n10375), .A3(n10374), .A4(n10373), .ZN(
        n10421) );
  AOI22_X1 U11421 ( .A1(n10378), .A2(keyinput78), .B1(n5298), .B2(keyinput37), 
        .ZN(n10377) );
  OAI221_X1 U11422 ( .B1(n10378), .B2(keyinput78), .C1(n5298), .C2(keyinput37), 
        .A(n10377), .ZN(n10388) );
  AOI22_X1 U11423 ( .A1(n10381), .A2(keyinput12), .B1(n10380), .B2(keyinput67), 
        .ZN(n10379) );
  OAI221_X1 U11424 ( .B1(n10381), .B2(keyinput12), .C1(n10380), .C2(keyinput67), .A(n10379), .ZN(n10387) );
  AOI22_X1 U11425 ( .A1(n7614), .A2(keyinput87), .B1(n10383), .B2(keyinput71), 
        .ZN(n10382) );
  OAI221_X1 U11426 ( .B1(n7614), .B2(keyinput87), .C1(n10383), .C2(keyinput71), 
        .A(n10382), .ZN(n10386) );
  AOI22_X1 U11427 ( .A1(n5971), .A2(keyinput20), .B1(n9695), .B2(keyinput111), 
        .ZN(n10384) );
  OAI221_X1 U11428 ( .B1(n5971), .B2(keyinput20), .C1(n9695), .C2(keyinput111), 
        .A(n10384), .ZN(n10385) );
  NOR4_X1 U11429 ( .A1(n10388), .A2(n10387), .A3(n10386), .A4(n10385), .ZN(
        n10420) );
  AOI22_X1 U11430 ( .A1(n10391), .A2(keyinput86), .B1(keyinput115), .B2(n10390), .ZN(n10389) );
  OAI221_X1 U11431 ( .B1(n10391), .B2(keyinput86), .C1(n10390), .C2(
        keyinput115), .A(n10389), .ZN(n10402) );
  AOI22_X1 U11432 ( .A1(n6768), .A2(keyinput103), .B1(keyinput8), .B2(n8909), 
        .ZN(n10392) );
  OAI221_X1 U11433 ( .B1(n6768), .B2(keyinput103), .C1(n8909), .C2(keyinput8), 
        .A(n10392), .ZN(n10401) );
  AOI22_X1 U11434 ( .A1(n10395), .A2(keyinput80), .B1(n10394), .B2(keyinput59), 
        .ZN(n10393) );
  OAI221_X1 U11435 ( .B1(n10395), .B2(keyinput80), .C1(n10394), .C2(keyinput59), .A(n10393), .ZN(n10400) );
  AOI22_X1 U11436 ( .A1(n10398), .A2(keyinput10), .B1(n10397), .B2(keyinput52), 
        .ZN(n10396) );
  OAI221_X1 U11437 ( .B1(n10398), .B2(keyinput10), .C1(n10397), .C2(keyinput52), .A(n10396), .ZN(n10399) );
  NOR4_X1 U11438 ( .A1(n10402), .A2(n10401), .A3(n10400), .A4(n10399), .ZN(
        n10419) );
  AOI22_X1 U11439 ( .A1(n10405), .A2(keyinput93), .B1(keyinput88), .B2(n10404), 
        .ZN(n10403) );
  OAI221_X1 U11440 ( .B1(n10405), .B2(keyinput93), .C1(n10404), .C2(keyinput88), .A(n10403), .ZN(n10417) );
  AOI22_X1 U11441 ( .A1(n10408), .A2(keyinput28), .B1(n10407), .B2(keyinput121), .ZN(n10406) );
  OAI221_X1 U11442 ( .B1(n10408), .B2(keyinput28), .C1(n10407), .C2(
        keyinput121), .A(n10406), .ZN(n10416) );
  AOI22_X1 U11443 ( .A1(n10410), .A2(keyinput14), .B1(keyinput39), .B2(n6038), 
        .ZN(n10409) );
  OAI221_X1 U11444 ( .B1(n10410), .B2(keyinput14), .C1(n6038), .C2(keyinput39), 
        .A(n10409), .ZN(n10415) );
  AOI22_X1 U11445 ( .A1(n10413), .A2(keyinput0), .B1(keyinput62), .B2(n10412), 
        .ZN(n10411) );
  OAI221_X1 U11446 ( .B1(n10413), .B2(keyinput0), .C1(n10412), .C2(keyinput62), 
        .A(n10411), .ZN(n10414) );
  NOR4_X1 U11447 ( .A1(n10417), .A2(n10416), .A3(n10415), .A4(n10414), .ZN(
        n10418) );
  NAND4_X1 U11448 ( .A1(n10421), .A2(n10420), .A3(n10419), .A4(n10418), .ZN(
        n10497) );
  OAI22_X1 U11449 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(keyinput74), .B1(
        P2_IR_REG_25__SCAN_IN), .B2(keyinput48), .ZN(n10422) );
  AOI221_X1 U11450 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(keyinput74), .C1(
        keyinput48), .C2(P2_IR_REG_25__SCAN_IN), .A(n10422), .ZN(n10429) );
  OAI22_X1 U11451 ( .A1(SI_27_), .A2(keyinput119), .B1(keyinput76), .B2(
        P1_DATAO_REG_23__SCAN_IN), .ZN(n10423) );
  AOI221_X1 U11452 ( .B1(SI_27_), .B2(keyinput119), .C1(
        P1_DATAO_REG_23__SCAN_IN), .C2(keyinput76), .A(n10423), .ZN(n10428) );
  OAI22_X1 U11453 ( .A1(P1_D_REG_5__SCAN_IN), .A2(keyinput21), .B1(
        P1_REG2_REG_16__SCAN_IN), .B2(keyinput1), .ZN(n10424) );
  AOI221_X1 U11454 ( .B1(P1_D_REG_5__SCAN_IN), .B2(keyinput21), .C1(keyinput1), 
        .C2(P1_REG2_REG_16__SCAN_IN), .A(n10424), .ZN(n10427) );
  OAI22_X1 U11455 ( .A1(P2_D_REG_10__SCAN_IN), .A2(keyinput47), .B1(
        P2_REG2_REG_16__SCAN_IN), .B2(keyinput57), .ZN(n10425) );
  AOI221_X1 U11456 ( .B1(P2_D_REG_10__SCAN_IN), .B2(keyinput47), .C1(
        keyinput57), .C2(P2_REG2_REG_16__SCAN_IN), .A(n10425), .ZN(n10426) );
  NAND4_X1 U11457 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10457) );
  OAI22_X1 U11458 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(keyinput25), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(keyinput3), .ZN(n10430) );
  AOI221_X1 U11459 ( .B1(P2_DATAO_REG_25__SCAN_IN), .B2(keyinput25), .C1(
        keyinput3), .C2(P1_DATAO_REG_19__SCAN_IN), .A(n10430), .ZN(n10437) );
  OAI22_X1 U11460 ( .A1(P1_REG1_REG_14__SCAN_IN), .A2(keyinput110), .B1(
        keyinput53), .B2(P1_REG2_REG_4__SCAN_IN), .ZN(n10431) );
  AOI221_X1 U11461 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(keyinput110), .C1(
        P1_REG2_REG_4__SCAN_IN), .C2(keyinput53), .A(n10431), .ZN(n10436) );
  OAI22_X1 U11462 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(keyinput4), .B1(
        keyinput117), .B2(P2_IR_REG_12__SCAN_IN), .ZN(n10432) );
  AOI221_X1 U11463 ( .B1(P1_DATAO_REG_4__SCAN_IN), .B2(keyinput4), .C1(
        P2_IR_REG_12__SCAN_IN), .C2(keyinput117), .A(n10432), .ZN(n10435) );
  OAI22_X1 U11464 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(keyinput96), .B1(
        keyinput79), .B2(P1_REG2_REG_23__SCAN_IN), .ZN(n10433) );
  AOI221_X1 U11465 ( .B1(P1_DATAO_REG_13__SCAN_IN), .B2(keyinput96), .C1(
        P1_REG2_REG_23__SCAN_IN), .C2(keyinput79), .A(n10433), .ZN(n10434) );
  NAND4_X1 U11466 ( .A1(n10437), .A2(n10436), .A3(n10435), .A4(n10434), .ZN(
        n10456) );
  OAI22_X1 U11467 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(keyinput23), .B1(
        keyinput118), .B2(P2_DATAO_REG_31__SCAN_IN), .ZN(n10438) );
  AOI221_X1 U11468 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(keyinput23), .C1(
        P2_DATAO_REG_31__SCAN_IN), .C2(keyinput118), .A(n10438), .ZN(n10445)
         );
  OAI22_X1 U11469 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput34), .B1(keyinput56), 
        .B2(P1_ADDR_REG_10__SCAN_IN), .ZN(n10439) );
  AOI221_X1 U11470 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput34), .C1(
        P1_ADDR_REG_10__SCAN_IN), .C2(keyinput56), .A(n10439), .ZN(n10444) );
  OAI22_X1 U11471 ( .A1(P1_D_REG_13__SCAN_IN), .A2(keyinput94), .B1(
        P2_REG0_REG_30__SCAN_IN), .B2(keyinput36), .ZN(n10440) );
  AOI221_X1 U11472 ( .B1(P1_D_REG_13__SCAN_IN), .B2(keyinput94), .C1(
        keyinput36), .C2(P2_REG0_REG_30__SCAN_IN), .A(n10440), .ZN(n10443) );
  OAI22_X1 U11473 ( .A1(P2_D_REG_9__SCAN_IN), .A2(keyinput116), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput35), .ZN(n10441) );
  AOI221_X1 U11474 ( .B1(P2_D_REG_9__SCAN_IN), .B2(keyinput116), .C1(
        keyinput35), .C2(P2_REG3_REG_26__SCAN_IN), .A(n10441), .ZN(n10442) );
  NAND4_X1 U11475 ( .A1(n10445), .A2(n10444), .A3(n10443), .A4(n10442), .ZN(
        n10455) );
  OAI22_X1 U11476 ( .A1(SI_10_), .A2(keyinput127), .B1(keyinput58), .B2(
        P1_REG3_REG_17__SCAN_IN), .ZN(n10446) );
  AOI221_X1 U11477 ( .B1(SI_10_), .B2(keyinput127), .C1(
        P1_REG3_REG_17__SCAN_IN), .C2(keyinput58), .A(n10446), .ZN(n10453) );
  OAI22_X1 U11478 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(keyinput7), .B1(
        keyinput18), .B2(P1_REG1_REG_2__SCAN_IN), .ZN(n10447) );
  AOI221_X1 U11479 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(keyinput7), .C1(
        P1_REG1_REG_2__SCAN_IN), .C2(keyinput18), .A(n10447), .ZN(n10452) );
  OAI22_X1 U11480 ( .A1(P1_D_REG_30__SCAN_IN), .A2(keyinput124), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(keyinput9), .ZN(n10448) );
  AOI221_X1 U11481 ( .B1(P1_D_REG_30__SCAN_IN), .B2(keyinput124), .C1(
        keyinput9), .C2(P1_DATAO_REG_1__SCAN_IN), .A(n10448), .ZN(n10451) );
  OAI22_X1 U11482 ( .A1(P2_D_REG_21__SCAN_IN), .A2(keyinput61), .B1(
        keyinput104), .B2(P2_D_REG_23__SCAN_IN), .ZN(n10449) );
  AOI221_X1 U11483 ( .B1(P2_D_REG_21__SCAN_IN), .B2(keyinput61), .C1(
        P2_D_REG_23__SCAN_IN), .C2(keyinput104), .A(n10449), .ZN(n10450) );
  NAND4_X1 U11484 ( .A1(n10453), .A2(n10452), .A3(n10451), .A4(n10450), .ZN(
        n10454) );
  NOR4_X1 U11485 ( .A1(n10457), .A2(n10456), .A3(n10455), .A4(n10454), .ZN(
        n10495) );
  OAI22_X1 U11486 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(keyinput70), .B1(
        keyinput45), .B2(P2_REG3_REG_28__SCAN_IN), .ZN(n10458) );
  AOI221_X1 U11487 ( .B1(P1_REG3_REG_15__SCAN_IN), .B2(keyinput70), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput45), .A(n10458), .ZN(n10465) );
  OAI22_X1 U11488 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(keyinput49), .B1(
        P2_REG0_REG_2__SCAN_IN), .B2(keyinput30), .ZN(n10459) );
  AOI221_X1 U11489 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(keyinput49), .C1(
        keyinput30), .C2(P2_REG0_REG_2__SCAN_IN), .A(n10459), .ZN(n10464) );
  OAI22_X1 U11490 ( .A1(P1_B_REG_SCAN_IN), .A2(keyinput91), .B1(
        P2_REG1_REG_21__SCAN_IN), .B2(keyinput100), .ZN(n10460) );
  AOI221_X1 U11491 ( .B1(P1_B_REG_SCAN_IN), .B2(keyinput91), .C1(keyinput100), 
        .C2(P2_REG1_REG_21__SCAN_IN), .A(n10460), .ZN(n10463) );
  OAI22_X1 U11492 ( .A1(P1_D_REG_6__SCAN_IN), .A2(keyinput101), .B1(keyinput83), .B2(P2_D_REG_7__SCAN_IN), .ZN(n10461) );
  AOI221_X1 U11493 ( .B1(P1_D_REG_6__SCAN_IN), .B2(keyinput101), .C1(
        P2_D_REG_7__SCAN_IN), .C2(keyinput83), .A(n10461), .ZN(n10462) );
  NAND4_X1 U11494 ( .A1(n10465), .A2(n10464), .A3(n10463), .A4(n10462), .ZN(
        n10493) );
  OAI22_X1 U11495 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(keyinput38), .B1(
        P2_REG2_REG_2__SCAN_IN), .B2(keyinput54), .ZN(n10466) );
  AOI221_X1 U11496 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(keyinput38), .C1(
        keyinput54), .C2(P2_REG2_REG_2__SCAN_IN), .A(n10466), .ZN(n10473) );
  OAI22_X1 U11497 ( .A1(SI_15_), .A2(keyinput120), .B1(keyinput50), .B2(
        P2_REG3_REG_17__SCAN_IN), .ZN(n10467) );
  AOI221_X1 U11498 ( .B1(SI_15_), .B2(keyinput120), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput50), .A(n10467), .ZN(n10472) );
  OAI22_X1 U11499 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput114), .B1(
        keyinput72), .B2(P2_D_REG_13__SCAN_IN), .ZN(n10468) );
  AOI221_X1 U11500 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput114), .C1(
        P2_D_REG_13__SCAN_IN), .C2(keyinput72), .A(n10468), .ZN(n10471) );
  OAI22_X1 U11501 ( .A1(SI_18_), .A2(keyinput102), .B1(keyinput63), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n10469) );
  AOI221_X1 U11502 ( .B1(SI_18_), .B2(keyinput102), .C1(
        P2_REG2_REG_25__SCAN_IN), .C2(keyinput63), .A(n10469), .ZN(n10470) );
  NAND4_X1 U11503 ( .A1(n10473), .A2(n10472), .A3(n10471), .A4(n10470), .ZN(
        n10492) );
  OAI22_X1 U11504 ( .A1(P1_D_REG_14__SCAN_IN), .A2(keyinput5), .B1(keyinput99), 
        .B2(P2_REG1_REG_3__SCAN_IN), .ZN(n10474) );
  AOI221_X1 U11505 ( .B1(P1_D_REG_14__SCAN_IN), .B2(keyinput5), .C1(
        P2_REG1_REG_3__SCAN_IN), .C2(keyinput99), .A(n10474), .ZN(n10481) );
  OAI22_X1 U11506 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(keyinput126), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(keyinput31), .ZN(n10475) );
  AOI221_X1 U11507 ( .B1(P1_REG3_REG_13__SCAN_IN), .B2(keyinput126), .C1(
        keyinput31), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10475), .ZN(n10480) );
  OAI22_X1 U11508 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput113), .B1(
        keyinput123), .B2(SI_17_), .ZN(n10476) );
  AOI221_X1 U11509 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput113), .C1(SI_17_), 
        .C2(keyinput123), .A(n10476), .ZN(n10479) );
  OAI22_X1 U11510 ( .A1(P1_D_REG_12__SCAN_IN), .A2(keyinput95), .B1(
        keyinput105), .B2(P2_REG1_REG_2__SCAN_IN), .ZN(n10477) );
  AOI221_X1 U11511 ( .B1(P1_D_REG_12__SCAN_IN), .B2(keyinput95), .C1(
        P2_REG1_REG_2__SCAN_IN), .C2(keyinput105), .A(n10477), .ZN(n10478) );
  NAND4_X1 U11512 ( .A1(n10481), .A2(n10480), .A3(n10479), .A4(n10478), .ZN(
        n10491) );
  OAI22_X1 U11513 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput97), .B1(keyinput60), .B2(P2_REG2_REG_26__SCAN_IN), .ZN(n10482) );
  AOI221_X1 U11514 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput97), .C1(
        P2_REG2_REG_26__SCAN_IN), .C2(keyinput60), .A(n10482), .ZN(n10489) );
  OAI22_X1 U11515 ( .A1(P1_REG0_REG_11__SCAN_IN), .A2(keyinput17), .B1(
        P2_REG1_REG_24__SCAN_IN), .B2(keyinput66), .ZN(n10483) );
  AOI221_X1 U11516 ( .B1(P1_REG0_REG_11__SCAN_IN), .B2(keyinput17), .C1(
        keyinput66), .C2(P2_REG1_REG_24__SCAN_IN), .A(n10483), .ZN(n10488) );
  OAI22_X1 U11517 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(keyinput64), .B1(
        keyinput107), .B2(P2_IR_REG_22__SCAN_IN), .ZN(n10484) );
  AOI221_X1 U11518 ( .B1(P1_DATAO_REG_17__SCAN_IN), .B2(keyinput64), .C1(
        P2_IR_REG_22__SCAN_IN), .C2(keyinput107), .A(n10484), .ZN(n10487) );
  OAI22_X1 U11519 ( .A1(P1_REG0_REG_8__SCAN_IN), .A2(keyinput108), .B1(
        keyinput81), .B2(P2_REG3_REG_22__SCAN_IN), .ZN(n10485) );
  AOI221_X1 U11520 ( .B1(P1_REG0_REG_8__SCAN_IN), .B2(keyinput108), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput81), .A(n10485), .ZN(n10486) );
  NAND4_X1 U11521 ( .A1(n10489), .A2(n10488), .A3(n10487), .A4(n10486), .ZN(
        n10490) );
  NOR4_X1 U11522 ( .A1(n10493), .A2(n10492), .A3(n10491), .A4(n10490), .ZN(
        n10494) );
  NAND2_X1 U11523 ( .A1(n10495), .A2(n10494), .ZN(n10496) );
  NOR4_X1 U11524 ( .A1(n10499), .A2(n10498), .A3(n10497), .A4(n10496), .ZN(
        n10500) );
  XNOR2_X1 U11525 ( .A(n10501), .B(n10500), .ZN(P2_U3307) );
  XOR2_X1 U11526 ( .A(n10502), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  XOR2_X1 U11527 ( .A(n10504), .B(n10503), .Z(ADD_1071_U54) );
  NOR2_X1 U11528 ( .A1(n10506), .A2(n10505), .ZN(n10507) );
  XOR2_X1 U11529 ( .A(n10507), .B(P1_ADDR_REG_5__SCAN_IN), .Z(ADD_1071_U51) );
  OAI21_X1 U11530 ( .B1(n10510), .B2(n10509), .A(n10508), .ZN(n10512) );
  XOR2_X1 U11531 ( .A(n10512), .B(n10511), .Z(ADD_1071_U55) );
  AOI21_X1 U11532 ( .B1(n10515), .B2(n10514), .A(n10513), .ZN(ADD_1071_U47) );
  XOR2_X1 U11533 ( .A(n10516), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11534 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10517), .Z(ADD_1071_U48) );
  XOR2_X1 U11535 ( .A(n10519), .B(n10518), .Z(ADD_1071_U53) );
  XNOR2_X1 U11536 ( .A(n10521), .B(n10520), .ZN(ADD_1071_U52) );
endmodule

