

module b15_C_AntiSAT_k_128_9 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695;

  NAND2_X1 U34450 ( .A1(n4029), .A2(n4028), .ZN(n4986) );
  CLKBUF_X1 U34460 ( .A(n3589), .Z(n3074) );
  CLKBUF_X1 U34470 ( .A(n4108), .Z(n4223) );
  INV_X1 U34480 ( .A(n4120), .ZN(n4117) );
  INV_X1 U3449 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6368) );
  BUF_X2 U3450 ( .A(n3204), .Z(n4062) );
  CLKBUF_X2 U34510 ( .A(n3182), .Z(n3978) );
  CLKBUF_X2 U34520 ( .A(n3264), .Z(n4071) );
  CLKBUF_X2 U34530 ( .A(n3278), .Z(n4060) );
  CLKBUF_X2 U3454 ( .A(n3160), .Z(n4058) );
  BUF_X2 U34550 ( .A(n3894), .Z(n4070) );
  CLKBUF_X2 U34560 ( .A(n3263), .Z(n4068) );
  AND2_X1 U3457 ( .A1(n4102), .A2(n3073), .ZN(n4356) );
  AND4_X1 U3458 ( .A1(n3173), .A2(n3172), .A3(n3171), .A4(n3170), .ZN(n3306)
         );
  AND4_X1 U34590 ( .A1(n3212), .A2(n3211), .A3(n3210), .A4(n3209), .ZN(n4102)
         );
  AND2_X4 U34600 ( .A1(n4433), .A2(n4458), .ZN(n3182) );
  CLKBUF_X2 U34610 ( .A(n3262), .Z(n4036) );
  NOR2_X1 U34620 ( .A1(n3247), .A2(n3215), .ZN(n3568) );
  NAND2_X1 U34630 ( .A1(n4289), .A2(n3419), .ZN(n3247) );
  AND2_X1 U34640 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3021) );
  NOR2_X2 U34650 ( .A1(n3247), .A2(n3061), .ZN(n3060) );
  NOR2_X1 U3466 ( .A1(n3331), .A2(n6368), .ZN(n3559) );
  NAND2_X1 U3467 ( .A1(n3060), .A2(n3249), .ZN(n4358) );
  NAND2_X2 U34690 ( .A1(n3103), .A2(n4427), .ZN(n3189) );
  NAND2_X1 U34700 ( .A1(n3566), .A2(n3565), .ZN(n4418) );
  INV_X1 U34710 ( .A(n3847), .ZN(n4954) );
  INV_X1 U34720 ( .A(n3575), .ZN(n3847) );
  INV_X2 U34730 ( .A(n3249), .ZN(n5787) );
  INV_X1 U34740 ( .A(n5724), .ZN(n5754) );
  AND2_X1 U3475 ( .A1(n3002), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4434)
         );
  INV_X1 U3476 ( .A(n5763), .ZN(n5738) );
  OR2_X1 U3477 ( .A1(n4216), .A2(n4219), .ZN(n2997) );
  XNOR2_X2 U3478 ( .A(n3449), .B(n3448), .ZN(n3032) );
  NAND2_X2 U3479 ( .A1(n3447), .A2(n3446), .ZN(n3449) );
  NOR2_X2 U3480 ( .A1(n4399), .A2(n4448), .ZN(n4447) );
  NAND2_X2 U3481 ( .A1(n3359), .A2(n3358), .ZN(n4608) );
  AND2_X4 U3482 ( .A1(n4458), .A2(n4434), .ZN(n3979) );
  NOR2_X4 U3483 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4458) );
  CLKBUF_X1 U3485 ( .A(n4985), .Z(n5058) );
  OR2_X1 U3486 ( .A1(n5069), .A2(n5070), .ZN(n5072) );
  INV_X1 U3488 ( .A(n3215), .ZN(n4101) );
  NAND2_X1 U3489 ( .A1(n3139), .A2(n3138), .ZN(n3573) );
  INV_X1 U3490 ( .A(n3189), .ZN(n3087) );
  CLKBUF_X2 U3491 ( .A(n3175), .Z(n4009) );
  INV_X4 U3492 ( .A(n3189), .ZN(n3984) );
  CLKBUF_X2 U3493 ( .A(n3176), .Z(n3072) );
  AND2_X2 U3494 ( .A1(n4428), .A2(n3021), .ZN(n3195) );
  INV_X1 U3495 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3090) );
  NAND2_X1 U3496 ( .A1(n3009), .A2(n2999), .ZN(n3008) );
  NOR2_X2 U3497 ( .A1(n5524), .A2(n3512), .ZN(n3514) );
  CLKBUF_X1 U3498 ( .A(n5063), .Z(n5076) );
  NOR2_X1 U3499 ( .A1(n4263), .A2(n5078), .ZN(n5073) );
  CLKBUF_X1 U3500 ( .A(n4263), .Z(n5079) );
  OAI211_X1 U3501 ( .C1(n5253), .C2(n3048), .A(n3045), .B(n5245), .ZN(n3049)
         );
  OR2_X1 U3502 ( .A1(n4888), .A2(n3729), .ZN(n5115) );
  NAND2_X1 U3503 ( .A1(n4218), .A2(n3000), .ZN(n3026) );
  AND3_X1 U3504 ( .A1(n5254), .A2(n5381), .A3(n3499), .ZN(n3084) );
  INV_X1 U3505 ( .A(n5695), .ZN(n2999) );
  AND2_X1 U3506 ( .A1(n4323), .A2(n4324), .ZN(n4322) );
  OR2_X1 U3507 ( .A1(n4478), .A2(n3014), .ZN(n4399) );
  AND2_X1 U3508 ( .A1(n4105), .A2(n4731), .ZN(n4402) );
  AND2_X1 U3509 ( .A1(n3150), .A2(n3229), .ZN(n4289) );
  CLKBUF_X3 U3510 ( .A(n4117), .Z(n5017) );
  AND2_X1 U3511 ( .A1(n4970), .A2(n3306), .ZN(n3572) );
  CLKBUF_X1 U3512 ( .A(n3169), .Z(n4597) );
  AND2_X1 U3513 ( .A1(n3059), .A2(n3217), .ZN(n4098) );
  NAND4_X1 U3514 ( .A1(n3112), .A2(n3111), .A3(n3110), .A4(n3109), .ZN(n3059)
         );
  NAND2_X2 U3515 ( .A1(n3149), .A2(n3148), .ZN(n3574) );
  AND4_X1 U3516 ( .A1(n3102), .A2(n3101), .A3(n3100), .A4(n3099), .ZN(n3110)
         );
  CLKBUF_X2 U3517 ( .A(n3195), .Z(n4069) );
  AND2_X2 U3518 ( .A1(n4434), .A2(n3021), .ZN(n3176) );
  CLKBUF_X2 U3519 ( .A(n3290), .Z(n4061) );
  AND2_X2 U3520 ( .A1(n4458), .A2(n4427), .ZN(n3177) );
  INV_X2 U3521 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3321) );
  INV_X1 U3522 ( .A(n4253), .ZN(n5197) );
  INV_X1 U3523 ( .A(n5130), .ZN(n3009) );
  XNOR2_X1 U3524 ( .A(n3515), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5285)
         );
  MUX2_X1 U3525 ( .A(n4940), .B(n4939), .S(INSTADDRPOINTER_REG_29__SCAN_IN), 
        .Z(n3515) );
  OR2_X1 U3526 ( .A1(n5198), .A2(n5199), .ZN(n4253) );
  NOR2_X1 U3527 ( .A1(n3514), .A2(n4901), .ZN(n4940) );
  NAND2_X1 U3528 ( .A1(n5204), .A2(n4252), .ZN(n5198) );
  NAND2_X1 U3529 ( .A1(n4250), .A2(n4249), .ZN(n5204) );
  AND2_X1 U3530 ( .A1(n3055), .A2(n3511), .ZN(n5526) );
  NAND2_X1 U3531 ( .A1(n3052), .A2(n3050), .ZN(n5524) );
  NAND2_X1 U3532 ( .A1(n5533), .A2(n3053), .ZN(n3052) );
  CLKBUF_X1 U3533 ( .A(n4254), .Z(n4255) );
  CLKBUF_X1 U3534 ( .A(n5227), .Z(n5240) );
  OAI21_X1 U3535 ( .B1(n3044), .B2(n3046), .A(n3047), .ZN(n5246) );
  NAND2_X1 U3536 ( .A1(n3049), .A2(n3502), .ZN(n5227) );
  NAND2_X1 U3537 ( .A1(n4894), .A2(n4218), .ZN(n3027) );
  NAND2_X1 U3538 ( .A1(n3026), .A2(n4894), .ZN(n4900) );
  NAND2_X1 U3539 ( .A1(n3047), .A2(n3046), .ZN(n3045) );
  INV_X1 U3540 ( .A(n3047), .ZN(n3048) );
  AND2_X1 U3541 ( .A1(n3007), .A2(n3501), .ZN(n3047) );
  NAND2_X1 U3542 ( .A1(n5066), .A2(n3022), .ZN(n4216) );
  NAND2_X1 U3543 ( .A1(n3084), .A2(n5255), .ZN(n3007) );
  AND2_X1 U3544 ( .A1(n5066), .A2(n5059), .ZN(n5061) );
  NAND2_X1 U3545 ( .A1(n3054), .A2(n3051), .ZN(n3050) );
  INV_X1 U3546 ( .A(n3084), .ZN(n3046) );
  OR2_X1 U3547 ( .A1(n4346), .A2(n4347), .ZN(n4348) );
  AND2_X1 U3548 ( .A1(n3054), .A2(n3078), .ZN(n3053) );
  INV_X1 U3549 ( .A(n3511), .ZN(n3051) );
  INV_X1 U3550 ( .A(n5525), .ZN(n3054) );
  NAND2_X1 U3551 ( .A1(n4322), .A2(n5081), .ZN(n5069) );
  OR2_X1 U3552 ( .A1(n5228), .A2(n5387), .ZN(n5381) );
  NAND2_X1 U3553 ( .A1(n5228), .A2(n4912), .ZN(n3511) );
  NAND2_X1 U3554 ( .A1(n3075), .A2(n3401), .ZN(n3078) );
  INV_X1 U3555 ( .A(n3497), .ZN(n3075) );
  AND2_X1 U3556 ( .A1(n4163), .A2(n3025), .ZN(n4323) );
  NAND2_X1 U3557 ( .A1(n3006), .A2(n3398), .ZN(n3478) );
  NOR2_X1 U3558 ( .A1(n5091), .A2(n5092), .ZN(n4163) );
  INV_X1 U3559 ( .A(n3466), .ZN(n3006) );
  NAND2_X1 U3560 ( .A1(n3596), .A2(n3595), .ZN(n4387) );
  NOR2_X1 U3561 ( .A1(n5000), .A2(n4154), .ZN(n4159) );
  OAI21_X1 U3562 ( .B1(n5908), .B2(n5904), .A(n5905), .ZN(n4437) );
  NOR2_X1 U3563 ( .A1(n3005), .A2(n3373), .ZN(n3453) );
  CLKBUF_X1 U3564 ( .A(n4971), .Z(n5784) );
  CLKBUF_X1 U3565 ( .A(n3597), .Z(n5957) );
  CLKBUF_X1 U3566 ( .A(n5015), .Z(n5357) );
  NOR2_X1 U3567 ( .A1(n5119), .A2(n5033), .ZN(n5111) );
  NAND2_X1 U3568 ( .A1(n3360), .A2(n4608), .ZN(n3005) );
  NOR2_X1 U3569 ( .A1(n5119), .A2(n3011), .ZN(n5015) );
  OR3_X1 U3570 ( .A1(n5119), .A2(n3013), .A3(n5033), .ZN(n3010) );
  NAND2_X1 U3571 ( .A1(n4281), .A2(n6361), .ZN(n4328) );
  NOR2_X1 U3572 ( .A1(n5042), .A2(n5043), .ZN(n5121) );
  NAND2_X1 U3573 ( .A1(n4875), .A2(n4891), .ZN(n5042) );
  OAI21_X1 U3574 ( .B1(n4529), .B2(STATE2_REG_0__SCAN_IN), .A(n3342), .ZN(
        n3426) );
  CLKBUF_X1 U3575 ( .A(n4529), .Z(n5420) );
  CLKBUF_X1 U3576 ( .A(n4450), .Z(n6101) );
  AOI21_X1 U3577 ( .B1(n3581), .B2(n4298), .A(n6367), .ZN(n4376) );
  NOR2_X2 U3578 ( .A1(n4876), .A2(n4877), .ZN(n4875) );
  NAND2_X1 U3579 ( .A1(n4754), .A2(n4862), .ZN(n4876) );
  XNOR2_X1 U3580 ( .A(n5406), .B(n4679), .ZN(n4450) );
  NOR2_X1 U3581 ( .A1(n4755), .A2(n4756), .ZN(n4754) );
  AOI21_X1 U3582 ( .B1(n3407), .B2(n3406), .A(n3405), .ZN(n4536) );
  NAND2_X1 U3583 ( .A1(n3030), .A2(n3028), .ZN(n4755) );
  AOI21_X1 U3584 ( .B1(n3402), .B2(n3310), .A(n3404), .ZN(n3068) );
  AOI21_X1 U3585 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6368), .A(n3561), 
        .ZN(n3562) );
  INV_X1 U3586 ( .A(n4565), .ZN(n3030) );
  NAND2_X1 U3587 ( .A1(n3347), .A2(n3346), .ZN(n4679) );
  NAND2_X1 U3588 ( .A1(n3036), .A2(n3035), .ZN(n3034) );
  NAND2_X1 U3589 ( .A1(n3039), .A2(n3040), .ZN(n3277) );
  AND2_X1 U3590 ( .A1(n3020), .A2(n3017), .ZN(n3016) );
  OR2_X1 U3591 ( .A1(n3244), .A2(n3321), .ZN(n3325) );
  AND2_X1 U3592 ( .A1(n3041), .A2(n3260), .ZN(n3035) );
  NAND2_X1 U3593 ( .A1(n3237), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3244) );
  AND2_X1 U3594 ( .A1(n5016), .A2(n4157), .ZN(n4158) );
  NAND2_X1 U3595 ( .A1(n3237), .A2(n3042), .ZN(n3041) );
  OAI211_X1 U3596 ( .C1(n4358), .C2(n3225), .A(n4283), .B(n4285), .ZN(n3004)
         );
  NAND2_X1 U3597 ( .A1(n5110), .A2(n3012), .ZN(n3011) );
  NOR2_X1 U3598 ( .A1(n4333), .A2(n4116), .ZN(n4561) );
  INV_X1 U3599 ( .A(n3060), .ZN(n4273) );
  NAND2_X1 U3600 ( .A1(n3015), .A2(n4400), .ZN(n3014) );
  CLKBUF_X1 U3601 ( .A(n4198), .Z(n4361) );
  NOR2_X1 U3602 ( .A1(n3024), .A2(n3023), .ZN(n3022) );
  NOR2_X1 U3603 ( .A1(n4566), .A2(n3029), .ZN(n3028) );
  INV_X1 U3604 ( .A(n4479), .ZN(n3015) );
  INV_X1 U3605 ( .A(n5110), .ZN(n3013) );
  OAI21_X1 U3606 ( .B1(n3031), .B2(n4303), .A(n5787), .ZN(n3259) );
  INV_X1 U3607 ( .A(n4895), .ZN(n3000) );
  INV_X1 U3608 ( .A(n4343), .ZN(n3029) );
  XNOR2_X1 U3609 ( .A(n4115), .B(n4486), .ZN(n4332) );
  NOR2_X1 U3610 ( .A1(n5033), .A2(n5358), .ZN(n3012) );
  NOR2_X1 U3611 ( .A1(n3224), .A2(n3031), .ZN(n4198) );
  AND2_X1 U3612 ( .A1(n3304), .A2(n3303), .ZN(n3403) );
  AOI22_X1 U3613 ( .A1(EBX_REG_0__SCAN_IN), .A2(n4123), .B1(n4117), .B2(n5760), 
        .ZN(n4486) );
  NOR2_X1 U3614 ( .A1(EBX_REG_2__SCAN_IN), .A2(n4897), .ZN(n4119) );
  AND2_X1 U3615 ( .A1(n3220), .A2(n3574), .ZN(n3229) );
  INV_X1 U3616 ( .A(n3169), .ZN(n4970) );
  AND2_X1 U3617 ( .A1(n5787), .A2(n4102), .ZN(n4731) );
  OR2_X1 U3618 ( .A1(n3288), .A2(n3287), .ZN(n3489) );
  INV_X1 U3619 ( .A(n3059), .ZN(n3169) );
  AND2_X1 U3620 ( .A1(n4303), .A2(n3249), .ZN(n4108) );
  INV_X1 U3621 ( .A(n4102), .ZN(n4303) );
  INV_X1 U3622 ( .A(n3419), .ZN(n4602) );
  OR2_X1 U3623 ( .A1(n3300), .A2(n3299), .ZN(n3418) );
  AND4_X1 U3624 ( .A1(n3125), .A2(n3124), .A3(n3123), .A4(n3122), .ZN(n3173)
         );
  AND2_X1 U3625 ( .A1(n3138), .A2(n3139), .ZN(n3217) );
  NAND2_X1 U3626 ( .A1(n3083), .A2(n3159), .ZN(n3419) );
  AND4_X1 U3627 ( .A1(n3116), .A2(n3115), .A3(n3114), .A4(n3113), .ZN(n3138)
         );
  AND4_X1 U3628 ( .A1(n3158), .A2(n3157), .A3(n3156), .A4(n3155), .ZN(n3159)
         );
  AND4_X1 U3629 ( .A1(n3194), .A2(n3193), .A3(n3192), .A4(n3191), .ZN(n3212)
         );
  AND4_X1 U3630 ( .A1(n3208), .A2(n3207), .A3(n3206), .A4(n3205), .ZN(n3209)
         );
  AND4_X1 U3631 ( .A1(n3199), .A2(n3198), .A3(n3197), .A4(n3196), .ZN(n3211)
         );
  AND4_X1 U3632 ( .A1(n3147), .A2(n3146), .A3(n3145), .A4(n3144), .ZN(n3148)
         );
  AND4_X1 U3633 ( .A1(n3129), .A2(n3128), .A3(n3127), .A4(n3126), .ZN(n3172)
         );
  AND4_X1 U3634 ( .A1(n3133), .A2(n3132), .A3(n3131), .A4(n3130), .ZN(n3171)
         );
  AND4_X1 U3635 ( .A1(n3098), .A2(n3097), .A3(n3096), .A4(n3095), .ZN(n3111)
         );
  AND4_X1 U3636 ( .A1(n3137), .A2(n3136), .A3(n3135), .A4(n3134), .ZN(n3170)
         );
  NOR2_X1 U3637 ( .A1(n6275), .A2(n4637), .ZN(n6283) );
  OR2_X1 U3638 ( .A1(n3189), .A2(n3190), .ZN(n3192) );
  AND4_X1 U3639 ( .A1(n3120), .A2(n3119), .A3(n3118), .A4(n3117), .ZN(n3139)
         );
  BUF_X2 U3640 ( .A(n4009), .Z(n4072) );
  AND4_X1 U3641 ( .A1(n3203), .A2(n3202), .A3(n3201), .A4(n3200), .ZN(n3210)
         );
  AND4_X1 U3642 ( .A1(n3143), .A2(n3142), .A3(n3141), .A4(n3140), .ZN(n3149)
         );
  BUF_X2 U3643 ( .A(n3700), .Z(n4057) );
  BUF_X2 U3644 ( .A(n3979), .Z(n3852) );
  BUF_X2 U3645 ( .A(n3177), .Z(n4059) );
  NOR2_X1 U3646 ( .A1(n3090), .A2(n3043), .ZN(n3042) );
  INV_X2 U3647 ( .A(n6491), .ZN(n6480) );
  AND2_X2 U3648 ( .A1(n4452), .A2(n4428), .ZN(n3700) );
  AND2_X2 U3649 ( .A1(n4428), .A2(n3103), .ZN(n3278) );
  AND2_X2 U3650 ( .A1(n4452), .A2(n4434), .ZN(n3894) );
  AND2_X1 U3651 ( .A1(n3001), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3103)
         );
  AND3_X2 U3652 ( .A1(n3090), .A2(n3104), .A3(n4451), .ZN(n3264) );
  AND2_X1 U3653 ( .A1(n3003), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4433)
         );
  AND2_X2 U3654 ( .A1(n3321), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4452)
         );
  AND2_X2 U3655 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4427) );
  AND2_X1 U3656 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4451) );
  INV_X1 U3657 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3001) );
  INV_X1 U3658 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3003) );
  INV_X1 U3659 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3002) );
  AND2_X2 U3660 ( .A1(n3003), .A2(n3002), .ZN(n4428) );
  INV_X1 U3661 ( .A(n3240), .ZN(n3228) );
  NAND2_X1 U3662 ( .A1(n3004), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3240) );
  NAND2_X1 U3663 ( .A1(n4402), .A2(n3216), .ZN(n4283) );
  NAND2_X1 U3664 ( .A1(n5533), .A2(n3078), .ZN(n3055) );
  AND2_X2 U3665 ( .A1(n3510), .A2(n3509), .ZN(n5533) );
  XNOR2_X1 U3666 ( .A(n3005), .B(n3444), .ZN(n3613) );
  NAND2_X2 U3667 ( .A1(n3478), .A2(n3400), .ZN(n3497) );
  NAND2_X1 U3668 ( .A1(n4984), .A2(n3008), .ZN(U2796) );
  NAND2_X1 U3669 ( .A1(n5015), .A2(n5100), .ZN(n5000) );
  OR2_X1 U3670 ( .A1(n4478), .A2(n4479), .ZN(n3020) );
  NAND2_X1 U3671 ( .A1(n4478), .A2(n4479), .ZN(n3017) );
  NAND2_X1 U3672 ( .A1(n4399), .A2(n3018), .ZN(n5729) );
  NAND2_X1 U3673 ( .A1(n3020), .A2(n3019), .ZN(n3018) );
  INV_X1 U3674 ( .A(n4400), .ZN(n3019) );
  INV_X1 U3675 ( .A(n3021), .ZN(n4461) );
  AND2_X2 U3676 ( .A1(n3021), .A2(n4427), .ZN(n3290) );
  AND2_X2 U3677 ( .A1(n4433), .A2(n3021), .ZN(n3204) );
  NAND2_X1 U3678 ( .A1(n5401), .A2(n3021), .ZN(n5402) );
  INV_X1 U3679 ( .A(n4991), .ZN(n3023) );
  INV_X1 U3680 ( .A(n5059), .ZN(n3024) );
  NOR2_X2 U3681 ( .A1(n5072), .A2(n5065), .ZN(n5066) );
  INV_X1 U3682 ( .A(n4163), .ZN(n5083) );
  INV_X1 U3683 ( .A(n5082), .ZN(n3025) );
  NAND2_X1 U3684 ( .A1(n3027), .A2(n4222), .ZN(n4946) );
  NOR2_X1 U3685 ( .A1(n4565), .A2(n4566), .ZN(n4564) );
  NAND3_X1 U3686 ( .A1(n3223), .A2(n3250), .A3(n3222), .ZN(n3031) );
  NAND2_X1 U3687 ( .A1(n3032), .A2(n4517), .ZN(n3451) );
  XNOR2_X1 U3688 ( .A(n4517), .B(n3032), .ZN(n4559) );
  NAND2_X1 U3689 ( .A1(n3034), .A2(n3277), .ZN(n3582) );
  NAND3_X1 U3690 ( .A1(n3034), .A2(n3277), .A3(n3033), .ZN(n3402) );
  INV_X1 U3691 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n3033) );
  NOR2_X1 U3692 ( .A1(n3038), .A2(n3037), .ZN(n3036) );
  INV_X1 U3693 ( .A(n3243), .ZN(n3037) );
  INV_X1 U3694 ( .A(n4295), .ZN(n3038) );
  NAND2_X1 U3695 ( .A1(n3260), .A2(n4295), .ZN(n3039) );
  NAND2_X1 U3696 ( .A1(n3041), .A2(n3243), .ZN(n3040) );
  INV_X1 U3697 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n3043) );
  INV_X1 U3698 ( .A(n5253), .ZN(n3044) );
  INV_X1 U3699 ( .A(n3055), .ZN(n5161) );
  OAI21_X1 U3700 ( .B1(n5285), .B2(n3056), .A(n4095), .ZN(U2956) );
  INV_X1 U3701 ( .A(n5916), .ZN(n3056) );
  INV_X1 U3702 ( .A(n3090), .ZN(n3057) );
  OAI21_X2 U3703 ( .B1(n3616), .B2(n3461), .A(n3460), .ZN(n3462) );
  CLKBUF_X1 U3704 ( .A(n4467), .Z(n3058) );
  NAND2_X1 U3705 ( .A1(n3451), .A2(n3450), .ZN(n4467) );
  NAND2_X1 U3706 ( .A1(n3473), .A2(n3472), .ZN(n4640) );
  NAND2_X1 U3707 ( .A1(n3326), .A2(n3327), .ZN(n5406) );
  INV_X1 U3708 ( .A(n3189), .ZN(n4067) );
  NAND2_X1 U3709 ( .A1(n4101), .A2(n3174), .ZN(n3061) );
  NAND2_X1 U3710 ( .A1(n4588), .A2(n4563), .ZN(n3062) );
  NOR2_X2 U3711 ( .A1(n3062), .A2(n3063), .ZN(n4860) );
  OR2_X1 U3712 ( .A1(n4799), .A2(n4347), .ZN(n3063) );
  XNOR2_X1 U3713 ( .A(n4888), .B(n3728), .ZN(n3064) );
  NOR2_X2 U3714 ( .A1(n4263), .A2(n3065), .ZN(n5063) );
  OR2_X1 U3715 ( .A1(n5078), .A2(n3066), .ZN(n3065) );
  INV_X1 U3716 ( .A(n5074), .ZN(n3066) );
  NOR2_X1 U3717 ( .A1(n4589), .A2(n4590), .ZN(n3067) );
  XNOR2_X1 U3718 ( .A(n4952), .B(n4951), .ZN(n3069) );
  XNOR2_X1 U3719 ( .A(n4888), .B(n3728), .ZN(n5038) );
  NOR2_X1 U3720 ( .A1(n4589), .A2(n4590), .ZN(n4588) );
  OR2_X1 U3721 ( .A1(n4395), .A2(n4445), .ZN(n4589) );
  AOI21_X1 U3722 ( .B1(n3402), .B2(n3310), .A(n3404), .ZN(n3414) );
  XNOR2_X1 U3723 ( .A(n4952), .B(n4951), .ZN(n4096) );
  CLKBUF_X1 U3724 ( .A(n4774), .Z(n3070) );
  CLKBUF_X1 U3725 ( .A(n4748), .Z(n3071) );
  OAI21_X2 U3726 ( .B1(n4437), .B2(n4438), .A(n3443), .ZN(n4517) );
  NAND2_X1 U3727 ( .A1(n3233), .A2(n3419), .ZN(n3250) );
  NAND2_X1 U3728 ( .A1(n5121), .A2(n5120), .ZN(n5119) );
  XNOR2_X1 U3729 ( .A(n3442), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4438)
         );
  NAND2_X1 U3730 ( .A1(n3441), .A2(n3440), .ZN(n3442) );
  OR2_X1 U3731 ( .A1(n3188), .A2(n3187), .ZN(n3073) );
  XNOR2_X1 U3732 ( .A(n3427), .B(n3426), .ZN(n3589) );
  AOI21_X1 U3733 ( .B1(n4196), .B2(n4986), .A(n4952), .ZN(n5157) );
  NOR2_X4 U3734 ( .A1(n4986), .A2(n4196), .ZN(n4952) );
  AND2_X1 U3735 ( .A1(n4100), .A2(n4294), .ZN(n4282) );
  INV_X1 U3736 ( .A(n3465), .ZN(n3398) );
  INV_X1 U3737 ( .A(n4025), .ZN(n4052) );
  AND2_X1 U3738 ( .A1(n3214), .A2(n4602), .ZN(n4105) );
  INV_X1 U3739 ( .A(n4328), .ZN(n4304) );
  NAND2_X1 U3740 ( .A1(n3169), .A2(n3573), .ZN(n3220) );
  NOR2_X1 U3742 ( .A1(n3305), .A2(n6368), .ZN(n3302) );
  INV_X1 U3743 ( .A(n5056), .ZN(n4005) );
  AND2_X1 U3744 ( .A1(n3849), .A2(n5012), .ZN(n4998) );
  OR2_X1 U3745 ( .A1(n4429), .A2(n6368), .ZN(n4046) );
  INV_X1 U3746 ( .A(n4397), .ZN(n3614) );
  NOR2_X1 U3747 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4025) );
  OR2_X1 U3748 ( .A1(n4597), .A2(n4550), .ZN(n3461) );
  AND2_X1 U3749 ( .A1(n5755), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4974) );
  AND3_X1 U3750 ( .A1(n3651), .A2(n3650), .A3(n3649), .ZN(n4347) );
  INV_X1 U3751 ( .A(n3997), .ZN(n3998) );
  NAND2_X1 U3752 ( .A1(n4394), .A2(n3592), .ZN(n4389) );
  AND2_X1 U3753 ( .A1(n4418), .A2(n6361), .ZN(n5840) );
  INV_X1 U3754 ( .A(n5598), .ZN(n5408) );
  OR2_X1 U3755 ( .A1(n4273), .A2(n6485), .ZN(n5839) );
  MUX2_X1 U3756 ( .A(n4279), .B(n4278), .S(n3215), .Z(n4280) );
  AND2_X1 U3757 ( .A1(n4422), .A2(n4421), .ZN(n6341) );
  NAND2_X1 U3758 ( .A1(n6368), .A2(n4523), .ZN(n5416) );
  INV_X2 U3759 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6367) );
  AND2_X1 U3760 ( .A1(n5755), .A2(n4235), .ZN(n5763) );
  NAND2_X1 U3761 ( .A1(n4107), .A2(n6361), .ZN(n5103) );
  INV_X2 U3762 ( .A(n5103), .ZN(n5776) );
  INV_X1 U3763 ( .A(n5909), .ZN(n5213) );
  INV_X1 U3764 ( .A(n5553), .ZN(n5919) );
  AND2_X1 U3765 ( .A1(n5840), .A2(n4357), .ZN(n5916) );
  XNOR2_X1 U3766 ( .A(n4260), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4288)
         );
  INV_X1 U3767 ( .A(n5944), .ZN(n6688) );
  OR2_X1 U3768 ( .A1(n4731), .A2(n3528), .ZN(n3554) );
  AND2_X1 U3769 ( .A1(n4200), .A2(n3541), .ZN(n3555) );
  NAND2_X1 U3770 ( .A1(n3229), .A2(n3306), .ZN(n4097) );
  OR2_X1 U3771 ( .A1(n3554), .A2(n3555), .ZN(n3535) );
  OR2_X1 U3772 ( .A1(n3395), .A2(n3394), .ZN(n3480) );
  OR2_X1 U3773 ( .A1(n3370), .A2(n3369), .ZN(n3455) );
  AND2_X1 U3774 ( .A1(n3256), .A2(n3255), .ZN(n3260) );
  NAND2_X1 U3775 ( .A1(n3249), .A2(n3305), .ZN(n3331) );
  INV_X1 U3776 ( .A(n3580), .ZN(n3218) );
  NOR2_X1 U3777 ( .A1(n3094), .A2(n3093), .ZN(n3112) );
  AOI22_X1 U3778 ( .A1(n3894), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3979), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3120) );
  AOI22_X1 U3779 ( .A1(n3087), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3700), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3116) );
  OR2_X1 U3780 ( .A1(n3357), .A2(n3356), .ZN(n3439) );
  OR3_X1 U3781 ( .A1(n3526), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(n3525), 
        .ZN(n4204) );
  AOI22_X1 U3782 ( .A1(n3894), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3186) );
  INV_X1 U3783 ( .A(n3541), .ZN(n3563) );
  NAND2_X1 U3784 ( .A1(n3524), .A2(n3523), .ZN(n4203) );
  OR2_X1 U3785 ( .A1(n3453), .A2(n3452), .ZN(n3454) );
  CLKBUF_X1 U3786 ( .A(n4996), .Z(n4997) );
  NAND2_X1 U3787 ( .A1(n3713), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3744)
         );
  AND2_X1 U3788 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n3617), .ZN(n3625)
         );
  AND2_X1 U3789 ( .A1(n4169), .A2(n4168), .ZN(n4324) );
  AND2_X1 U3790 ( .A1(n4155), .A2(n5004), .ZN(n4154) );
  AND2_X1 U3791 ( .A1(n5228), .A2(n5387), .ZN(n5255) );
  NOR2_X1 U3792 ( .A1(n3571), .A2(n3570), .ZN(n4100) );
  OR2_X1 U3793 ( .A1(n3341), .A2(n3340), .ZN(n3428) );
  AND2_X1 U3794 ( .A1(n3331), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3541) );
  OR2_X1 U3795 ( .A1(n3244), .A2(n3104), .ZN(n3347) );
  OAI21_X1 U3796 ( .B1(n6486), .B2(n6462), .A(n4931), .ZN(n4523) );
  INV_X1 U3797 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6344) );
  INV_X1 U3798 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6337) );
  AND2_X1 U3799 ( .A1(n4282), .A2(n4731), .ZN(n4381) );
  AND2_X1 U3800 ( .A1(n3798), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3794)
         );
  NAND2_X1 U3801 ( .A1(n4114), .A2(n4113), .ZN(n4115) );
  NAND2_X1 U3802 ( .A1(n4217), .A2(n4291), .ZN(n4218) );
  AND2_X1 U3803 ( .A1(n4166), .A2(n4165), .ZN(n5082) );
  AND2_X1 U3804 ( .A1(n3850), .A2(n4998), .ZN(n3851) );
  INV_X1 U3805 ( .A(n4896), .ZN(n4487) );
  NAND2_X1 U3806 ( .A1(n5840), .A2(n4197), .ZN(n5842) );
  AND2_X1 U3807 ( .A1(n6367), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4953) );
  OR2_X1 U3808 ( .A1(n5155), .A2(n4052), .ZN(n4053) );
  INV_X1 U3809 ( .A(n4985), .ZN(n4029) );
  OR2_X1 U3810 ( .A1(n5442), .A2(n4052), .ZN(n4003) );
  AND2_X1 U3811 ( .A1(n5447), .A2(n4207), .ZN(n3975) );
  NOR2_X1 U3812 ( .A1(n3955), .A2(n3954), .ZN(n3956) );
  AND2_X1 U3813 ( .A1(n3959), .A2(n3958), .ZN(n5074) );
  OR2_X1 U3814 ( .A1(n5531), .A2(n4052), .ZN(n3958) );
  CLKBUF_X1 U3815 ( .A(n4261), .Z(n4262) );
  AND2_X1 U3816 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n3867), .ZN(n3868)
         );
  INV_X1 U3817 ( .A(n3866), .ZN(n3867) );
  NOR2_X1 U3818 ( .A1(n3793), .A2(n3745), .ZN(n3748) );
  NAND2_X1 U3819 ( .A1(n3748), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3866)
         );
  NOR2_X1 U3820 ( .A1(n3814), .A2(n5029), .ZN(n3798) );
  NOR2_X1 U3821 ( .A1(n3744), .A2(n5247), .ZN(n3843) );
  NOR2_X1 U3822 ( .A1(n3696), .A2(n3692), .ZN(n3713) );
  NAND2_X1 U3823 ( .A1(n3691), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3696)
         );
  NOR2_X1 U3824 ( .A1(n3667), .A2(n5682), .ZN(n3691) );
  NAND2_X1 U3825 ( .A1(n3635), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3652)
         );
  AND2_X1 U3826 ( .A1(n3625), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3635)
         );
  AOI21_X1 U3827 ( .B1(n3633), .B2(n3842), .A(n3632), .ZN(n4590) );
  INV_X1 U3828 ( .A(n3598), .ZN(n3599) );
  NAND2_X1 U3829 ( .A1(n3599), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3608)
         );
  INV_X1 U3830 ( .A(n4394), .ZN(n3593) );
  INV_X1 U3831 ( .A(n5563), .ZN(n4911) );
  INV_X1 U3832 ( .A(n5207), .ZN(n4249) );
  INV_X1 U3833 ( .A(n5343), .ZN(n5572) );
  NOR2_X1 U3834 ( .A1(n5948), .A2(n5365), .ZN(n5341) );
  OR2_X1 U3835 ( .A1(n4273), .A2(n4897), .ZN(n4413) );
  AND2_X1 U3836 ( .A1(n4100), .A2(n3572), .ZN(n4357) );
  AND2_X1 U3837 ( .A1(n5371), .A2(n5366), .ZN(n5948) );
  NAND2_X1 U3838 ( .A1(n3402), .A2(n3403), .ZN(n3407) );
  CLKBUF_X1 U3839 ( .A(n4425), .Z(n4426) );
  NAND2_X1 U3840 ( .A1(n3569), .A2(n4970), .ZN(n4429) );
  INV_X1 U3841 ( .A(n3248), .ZN(n3569) );
  NOR2_X1 U3842 ( .A1(n5957), .A2(n5956), .ZN(n5987) );
  AND2_X1 U3843 ( .A1(n4651), .A2(n5957), .ZN(n6103) );
  AND2_X1 U3844 ( .A1(n6276), .A2(n4609), .ZN(n6185) );
  OR2_X1 U3845 ( .A1(n5413), .A2(n5412), .ZN(n6356) );
  NAND2_X1 U3846 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4418), .ZN(n4931) );
  INV_X1 U3847 ( .A(n6374), .ZN(n6361) );
  INV_X1 U3848 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U3849 ( .A1(n5842), .A2(n5432), .ZN(n6481) );
  INV_X1 U3850 ( .A(n5764), .ZN(n5683) );
  AND2_X1 U3851 ( .A1(n4974), .A2(n4231), .ZN(n5724) );
  AND2_X1 U3852 ( .A1(n4732), .A2(n5695), .ZN(n5767) );
  AND2_X1 U3853 ( .A1(n5755), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5764) );
  AND2_X1 U3854 ( .A1(n4974), .A2(n4224), .ZN(n5758) );
  INV_X1 U3855 ( .A(n5630), .ZN(n5777) );
  INV_X1 U3856 ( .A(n5507), .ZN(n5781) );
  AND2_X1 U3857 ( .A1(n5151), .A2(n3216), .ZN(n5780) );
  INV_X1 U3858 ( .A(n5148), .ZN(n5152) );
  AND2_X1 U3859 ( .A1(n5840), .A2(n5430), .ZN(n5814) );
  AND2_X1 U3860 ( .A1(n5840), .A2(n4377), .ZN(n5893) );
  NOR2_X1 U3861 ( .A1(n4413), .A2(READY_N), .ZN(n4377) );
  INV_X1 U3862 ( .A(n5887), .ZN(n5895) );
  OR2_X1 U3863 ( .A1(n4212), .A2(n4211), .ZN(n4214) );
  AND2_X1 U3864 ( .A1(n4050), .A2(n4024), .ZN(n5164) );
  INV_X1 U3865 ( .A(n5200), .ZN(n5514) );
  OR2_X1 U3866 ( .A1(n5916), .A2(n4087), .ZN(n5553) );
  NAND2_X1 U3867 ( .A1(n5553), .A2(n5918), .ZN(n5914) );
  INV_X1 U3868 ( .A(n6275), .ZN(n5909) );
  AOI21_X1 U3869 ( .B1(n4941), .B2(n5572), .A(n4943), .ZN(n5282) );
  AOI21_X1 U3870 ( .B1(n5572), .B2(n5306), .A(n5558), .ZN(n5300) );
  AOI211_X1 U3871 ( .C1(n4313), .C2(n4308), .A(n4306), .B(n4307), .ZN(n5939)
         );
  NOR2_X2 U3872 ( .A1(n4328), .A2(n4327), .ZN(n5944) );
  AND2_X1 U3873 ( .A1(n5839), .A2(n4326), .ZN(n4327) );
  NAND2_X1 U3874 ( .A1(n4304), .A2(n4362), .ZN(n5940) );
  AND2_X1 U3875 ( .A1(n5375), .A2(n5371), .ZN(n5343) );
  NAND2_X1 U3876 ( .A1(n4304), .A2(n5429), .ZN(n5371) );
  CLKBUF_X1 U3877 ( .A(n4536), .Z(n6465) );
  CLKBUF_X1 U3878 ( .A(n4525), .Z(n4526) );
  INV_X1 U3879 ( .A(n4426), .ZN(n5396) );
  NOR2_X2 U3880 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6464) );
  AND2_X1 U3881 ( .A1(n4361), .A2(n4303), .ZN(n5429) );
  NOR2_X1 U3882 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n5597) );
  INV_X1 U3883 ( .A(n6049), .ZN(n6023) );
  NOR2_X1 U3884 ( .A1(n4537), .A2(n3581), .ZN(n4801) );
  OR3_X1 U3885 ( .A1(n4656), .A2(n4655), .A3(n4654), .ZN(n6098) );
  AND2_X1 U3886 ( .A1(n4571), .A2(n5957), .ZN(n6156) );
  AND2_X1 U3887 ( .A1(n4616), .A2(n5957), .ZN(n6181) );
  INV_X1 U3888 ( .A(n6211), .ZN(n6212) );
  OAI21_X1 U3889 ( .B1(n6262), .B2(n6458), .A(n6232), .ZN(n6265) );
  INV_X1 U3890 ( .A(n5979), .ZN(n6327) );
  INV_X1 U3891 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U3892 ( .A1(n3567), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6374) );
  AOI21_X1 U3893 ( .B1(n3086), .B2(n4194), .A(n4193), .ZN(n4195) );
  NOR2_X1 U3894 ( .A1(n5776), .A2(n6647), .ZN(n4193) );
  INV_X1 U3895 ( .A(n4268), .ZN(n4269) );
  OAI21_X1 U3896 ( .B1(n5472), .B2(n5213), .A(n4267), .ZN(n4268) );
  OAI211_X1 U3897 ( .C1(n4941), .C2(n4948), .A(n4947), .B(n3082), .ZN(n4949)
         );
  OR2_X1 U3898 ( .A1(n3239), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3076)
         );
  NAND2_X1 U3899 ( .A1(n3217), .A2(n3574), .ZN(n3580) );
  AND2_X1 U3900 ( .A1(n3919), .A2(n3918), .ZN(n3077) );
  OR2_X1 U3901 ( .A1(n3074), .A2(n6218), .ZN(n4617) );
  AND2_X1 U3902 ( .A1(n3074), .A2(n4608), .ZN(n6276) );
  INV_X1 U3903 ( .A(n3277), .ZN(n3317) );
  OR2_X1 U3904 ( .A1(n6383), .A2(n6271), .ZN(n6275) );
  INV_X1 U3905 ( .A(n4536), .ZN(n3581) );
  NOR2_X1 U3906 ( .A1(n5170), .A2(n4914), .ZN(n4939) );
  AND4_X1 U3907 ( .A1(n3164), .A2(n3163), .A3(n3162), .A4(n3161), .ZN(n3079)
         );
  OR2_X1 U3908 ( .A1(n4946), .A2(n5671), .ZN(n3080) );
  OR2_X1 U3909 ( .A1(n5473), .A2(n6688), .ZN(n3081) );
  OR2_X1 U3910 ( .A1(n4946), .A2(n6688), .ZN(n3082) );
  AND4_X1 U3911 ( .A1(n3154), .A2(n3153), .A3(n3152), .A4(n3151), .ZN(n3083)
         );
  AND4_X1 U3912 ( .A1(n3168), .A2(n3167), .A3(n3166), .A4(n3165), .ZN(n3085)
         );
  INV_X1 U3913 ( .A(n5122), .ZN(n4194) );
  INV_X1 U3914 ( .A(n5126), .ZN(n5772) );
  NAND4_X1 U3915 ( .A1(n3173), .A2(n3172), .A3(n3171), .A4(n3170), .ZN(n3305)
         );
  AND2_X1 U3916 ( .A1(n4192), .A2(n4191), .ZN(n3086) );
  NAND2_X2 U3917 ( .A1(n5151), .A2(n4385), .ZN(n5507) );
  OR2_X1 U3918 ( .A1(n3552), .A2(n3551), .ZN(n3553) );
  AND2_X1 U3919 ( .A1(n6468), .A2(n3057), .ZN(n3538) );
  NAND2_X1 U3920 ( .A1(n3518), .A2(n3517), .ZN(n3532) );
  NOR2_X1 U3921 ( .A1(n4970), .A2(n3305), .ZN(n3174) );
  INV_X1 U3922 ( .A(n3239), .ZN(n3241) );
  AND2_X1 U3923 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n3525), .ZN(n3521)
         );
  INV_X1 U3924 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4109) );
  OR2_X1 U3925 ( .A1(n3274), .A2(n3273), .ZN(n3417) );
  NAND2_X1 U3926 ( .A1(n3092), .A2(n3091), .ZN(n3093) );
  INV_X1 U3927 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3525) );
  OR2_X1 U3928 ( .A1(n3526), .A2(n3521), .ZN(n3524) );
  NAND2_X1 U3929 ( .A1(n3594), .A2(n3593), .ZN(n3595) );
  OR2_X1 U3930 ( .A1(n5476), .A2(n4052), .ZN(n3918) );
  NAND2_X1 U3931 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3503) );
  OR2_X1 U3932 ( .A1(n3311), .A2(n3301), .ZN(n3304) );
  OR2_X1 U3933 ( .A1(n3189), .A2(n3121), .ZN(n3123) );
  AND4_X1 U3934 ( .A1(n3108), .A2(n3107), .A3(n3106), .A4(n3105), .ZN(n3109)
         );
  NAND2_X1 U3935 ( .A1(n3559), .A2(n3527), .ZN(n3564) );
  NOR2_X1 U3936 ( .A1(n4023), .A2(n6650), .ZN(n4048) );
  AND2_X1 U3937 ( .A1(n3397), .A2(n3396), .ZN(n3465) );
  OR2_X1 U3938 ( .A1(n3383), .A2(n3382), .ZN(n3458) );
  INV_X1 U3939 ( .A(n3461), .ZN(n3527) );
  NAND2_X1 U3940 ( .A1(n3325), .A2(n3324), .ZN(n3327) );
  XNOR2_X1 U3941 ( .A(n3437), .B(n4608), .ZN(n3597) );
  OR2_X1 U3942 ( .A1(n3564), .A2(n4203), .ZN(n3565) );
  INV_X1 U3943 ( .A(n4123), .ZN(n4182) );
  NAND2_X1 U3944 ( .A1(n3249), .A2(n4602), .ZN(n4123) );
  INV_X1 U3945 ( .A(n4988), .ZN(n4028) );
  OR2_X1 U3946 ( .A1(n3652), .A2(n4342), .ZN(n3667) );
  NOR2_X1 U3947 ( .A1(n3608), .A2(n4555), .ZN(n3617) );
  AND2_X1 U3948 ( .A1(n5228), .A2(n5559), .ZN(n3512) );
  NAND2_X1 U3949 ( .A1(n3410), .A2(n3409), .ZN(n4481) );
  AND2_X1 U3950 ( .A1(n3404), .A2(n3403), .ZN(n3405) );
  INV_X1 U3951 ( .A(n5416), .ZN(n4803) );
  AND2_X1 U3952 ( .A1(n5399), .A2(n5398), .ZN(n6343) );
  INV_X1 U3953 ( .A(n4356), .ZN(n6485) );
  AND2_X1 U3954 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n3998), .ZN(n3999)
         );
  NOR2_X1 U3955 ( .A1(n3915), .A2(n5477), .ZN(n3916) );
  INV_X1 U3956 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5029) );
  INV_X1 U3957 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U3958 ( .A1(n3868), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3915)
         );
  AND2_X1 U3959 ( .A1(n5013), .A2(n5011), .ZN(n5012) );
  NAND2_X1 U3960 ( .A1(n3843), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3814)
         );
  INV_X1 U3961 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5247) );
  INV_X1 U3962 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4555) );
  INV_X1 U3963 ( .A(n4898), .ZN(n4899) );
  AOI21_X1 U3964 ( .B1(n5323), .B2(n5572), .A(n5332), .ZN(n4906) );
  OR2_X1 U3965 ( .A1(n5929), .A2(n4317), .ZN(n5563) );
  INV_X1 U3966 ( .A(n5925), .ZN(n5385) );
  INV_X1 U3967 ( .A(n5917), .ZN(n6684) );
  OR2_X1 U3968 ( .A1(n3074), .A2(n4526), .ZN(n5956) );
  OR2_X1 U3969 ( .A1(n5424), .A2(n4526), .ZN(n4537) );
  INV_X1 U3970 ( .A(n4801), .ZN(n4838) );
  NAND2_X1 U3971 ( .A1(n3074), .A2(n4524), .ZN(n5424) );
  OAI21_X1 U3972 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6458), .A(n4803), 
        .ZN(n6191) );
  INV_X1 U3973 ( .A(n4526), .ZN(n4609) );
  NAND3_X1 U3975 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6368), .A3(n4523), .ZN(
        n4740) );
  INV_X1 U3976 ( .A(n4052), .ZN(n4207) );
  OR2_X1 U3977 ( .A1(n4354), .A2(n6374), .ZN(n5432) );
  INV_X1 U3978 ( .A(n6382), .ZN(n6486) );
  NOR2_X1 U3979 ( .A1(n4239), .A2(n4243), .ZN(n4244) );
  NAND2_X1 U3980 ( .A1(n3999), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4023)
         );
  NAND2_X1 U3981 ( .A1(n3916), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3955)
         );
  NAND2_X1 U3982 ( .A1(n3794), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3793)
         );
  INV_X1 U3983 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4342) );
  OR2_X1 U3984 ( .A1(n6481), .A2(n4210), .ZN(n5755) );
  AND2_X1 U3985 ( .A1(n4974), .A2(n4228), .ZN(n5743) );
  INV_X2 U3986 ( .A(n4108), .ZN(n4897) );
  AND2_X1 U3987 ( .A1(n5098), .A2(n5097), .ZN(n5534) );
  INV_X1 U3988 ( .A(n5151), .ZN(n5783) );
  AND2_X1 U3989 ( .A1(n5151), .A2(n4386), .ZN(n5148) );
  NOR2_X1 U3990 ( .A1(n5787), .A2(n5837), .ZN(n5805) );
  NAND2_X1 U3991 ( .A1(n4092), .A2(n4091), .ZN(n4093) );
  NAND2_X1 U3992 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n3956), .ZN(n3997)
         );
  AND2_X1 U3993 ( .A1(n3779), .A2(n3778), .ZN(n5013) );
  AND2_X1 U3994 ( .A1(n5118), .A2(n5117), .ZN(n5654) );
  INV_X1 U3995 ( .A(n5914), .ZN(n5897) );
  XNOR2_X1 U3996 ( .A(n4900), .B(n4899), .ZN(n4983) );
  AOI21_X1 U3997 ( .B1(n5228), .B2(n5183), .A(n5197), .ZN(n5193) );
  INV_X1 U3998 ( .A(n5940), .ZN(n5342) );
  NOR3_X1 U3999 ( .A1(n4316), .A2(n4315), .A3(n4470), .ZN(n5368) );
  INV_X1 U4000 ( .A(n5394), .ZN(n5951) );
  INV_X1 U4001 ( .A(n6464), .ZN(n6271) );
  OAI21_X1 U4002 ( .B1(n5989), .B2(n5966), .A(n5965), .ZN(n5984) );
  INV_X1 U4003 ( .A(n6017), .ZN(n6001) );
  OAI21_X1 U4004 ( .B1(n6044), .B2(n6028), .A(n6136), .ZN(n6046) );
  INV_X1 U4005 ( .A(n4714), .ZN(n4793) );
  INV_X1 U4006 ( .A(n4808), .ZN(n6080) );
  OR2_X1 U4007 ( .A1(n6191), .A2(n4570), .ZN(n6171) );
  AND2_X1 U4008 ( .A1(n6185), .A2(n6465), .ZN(n6263) );
  AND2_X1 U4009 ( .A1(n6376), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3567) );
  NOR2_X1 U4010 ( .A1(n6376), .A2(n6367), .ZN(n6462) );
  INV_X1 U4011 ( .A(n6449), .ZN(n6443) );
  INV_X1 U4012 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6224) );
  AND2_X1 U4013 ( .A1(n3080), .A2(n4244), .ZN(n4245) );
  INV_X1 U4014 ( .A(n5743), .ZN(n5761) );
  INV_X1 U4015 ( .A(n5758), .ZN(n5671) );
  NAND2_X1 U4016 ( .A1(n5755), .A2(n4215), .ZN(n5695) );
  OR2_X1 U4017 ( .A1(n5543), .A2(n5109), .ZN(n5641) );
  NAND2_X1 U4018 ( .A1(n5776), .A2(n5127), .ZN(n5122) );
  OR2_X1 U4019 ( .A1(n5893), .A2(n4384), .ZN(n5151) );
  INV_X1 U4020 ( .A(n5805), .ZN(n5809) );
  OR2_X1 U4021 ( .A1(n5816), .A2(n5814), .ZN(n5824) );
  INV_X1 U4022 ( .A(n5814), .ZN(n5837) );
  INV_X1 U4023 ( .A(n5893), .ZN(n5890) );
  NOR2_X1 U4024 ( .A1(n4094), .A2(n4093), .ZN(n4095) );
  OAI21_X1 U4025 ( .B1(n5014), .B2(n5013), .A(n5096), .ZN(n5222) );
  AND2_X1 U4026 ( .A1(n4329), .A2(n3081), .ZN(n4330) );
  NOR2_X1 U4027 ( .A1(n5341), .A2(n5368), .ZN(n5929) );
  NAND2_X1 U4028 ( .A1(n4304), .A2(n4287), .ZN(n5394) );
  INV_X1 U4029 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U4030 ( .A1(n6276), .A2(n5961), .ZN(n5979) );
  NAND2_X1 U4031 ( .A1(n5987), .A2(n3581), .ZN(n6017) );
  NAND2_X1 U4032 ( .A1(n5987), .A2(n6465), .ZN(n6049) );
  INV_X1 U4033 ( .A(n4704), .ZN(n4798) );
  INV_X1 U4034 ( .A(n4806), .ZN(n4843) );
  NAND2_X1 U4035 ( .A1(n6103), .A2(n3581), .ZN(n6125) );
  NAND2_X1 U4036 ( .A1(n6103), .A2(n6465), .ZN(n6162) );
  INV_X1 U4037 ( .A(n6156), .ZN(n6174) );
  INV_X1 U4038 ( .A(n6182), .ZN(n4773) );
  INV_X1 U4039 ( .A(n6263), .ZN(n6225) );
  NAND2_X1 U4040 ( .A1(n6276), .A2(n6219), .ZN(n6332) );
  INV_X1 U4041 ( .A(n6365), .ZN(n6457) );
  INV_X1 U4042 ( .A(n6455), .ZN(n6452) );
  INV_X1 U4043 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6392) );
  OAI21_X1 U4044 ( .B1(n5133), .B2(n5695), .A(n4245), .ZN(U2798) );
  OAI21_X1 U4045 ( .B1(n3069), .B2(n5126), .A(n4195), .ZN(U2829) );
  NAND2_X1 U4046 ( .A1(n3700), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3089) );
  NAND2_X1 U4047 ( .A1(n3087), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3088) );
  NAND2_X1 U4048 ( .A1(n3089), .A2(n3088), .ZN(n3094) );
  AND2_X2 U4049 ( .A1(n4452), .A2(n4427), .ZN(n3160) );
  NAND2_X1 U4050 ( .A1(n3160), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3092)
         );
  NAND2_X1 U4051 ( .A1(n3176), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3091)
         );
  NAND2_X1 U4052 ( .A1(n3204), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3098)
         );
  NAND2_X1 U4053 ( .A1(n3182), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3097) );
  AND2_X2 U4054 ( .A1(n4458), .A2(n4428), .ZN(n3263) );
  NAND2_X1 U4055 ( .A1(n3263), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3096) );
  NAND2_X1 U4056 ( .A1(n3290), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3095)
         );
  AND2_X2 U4057 ( .A1(n3103), .A2(n4433), .ZN(n3262) );
  NAND2_X1 U4058 ( .A1(n3262), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3102) );
  NAND2_X1 U4059 ( .A1(n3979), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3101) );
  NAND2_X1 U4060 ( .A1(n3894), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3100)
         );
  NAND2_X1 U4061 ( .A1(n3195), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3099)
         );
  AND2_X2 U4062 ( .A1(n4452), .A2(n4433), .ZN(n3175) );
  NAND2_X1 U4063 ( .A1(n3175), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3108) );
  NAND2_X1 U4064 ( .A1(n3278), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3107) );
  NAND2_X1 U4065 ( .A1(n3177), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3106) );
  INV_X1 U4066 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3104) );
  NAND2_X1 U4067 ( .A1(n3264), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3105) );
  AOI22_X1 U4068 ( .A1(n3176), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3160), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3115) );
  AOI22_X1 U4069 ( .A1(n3175), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3278), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3114) );
  AOI22_X1 U4070 ( .A1(n3177), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3264), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3113) );
  AOI22_X1 U4071 ( .A1(n3204), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3263), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3119) );
  AOI22_X1 U4072 ( .A1(n3262), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3118) );
  AOI22_X1 U4073 ( .A1(n3182), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3117) );
  NAND2_X1 U4074 ( .A1(n3176), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3125)
         );
  NAND2_X1 U4075 ( .A1(n3160), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3124)
         );
  INV_X1 U4076 ( .A(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3121) );
  NAND2_X1 U4077 ( .A1(n3700), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3122) );
  NAND2_X1 U4078 ( .A1(n3894), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3129)
         );
  NAND2_X1 U4079 ( .A1(n3262), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3128) );
  NAND2_X1 U4080 ( .A1(n3979), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3127) );
  NAND2_X1 U4081 ( .A1(n3195), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3126)
         );
  NAND2_X1 U4082 ( .A1(n3175), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3133) );
  NAND2_X1 U4083 ( .A1(n3278), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3132) );
  NAND2_X1 U4084 ( .A1(n3177), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3131) );
  NAND2_X1 U4085 ( .A1(n3264), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3130) );
  NAND2_X1 U4086 ( .A1(n3182), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3137) );
  NAND2_X1 U4087 ( .A1(n3204), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3136)
         );
  NAND2_X1 U4088 ( .A1(n3263), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3135) );
  NAND2_X1 U4089 ( .A1(n3290), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3134)
         );
  NAND2_X1 U4090 ( .A1(n4098), .A2(n3306), .ZN(n3150) );
  AOI22_X1 U4091 ( .A1(n3894), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3979), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3143) );
  AOI22_X1 U4092 ( .A1(n3262), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3142) );
  AOI22_X1 U4093 ( .A1(n3204), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3263), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3141) );
  AOI22_X1 U4094 ( .A1(n3182), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3140) );
  AOI22_X1 U4095 ( .A1(n3087), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3700), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3147) );
  AOI22_X1 U4096 ( .A1(n3176), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3160), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3146) );
  AOI22_X1 U4097 ( .A1(n3175), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3278), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3145) );
  AOI22_X1 U4098 ( .A1(n3177), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3264), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3144) );
  AOI22_X1 U4099 ( .A1(n3176), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3177), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3154) );
  AOI22_X1 U4100 ( .A1(n3700), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3263), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3153) );
  AOI22_X1 U4101 ( .A1(n3262), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3152) );
  AOI22_X1 U4102 ( .A1(n3204), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U4103 ( .A1(n4009), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3160), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3158) );
  AOI22_X1 U4104 ( .A1(n3984), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3157) );
  AOI22_X1 U4105 ( .A1(n3894), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3979), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3156) );
  AOI22_X1 U4106 ( .A1(n3278), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3264), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3155) );
  AOI22_X1 U4107 ( .A1(n4009), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3278), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3164) );
  AOI22_X1 U4108 ( .A1(n3176), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3160), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3163) );
  AOI22_X1 U4109 ( .A1(n3984), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3700), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3162) );
  AOI22_X1 U4110 ( .A1(n3177), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3264), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3161) );
  AOI22_X1 U4111 ( .A1(n3204), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3263), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3168) );
  AOI22_X1 U4112 ( .A1(n3894), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3979), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3167) );
  AOI22_X1 U4113 ( .A1(n3290), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        INSTQUEUE_REG_1__2__SCAN_IN), .B2(n3182), .ZN(n3166) );
  AOI22_X1 U4114 ( .A1(n3262), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3165) );
  NAND2_X2 U4115 ( .A1(n3079), .A2(n3085), .ZN(n3215) );
  AOI22_X1 U4116 ( .A1(n3204), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3979), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U4117 ( .A1(n3175), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3176), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3180) );
  AOI22_X1 U4118 ( .A1(n3700), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3263), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3179) );
  AOI22_X1 U4119 ( .A1(n3278), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3177), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3178) );
  NAND4_X1 U4120 ( .A1(n3181), .A2(n3180), .A3(n3179), .A4(n3178), .ZN(n3188)
         );
  AOI22_X1 U4121 ( .A1(n4067), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3185) );
  AOI22_X1 U4122 ( .A1(n3160), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3264), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3184) );
  AOI22_X1 U4123 ( .A1(n3262), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3183) );
  NAND4_X1 U4124 ( .A1(n3186), .A2(n3185), .A3(n3184), .A4(n3183), .ZN(n3187)
         );
  OR2_X2 U4125 ( .A1(n3188), .A2(n3187), .ZN(n3249) );
  NAND2_X1 U4126 ( .A1(n3176), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3194)
         );
  NAND2_X1 U4127 ( .A1(n3160), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3193)
         );
  INV_X1 U4128 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3190) );
  NAND2_X1 U4129 ( .A1(n3700), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3191) );
  NAND2_X1 U4130 ( .A1(n3894), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3199)
         );
  NAND2_X1 U4131 ( .A1(n3262), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3198) );
  NAND2_X1 U4132 ( .A1(n3979), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3197) );
  NAND2_X1 U4133 ( .A1(n3195), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3196)
         );
  NAND2_X1 U4134 ( .A1(n3278), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3203) );
  NAND2_X1 U4135 ( .A1(n3175), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3202) );
  NAND2_X1 U4136 ( .A1(n3177), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3201) );
  NAND2_X1 U4137 ( .A1(n3264), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3200) );
  NAND2_X1 U4138 ( .A1(n3182), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3208) );
  NAND2_X1 U4139 ( .A1(n3204), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3207)
         );
  NAND2_X1 U4140 ( .A1(n3263), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3206) );
  NAND2_X1 U4141 ( .A1(n3290), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3205)
         );
  NOR2_X1 U4142 ( .A1(n6529), .A2(n6392), .ZN(n6395) );
  INV_X1 U4143 ( .A(n6395), .ZN(n3213) );
  OAI21_X1 U4144 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n3213), .ZN(n4225) );
  NAND2_X1 U4145 ( .A1(n4102), .A2(n4225), .ZN(n3232) );
  INV_X1 U4146 ( .A(n3232), .ZN(n3225) );
  NOR2_X1 U4147 ( .A1(n3215), .A2(n4970), .ZN(n3214) );
  AND2_X2 U4148 ( .A1(n3574), .A2(n3573), .ZN(n3216) );
  INV_X1 U4149 ( .A(n3216), .ZN(n4275) );
  AOI22_X1 U4150 ( .A1(n3216), .A2(n3169), .B1(n3574), .B2(n3215), .ZN(n3219)
         );
  NAND2_X1 U4151 ( .A1(n3218), .A2(n3305), .ZN(n3248) );
  NAND2_X1 U4152 ( .A1(n3219), .A2(n3248), .ZN(n3223) );
  NAND3_X1 U4153 ( .A1(n3580), .A2(n3306), .A3(n3220), .ZN(n3221) );
  NAND2_X1 U4154 ( .A1(n3221), .A2(n3215), .ZN(n3222) );
  INV_X1 U4155 ( .A(n4098), .ZN(n3233) );
  NAND2_X1 U4156 ( .A1(n3572), .A2(n5787), .ZN(n3224) );
  NAND2_X1 U4157 ( .A1(n4198), .A2(n4550), .ZN(n4285) );
  NAND2_X1 U4158 ( .A1(n5597), .A2(n6368), .ZN(n4086) );
  INV_X1 U4159 ( .A(n4086), .ZN(n3345) );
  XNOR2_X1 U4160 ( .A(n6468), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6138)
         );
  NAND2_X1 U4161 ( .A1(n3345), .A2(n6138), .ZN(n3227) );
  INV_X1 U4162 ( .A(n3567), .ZN(n3344) );
  NAND2_X1 U4163 ( .A1(n3344), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3226) );
  NAND2_X1 U4164 ( .A1(n3227), .A2(n3226), .ZN(n3239) );
  NAND2_X1 U4165 ( .A1(n3228), .A2(n3076), .ZN(n3319) );
  NAND2_X1 U4166 ( .A1(n4097), .A2(n4356), .ZN(n3231) );
  AND2_X2 U4167 ( .A1(n4303), .A2(n3419), .ZN(n4120) );
  NAND2_X1 U4168 ( .A1(n4120), .A2(n3572), .ZN(n4297) );
  NAND2_X1 U4169 ( .A1(n3231), .A2(n4297), .ZN(n3253) );
  NAND2_X1 U4170 ( .A1(n3232), .A2(n4597), .ZN(n3234) );
  NAND2_X1 U4171 ( .A1(n3233), .A2(n3305), .ZN(n3245) );
  NAND2_X1 U4172 ( .A1(n3234), .A2(n3245), .ZN(n3235) );
  NOR2_X1 U4173 ( .A1(n3253), .A2(n3235), .ZN(n3236) );
  NAND3_X1 U4174 ( .A1(n3236), .A2(n3259), .A3(n3568), .ZN(n3237) );
  INV_X1 U4175 ( .A(n3244), .ZN(n3238) );
  NAND2_X1 U4176 ( .A1(n3238), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3242) );
  NAND3_X1 U4177 ( .A1(n3242), .A2(n3241), .A3(n3240), .ZN(n3318) );
  NAND2_X1 U4178 ( .A1(n3319), .A2(n3318), .ZN(n3261) );
  MUX2_X1 U4179 ( .A(n3567), .B(n4086), .S(n6468), .Z(n3243) );
  INV_X1 U4180 ( .A(n3245), .ZN(n3246) );
  OAI21_X1 U4181 ( .B1(n3247), .B2(n3246), .A(n4303), .ZN(n3256) );
  NAND3_X1 U4182 ( .A1(n4602), .A2(n5787), .A3(n4101), .ZN(n4300) );
  NAND2_X1 U4183 ( .A1(n5597), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6375) );
  AOI21_X1 U4184 ( .B1(n3215), .B2(n3249), .A(n6375), .ZN(n3252) );
  NAND2_X1 U4185 ( .A1(n3250), .A2(n4356), .ZN(n3251) );
  OAI211_X1 U4186 ( .C1(n3248), .C2(n4300), .A(n3252), .B(n3251), .ZN(n3254)
         );
  NOR2_X1 U4187 ( .A1(n3254), .A2(n3253), .ZN(n3255) );
  INV_X1 U4188 ( .A(n3572), .ZN(n3257) );
  NOR2_X1 U4189 ( .A1(n3257), .A2(n4550), .ZN(n3258) );
  OR2_X1 U4190 ( .A1(n3259), .A2(n3258), .ZN(n4295) );
  XNOR2_X1 U4191 ( .A(n3261), .B(n3317), .ZN(n4425) );
  NAND2_X1 U4192 ( .A1(n4425), .A2(n6368), .ZN(n3276) );
  AOI22_X1 U4193 ( .A1(n4060), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U4194 ( .A1(n3072), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3267) );
  AOI22_X1 U4195 ( .A1(n4036), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3266) );
  AOI22_X1 U4196 ( .A1(n4058), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3265) );
  NAND4_X1 U4197 ( .A1(n3268), .A2(n3267), .A3(n3266), .A4(n3265), .ZN(n3274)
         );
  AOI22_X1 U4198 ( .A1(n4072), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3272) );
  AOI22_X1 U4199 ( .A1(n3852), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4059), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3271) );
  AOI22_X1 U4200 ( .A1(n4070), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3270) );
  AOI22_X1 U4201 ( .A1(n4062), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3269) );
  NAND4_X1 U4202 ( .A1(n3272), .A2(n3271), .A3(n3270), .A4(n3269), .ZN(n3273)
         );
  NAND2_X1 U4203 ( .A1(n3302), .A2(n3417), .ZN(n3275) );
  NAND2_X1 U4204 ( .A1(n3276), .A2(n3275), .ZN(n3416) );
  AOI22_X1 U4205 ( .A1(n4009), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3282) );
  AOI22_X1 U4206 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n3984), .B1(n4058), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3281) );
  AOI22_X1 U4207 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n4070), .B1(n4057), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U4208 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n3852), .B1(n3195), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3279) );
  NAND4_X1 U4209 ( .A1(n3282), .A2(n3281), .A3(n3280), .A4(n3279), .ZN(n3288)
         );
  AOI22_X1 U4210 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n4062), .B1(n3978), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4211 ( .A1(n3072), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4212 ( .A1(n4059), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4213 ( .A1(n4036), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3283) );
  NAND4_X1 U4214 ( .A1(n3286), .A2(n3285), .A3(n3284), .A4(n3283), .ZN(n3287)
         );
  INV_X1 U4215 ( .A(n3489), .ZN(n3289) );
  NAND2_X1 U4216 ( .A1(n3302), .A2(n3289), .ZN(n3311) );
  AOI22_X1 U4217 ( .A1(n3894), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4036), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3294) );
  AOI22_X1 U4218 ( .A1(n3072), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3293) );
  AOI22_X1 U4219 ( .A1(n4072), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U4220 ( .A1(n3978), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3291) );
  NAND4_X1 U4221 ( .A1(n3294), .A2(n3293), .A3(n3292), .A4(n3291), .ZN(n3300)
         );
  AOI22_X1 U4222 ( .A1(n3984), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4223 ( .A1(n4060), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4059), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4224 ( .A1(n3700), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4225 ( .A1(n3852), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3295) );
  NAND4_X1 U4226 ( .A1(n3298), .A2(n3297), .A3(n3296), .A4(n3295), .ZN(n3299)
         );
  INV_X1 U4227 ( .A(n3418), .ZN(n3301) );
  NAND2_X1 U4228 ( .A1(n3302), .A2(n3489), .ZN(n3399) );
  OR2_X1 U4229 ( .A1(n3418), .A2(n3399), .ZN(n3303) );
  AND2_X1 U4230 ( .A1(n3403), .A2(n3399), .ZN(n3310) );
  NAND2_X1 U4231 ( .A1(n3306), .A2(n3489), .ZN(n3308) );
  NAND2_X1 U4232 ( .A1(n5787), .A2(n3418), .ZN(n3307) );
  NAND3_X1 U4233 ( .A1(n3308), .A2(n3307), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3309) );
  AOI21_X1 U4234 ( .B1(n3559), .B2(INSTQUEUE_REG_0__0__SCAN_IN), .A(n3309), 
        .ZN(n3404) );
  INV_X1 U4235 ( .A(n3414), .ZN(n3315) );
  NAND2_X1 U4236 ( .A1(n3417), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3313) );
  NAND2_X1 U4237 ( .A1(n3559), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3312) );
  OAI211_X1 U4238 ( .C1(n3249), .C2(n3313), .A(n3312), .B(n3311), .ZN(n3413)
         );
  INV_X1 U4239 ( .A(n3413), .ZN(n3314) );
  NAND2_X1 U4240 ( .A1(n3315), .A2(n3314), .ZN(n3316) );
  NAND2_X1 U4241 ( .A1(n3416), .A2(n3316), .ZN(n3427) );
  INV_X1 U4242 ( .A(n3427), .ZN(n3343) );
  NAND2_X1 U4243 ( .A1(n3318), .A2(n3317), .ZN(n3320) );
  NAND2_X1 U4244 ( .A1(n3320), .A2(n3319), .ZN(n3326) );
  NOR2_X1 U4245 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6337), .ZN(n4611)
         );
  NAND2_X1 U4246 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4611), .ZN(n4606) );
  NAND2_X1 U4247 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3322) );
  NAND2_X1 U4248 ( .A1(n3322), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3323) );
  NAND2_X1 U4249 ( .A1(n4606), .A2(n3323), .ZN(n4657) );
  AOI22_X1 U4250 ( .A1(n4657), .A2(n3345), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3344), .ZN(n3324) );
  INV_X1 U4251 ( .A(n3326), .ZN(n3329) );
  INV_X1 U4252 ( .A(n3327), .ZN(n3328) );
  NAND2_X1 U4253 ( .A1(n3329), .A2(n3328), .ZN(n3330) );
  NAND2_X1 U4254 ( .A1(n5406), .A2(n3330), .ZN(n4529) );
  AOI22_X1 U4255 ( .A1(n4058), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4256 ( .A1(n4062), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4257 ( .A1(n4072), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4258 ( .A1(n3979), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3332) );
  NAND4_X1 U4259 ( .A1(n3335), .A2(n3334), .A3(n3333), .A4(n3332), .ZN(n3341)
         );
  AOI22_X1 U4260 ( .A1(n3984), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3072), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4261 ( .A1(n4060), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4059), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4262 ( .A1(n4070), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3337) );
  AOI22_X1 U4263 ( .A1(n4036), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3336) );
  NAND4_X1 U4264 ( .A1(n3339), .A2(n3338), .A3(n3337), .A4(n3336), .ZN(n3340)
         );
  AOI22_X1 U4265 ( .A1(n3559), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3541), 
        .B2(n3428), .ZN(n3342) );
  NAND2_X1 U4266 ( .A1(n3343), .A2(n3426), .ZN(n3437) );
  INV_X1 U4267 ( .A(n3437), .ZN(n3360) );
  NOR3_X1 U4268 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6344), .A3(n6337), 
        .ZN(n6058) );
  NAND2_X1 U4269 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6058), .ZN(n6053) );
  NAND3_X1 U4270 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6274) );
  NOR2_X1 U4271 ( .A1(n6468), .A2(n6274), .ZN(n6325) );
  AOI21_X1 U4272 ( .B1(n6231), .B2(n6053), .A(n6325), .ZN(n4700) );
  AOI22_X1 U4273 ( .A1(n3345), .A2(n4700), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3344), .ZN(n3346) );
  NAND2_X1 U4274 ( .A1(n4450), .A2(n6368), .ZN(n3359) );
  AOI22_X1 U4275 ( .A1(n4072), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3351) );
  AOI22_X1 U4276 ( .A1(n3072), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3350) );
  AOI22_X1 U4277 ( .A1(n3984), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3349) );
  AOI22_X1 U4278 ( .A1(n4059), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3348) );
  NAND4_X1 U4279 ( .A1(n3351), .A2(n3350), .A3(n3349), .A4(n3348), .ZN(n3357)
         );
  AOI22_X1 U4280 ( .A1(n4070), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4281 ( .A1(n4062), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4282 ( .A1(n4036), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4283 ( .A1(n3978), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3352) );
  NAND4_X1 U4284 ( .A1(n3355), .A2(n3354), .A3(n3353), .A4(n3352), .ZN(n3356)
         );
  AOI22_X1 U4285 ( .A1(n3559), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3541), 
        .B2(n3439), .ZN(n3358) );
  NAND2_X1 U4286 ( .A1(n3559), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4287 ( .A1(n4060), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4288 ( .A1(n4036), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3363) );
  AOI22_X1 U4289 ( .A1(n4072), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4290 ( .A1(n4058), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3361) );
  NAND4_X1 U4291 ( .A1(n3364), .A2(n3363), .A3(n3362), .A4(n3361), .ZN(n3370)
         );
  AOI22_X1 U4292 ( .A1(n3984), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3072), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4293 ( .A1(n3852), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4059), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4294 ( .A1(n4062), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4295 ( .A1(n4070), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3365) );
  NAND4_X1 U4296 ( .A1(n3368), .A2(n3367), .A3(n3366), .A4(n3365), .ZN(n3369)
         );
  NAND2_X1 U4297 ( .A1(n3541), .A2(n3455), .ZN(n3371) );
  NAND2_X1 U4298 ( .A1(n3372), .A2(n3371), .ZN(n3444) );
  INV_X1 U4299 ( .A(n3444), .ZN(n3373) );
  NAND2_X1 U4300 ( .A1(n3559), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3385) );
  AOI22_X1 U4301 ( .A1(n4072), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4302 ( .A1(n3072), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4303 ( .A1(n3984), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U4304 ( .A1(n4059), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3374) );
  NAND4_X1 U4305 ( .A1(n3377), .A2(n3376), .A3(n3375), .A4(n3374), .ZN(n3383)
         );
  INV_X1 U4306 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n6517) );
  AOI22_X1 U4307 ( .A1(n4070), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4308 ( .A1(n4062), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3380) );
  AOI22_X1 U4309 ( .A1(n4036), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3379) );
  AOI22_X1 U4310 ( .A1(n3978), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3378) );
  NAND4_X1 U4311 ( .A1(n3381), .A2(n3380), .A3(n3379), .A4(n3378), .ZN(n3382)
         );
  NAND2_X1 U4312 ( .A1(n3541), .A2(n3458), .ZN(n3384) );
  NAND2_X1 U4313 ( .A1(n3385), .A2(n3384), .ZN(n3452) );
  NAND2_X1 U4314 ( .A1(n3453), .A2(n3452), .ZN(n3466) );
  NAND2_X1 U4315 ( .A1(n3559), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3397) );
  AOI22_X1 U4316 ( .A1(n3072), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4317 ( .A1(n3700), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4318 ( .A1(n4070), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3387) );
  AOI22_X1 U4319 ( .A1(n4072), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3386) );
  NAND4_X1 U4320 ( .A1(n3389), .A2(n3388), .A3(n3387), .A4(n3386), .ZN(n3395)
         );
  AOI22_X1 U4321 ( .A1(n4060), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4059), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4322 ( .A1(n3984), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3392) );
  AOI22_X1 U4323 ( .A1(n4036), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3391) );
  AOI22_X1 U4324 ( .A1(n3852), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3390) );
  NAND4_X1 U4325 ( .A1(n3393), .A2(n3392), .A3(n3391), .A4(n3390), .ZN(n3394)
         );
  NAND2_X1 U4326 ( .A1(n3541), .A2(n3480), .ZN(n3396) );
  NOR2_X1 U4327 ( .A1(n3399), .A2(n3461), .ZN(n3400) );
  NOR2_X1 U4328 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5344) );
  NOR2_X1 U4329 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5325) );
  INV_X1 U4330 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5315) );
  INV_X1 U4331 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6606) );
  NAND4_X1 U4332 ( .A1(n5344), .A2(n5325), .A3(n5315), .A4(n6606), .ZN(n3401)
         );
  INV_X1 U4333 ( .A(n3404), .ZN(n3406) );
  NAND2_X1 U4334 ( .A1(n4536), .A2(n3527), .ZN(n3410) );
  NAND2_X1 U4335 ( .A1(n5787), .A2(n3419), .ZN(n3431) );
  OAI21_X1 U4336 ( .B1(n6485), .B2(n3418), .A(n3431), .ZN(n3408) );
  INV_X1 U4337 ( .A(n3408), .ZN(n3409) );
  INV_X1 U4338 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4930) );
  NAND2_X1 U4339 ( .A1(n4481), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4482)
         );
  NAND2_X1 U4340 ( .A1(n4482), .A2(n4109), .ZN(n3412) );
  NAND2_X1 U4341 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5941) );
  INV_X1 U4342 ( .A(n5941), .ZN(n3411) );
  NAND2_X1 U4343 ( .A1(n4481), .A2(n3411), .ZN(n3425) );
  AND2_X1 U4344 ( .A1(n3412), .A2(n3425), .ZN(n4336) );
  XNOR2_X1 U4345 ( .A(n3068), .B(n3413), .ZN(n3415) );
  XNOR2_X1 U4346 ( .A(n3416), .B(n3415), .ZN(n4525) );
  NAND2_X1 U4347 ( .A1(n4525), .A2(n3527), .ZN(n3424) );
  NAND2_X1 U4348 ( .A1(n3418), .A2(n3417), .ZN(n3429) );
  OAI21_X1 U4349 ( .B1(n3418), .B2(n3417), .A(n3429), .ZN(n3421) );
  NOR2_X1 U4350 ( .A1(n4597), .A2(n3215), .ZN(n3420) );
  OAI211_X1 U4351 ( .C1(n3421), .C2(n6485), .A(n3420), .B(n3419), .ZN(n3422)
         );
  INV_X1 U4352 ( .A(n3422), .ZN(n3423) );
  NAND2_X1 U4353 ( .A1(n3424), .A2(n3423), .ZN(n4335) );
  NAND2_X1 U4354 ( .A1(n4336), .A2(n4335), .ZN(n4334) );
  NAND2_X1 U4355 ( .A1(n4334), .A2(n3425), .ZN(n5908) );
  NAND2_X1 U4356 ( .A1(n3589), .A2(n3527), .ZN(n3435) );
  INV_X1 U4357 ( .A(n3428), .ZN(n3430) );
  NAND2_X1 U4358 ( .A1(n3429), .A2(n3430), .ZN(n3438) );
  OAI21_X1 U4359 ( .B1(n3430), .B2(n3429), .A(n3438), .ZN(n3433) );
  INV_X1 U4360 ( .A(n3431), .ZN(n3432) );
  AOI21_X1 U4361 ( .B1(n3433), .B2(n4356), .A(n3432), .ZN(n3434) );
  NAND2_X1 U4362 ( .A1(n3435), .A2(n3434), .ZN(n3436) );
  AND2_X1 U4363 ( .A1(n3436), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n5904)
         );
  OR2_X1 U4364 ( .A1(n3436), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n5905)
         );
  NAND2_X1 U4365 ( .A1(n3597), .A2(n3527), .ZN(n3441) );
  NAND2_X1 U4366 ( .A1(n3438), .A2(n3439), .ZN(n3457) );
  OAI211_X1 U4367 ( .C1(n3439), .C2(n3438), .A(n3457), .B(n4356), .ZN(n3440)
         );
  NAND2_X1 U4368 ( .A1(n3442), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3443)
         );
  NAND2_X1 U4369 ( .A1(n3613), .A2(n3527), .ZN(n3447) );
  XNOR2_X1 U4370 ( .A(n3457), .B(n3455), .ZN(n3445) );
  NAND2_X1 U4371 ( .A1(n3445), .A2(n4356), .ZN(n3446) );
  INV_X1 U4372 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3448) );
  NAND2_X1 U4373 ( .A1(n3449), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3450)
         );
  NAND2_X1 U4374 ( .A1(n3466), .A2(n3454), .ZN(n3616) );
  INV_X1 U4375 ( .A(n3455), .ZN(n3456) );
  NOR2_X1 U4376 ( .A1(n3457), .A2(n3456), .ZN(n3459) );
  NAND2_X1 U4377 ( .A1(n3459), .A2(n3458), .ZN(n3479) );
  OAI211_X1 U4378 ( .C1(n3459), .C2(n3458), .A(n3479), .B(n4356), .ZN(n3460)
         );
  INV_X1 U4379 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4471) );
  XNOR2_X1 U4380 ( .A(n3462), .B(n4471), .ZN(n4468) );
  NAND2_X1 U4381 ( .A1(n4467), .A2(n4468), .ZN(n3464) );
  NAND2_X1 U4382 ( .A1(n3462), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3463)
         );
  NAND2_X1 U4383 ( .A1(n3464), .A2(n3463), .ZN(n4494) );
  NAND2_X1 U4384 ( .A1(n3466), .A2(n3465), .ZN(n3633) );
  NAND3_X1 U4385 ( .A1(n3478), .A2(n3633), .A3(n3527), .ZN(n3469) );
  XNOR2_X1 U4386 ( .A(n3479), .B(n3480), .ZN(n3467) );
  NAND2_X1 U4387 ( .A1(n3467), .A2(n4356), .ZN(n3468) );
  NAND2_X1 U4388 ( .A1(n3469), .A2(n3468), .ZN(n3471) );
  INV_X1 U4389 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3470) );
  XNOR2_X1 U4390 ( .A(n3471), .B(n3470), .ZN(n4495) );
  NAND2_X1 U4391 ( .A1(n4494), .A2(n4495), .ZN(n3473) );
  NAND2_X1 U4392 ( .A1(n3471), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3472)
         );
  INV_X1 U4393 ( .A(n3559), .ZN(n3476) );
  INV_X1 U4394 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3475) );
  NAND2_X1 U4395 ( .A1(n3541), .A2(n3489), .ZN(n3474) );
  OAI21_X1 U4396 ( .B1(n3476), .B2(n3475), .A(n3474), .ZN(n3477) );
  XNOR2_X1 U4397 ( .A(n3478), .B(n3477), .ZN(n3634) );
  NAND2_X1 U4398 ( .A1(n3634), .A2(n3527), .ZN(n3484) );
  INV_X1 U4399 ( .A(n3479), .ZN(n3481) );
  NAND2_X1 U4400 ( .A1(n3481), .A2(n3480), .ZN(n3488) );
  XNOR2_X1 U4401 ( .A(n3488), .B(n3489), .ZN(n3482) );
  NAND2_X1 U4402 ( .A1(n3482), .A2(n4356), .ZN(n3483) );
  NAND2_X1 U4403 ( .A1(n3484), .A2(n3483), .ZN(n3485) );
  INV_X1 U4404 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5938) );
  XNOR2_X1 U4405 ( .A(n3485), .B(n5938), .ZN(n4641) );
  NAND2_X1 U4406 ( .A1(n4640), .A2(n4641), .ZN(n3487) );
  NAND2_X1 U4407 ( .A1(n3485), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3486)
         );
  NAND2_X1 U4408 ( .A1(n3487), .A2(n3486), .ZN(n4774) );
  INV_X1 U4409 ( .A(n3488), .ZN(n3490) );
  NAND3_X1 U4410 ( .A1(n3490), .A2(n4356), .A3(n3489), .ZN(n3491) );
  NAND2_X1 U4411 ( .A1(n3497), .A2(n3491), .ZN(n3492) );
  INV_X1 U4412 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4780) );
  XNOR2_X1 U4413 ( .A(n3492), .B(n4780), .ZN(n4775) );
  NAND2_X1 U4414 ( .A1(n4774), .A2(n4775), .ZN(n3494) );
  NAND2_X1 U4415 ( .A1(n3492), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3493)
         );
  NAND2_X1 U4416 ( .A1(n3494), .A2(n3493), .ZN(n4748) );
  XNOR2_X1 U4417 ( .A(n5228), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4749)
         );
  NAND2_X1 U4418 ( .A1(n4748), .A2(n4749), .ZN(n3496) );
  NAND2_X1 U4419 ( .A1(n3075), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3495)
         );
  NAND2_X1 U4420 ( .A1(n3496), .A2(n3495), .ZN(n4865) );
  CLKBUF_X3 U4421 ( .A(n3497), .Z(n5228) );
  INV_X1 U4422 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3498) );
  NAND2_X1 U4423 ( .A1(n5228), .A2(n3498), .ZN(n4864) );
  NAND2_X1 U4424 ( .A1(n4865), .A2(n4864), .ZN(n5253) );
  INV_X1 U4425 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U4426 ( .A1(n3075), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U4427 ( .A1(n3075), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3499) );
  INV_X1 U4428 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3500) );
  NAND2_X1 U4429 ( .A1(n5228), .A2(n3500), .ZN(n3501) );
  XNOR2_X1 U4430 ( .A(n5228), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5245)
         );
  INV_X1 U4431 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U4432 ( .A1(n5228), .A2(n5373), .ZN(n3502) );
  INV_X1 U4433 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5238) );
  OAI21_X1 U4434 ( .B1(n5227), .B2(n3503), .A(n5228), .ZN(n3507) );
  NOR2_X1 U4435 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3504) );
  NAND2_X1 U4436 ( .A1(n5227), .A2(n3504), .ZN(n3505) );
  NAND2_X1 U4437 ( .A1(n3507), .A2(n3505), .ZN(n4254) );
  NOR2_X1 U4438 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3506) );
  NAND2_X1 U4439 ( .A1(n4254), .A2(n3506), .ZN(n5215) );
  OAI21_X1 U4440 ( .B1(n5215), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n3075), 
        .ZN(n3510) );
  NAND2_X1 U4441 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4909) );
  INV_X1 U4442 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5574) );
  NOR2_X1 U4443 ( .A1(n4909), .A2(n5574), .ZN(n3508) );
  NAND2_X1 U4444 ( .A1(n3507), .A2(n3508), .ZN(n3509) );
  NAND2_X1 U4445 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U4446 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5346) );
  NOR2_X1 U4447 ( .A1(n5323), .A2(n5346), .ZN(n4256) );
  AND2_X1 U4448 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4907) );
  NAND2_X1 U4449 ( .A1(n4256), .A2(n4907), .ZN(n4912) );
  XOR2_X1 U4450 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(n5228), .Z(n5525) );
  INV_X1 U4451 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5559) );
  NOR2_X1 U4452 ( .A1(n5228), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5177)
         );
  NOR2_X1 U4453 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3513) );
  NAND2_X1 U4454 ( .A1(n5177), .A2(n3513), .ZN(n4901) );
  AND2_X1 U4455 ( .A1(n5228), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5176)
         );
  NAND2_X1 U4456 ( .A1(n3514), .A2(n5176), .ZN(n5170) );
  NAND2_X1 U4457 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4914) );
  XNOR2_X1 U4458 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3537) );
  NAND2_X1 U4459 ( .A1(n3537), .A2(n3538), .ZN(n3536) );
  NAND2_X1 U4460 ( .A1(n6337), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3516) );
  NAND2_X1 U4461 ( .A1(n3536), .A2(n3516), .ZN(n3531) );
  XNOR2_X1 U4462 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3529) );
  NAND2_X1 U4463 ( .A1(n3531), .A2(n3529), .ZN(n3518) );
  NAND2_X1 U4464 ( .A1(n6344), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3517) );
  XNOR2_X1 U4465 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3533) );
  NAND2_X1 U4466 ( .A1(n3532), .A2(n3533), .ZN(n3520) );
  NAND2_X1 U4467 ( .A1(n6231), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3519) );
  NAND2_X1 U4468 ( .A1(n3520), .A2(n3519), .ZN(n3526) );
  INV_X1 U4469 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3522) );
  NAND2_X1 U4470 ( .A1(n3522), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3523) );
  AND2_X1 U4471 ( .A1(n4970), .A2(n4550), .ZN(n3528) );
  INV_X1 U4472 ( .A(n3529), .ZN(n3530) );
  XNOR2_X1 U4473 ( .A(n3531), .B(n3530), .ZN(n4200) );
  XOR2_X1 U4474 ( .A(n3533), .B(n3532), .Z(n4201) );
  INV_X1 U4475 ( .A(n4200), .ZN(n3534) );
  AOI22_X1 U4476 ( .A1(n3535), .A2(n4201), .B1(n3559), .B2(n3534), .ZN(n3557)
         );
  OAI21_X1 U4477 ( .B1(n3538), .B2(n3537), .A(n3536), .ZN(n3549) );
  INV_X1 U4478 ( .A(n3549), .ZN(n4199) );
  INV_X1 U4479 ( .A(n3554), .ZN(n3540) );
  XNOR2_X1 U4480 ( .A(n3057), .B(n6468), .ZN(n3543) );
  OAI21_X1 U4481 ( .B1(n3572), .B2(n3543), .A(n3249), .ZN(n3539) );
  NAND2_X1 U4482 ( .A1(n3540), .A2(n3539), .ZN(n3544) );
  INV_X1 U4483 ( .A(n3544), .ZN(n3547) );
  NAND2_X1 U4484 ( .A1(n3541), .A2(n4303), .ZN(n3542) );
  NAND2_X1 U4485 ( .A1(n3542), .A2(n4970), .ZN(n3548) );
  NOR2_X1 U4486 ( .A1(n3563), .A2(n3543), .ZN(n3545) );
  OAI211_X1 U4487 ( .C1(n4199), .C2(n3548), .A(n3545), .B(n3544), .ZN(n3546)
         );
  AOI22_X1 U4488 ( .A1(n4199), .A2(n3547), .B1(n3564), .B2(n3546), .ZN(n3552)
         );
  INV_X1 U4489 ( .A(n3548), .ZN(n3550) );
  NOR3_X1 U4490 ( .A1(n3550), .A2(n6368), .A3(n3549), .ZN(n3551) );
  AOI21_X1 U4491 ( .B1(n3555), .B2(n3554), .A(n3553), .ZN(n3556) );
  OAI22_X1 U4492 ( .A1(n3557), .A2(n3556), .B1(n4201), .B2(n3564), .ZN(n3558)
         );
  OAI21_X1 U4493 ( .B1(n3559), .B2(n4204), .A(n3558), .ZN(n3560) );
  OAI21_X1 U4494 ( .B1(n4204), .B2(n3564), .A(n3560), .ZN(n3561) );
  OAI21_X1 U4495 ( .B1(n4203), .B2(n3563), .A(n3562), .ZN(n3566) );
  INV_X1 U4496 ( .A(n3568), .ZN(n3571) );
  AND2_X1 U4497 ( .A1(n4429), .A2(n5787), .ZN(n3570) );
  NOR2_X2 U4498 ( .A1(n3573), .A2(n6367), .ZN(n3842) );
  NAND2_X1 U4499 ( .A1(n4525), .A2(n3842), .ZN(n3579) );
  AND2_X1 U4500 ( .A1(n3216), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3606) );
  NAND2_X1 U4501 ( .A1(n3606), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3577) );
  NOR2_X2 U4502 ( .A1(n3574), .A2(n6367), .ZN(n3575) );
  AOI22_X1 U4503 ( .A1(n4954), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6367), .ZN(n3576) );
  AND2_X1 U4504 ( .A1(n3577), .A2(n3576), .ZN(n3578) );
  NAND2_X1 U4505 ( .A1(n3579), .A2(n3578), .ZN(n4392) );
  INV_X1 U4506 ( .A(n3580), .ZN(n4298) );
  INV_X1 U4507 ( .A(n3842), .ZN(n3828) );
  OR2_X1 U4508 ( .A1(n3582), .A2(n3828), .ZN(n3586) );
  NAND2_X1 U4509 ( .A1(n3606), .A2(n3057), .ZN(n3584) );
  AOI22_X1 U4510 ( .A1(n4954), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6367), .ZN(n3583) );
  AND2_X1 U4511 ( .A1(n3584), .A2(n3583), .ZN(n3585) );
  NAND2_X1 U4512 ( .A1(n3586), .A2(n3585), .ZN(n4375) );
  NAND2_X1 U4513 ( .A1(n4376), .A2(n4375), .ZN(n4374) );
  INV_X1 U4514 ( .A(n4375), .ZN(n3587) );
  NAND2_X1 U4515 ( .A1(n3587), .A2(n4025), .ZN(n3588) );
  NAND2_X1 U4516 ( .A1(n4374), .A2(n3588), .ZN(n4391) );
  NAND2_X1 U4517 ( .A1(n4392), .A2(n4391), .ZN(n4394) );
  AOI21_X1 U4518 ( .B1(n3589), .B2(n3842), .A(n4953), .ZN(n3592) );
  INV_X1 U4519 ( .A(n3606), .ZN(n3602) );
  NAND2_X1 U4520 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3598) );
  OAI21_X1 U4521 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3598), .ZN(n5913) );
  AOI22_X1 U4522 ( .A1(n4953), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n4207), 
        .B2(n5913), .ZN(n3591) );
  NAND2_X1 U4523 ( .A1(n4954), .A2(EAX_REG_2__SCAN_IN), .ZN(n3590) );
  OAI211_X1 U4524 ( .C1(n3602), .C2(n3321), .A(n3591), .B(n3590), .ZN(n4390)
         );
  NAND2_X1 U4525 ( .A1(n4389), .A2(n4390), .ZN(n3596) );
  INV_X1 U4526 ( .A(n3592), .ZN(n3594) );
  NAND2_X1 U4527 ( .A1(n3597), .A2(n3842), .ZN(n3605) );
  OAI21_X1 U4528 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3599), .A(n3608), 
        .ZN(n5741) );
  AOI22_X1 U4529 ( .A1(n4207), .A2(n5741), .B1(n4953), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3601) );
  NAND2_X1 U4530 ( .A1(n4954), .A2(EAX_REG_3__SCAN_IN), .ZN(n3600) );
  OAI211_X1 U4531 ( .C1(n3602), .C2(n3104), .A(n3601), .B(n3600), .ZN(n3603)
         );
  INV_X1 U4532 ( .A(n3603), .ZN(n3604) );
  NAND2_X1 U4533 ( .A1(n3605), .A2(n3604), .ZN(n4439) );
  NAND2_X1 U4534 ( .A1(n4387), .A2(n4439), .ZN(n4396) );
  INV_X1 U4535 ( .A(n4396), .ZN(n3615) );
  NAND2_X1 U4536 ( .A1(n3606), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3611) );
  AOI21_X1 U4537 ( .B1(n4555), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3607) );
  AOI21_X1 U4538 ( .B1(n3575), .B2(EAX_REG_4__SCAN_IN), .A(n3607), .ZN(n3610)
         );
  NAND2_X1 U4539 ( .A1(n4555), .A2(n3608), .ZN(n3609) );
  INV_X1 U4540 ( .A(n3617), .ZN(n3618) );
  AND2_X1 U4541 ( .A1(n3609), .A2(n3618), .ZN(n5722) );
  AOI22_X1 U4542 ( .A1(n3611), .A2(n3610), .B1(n4207), .B2(n5722), .ZN(n3612)
         );
  AOI21_X1 U4543 ( .B1(n3613), .B2(n3842), .A(n3612), .ZN(n4397) );
  NAND2_X1 U4544 ( .A1(n3615), .A2(n3614), .ZN(n4395) );
  INV_X1 U4545 ( .A(n3616), .ZN(n3624) );
  INV_X1 U4546 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3622) );
  INV_X1 U4547 ( .A(n3625), .ZN(n3626) );
  INV_X1 U4548 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3619) );
  NAND2_X1 U4549 ( .A1(n3619), .A2(n3618), .ZN(n3620) );
  NAND2_X1 U4550 ( .A1(n3626), .A2(n3620), .ZN(n5721) );
  AOI22_X1 U4551 ( .A1(n5721), .A2(n4025), .B1(n4953), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3621) );
  OAI21_X1 U4552 ( .B1(n3847), .B2(n3622), .A(n3621), .ZN(n3623) );
  AOI21_X1 U4553 ( .B1(n3624), .B2(n3842), .A(n3623), .ZN(n4445) );
  INV_X1 U4554 ( .A(n3635), .ZN(n3628) );
  INV_X1 U4555 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3629) );
  NAND2_X1 U4556 ( .A1(n3626), .A2(n3629), .ZN(n3627) );
  NAND2_X1 U4557 ( .A1(n3628), .A2(n3627), .ZN(n5705) );
  INV_X1 U4558 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3630) );
  OAI22_X1 U4559 ( .A1(n3847), .A2(n3630), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3629), .ZN(n3631) );
  MUX2_X1 U4560 ( .A(n5705), .B(n3631), .S(n4052), .Z(n3632) );
  INV_X1 U4561 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3638) );
  NAND2_X1 U4562 ( .A1(n3634), .A2(n3842), .ZN(n3637) );
  OAI21_X1 U4563 ( .B1(n3635), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3652), 
        .ZN(n5694) );
  AOI22_X1 U4564 ( .A1(n5694), .A2(n4025), .B1(n4953), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3636) );
  OAI211_X1 U4565 ( .C1(n3847), .C2(n3638), .A(n3637), .B(n3636), .ZN(n4563)
         );
  NAND2_X1 U4566 ( .A1(n3067), .A2(n4563), .ZN(n4346) );
  AOI22_X1 U4567 ( .A1(n3984), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3072), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4568 ( .A1(n4057), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4569 ( .A1(n4060), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4570 ( .A1(n4070), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3639) );
  NAND4_X1 U4571 ( .A1(n3642), .A2(n3641), .A3(n3640), .A4(n3639), .ZN(n3648)
         );
  AOI22_X1 U4572 ( .A1(n4036), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4573 ( .A1(n4058), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4574 ( .A1(n4072), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4059), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4575 ( .A1(n3978), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3643) );
  NAND4_X1 U4576 ( .A1(n3646), .A2(n3645), .A3(n3644), .A4(n3643), .ZN(n3647)
         );
  OAI21_X1 U4577 ( .B1(n3648), .B2(n3647), .A(n3842), .ZN(n3651) );
  XOR2_X1 U4578 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3652), .Z(n4847) );
  AOI22_X1 U4579 ( .A1(n4953), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n4207), 
        .B2(n4847), .ZN(n3650) );
  NAND2_X1 U4580 ( .A1(n4954), .A2(EAX_REG_8__SCAN_IN), .ZN(n3649) );
  XNOR2_X1 U4581 ( .A(n3667), .B(n5682), .ZN(n5687) );
  AOI22_X1 U4582 ( .A1(n3072), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4583 ( .A1(n4070), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3655) );
  AOI22_X1 U4584 ( .A1(n4062), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4585 ( .A1(n4060), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4059), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3653) );
  NAND4_X1 U4586 ( .A1(n3656), .A2(n3655), .A3(n3654), .A4(n3653), .ZN(n3662)
         );
  AOI22_X1 U4587 ( .A1(n3984), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4588 ( .A1(n4036), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3659) );
  AOI22_X1 U4589 ( .A1(n4072), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4590 ( .A1(n3978), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3657) );
  NAND4_X1 U4591 ( .A1(n3660), .A2(n3659), .A3(n3658), .A4(n3657), .ZN(n3661)
         );
  NOR2_X1 U4592 ( .A1(n3662), .A2(n3661), .ZN(n3665) );
  NAND2_X1 U4593 ( .A1(n4954), .A2(EAX_REG_9__SCAN_IN), .ZN(n3664) );
  NAND2_X1 U4594 ( .A1(n4953), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3663)
         );
  OAI211_X1 U4595 ( .C1(n3828), .C2(n3665), .A(n3664), .B(n3663), .ZN(n3666)
         );
  AOI21_X1 U4596 ( .B1(n4207), .B2(n5687), .A(n3666), .ZN(n4799) );
  XOR2_X1 U4597 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3691), .Z(n5674) );
  AOI22_X1 U4598 ( .A1(n4058), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4599 ( .A1(n4070), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4600 ( .A1(n3177), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4601 ( .A1(n4062), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3668) );
  NAND4_X1 U4602 ( .A1(n3671), .A2(n3670), .A3(n3669), .A4(n3668), .ZN(n3677)
         );
  AOI22_X1 U4603 ( .A1(n4072), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3675) );
  AOI22_X1 U4604 ( .A1(n3984), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3072), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3674) );
  AOI22_X1 U4605 ( .A1(n3978), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3673) );
  AOI22_X1 U4606 ( .A1(n4036), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3672) );
  NAND4_X1 U4607 ( .A1(n3675), .A2(n3674), .A3(n3673), .A4(n3672), .ZN(n3676)
         );
  OR2_X1 U4608 ( .A1(n3677), .A2(n3676), .ZN(n3678) );
  AOI22_X1 U4609 ( .A1(n3842), .A2(n3678), .B1(n4953), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3680) );
  NAND2_X1 U4610 ( .A1(n3575), .A2(EAX_REG_10__SCAN_IN), .ZN(n3679) );
  OAI211_X1 U4611 ( .C1(n5674), .C2(n4052), .A(n3680), .B(n3679), .ZN(n4859)
         );
  AND2_X2 U4612 ( .A1(n4860), .A2(n4859), .ZN(n4858) );
  AOI22_X1 U4613 ( .A1(n3984), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4614 ( .A1(n4036), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4615 ( .A1(n4058), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4616 ( .A1(n4068), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4059), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3681) );
  NAND4_X1 U4617 ( .A1(n3684), .A2(n3683), .A3(n3682), .A4(n3681), .ZN(n3690)
         );
  AOI22_X1 U4618 ( .A1(n4070), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4619 ( .A1(n4072), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3072), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4620 ( .A1(n4057), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4621 ( .A1(n3979), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3685) );
  NAND4_X1 U4622 ( .A1(n3688), .A2(n3687), .A3(n3686), .A4(n3685), .ZN(n3689)
         );
  NOR2_X1 U4623 ( .A1(n3690), .A2(n3689), .ZN(n3695) );
  INV_X1 U4624 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3692) );
  XNOR2_X1 U4625 ( .A(n3696), .B(n3692), .ZN(n5260) );
  NAND2_X1 U4626 ( .A1(n5260), .A2(n4025), .ZN(n3694) );
  AOI22_X1 U4627 ( .A1(n4954), .A2(EAX_REG_11__SCAN_IN), .B1(n4953), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3693) );
  OAI211_X1 U4628 ( .C1(n3695), .C2(n3828), .A(n3694), .B(n3693), .ZN(n4873)
         );
  AND2_X2 U4629 ( .A1(n4858), .A2(n4873), .ZN(n4890) );
  XOR2_X1 U4630 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3713), .Z(n5898) );
  NAND2_X1 U4631 ( .A1(n5898), .A2(n4025), .ZN(n3699) );
  INV_X1 U4632 ( .A(EAX_REG_12__SCAN_IN), .ZN(n4893) );
  OAI21_X1 U4633 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6224), .A(n6367), 
        .ZN(n3697) );
  OAI21_X1 U4634 ( .B1(n3847), .B2(n4893), .A(n3697), .ZN(n3698) );
  NAND2_X1 U4635 ( .A1(n3699), .A2(n3698), .ZN(n3712) );
  AOI22_X1 U4636 ( .A1(n3072), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4637 ( .A1(n4070), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4638 ( .A1(n3700), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4639 ( .A1(n4036), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3701) );
  NAND4_X1 U4640 ( .A1(n3704), .A2(n3703), .A3(n3702), .A4(n3701), .ZN(n3710)
         );
  AOI22_X1 U4641 ( .A1(n4072), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3708) );
  AOI22_X1 U4642 ( .A1(n3984), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3707) );
  AOI22_X1 U4643 ( .A1(n3852), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4059), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4644 ( .A1(n3978), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3705) );
  NAND4_X1 U4645 ( .A1(n3708), .A2(n3707), .A3(n3706), .A4(n3705), .ZN(n3709)
         );
  OAI21_X1 U4646 ( .B1(n3710), .B2(n3709), .A(n3842), .ZN(n3711) );
  NAND2_X1 U4647 ( .A1(n3712), .A2(n3711), .ZN(n4889) );
  XNOR2_X1 U4649 ( .A(n3744), .B(n5247), .ZN(n5041) );
  NAND2_X1 U4650 ( .A1(n5041), .A2(n4025), .ZN(n3716) );
  INV_X1 U4651 ( .A(n4953), .ZN(n3809) );
  NOR2_X1 U4652 ( .A1(n3809), .A2(n5247), .ZN(n3714) );
  AOI21_X1 U4653 ( .B1(n3575), .B2(EAX_REG_13__SCAN_IN), .A(n3714), .ZN(n3715)
         );
  NAND2_X1 U4654 ( .A1(n3716), .A2(n3715), .ZN(n3728) );
  AOI22_X1 U4655 ( .A1(n3984), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3072), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4656 ( .A1(n4072), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3979), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4657 ( .A1(n4036), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4658 ( .A1(n4060), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3717) );
  NAND4_X1 U4659 ( .A1(n3720), .A2(n3719), .A3(n3718), .A4(n3717), .ZN(n3726)
         );
  AOI22_X1 U4660 ( .A1(n4070), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4661 ( .A1(n4057), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4662 ( .A1(n4062), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4059), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4663 ( .A1(n4058), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3721) );
  NAND4_X1 U4664 ( .A1(n3724), .A2(n3723), .A3(n3722), .A4(n3721), .ZN(n3725)
         );
  OR2_X1 U4665 ( .A1(n3726), .A2(n3725), .ZN(n3727) );
  AND2_X1 U4666 ( .A1(n3842), .A2(n3727), .ZN(n5037) );
  NAND2_X1 U4667 ( .A1(n5038), .A2(n5037), .ZN(n5036) );
  INV_X1 U4668 ( .A(n3728), .ZN(n3729) );
  NAND2_X1 U4669 ( .A1(n5036), .A2(n5115), .ZN(n4996) );
  AOI22_X1 U4670 ( .A1(n4072), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4671 ( .A1(n4060), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3177), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3732) );
  AOI22_X1 U4672 ( .A1(n3984), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4673 ( .A1(n4062), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3730) );
  NAND4_X1 U4674 ( .A1(n3733), .A2(n3732), .A3(n3731), .A4(n3730), .ZN(n3741)
         );
  AOI22_X1 U4675 ( .A1(n3072), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4676 ( .A1(n4070), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4677 ( .A1(n3852), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3737) );
  NAND2_X1 U4678 ( .A1(n4036), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3735) );
  AOI21_X1 U4679 ( .B1(n4071), .B2(INSTQUEUE_REG_9__4__SCAN_IN), .A(n4207), 
        .ZN(n3734) );
  AND2_X1 U4680 ( .A1(n3735), .A2(n3734), .ZN(n3736) );
  NAND4_X1 U4681 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3740)
         );
  NAND2_X1 U4682 ( .A1(n4046), .A2(n4052), .ZN(n3886) );
  OAI21_X1 U4683 ( .B1(n3741), .B2(n3740), .A(n3886), .ZN(n3743) );
  AOI22_X1 U4684 ( .A1(n4954), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6367), .ZN(n3742) );
  NAND2_X1 U4685 ( .A1(n3743), .A2(n3742), .ZN(n3747) );
  INV_X1 U4686 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3745) );
  XNOR2_X1 U4687 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n3866), .ZN(n5210)
         );
  NAND2_X1 U4688 ( .A1(n4207), .A2(n5210), .ZN(n3746) );
  NAND2_X1 U4689 ( .A1(n3747), .A2(n3746), .ZN(n4999) );
  INV_X1 U4690 ( .A(n4999), .ZN(n3850) );
  OR2_X1 U4691 ( .A1(n3748), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3749)
         );
  NAND2_X1 U4692 ( .A1(n3749), .A2(n3866), .ZN(n5537) );
  AOI22_X1 U4693 ( .A1(n3072), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4694 ( .A1(n3978), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4695 ( .A1(n4072), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4696 ( .A1(n4036), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3750) );
  NAND4_X1 U4697 ( .A1(n3753), .A2(n3752), .A3(n3751), .A4(n3750), .ZN(n3759)
         );
  AOI22_X1 U4698 ( .A1(n4070), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4699 ( .A1(n4058), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4700 ( .A1(n3984), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3177), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4701 ( .A1(n4060), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3754) );
  NAND4_X1 U4702 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3758)
         );
  NOR2_X1 U4703 ( .A1(n3759), .A2(n3758), .ZN(n3762) );
  OAI21_X1 U4704 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6224), .A(n6367), 
        .ZN(n3761) );
  NAND2_X1 U4705 ( .A1(n4954), .A2(EAX_REG_19__SCAN_IN), .ZN(n3760) );
  OAI211_X1 U4706 ( .C1(n4046), .C2(n3762), .A(n3761), .B(n3760), .ZN(n3763)
         );
  OAI21_X1 U4707 ( .B1(n5537), .B2(n4052), .A(n3763), .ZN(n5095) );
  INV_X1 U4708 ( .A(n5095), .ZN(n3849) );
  AOI22_X1 U4709 ( .A1(n3072), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4710 ( .A1(n4036), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4711 ( .A1(n4062), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4712 ( .A1(n4060), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3177), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3764) );
  NAND4_X1 U4713 ( .A1(n3767), .A2(n3766), .A3(n3765), .A4(n3764), .ZN(n3775)
         );
  AOI22_X1 U4714 ( .A1(n4072), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4715 ( .A1(n4070), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4716 ( .A1(n3852), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3771) );
  AOI21_X1 U4717 ( .B1(n4071), .B2(INSTQUEUE_REG_9__2__SCAN_IN), .A(n4207), 
        .ZN(n3769) );
  NAND2_X1 U4718 ( .A1(n4069), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3768)
         );
  AND2_X1 U4719 ( .A1(n3769), .A2(n3768), .ZN(n3770) );
  NAND4_X1 U4720 ( .A1(n3773), .A2(n3772), .A3(n3771), .A4(n3770), .ZN(n3774)
         );
  OAI21_X1 U4721 ( .B1(n3775), .B2(n3774), .A(n3886), .ZN(n3777) );
  AOI22_X1 U4722 ( .A1(n4954), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6367), .ZN(n3776) );
  NAND2_X1 U4723 ( .A1(n3777), .A2(n3776), .ZN(n3779) );
  XNOR2_X1 U4724 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3793), .ZN(n5219)
         );
  NAND2_X1 U4725 ( .A1(n4207), .A2(n5219), .ZN(n3778) );
  AOI22_X1 U4726 ( .A1(n4060), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4727 ( .A1(n3984), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3072), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4728 ( .A1(n3978), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3979), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4729 ( .A1(n4057), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3780) );
  NAND4_X1 U4730 ( .A1(n3783), .A2(n3782), .A3(n3781), .A4(n3780), .ZN(n3789)
         );
  AOI22_X1 U4731 ( .A1(n4072), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4732 ( .A1(n4036), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4733 ( .A1(n4059), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4734 ( .A1(n4070), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3784) );
  NAND4_X1 U4735 ( .A1(n3787), .A2(n3786), .A3(n3785), .A4(n3784), .ZN(n3788)
         );
  NOR2_X1 U4736 ( .A1(n3789), .A2(n3788), .ZN(n3790) );
  OR2_X1 U4737 ( .A1(n4046), .A2(n3790), .ZN(n3797) );
  NAND2_X1 U4738 ( .A1(n6367), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3791)
         );
  NAND2_X1 U4739 ( .A1(n4052), .A2(n3791), .ZN(n3792) );
  AOI21_X1 U4740 ( .B1(n3575), .B2(EAX_REG_17__SCAN_IN), .A(n3792), .ZN(n3796)
         );
  OAI21_X1 U4741 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3794), .A(n3793), 
        .ZN(n5633) );
  NOR2_X1 U4742 ( .A1(n5633), .A2(n4052), .ZN(n3795) );
  AOI21_X1 U4743 ( .B1(n3797), .B2(n3796), .A(n3795), .ZN(n5542) );
  XNOR2_X1 U4744 ( .A(n3798), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5640)
         );
  AOI22_X1 U4745 ( .A1(n4072), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4746 ( .A1(n4070), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4747 ( .A1(n4057), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4748 ( .A1(n4069), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3799) );
  NAND4_X1 U4749 ( .A1(n3802), .A2(n3801), .A3(n3800), .A4(n3799), .ZN(n3808)
         );
  AOI22_X1 U4750 ( .A1(n4060), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4751 ( .A1(n3984), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3072), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4752 ( .A1(n3852), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4753 ( .A1(n4036), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3177), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3803) );
  NAND4_X1 U4754 ( .A1(n3806), .A2(n3805), .A3(n3804), .A4(n3803), .ZN(n3807)
         );
  NOR2_X1 U4755 ( .A1(n3808), .A2(n3807), .ZN(n3812) );
  INV_X1 U4756 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5638) );
  NOR2_X1 U4757 ( .A1(n3809), .A2(n5638), .ZN(n3810) );
  AOI21_X1 U4758 ( .B1(n3575), .B2(EAX_REG_16__SCAN_IN), .A(n3810), .ZN(n3811)
         );
  OAI21_X1 U4759 ( .B1(n4046), .B2(n3812), .A(n3811), .ZN(n3813) );
  AOI21_X1 U4760 ( .B1(n5640), .B2(n4025), .A(n3813), .ZN(n5107) );
  XNOR2_X1 U4761 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3814), .ZN(n5234)
         );
  INV_X1 U4762 ( .A(n5234), .ZN(n3830) );
  AOI22_X1 U4763 ( .A1(n4072), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4764 ( .A1(n3072), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4765 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n3978), .B1(n4062), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4766 ( .A1(n3852), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3815) );
  NAND4_X1 U4767 ( .A1(n3818), .A2(n3817), .A3(n3816), .A4(n3815), .ZN(n3824)
         );
  AOI22_X1 U4768 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n4060), .B1(n3984), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4769 ( .A1(n4070), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4770 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n4036), .B1(n4069), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4771 ( .A1(n4059), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3819) );
  NAND4_X1 U4772 ( .A1(n3822), .A2(n3821), .A3(n3820), .A4(n3819), .ZN(n3823)
         );
  NOR2_X1 U4773 ( .A1(n3824), .A2(n3823), .ZN(n3827) );
  NAND2_X1 U4774 ( .A1(n3575), .A2(EAX_REG_15__SCAN_IN), .ZN(n3826) );
  NAND2_X1 U4775 ( .A1(n4953), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3825)
         );
  OAI211_X1 U4776 ( .C1(n3828), .C2(n3827), .A(n3826), .B(n3825), .ZN(n3829)
         );
  AOI21_X1 U4777 ( .B1(n3830), .B2(n4025), .A(n3829), .ZN(n5106) );
  NOR2_X1 U4778 ( .A1(n5107), .A2(n5106), .ZN(n3848) );
  INV_X1 U4779 ( .A(EAX_REG_14__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4780 ( .A1(n4060), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4781 ( .A1(n3984), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3072), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4782 ( .A1(n4070), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4783 ( .A1(n3852), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3831) );
  NAND4_X1 U4784 ( .A1(n3834), .A2(n3833), .A3(n3832), .A4(n3831), .ZN(n3840)
         );
  AOI22_X1 U4785 ( .A1(n4072), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4786 ( .A1(n3978), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4787 ( .A1(n4059), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4788 ( .A1(n4036), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3835) );
  NAND4_X1 U4789 ( .A1(n3838), .A2(n3837), .A3(n3836), .A4(n3835), .ZN(n3839)
         );
  OR2_X1 U4790 ( .A1(n3840), .A2(n3839), .ZN(n3841) );
  NAND2_X1 U4791 ( .A1(n3842), .A2(n3841), .ZN(n3845) );
  XNOR2_X1 U4792 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3843), .ZN(n5652)
         );
  AOI22_X1 U4793 ( .A1(n4207), .A2(n5652), .B1(n4953), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3844) );
  OAI211_X1 U4794 ( .C1(n3847), .C2(n3846), .A(n3845), .B(n3844), .ZN(n5114)
         );
  AND2_X1 U4795 ( .A1(n3848), .A2(n5114), .ZN(n5105) );
  AND2_X1 U4796 ( .A1(n5542), .A2(n5105), .ZN(n5011) );
  AND2_X2 U4797 ( .A1(n4996), .A2(n3851), .ZN(n5089) );
  AOI22_X1 U4798 ( .A1(n4067), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3072), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4799 ( .A1(n4062), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4800 ( .A1(n4058), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3177), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4801 ( .A1(n3852), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3853) );
  NAND4_X1 U4802 ( .A1(n3856), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(n3862)
         );
  AOI22_X1 U4803 ( .A1(n4072), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4804 ( .A1(n4070), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4805 ( .A1(n4036), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4806 ( .A1(n4060), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3857) );
  NAND4_X1 U4807 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3861)
         );
  NOR2_X1 U4808 ( .A1(n3862), .A2(n3861), .ZN(n3863) );
  OR2_X1 U4809 ( .A1(n4046), .A2(n3863), .ZN(n3871) );
  NAND2_X1 U4810 ( .A1(n6367), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3864)
         );
  NAND2_X1 U4811 ( .A1(n4052), .A2(n3864), .ZN(n3865) );
  AOI21_X1 U4812 ( .B1(n3575), .B2(EAX_REG_21__SCAN_IN), .A(n3865), .ZN(n3870)
         );
  OAI21_X1 U4813 ( .B1(n3868), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n3915), 
        .ZN(n5491) );
  NOR2_X1 U4814 ( .A1(n5491), .A2(n4052), .ZN(n3869) );
  AOI21_X1 U4815 ( .B1(n3871), .B2(n3870), .A(n3869), .ZN(n5088) );
  AND2_X2 U4816 ( .A1(n5089), .A2(n5088), .ZN(n5085) );
  AOI22_X1 U4817 ( .A1(n4072), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4818 ( .A1(n3984), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4819 ( .A1(n4036), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3875) );
  AOI21_X1 U4820 ( .B1(n4071), .B2(INSTQUEUE_REG_9__6__SCAN_IN), .A(n4025), 
        .ZN(n3873) );
  NAND2_X1 U4821 ( .A1(n3195), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3872)
         );
  AND2_X1 U4822 ( .A1(n3873), .A2(n3872), .ZN(n3874) );
  NAND4_X1 U4823 ( .A1(n3877), .A2(n3876), .A3(n3875), .A4(n3874), .ZN(n3884)
         );
  AOI22_X1 U4824 ( .A1(n4060), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4825 ( .A1(n3072), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4826 ( .A1(n4070), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4827 ( .A1(n4058), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4059), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3879) );
  NAND4_X1 U4828 ( .A1(n3882), .A2(n3881), .A3(n3880), .A4(n3879), .ZN(n3883)
         );
  OR2_X1 U4829 ( .A1(n3884), .A2(n3883), .ZN(n3885) );
  NAND2_X1 U4830 ( .A1(n3886), .A2(n3885), .ZN(n3889) );
  AOI22_X1 U4831 ( .A1(n4954), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6367), .ZN(n3888) );
  XNOR2_X1 U4832 ( .A(n3915), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5483)
         );
  AND2_X1 U4833 ( .A1(n5483), .A2(n4207), .ZN(n3887) );
  AOI21_X1 U4834 ( .B1(n3889), .B2(n3888), .A(n3887), .ZN(n5086) );
  NAND2_X1 U4835 ( .A1(n5085), .A2(n5086), .ZN(n4261) );
  INV_X1 U4836 ( .A(n4261), .ZN(n3920) );
  AOI22_X1 U4837 ( .A1(n3072), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4838 ( .A1(n3984), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4839 ( .A1(n4060), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4840 ( .A1(n4036), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3890) );
  NAND4_X1 U4841 ( .A1(n3893), .A2(n3892), .A3(n3891), .A4(n3890), .ZN(n3900)
         );
  AOI22_X1 U4842 ( .A1(n3894), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4843 ( .A1(n4057), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4844 ( .A1(n4009), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4059), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4845 ( .A1(n4062), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3895) );
  NAND4_X1 U4846 ( .A1(n3898), .A2(n3897), .A3(n3896), .A4(n3895), .ZN(n3899)
         );
  NOR2_X1 U4847 ( .A1(n3900), .A2(n3899), .ZN(n3921) );
  AOI22_X1 U4848 ( .A1(n3072), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4849 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n4057), .B1(n4062), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4850 ( .A1(n4060), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4851 ( .A1(n4070), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3901) );
  NAND4_X1 U4852 ( .A1(n3904), .A2(n3903), .A3(n3902), .A4(n3901), .ZN(n3910)
         );
  AOI22_X1 U4853 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(n3978), .B1(n3852), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4854 ( .A1(n4009), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4059), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4855 ( .A1(n3087), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4856 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n4036), .B1(n4069), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3905) );
  NAND4_X1 U4857 ( .A1(n3908), .A2(n3907), .A3(n3906), .A4(n3905), .ZN(n3909)
         );
  NOR2_X1 U4858 ( .A1(n3910), .A2(n3909), .ZN(n3922) );
  XNOR2_X1 U4859 ( .A(n3921), .B(n3922), .ZN(n3914) );
  NAND2_X1 U4860 ( .A1(n6367), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3911)
         );
  NAND2_X1 U4861 ( .A1(n4052), .A2(n3911), .ZN(n3912) );
  AOI21_X1 U4862 ( .B1(n3575), .B2(EAX_REG_23__SCAN_IN), .A(n3912), .ZN(n3913)
         );
  OAI21_X1 U4863 ( .B1(n4046), .B2(n3914), .A(n3913), .ZN(n3919) );
  INV_X1 U4864 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5477) );
  OR2_X1 U4865 ( .A1(n3916), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3917)
         );
  NAND2_X1 U4866 ( .A1(n3955), .A2(n3917), .ZN(n5476) );
  NAND2_X1 U4867 ( .A1(n3920), .A2(n3077), .ZN(n4263) );
  NOR2_X1 U4868 ( .A1(n3922), .A2(n3921), .ZN(n3939) );
  AOI22_X1 U4869 ( .A1(n4009), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4870 ( .A1(n3072), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4871 ( .A1(n4067), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4872 ( .A1(n4059), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3923) );
  NAND4_X1 U4873 ( .A1(n3926), .A2(n3925), .A3(n3924), .A4(n3923), .ZN(n3932)
         );
  AOI22_X1 U4874 ( .A1(n4070), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4875 ( .A1(n4062), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4876 ( .A1(n4036), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4877 ( .A1(n3978), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3927) );
  NAND4_X1 U4878 ( .A1(n3930), .A2(n3929), .A3(n3928), .A4(n3927), .ZN(n3931)
         );
  OR2_X1 U4879 ( .A1(n3932), .A2(n3931), .ZN(n3938) );
  INV_X1 U4880 ( .A(n3938), .ZN(n3933) );
  XNOR2_X1 U4881 ( .A(n3939), .B(n3933), .ZN(n3937) );
  INV_X1 U4882 ( .A(n4046), .ZN(n4081) );
  XNOR2_X1 U4883 ( .A(n3955), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5463)
         );
  NAND2_X1 U4884 ( .A1(n4954), .A2(EAX_REG_24__SCAN_IN), .ZN(n3935) );
  NAND2_X1 U4885 ( .A1(n4953), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3934)
         );
  OAI211_X1 U4886 ( .C1(n5463), .C2(n4052), .A(n3935), .B(n3934), .ZN(n3936)
         );
  AOI21_X1 U4887 ( .B1(n3937), .B2(n4081), .A(n3936), .ZN(n5078) );
  NAND2_X1 U4888 ( .A1(n3939), .A2(n3938), .ZN(n3960) );
  AOI22_X1 U4889 ( .A1(n4070), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4890 ( .A1(n4036), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4891 ( .A1(n3072), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4892 ( .A1(n4058), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4059), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3940) );
  NAND4_X1 U4893 ( .A1(n3943), .A2(n3942), .A3(n3941), .A4(n3940), .ZN(n3949)
         );
  AOI22_X1 U4894 ( .A1(n4009), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4895 ( .A1(n4057), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4896 ( .A1(n4060), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4897 ( .A1(n4069), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3944) );
  NAND4_X1 U4898 ( .A1(n3947), .A2(n3946), .A3(n3945), .A4(n3944), .ZN(n3948)
         );
  NOR2_X1 U4899 ( .A1(n3949), .A2(n3948), .ZN(n3961) );
  XNOR2_X1 U4900 ( .A(n3960), .B(n3961), .ZN(n3953) );
  INV_X1 U4901 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3950) );
  OAI21_X1 U4902 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n3950), .A(n4052), .ZN(
        n3951) );
  AOI21_X1 U4903 ( .B1(n3575), .B2(EAX_REG_25__SCAN_IN), .A(n3951), .ZN(n3952)
         );
  OAI21_X1 U4904 ( .B1(n3953), .B2(n4046), .A(n3952), .ZN(n3959) );
  INV_X1 U4905 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3954) );
  OR2_X1 U4906 ( .A1(n3956), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3957)
         );
  NAND2_X1 U4907 ( .A1(n3957), .A2(n3997), .ZN(n5531) );
  NOR2_X1 U4908 ( .A1(n3961), .A2(n3960), .ZN(n3992) );
  AOI22_X1 U4909 ( .A1(n4009), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4910 ( .A1(n3072), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4911 ( .A1(n3984), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4912 ( .A1(n4059), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3962) );
  NAND4_X1 U4913 ( .A1(n3965), .A2(n3964), .A3(n3963), .A4(n3962), .ZN(n3971)
         );
  AOI22_X1 U4914 ( .A1(n4070), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U4915 ( .A1(n4062), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4916 ( .A1(n4036), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4917 ( .A1(n3978), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3966) );
  NAND4_X1 U4918 ( .A1(n3969), .A2(n3968), .A3(n3967), .A4(n3966), .ZN(n3970)
         );
  OR2_X1 U4919 ( .A1(n3971), .A2(n3970), .ZN(n3991) );
  INV_X1 U4920 ( .A(n3991), .ZN(n3972) );
  XNOR2_X1 U4921 ( .A(n3992), .B(n3972), .ZN(n3973) );
  NAND2_X1 U4922 ( .A1(n3973), .A2(n4081), .ZN(n3977) );
  INV_X1 U4923 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5179) );
  AOI21_X1 U4924 ( .B1(n5179), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3974) );
  AOI21_X1 U4925 ( .B1(n3575), .B2(EAX_REG_26__SCAN_IN), .A(n3974), .ZN(n3976)
         );
  XNOR2_X1 U4926 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .B(n3997), .ZN(n5447)
         );
  AOI21_X1 U4927 ( .B1(n3977), .B2(n3976), .A(n3975), .ZN(n5064) );
  NAND2_X1 U4928 ( .A1(n5063), .A2(n5064), .ZN(n5055) );
  INV_X1 U4929 ( .A(n5055), .ZN(n4006) );
  AOI22_X1 U4930 ( .A1(n4070), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4931 ( .A1(n4058), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4059), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4932 ( .A1(n3072), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4933 ( .A1(n3979), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3980) );
  NAND4_X1 U4934 ( .A1(n3983), .A2(n3982), .A3(n3981), .A4(n3980), .ZN(n3990)
         );
  AOI22_X1 U4935 ( .A1(n4009), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U4936 ( .A1(n4057), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U4937 ( .A1(n4060), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U4938 ( .A1(n4036), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3985) );
  NAND4_X1 U4939 ( .A1(n3988), .A2(n3987), .A3(n3986), .A4(n3985), .ZN(n3989)
         );
  NOR2_X1 U4940 ( .A1(n3990), .A2(n3989), .ZN(n4008) );
  NAND2_X1 U4941 ( .A1(n3992), .A2(n3991), .ZN(n4007) );
  XNOR2_X1 U4942 ( .A(n4008), .B(n4007), .ZN(n3996) );
  NAND2_X1 U4943 ( .A1(n6367), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3993)
         );
  NAND2_X1 U4944 ( .A1(n4052), .A2(n3993), .ZN(n3994) );
  AOI21_X1 U4945 ( .B1(n3575), .B2(EAX_REG_27__SCAN_IN), .A(n3994), .ZN(n3995)
         );
  OAI21_X1 U4946 ( .B1(n3996), .B2(n4046), .A(n3995), .ZN(n4004) );
  INV_X1 U4947 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4001) );
  INV_X1 U4948 ( .A(n3999), .ZN(n4000) );
  NAND2_X1 U4949 ( .A1(n4001), .A2(n4000), .ZN(n4002) );
  NAND2_X1 U4950 ( .A1(n4023), .A2(n4002), .ZN(n5442) );
  NAND2_X1 U4951 ( .A1(n4004), .A2(n4003), .ZN(n5056) );
  NAND2_X1 U4952 ( .A1(n4006), .A2(n4005), .ZN(n4985) );
  NOR2_X1 U4953 ( .A1(n4008), .A2(n4007), .ZN(n4031) );
  AOI22_X1 U4954 ( .A1(n4009), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4955 ( .A1(n3072), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4956 ( .A1(n3984), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4957 ( .A1(n4059), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4010) );
  NAND4_X1 U4958 ( .A1(n4013), .A2(n4012), .A3(n4011), .A4(n4010), .ZN(n4019)
         );
  AOI22_X1 U4959 ( .A1(n4070), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3852), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4960 ( .A1(n4062), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U4961 ( .A1(n4036), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U4962 ( .A1(n3978), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4014) );
  NAND4_X1 U4963 ( .A1(n4017), .A2(n4016), .A3(n4015), .A4(n4014), .ZN(n4018)
         );
  OR2_X1 U4964 ( .A1(n4019), .A2(n4018), .ZN(n4030) );
  XNOR2_X1 U4965 ( .A(n4031), .B(n4030), .ZN(n4022) );
  INV_X1 U4966 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6650) );
  OAI21_X1 U4967 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6650), .A(n4052), .ZN(
        n4020) );
  AOI21_X1 U4968 ( .B1(n3575), .B2(EAX_REG_28__SCAN_IN), .A(n4020), .ZN(n4021)
         );
  OAI21_X1 U4969 ( .B1(n4022), .B2(n4046), .A(n4021), .ZN(n4027) );
  INV_X1 U4970 ( .A(n4048), .ZN(n4050) );
  NAND2_X1 U4971 ( .A1(n4023), .A2(n6650), .ZN(n4024) );
  NAND2_X1 U4972 ( .A1(n5164), .A2(n4025), .ZN(n4026) );
  NAND2_X1 U4973 ( .A1(n4027), .A2(n4026), .ZN(n4988) );
  NAND2_X1 U4974 ( .A1(n4031), .A2(n4030), .ZN(n4055) );
  AOI22_X1 U4975 ( .A1(n4062), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U4976 ( .A1(n4070), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U4977 ( .A1(n3087), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U4978 ( .A1(n3182), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4032) );
  NAND4_X1 U4979 ( .A1(n4035), .A2(n4034), .A3(n4033), .A4(n4032), .ZN(n4042)
         );
  AOI22_X1 U4980 ( .A1(n4072), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U4981 ( .A1(n3072), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U4982 ( .A1(n4036), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3979), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U4983 ( .A1(n4060), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4059), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4037) );
  NAND4_X1 U4984 ( .A1(n4040), .A2(n4039), .A3(n4038), .A4(n4037), .ZN(n4041)
         );
  NOR2_X1 U4985 ( .A1(n4042), .A2(n4041), .ZN(n4056) );
  XNOR2_X1 U4986 ( .A(n4055), .B(n4056), .ZN(n4047) );
  NAND2_X1 U4987 ( .A1(n6367), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4043)
         );
  NAND2_X1 U4988 ( .A1(n4052), .A2(n4043), .ZN(n4044) );
  AOI21_X1 U4989 ( .B1(n3575), .B2(EAX_REG_29__SCAN_IN), .A(n4044), .ZN(n4045)
         );
  OAI21_X1 U4990 ( .B1(n4047), .B2(n4046), .A(n4045), .ZN(n4054) );
  NAND2_X1 U4991 ( .A1(n4048), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4212)
         );
  INV_X1 U4992 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4049) );
  NAND2_X1 U4993 ( .A1(n4050), .A2(n4049), .ZN(n4051) );
  NAND2_X1 U4994 ( .A1(n4212), .A2(n4051), .ZN(n5155) );
  NAND2_X1 U4995 ( .A1(n4054), .A2(n4053), .ZN(n4196) );
  NOR2_X1 U4996 ( .A1(n4056), .A2(n4055), .ZN(n4080) );
  AOI22_X1 U4997 ( .A1(n4058), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U4998 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4036), .B1(n3979), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U4999 ( .A1(n4060), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4059), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5000 ( .A1(n4062), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4061), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4063) );
  NAND4_X1 U5001 ( .A1(n4066), .A2(n4065), .A3(n4064), .A4(n4063), .ZN(n4078)
         );
  AOI22_X1 U5002 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n3984), .B1(n3072), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5003 ( .A1(n3182), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4075) );
  AOI22_X1 U5004 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n4070), .B1(n4069), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4074) );
  AOI22_X1 U5005 ( .A1(n4072), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4073) );
  NAND4_X1 U5006 ( .A1(n4076), .A2(n4075), .A3(n4074), .A4(n4073), .ZN(n4077)
         );
  NOR2_X1 U5007 ( .A1(n4078), .A2(n4077), .ZN(n4079) );
  XNOR2_X1 U5008 ( .A(n4080), .B(n4079), .ZN(n4082) );
  NAND2_X1 U5009 ( .A1(n4082), .A2(n4081), .ZN(n4085) );
  INV_X1 U5010 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4211) );
  NOR2_X1 U5011 ( .A1(n4211), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4083) );
  AOI211_X1 U5012 ( .C1(n3575), .C2(EAX_REG_30__SCAN_IN), .A(n4083), .B(n4207), 
        .ZN(n4084) );
  XNOR2_X1 U5013 ( .A(n4212), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4964)
         );
  AOI22_X1 U5014 ( .A1(n4085), .A2(n4084), .B1(n4964), .B2(n4207), .ZN(n4951)
         );
  AND2_X1 U5015 ( .A1(n6368), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4208) );
  NAND2_X1 U5016 ( .A1(n4208), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6383) );
  NOR2_X1 U5017 ( .A1(n4096), .A2(n6275), .ZN(n4094) );
  NAND2_X1 U5018 ( .A1(n6271), .A2(n4086), .ZN(n6482) );
  AND2_X1 U5019 ( .A1(n6482), .A2(n6368), .ZN(n4087) );
  NAND2_X1 U5020 ( .A1(n6368), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4089) );
  NAND2_X1 U5021 ( .A1(n6224), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4088) );
  NAND2_X1 U5022 ( .A1(n4089), .A2(n4088), .ZN(n5918) );
  NAND2_X1 U5023 ( .A1(n5897), .A2(n4964), .ZN(n4092) );
  NOR2_X1 U5024 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6385) );
  AND2_X2 U5025 ( .A1(n5597), .A2(n6385), .ZN(n5917) );
  NAND2_X1 U5026 ( .A1(n5917), .A2(REIP_REG_30__SCAN_IN), .ZN(n5280) );
  OAI21_X1 U5027 ( .B1(n5553), .B2(n4211), .A(n5280), .ZN(n4090) );
  INV_X1 U5028 ( .A(n4090), .ZN(n4091) );
  NAND2_X1 U5029 ( .A1(n4097), .A2(n3249), .ZN(n4099) );
  MUX2_X1 U5030 ( .A(n4099), .B(n6485), .S(n4098), .Z(n4294) );
  NOR2_X1 U5031 ( .A1(n4550), .A2(n3249), .ZN(n4735) );
  NAND2_X1 U5032 ( .A1(n4735), .A2(n4101), .ZN(n4415) );
  NAND2_X1 U5033 ( .A1(n4415), .A2(n4303), .ZN(n4103) );
  NOR2_X1 U5034 ( .A1(n4429), .A2(n4103), .ZN(n4104) );
  NAND2_X1 U5035 ( .A1(n4282), .A2(n4104), .ZN(n4456) );
  INV_X1 U5036 ( .A(n3574), .ZN(n5127) );
  AND3_X1 U5037 ( .A1(n5127), .A2(n3306), .A3(n3573), .ZN(n4382) );
  NAND3_X1 U5038 ( .A1(n4223), .A2(n4105), .A3(n4382), .ZN(n4106) );
  OAI21_X1 U5039 ( .B1(n4418), .B2(n4456), .A(n4106), .ZN(n4107) );
  NAND2_X2 U5040 ( .A1(n5776), .A2(n3574), .ZN(n5126) );
  INV_X1 U5041 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4736) );
  NAND2_X1 U5042 ( .A1(n4108), .A2(n4736), .ZN(n4111) );
  NAND2_X1 U5043 ( .A1(n4123), .A2(n4109), .ZN(n4110) );
  NAND3_X1 U5044 ( .A1(n4117), .A2(n4111), .A3(n4110), .ZN(n4114) );
  INV_X1 U5045 ( .A(n4111), .ZN(n4112) );
  NAND2_X1 U5046 ( .A1(n4112), .A2(n4120), .ZN(n4113) );
  INV_X1 U5047 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5760) );
  NOR2_X1 U5048 ( .A1(n4897), .A2(n4332), .ZN(n4333) );
  INV_X1 U5049 ( .A(n4115), .ZN(n4116) );
  AOI21_X1 U5050 ( .B1(n5017), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(n4119), 
        .ZN(n4118) );
  AOI22_X1 U5051 ( .A1(n5017), .A2(n4119), .B1(n4178), .B2(n4118), .ZN(n4560)
         );
  NAND2_X1 U5052 ( .A1(n4561), .A2(n4560), .ZN(n4478) );
  NOR2_X1 U5053 ( .A1(EBX_REG_3__SCAN_IN), .A2(n4897), .ZN(n4122) );
  INV_X1 U5054 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4505) );
  AOI21_X1 U5055 ( .B1(n4505), .B2(n4178), .A(n4122), .ZN(n4121) );
  OAI22_X1 U5056 ( .A1(n4122), .A2(n5017), .B1(n4291), .B2(n4121), .ZN(n4479)
         );
  INV_X1 U5057 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4401) );
  NAND2_X1 U5058 ( .A1(n4223), .A2(n4401), .ZN(n4125) );
  OAI211_X1 U5059 ( .C1(n4182), .C2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n5017), 
        .B(n4125), .ZN(n4124) );
  OAI21_X1 U5060 ( .B1(n5017), .B2(n4125), .A(n4124), .ZN(n4400) );
  INV_X1 U5061 ( .A(EBX_REG_5__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U5062 ( .A1(n4223), .A2(n5713), .ZN(n4127) );
  OAI211_X1 U5063 ( .C1(n4291), .C2(n4471), .A(n4178), .B(n4127), .ZN(n4126)
         );
  OAI21_X1 U5064 ( .B1(n4291), .B2(n4127), .A(n4126), .ZN(n4448) );
  INV_X1 U5065 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5775) );
  NAND2_X1 U5066 ( .A1(n4223), .A2(n5775), .ZN(n4129) );
  OAI211_X1 U5067 ( .C1(n4182), .C2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n5017), 
        .B(n4129), .ZN(n4128) );
  OAI21_X1 U5068 ( .B1(n5017), .B2(n4129), .A(n4128), .ZN(n4500) );
  NAND2_X1 U5069 ( .A1(n4447), .A2(n4500), .ZN(n4565) );
  NOR2_X1 U5070 ( .A1(EBX_REG_7__SCAN_IN), .A2(n4897), .ZN(n4131) );
  AOI21_X1 U5071 ( .B1(n5938), .B2(n4178), .A(n4131), .ZN(n4130) );
  OAI22_X1 U5072 ( .A1(n4131), .A2(n5017), .B1(n4291), .B2(n4130), .ZN(n4566)
         );
  NOR2_X1 U5073 ( .A1(EBX_REG_8__SCAN_IN), .A2(n4897), .ZN(n4133) );
  AOI21_X1 U5074 ( .B1(n5017), .B2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n4133), 
        .ZN(n4132) );
  AOI22_X1 U5075 ( .A1(n5017), .A2(n4133), .B1(n4178), .B2(n4132), .ZN(n4343)
         );
  NOR2_X1 U5076 ( .A1(EBX_REG_9__SCAN_IN), .A2(n4897), .ZN(n4135) );
  INV_X1 U5077 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4753) );
  AOI21_X1 U5078 ( .B1(n4753), .B2(n4178), .A(n4135), .ZN(n4134) );
  OAI22_X1 U5079 ( .A1(n4135), .A2(n5017), .B1(n4291), .B2(n4134), .ZN(n4756)
         );
  INV_X1 U5080 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4863) );
  NAND2_X1 U5081 ( .A1(n4223), .A2(n4863), .ZN(n4137) );
  OAI211_X1 U5082 ( .C1(n4182), .C2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5017), .B(n4137), .ZN(n4136) );
  OAI21_X1 U5083 ( .B1(n5017), .B2(n4137), .A(n4136), .ZN(n4862) );
  NOR2_X1 U5084 ( .A1(EBX_REG_11__SCAN_IN), .A2(n4897), .ZN(n4139) );
  AOI21_X1 U5085 ( .B1(n5387), .B2(n4178), .A(n4139), .ZN(n4138) );
  OAI22_X1 U5086 ( .A1(n4139), .A2(n5017), .B1(n4291), .B2(n4138), .ZN(n4877)
         );
  INV_X1 U5087 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U5088 ( .A1(n4223), .A2(n5661), .ZN(n4141) );
  OAI211_X1 U5089 ( .C1(n4182), .C2(INSTADDRPOINTER_REG_12__SCAN_IN), .A(n5017), .B(n4141), .ZN(n4140) );
  OAI21_X1 U5090 ( .B1(n5017), .B2(n4141), .A(n4140), .ZN(n4891) );
  INV_X1 U5091 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U5092 ( .A1(n4223), .A2(n5125), .ZN(n4143) );
  OAI211_X1 U5093 ( .C1(n4291), .C2(n5373), .A(n4178), .B(n4143), .ZN(n4142)
         );
  OAI21_X1 U5094 ( .B1(n4291), .B2(n4143), .A(n4142), .ZN(n5043) );
  NOR2_X1 U5095 ( .A1(EBX_REG_14__SCAN_IN), .A2(n4897), .ZN(n4145) );
  AOI21_X1 U5096 ( .B1(n5017), .B2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n4145), 
        .ZN(n4144) );
  AOI22_X1 U5097 ( .A1(n5017), .A2(n4145), .B1(n4178), .B2(n4144), .ZN(n5120)
         );
  INV_X1 U5098 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6671) );
  NAND2_X1 U5099 ( .A1(n4223), .A2(n6671), .ZN(n4147) );
  INV_X1 U5100 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4305) );
  OAI211_X1 U5101 ( .C1(n4291), .C2(n4305), .A(n4178), .B(n4147), .ZN(n4146)
         );
  OAI21_X1 U5102 ( .B1(n4291), .B2(n4147), .A(n4146), .ZN(n5033) );
  NOR2_X1 U5103 ( .A1(EBX_REG_16__SCAN_IN), .A2(n4897), .ZN(n4149) );
  AOI21_X1 U5104 ( .B1(n5017), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n4149), 
        .ZN(n4148) );
  AOI22_X1 U5105 ( .A1(n5017), .A2(n4149), .B1(n4178), .B2(n4148), .ZN(n5110)
         );
  INV_X1 U5106 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U5107 ( .A1(n4223), .A2(n5770), .ZN(n4151) );
  INV_X1 U5108 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5564) );
  OAI211_X1 U5109 ( .C1(n4291), .C2(n5564), .A(n4178), .B(n4151), .ZN(n4150)
         );
  OAI21_X1 U5110 ( .B1(n4291), .B2(n4151), .A(n4150), .ZN(n5358) );
  NOR2_X1 U5111 ( .A1(EBX_REG_19__SCAN_IN), .A2(n4897), .ZN(n4153) );
  AOI21_X1 U5112 ( .B1(n5017), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n4153), 
        .ZN(n4152) );
  AOI22_X1 U5113 ( .A1(n5017), .A2(n4153), .B1(n4178), .B2(n4152), .ZN(n5100)
         );
  NAND2_X1 U5114 ( .A1(n5017), .A2(n4178), .ZN(n4896) );
  INV_X1 U5115 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6626) );
  NOR2_X1 U5116 ( .A1(EBX_REG_18__SCAN_IN), .A2(n4897), .ZN(n5018) );
  AOI21_X1 U5117 ( .B1(n4487), .B2(n6626), .A(n5018), .ZN(n4155) );
  OAI22_X1 U5118 ( .A1(EBX_REG_20__SCAN_IN), .A2(n4897), .B1(
        INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n4896), .ZN(n5004) );
  INV_X1 U5119 ( .A(n4155), .ZN(n5001) );
  NAND2_X1 U5120 ( .A1(n5017), .A2(n5001), .ZN(n5016) );
  INV_X1 U5121 ( .A(EBX_REG_20__SCAN_IN), .ZN(n4156) );
  NAND2_X1 U5122 ( .A1(EBX_REG_20__SCAN_IN), .A2(n4291), .ZN(n4157) );
  NAND2_X1 U5123 ( .A1(n4159), .A2(n4158), .ZN(n5091) );
  INV_X1 U5124 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U5125 ( .A1(n4223), .A2(n5496), .ZN(n4160) );
  OR2_X1 U5126 ( .A1(n4160), .A2(n4291), .ZN(n4162) );
  INV_X1 U5127 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5183) );
  OAI211_X1 U5128 ( .C1(n4291), .C2(n5183), .A(n4178), .B(n4160), .ZN(n4161)
         );
  NAND2_X1 U5129 ( .A1(n4162), .A2(n4161), .ZN(n5092) );
  INV_X1 U5130 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U5131 ( .A1(n4223), .A2(n5478), .ZN(n4164) );
  OR2_X1 U5132 ( .A1(n4164), .A2(n5017), .ZN(n4166) );
  OAI211_X1 U5133 ( .C1(n4182), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5017), .B(n4164), .ZN(n4165) );
  INV_X1 U5134 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U5135 ( .A1(n4223), .A2(n5506), .ZN(n4167) );
  OR2_X1 U5136 ( .A1(n4167), .A2(n4291), .ZN(n4169) );
  OAI211_X1 U5137 ( .C1(n4291), .C2(n5315), .A(n4178), .B(n4167), .ZN(n4168)
         );
  INV_X1 U5138 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U5139 ( .A1(n4223), .A2(n5460), .ZN(n4170) );
  OR2_X1 U5140 ( .A1(n4170), .A2(n5017), .ZN(n4172) );
  OAI211_X1 U5141 ( .C1(n4182), .C2(INSTADDRPOINTER_REG_24__SCAN_IN), .A(n5017), .B(n4170), .ZN(n4171) );
  NAND2_X1 U5142 ( .A1(n4172), .A2(n4171), .ZN(n5081) );
  NOR2_X1 U5143 ( .A1(EBX_REG_25__SCAN_IN), .A2(n4897), .ZN(n4174) );
  AOI21_X1 U5144 ( .B1(n5559), .B2(n4178), .A(n4174), .ZN(n4173) );
  OAI22_X1 U5145 ( .A1(n4174), .A2(n5017), .B1(n4291), .B2(n4173), .ZN(n5070)
         );
  INV_X1 U5146 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5068) );
  NAND2_X1 U5147 ( .A1(n4223), .A2(n5068), .ZN(n4176) );
  OAI211_X1 U5148 ( .C1(n4182), .C2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5017), .B(n4176), .ZN(n4175) );
  OAI21_X1 U5149 ( .B1(n5017), .B2(n4176), .A(n4175), .ZN(n4177) );
  INV_X1 U5150 ( .A(n4177), .ZN(n5065) );
  INV_X1 U5151 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5299) );
  INV_X1 U5152 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5062) );
  AND2_X1 U5153 ( .A1(n4223), .A2(n5062), .ZN(n4179) );
  AOI21_X1 U5154 ( .B1(n5299), .B2(n4178), .A(n4179), .ZN(n4180) );
  MUX2_X1 U5155 ( .A(n4180), .B(n4179), .S(n4291), .Z(n5059) );
  INV_X1 U5156 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5054) );
  NAND2_X1 U5157 ( .A1(n4223), .A2(n5054), .ZN(n4181) );
  OR2_X1 U5158 ( .A1(n4181), .A2(n5017), .ZN(n4184) );
  OAI211_X1 U5159 ( .C1(n4182), .C2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n4117), .B(n4181), .ZN(n4183) );
  NAND2_X1 U5160 ( .A1(n4184), .A2(n4183), .ZN(n4991) );
  INV_X1 U5161 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4938) );
  NAND2_X1 U5162 ( .A1(n4223), .A2(n4938), .ZN(n4220) );
  INV_X1 U5163 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4941) );
  NAND2_X1 U5164 ( .A1(n4941), .A2(n4487), .ZN(n4185) );
  NAND2_X1 U5165 ( .A1(n4220), .A2(n4185), .ZN(n4219) );
  NAND2_X1 U5166 ( .A1(n2997), .A2(n4117), .ZN(n4894) );
  INV_X1 U5167 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5281) );
  OR2_X1 U5168 ( .A1(n4223), .A2(n5281), .ZN(n4187) );
  NAND2_X1 U5169 ( .A1(EBX_REG_30__SCAN_IN), .A2(n4896), .ZN(n4186) );
  NAND2_X1 U5170 ( .A1(n4187), .A2(n4186), .ZN(n4895) );
  INV_X1 U5171 ( .A(n4216), .ZN(n4188) );
  NAND2_X1 U5172 ( .A1(n2997), .A2(n4188), .ZN(n4189) );
  NAND3_X1 U5173 ( .A1(n4894), .A2(n4895), .A3(n4189), .ZN(n4192) );
  NAND2_X1 U5174 ( .A1(n4216), .A2(n4291), .ZN(n4190) );
  NAND3_X1 U5175 ( .A1(n2997), .A2(n3000), .A3(n4190), .ZN(n4191) );
  INV_X1 U5176 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6647) );
  INV_X1 U5177 ( .A(n5157), .ZN(n5133) );
  INV_X1 U5178 ( .A(n4358), .ZN(n4197) );
  NAND3_X1 U5179 ( .A1(n4201), .A2(n4200), .A3(n4199), .ZN(n4202) );
  NAND2_X1 U5180 ( .A1(n4203), .A2(n4202), .ZN(n4205) );
  AND2_X1 U5181 ( .A1(n4205), .A2(n4204), .ZN(n4360) );
  INV_X1 U5182 ( .A(n4360), .ZN(n4206) );
  NAND2_X1 U5183 ( .A1(n4361), .A2(n4206), .ZN(n4354) );
  AND2_X1 U5184 ( .A1(n4208), .A2(n4207), .ZN(n6378) );
  OR2_X1 U5185 ( .A1(n6378), .A2(n5917), .ZN(n4209) );
  INV_X1 U5186 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U5187 ( .A1(n6376), .A2(n6367), .ZN(n6382) );
  NOR3_X1 U5188 ( .A1(n6368), .A2(n6458), .A3(n6382), .ZN(n6359) );
  OR2_X1 U5189 ( .A1(n4209), .A2(n6359), .ZN(n4210) );
  INV_X1 U5190 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4213) );
  XNOR2_X1 U5191 ( .A(n4214), .B(n4213), .ZN(n4959) );
  NOR2_X1 U5192 ( .A1(n4959), .A2(n6376), .ZN(n4215) );
  OR2_X1 U5193 ( .A1(n4216), .A2(n4220), .ZN(n4217) );
  MUX2_X1 U5194 ( .A(n4220), .B(n4219), .S(n4117), .Z(n4221) );
  NAND2_X1 U5195 ( .A1(n4216), .A2(n4221), .ZN(n4222) );
  INV_X1 U5196 ( .A(READY_N), .ZN(n6483) );
  NAND2_X1 U5197 ( .A1(n6483), .A2(n6224), .ZN(n4229) );
  AND3_X1 U5198 ( .A1(n4223), .A2(EBX_REG_31__SCAN_IN), .A3(n4229), .ZN(n4224)
         );
  INV_X1 U5199 ( .A(n4225), .ZN(n4226) );
  INV_X1 U5200 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U5201 ( .A1(n4226), .A2(n6393), .ZN(n6391) );
  NOR2_X1 U5202 ( .A1(n6391), .A2(n4229), .ZN(n6363) );
  INV_X1 U5203 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5052) );
  NAND3_X1 U5204 ( .A1(n3249), .A2(n4229), .A3(n5052), .ZN(n4227) );
  OAI21_X1 U5205 ( .B1(n6485), .B2(n6363), .A(n4227), .ZN(n4228) );
  INV_X1 U5206 ( .A(n6391), .ZN(n4412) );
  NAND2_X1 U5207 ( .A1(n3249), .A2(n4412), .ZN(n4230) );
  AOI21_X1 U5208 ( .B1(n4897), .B2(n4230), .A(n4229), .ZN(n4231) );
  NAND3_X1 U5209 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4233) );
  INV_X1 U5210 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6433) );
  INV_X1 U5211 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6424) );
  INV_X1 U5212 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6421) );
  INV_X1 U5213 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6415) );
  INV_X1 U5214 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6411) );
  INV_X1 U5215 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6505) );
  NAND3_X1 U5216 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5728) );
  NOR2_X1 U5217 ( .A1(n6505), .A2(n5728), .ZN(n5718) );
  NAND2_X1 U5218 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5718), .ZN(n5693) );
  NOR2_X1 U5219 ( .A1(n6411), .A2(n5693), .ZN(n5698) );
  NAND2_X1 U5220 ( .A1(REIP_REG_7__SCAN_IN), .A2(n5698), .ZN(n4345) );
  NOR2_X1 U5221 ( .A1(n6415), .A2(n4345), .ZN(n4880) );
  NAND4_X1 U5222 ( .A1(n4880), .A2(REIP_REG_11__SCAN_IN), .A3(
        REIP_REG_10__SCAN_IN), .A4(REIP_REG_9__SCAN_IN), .ZN(n4881) );
  NOR2_X1 U5223 ( .A1(n6421), .A2(n4881), .ZN(n5045) );
  NAND2_X1 U5224 ( .A1(REIP_REG_13__SCAN_IN), .A2(n5045), .ZN(n5650) );
  NOR2_X1 U5225 ( .A1(n6424), .A2(n5650), .ZN(n5646) );
  NAND4_X1 U5226 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .A4(n5646), .ZN(n5022) );
  NAND2_X1 U5227 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5497) );
  NOR2_X1 U5228 ( .A1(n5022), .A2(n5497), .ZN(n5005) );
  NAND2_X1 U5229 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5005), .ZN(n5488) );
  NOR2_X1 U5230 ( .A1(n6433), .A2(n5488), .ZN(n5468) );
  NAND3_X1 U5231 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        n5468), .ZN(n4240) );
  INV_X1 U5232 ( .A(n5755), .ZN(n5723) );
  AOI21_X1 U5233 ( .B1(n4240), .B2(n5724), .A(n5723), .ZN(n5470) );
  INV_X1 U5234 ( .A(n5470), .ZN(n4232) );
  AOI21_X1 U5235 ( .B1(n5724), .B2(n4233), .A(n4232), .ZN(n5451) );
  NAND2_X1 U5236 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4241) );
  NAND2_X1 U5237 ( .A1(n5724), .A2(n4241), .ZN(n4234) );
  NAND2_X1 U5238 ( .A1(n5451), .A2(n4234), .ZN(n4994) );
  NAND2_X1 U5239 ( .A1(n4994), .A2(REIP_REG_29__SCAN_IN), .ZN(n4238) );
  AND2_X1 U5240 ( .A1(n4959), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4235) );
  INV_X1 U5241 ( .A(n5155), .ZN(n4236) );
  AOI22_X1 U5242 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n5764), .B1(n5763), 
        .B2(n4236), .ZN(n4237) );
  OAI211_X1 U5243 ( .C1(n4938), .C2(n5761), .A(n4238), .B(n4237), .ZN(n4239)
         );
  INV_X1 U5244 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6438) );
  NOR2_X1 U5245 ( .A1(n5754), .A2(n4240), .ZN(n5452) );
  NAND2_X1 U5246 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5452), .ZN(n5453) );
  NOR2_X1 U5247 ( .A1(n6438), .A2(n5453), .ZN(n5443) );
  AND2_X1 U5248 ( .A1(n5443), .A2(REIP_REG_26__SCAN_IN), .ZN(n5438) );
  INV_X1 U5249 ( .A(n4241), .ZN(n4242) );
  NAND2_X1 U5250 ( .A1(n5438), .A2(n4242), .ZN(n4977) );
  NOR2_X1 U5251 ( .A1(n4977), .A2(REIP_REG_29__SCAN_IN), .ZN(n4243) );
  XNOR2_X1 U5252 ( .A(n5228), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5532)
         );
  NAND2_X1 U5253 ( .A1(n5533), .A2(n5532), .ZN(n4248) );
  INV_X1 U5254 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4246) );
  NAND2_X1 U5255 ( .A1(n5228), .A2(n4246), .ZN(n4247) );
  NAND2_X1 U5256 ( .A1(n4248), .A2(n4247), .ZN(n5206) );
  INV_X1 U5257 ( .A(n5206), .ZN(n4250) );
  INV_X1 U5258 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4251) );
  XNOR2_X1 U5259 ( .A(n5228), .B(n4251), .ZN(n5207) );
  OR2_X1 U5260 ( .A1(n5228), .A2(n4251), .ZN(n4252) );
  XNOR2_X1 U5261 ( .A(n5228), .B(n5183), .ZN(n5199) );
  NOR3_X1 U5262 ( .A1(n4253), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n5228), 
        .ZN(n5185) );
  OR2_X1 U5263 ( .A1(n4255), .A2(n5574), .ZN(n5214) );
  OR2_X1 U5264 ( .A1(n5214), .A2(n4909), .ZN(n4258) );
  INV_X1 U5265 ( .A(n4256), .ZN(n4257) );
  NOR3_X1 U5266 ( .A1(n4258), .A2(n3075), .A3(n4257), .ZN(n4259) );
  NOR2_X1 U5267 ( .A1(n5185), .A2(n4259), .ZN(n4260) );
  NAND2_X1 U5268 ( .A1(n4288), .A2(n5916), .ZN(n4270) );
  INV_X1 U5269 ( .A(n4262), .ZN(n4264) );
  OAI21_X1 U5270 ( .B1(n4264), .B2(n3077), .A(n5079), .ZN(n5472) );
  INV_X1 U5271 ( .A(REIP_REG_23__SCAN_IN), .ZN(n4265) );
  NOR2_X1 U5272 ( .A1(n6684), .A2(n4265), .ZN(n4320) );
  NOR2_X1 U5273 ( .A1(n5914), .A2(n5476), .ZN(n4266) );
  AOI211_X1 U5274 ( .C1(n5919), .C2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n4320), 
        .B(n4266), .ZN(n4267) );
  NAND2_X1 U5275 ( .A1(n4270), .A2(n4269), .ZN(U2963) );
  OR2_X1 U5276 ( .A1(n4429), .A2(n4550), .ZN(n4271) );
  OAI22_X1 U5277 ( .A1(n4418), .A2(n4271), .B1(n4361), .B2(n4282), .ZN(n4272)
         );
  INV_X1 U5278 ( .A(n4272), .ZN(n4421) );
  OAI21_X1 U5279 ( .B1(n4273), .B2(READY_N), .A(n3249), .ZN(n4274) );
  OAI21_X1 U5280 ( .B1(n4412), .B2(n6485), .A(n4274), .ZN(n4276) );
  NAND2_X1 U5281 ( .A1(n4276), .A2(n4275), .ZN(n4277) );
  NAND2_X1 U5282 ( .A1(n4418), .A2(n4277), .ZN(n4279) );
  NOR2_X1 U5283 ( .A1(READY_N), .A2(n4360), .ZN(n4378) );
  OAI21_X1 U5284 ( .B1(n4550), .B2(n4412), .A(n4378), .ZN(n4278) );
  NAND2_X1 U5285 ( .A1(n4421), .A2(n4280), .ZN(n4281) );
  INV_X1 U5286 ( .A(n4381), .ZN(n4457) );
  NOR2_X1 U5287 ( .A1(n4283), .A2(n3306), .ZN(n4284) );
  NOR2_X1 U5288 ( .A1(n4357), .A2(n4284), .ZN(n4286) );
  INV_X1 U5289 ( .A(n4285), .ZN(n5598) );
  NAND4_X1 U5290 ( .A1(n4457), .A2(n4286), .A3(n5408), .A4(n4413), .ZN(n4287)
         );
  NAND2_X1 U5291 ( .A1(n4288), .A2(n5951), .ZN(n4331) );
  INV_X1 U5292 ( .A(n4456), .ZN(n4362) );
  INV_X1 U5293 ( .A(n4289), .ZN(n4292) );
  AOI21_X1 U5294 ( .B1(n3216), .B2(n5787), .A(n4101), .ZN(n4290) );
  AOI21_X1 U5295 ( .B1(n4292), .B2(n4291), .A(n4290), .ZN(n4293) );
  AND2_X1 U5296 ( .A1(n4294), .A2(n4293), .ZN(n4296) );
  AND2_X1 U5297 ( .A1(n4296), .A2(n4295), .ZN(n4407) );
  INV_X1 U5298 ( .A(n4297), .ZN(n4403) );
  AOI22_X1 U5299 ( .A1(n4403), .A2(n5787), .B1(n4402), .B2(n4298), .ZN(n4301)
         );
  NAND2_X1 U5300 ( .A1(n4415), .A2(n4487), .ZN(n4299) );
  NAND2_X1 U5301 ( .A1(n4299), .A2(n4602), .ZN(n4404) );
  OR2_X1 U5302 ( .A1(n4429), .A2(n4300), .ZN(n4923) );
  NAND4_X1 U5303 ( .A1(n4407), .A2(n4301), .A3(n4404), .A4(n4923), .ZN(n4302)
         );
  NAND2_X1 U5304 ( .A1(n4304), .A2(n4302), .ZN(n4310) );
  AND2_X1 U5305 ( .A1(n5940), .A2(n4310), .ZN(n5375) );
  NOR2_X1 U5306 ( .A1(n4909), .A2(n5346), .ZN(n4318) );
  NOR2_X1 U5307 ( .A1(n3500), .A2(n5387), .ZN(n5374) );
  NAND3_X1 U5308 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n5374), .ZN(n5573) );
  NOR2_X1 U5309 ( .A1(n4305), .A2(n5573), .ZN(n5571) );
  NAND2_X1 U5310 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n5571), .ZN(n4317) );
  INV_X1 U5311 ( .A(n4317), .ZN(n4309) );
  NAND2_X1 U5312 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4315) );
  NAND2_X1 U5313 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4520) );
  NOR2_X1 U5314 ( .A1(n4315), .A2(n4520), .ZN(n4751) );
  NAND3_X1 U5315 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4751), .ZN(n4313) );
  NAND2_X1 U5316 ( .A1(n5371), .A2(n4310), .ZN(n4308) );
  INV_X1 U5317 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U5318 ( .A1(n5954), .A2(n5941), .ZN(n5942) );
  INV_X1 U5319 ( .A(n5942), .ZN(n4504) );
  NOR2_X1 U5320 ( .A1(n4520), .A2(n4504), .ZN(n4314) );
  AND2_X1 U5321 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4314), .ZN(n4498)
         );
  AOI21_X1 U5322 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n4498), .A(n5940), 
        .ZN(n4306) );
  NAND2_X1 U5323 ( .A1(n4328), .A2(n6684), .ZN(n4485) );
  OAI21_X1 U5324 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n4310), .A(n4485), 
        .ZN(n4307) );
  NAND2_X1 U5325 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4752) );
  NAND2_X1 U5326 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4867) );
  NOR2_X1 U5327 ( .A1(n4752), .A2(n4867), .ZN(n4312) );
  NAND2_X1 U5328 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4469) );
  AOI21_X1 U5329 ( .B1(n4469), .B2(n4308), .A(n4307), .ZN(n5955) );
  AOI22_X1 U5330 ( .A1(n2998), .A2(n4312), .B1(n5343), .B2(n5955), .ZN(n5925)
         );
  OAI21_X1 U5331 ( .B1(n5343), .B2(n4309), .A(n5385), .ZN(n5340) );
  INV_X1 U5332 ( .A(n5340), .ZN(n5362) );
  OAI21_X1 U5333 ( .B1(n5343), .B2(n4318), .A(n5362), .ZN(n5332) );
  INV_X1 U5334 ( .A(n4906), .ZN(n4321) );
  INV_X1 U5335 ( .A(n4310), .ZN(n4311) );
  NAND2_X1 U5336 ( .A1(n4311), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5366)
         );
  INV_X1 U5337 ( .A(n4312), .ZN(n4316) );
  NOR2_X1 U5338 ( .A1(n4316), .A2(n4313), .ZN(n5370) );
  INV_X1 U5339 ( .A(n5370), .ZN(n5365) );
  NAND2_X1 U5340 ( .A1(n5342), .A2(n4314), .ZN(n4470) );
  NAND2_X1 U5341 ( .A1(n4911), .A2(n4318), .ZN(n5335) );
  NOR3_X1 U5342 ( .A1(n5335), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n5323), 
        .ZN(n4319) );
  AOI211_X1 U5343 ( .C1(n4321), .C2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n4320), .B(n4319), .ZN(n4329) );
  NOR2_X1 U5344 ( .A1(n4323), .A2(n4324), .ZN(n4325) );
  OR2_X1 U5345 ( .A1(n4322), .A2(n4325), .ZN(n5473) );
  NAND3_X1 U5346 ( .A1(n4402), .A2(n3306), .A3(n3216), .ZN(n4326) );
  NAND2_X1 U5347 ( .A1(n4331), .A2(n4330), .ZN(U2995) );
  OR2_X1 U5348 ( .A1(n5375), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4488)
         );
  AOI21_X1 U5349 ( .B1(n4485), .B2(n4488), .A(n4109), .ZN(n4340) );
  AOI211_X1 U5350 ( .C1(n4930), .C2(n5371), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .B(n5343), .ZN(n4339) );
  AOI21_X1 U5351 ( .B1(n4332), .B2(n4897), .A(n4333), .ZN(n4476) );
  NOR2_X1 U5352 ( .A1(n6688), .A2(n4476), .ZN(n4338) );
  OAI21_X1 U5353 ( .B1(n4336), .B2(n4335), .A(n4334), .ZN(n5271) );
  NAND2_X1 U5354 ( .A1(n5917), .A2(REIP_REG_1__SCAN_IN), .ZN(n5275) );
  OAI21_X1 U5355 ( .B1(n5394), .B2(n5271), .A(n5275), .ZN(n4337) );
  OR4_X1 U5356 ( .A1(n4340), .A2(n4339), .A3(n4338), .A4(n4337), .ZN(U3017) );
  OAI21_X1 U5357 ( .B1(n4880), .B2(n5754), .A(n5755), .ZN(n5680) );
  AOI22_X1 U5358 ( .A1(EBX_REG_8__SCAN_IN), .A2(n5743), .B1(
        REIP_REG_8__SCAN_IN), .B2(n5680), .ZN(n4341) );
  NAND3_X1 U5359 ( .A1(n6464), .A2(n6376), .A3(n5755), .ZN(n5712) );
  OAI211_X1 U5360 ( .C1(n5683), .C2(n4342), .A(n4341), .B(n5712), .ZN(n4353)
         );
  OAI21_X1 U5361 ( .B1(n4564), .B2(n4343), .A(n4755), .ZN(n4778) );
  OR2_X1 U5362 ( .A1(n5754), .A2(n4880), .ZN(n4344) );
  OAI22_X1 U5363 ( .A1(n5671), .A2(n4778), .B1(n4345), .B2(n4344), .ZN(n4352)
         );
  INV_X1 U5364 ( .A(n4346), .ZN(n4350) );
  INV_X1 U5365 ( .A(n4347), .ZN(n4349) );
  OAI21_X1 U5366 ( .B1(n4350), .B2(n4349), .A(n4348), .ZN(n4845) );
  OAI22_X1 U5367 ( .A1(n4845), .A2(n5695), .B1(n5738), .B2(n4847), .ZN(n4351)
         );
  OR3_X1 U5368 ( .A1(n4353), .A2(n4352), .A3(n4351), .ZN(U2819) );
  NAND2_X1 U5369 ( .A1(n4358), .A2(n4354), .ZN(n4355) );
  OAI21_X1 U5370 ( .B1(n4418), .B2(n4731), .A(n4355), .ZN(n5603) );
  OR2_X1 U5371 ( .A1(n4356), .A2(n4735), .ZN(n4370) );
  AOI21_X1 U5372 ( .B1(n6391), .B2(n4370), .A(READY_N), .ZN(n6484) );
  NOR2_X1 U5373 ( .A1(n5603), .A2(n6484), .ZN(n6350) );
  NOR2_X1 U5374 ( .A1(n6350), .A2(n6374), .ZN(n5610) );
  INV_X1 U5375 ( .A(MORE_REG_SCAN_IN), .ZN(n4367) );
  INV_X1 U5376 ( .A(n4357), .ZN(n6352) );
  NAND2_X1 U5377 ( .A1(n6352), .A2(n4358), .ZN(n4359) );
  NOR2_X1 U5378 ( .A1(n4359), .A2(n4381), .ZN(n4365) );
  NAND2_X1 U5379 ( .A1(n4361), .A2(n4360), .ZN(n4364) );
  NAND2_X1 U5380 ( .A1(n4418), .A2(n4362), .ZN(n4363) );
  OAI211_X1 U5381 ( .C1(n4418), .C2(n4365), .A(n4364), .B(n4363), .ZN(n6349)
         );
  NAND2_X1 U5382 ( .A1(n5610), .A2(n6349), .ZN(n4366) );
  OAI21_X1 U5383 ( .B1(n5610), .B2(n4367), .A(n4366), .ZN(U3471) );
  NAND2_X1 U5384 ( .A1(n6464), .A2(n6376), .ZN(n4368) );
  NAND2_X1 U5385 ( .A1(n5842), .A2(n4368), .ZN(n5431) );
  INV_X1 U5386 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n4369) );
  NAND2_X1 U5387 ( .A1(n5432), .A2(n4369), .ZN(n4372) );
  NAND2_X1 U5388 ( .A1(n6481), .A2(n4370), .ZN(n4371) );
  OAI21_X1 U5389 ( .B1(n5431), .B2(n4372), .A(n4371), .ZN(n4373) );
  INV_X1 U5390 ( .A(n4373), .ZN(U3474) );
  OAI21_X1 U5391 ( .B1(n4376), .B2(n4375), .A(n4374), .ZN(n5922) );
  INV_X1 U5392 ( .A(n4378), .ZN(n4379) );
  NOR2_X1 U5393 ( .A1(n5408), .A2(n4379), .ZN(n4380) );
  AOI21_X1 U5394 ( .B1(n4418), .B2(n4381), .A(n4380), .ZN(n4420) );
  NAND2_X1 U5395 ( .A1(n4402), .A2(n4382), .ZN(n4383) );
  AOI21_X1 U5396 ( .B1(n4420), .B2(n4383), .A(n6374), .ZN(n4384) );
  OR2_X1 U5397 ( .A1(n4098), .A2(n5127), .ZN(n4385) );
  INV_X1 U5398 ( .A(n4385), .ZN(n4386) );
  INV_X1 U5399 ( .A(DATAI_0_), .ZN(n6603) );
  INV_X1 U5400 ( .A(EAX_REG_0__SCAN_IN), .ZN(n5838) );
  OAI222_X1 U5401 ( .A1(n5922), .A2(n5507), .B1(n5152), .B2(n6603), .C1(n5151), 
        .C2(n5838), .ZN(U2891) );
  INV_X1 U5402 ( .A(n4387), .ZN(n4388) );
  OAI21_X1 U5403 ( .B1(n4390), .B2(n4389), .A(n4388), .ZN(n5903) );
  INV_X1 U5404 ( .A(DATAI_2_), .ZN(n5866) );
  INV_X1 U5405 ( .A(EAX_REG_2__SCAN_IN), .ZN(n5832) );
  OAI222_X1 U5406 ( .A1(n5903), .A2(n5507), .B1(n5152), .B2(n5866), .C1(n5151), 
        .C2(n5832), .ZN(U2889) );
  OR2_X1 U5407 ( .A1(n4392), .A2(n4391), .ZN(n4393) );
  AND2_X1 U5408 ( .A1(n4394), .A2(n4393), .ZN(n5272) );
  INV_X1 U5409 ( .A(n5272), .ZN(n4477) );
  INV_X1 U5410 ( .A(DATAI_1_), .ZN(n5864) );
  INV_X1 U5411 ( .A(EAX_REG_1__SCAN_IN), .ZN(n5834) );
  OAI222_X1 U5412 ( .A1(n4477), .A2(n5507), .B1(n5152), .B2(n5864), .C1(n5151), 
        .C2(n5834), .ZN(U2890) );
  NAND2_X1 U5413 ( .A1(n4396), .A2(n4397), .ZN(n4398) );
  NAND2_X1 U5414 ( .A1(n4395), .A2(n4398), .ZN(n5733) );
  OAI222_X1 U5415 ( .A1(n5733), .A2(n5126), .B1(n5776), .B2(n4401), .C1(n5122), 
        .C2(n5729), .ZN(U2855) );
  INV_X1 U5416 ( .A(DATAI_4_), .ZN(n5870) );
  INV_X1 U5417 ( .A(EAX_REG_4__SCAN_IN), .ZN(n5828) );
  OAI222_X1 U5418 ( .A1(n5733), .A2(n5507), .B1(n5152), .B2(n5870), .C1(n5151), 
        .C2(n5828), .ZN(U2887) );
  INV_X1 U5419 ( .A(n3582), .ZN(n6461) );
  NOR2_X1 U5420 ( .A1(n4403), .A2(n4402), .ZN(n4405) );
  AND4_X1 U5421 ( .A1(n5408), .A2(n4273), .A3(n4405), .A4(n4404), .ZN(n4406)
         );
  AND2_X1 U5422 ( .A1(n4407), .A2(n4406), .ZN(n4928) );
  INV_X1 U5423 ( .A(n4928), .ZN(n4409) );
  INV_X1 U5424 ( .A(n4429), .ZN(n4408) );
  AOI22_X1 U5425 ( .A1(n6461), .A2(n4409), .B1(n4408), .B2(n3090), .ZN(n6334)
         );
  INV_X1 U5426 ( .A(n6334), .ZN(n4411) );
  OAI22_X1 U5427 ( .A1(n6376), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(n3057), 
        .B2(n4931), .ZN(n4410) );
  AOI21_X1 U5428 ( .B1(n4411), .B2(n5597), .A(n4410), .ZN(n4424) );
  OAI21_X1 U5429 ( .B1(n3060), .B2(n5429), .A(n4412), .ZN(n4414) );
  AOI21_X1 U5430 ( .B1(n4414), .B2(n4413), .A(READY_N), .ZN(n4417) );
  INV_X1 U5431 ( .A(n4415), .ZN(n4416) );
  AOI21_X1 U5432 ( .B1(n4418), .B2(n4417), .A(n4416), .ZN(n4419) );
  AND2_X1 U5433 ( .A1(n4420), .A2(n4419), .ZN(n4422) );
  NAND2_X1 U5434 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6462), .ZN(n6456) );
  INV_X1 U5435 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5609) );
  OAI22_X1 U5436 ( .A1(n6341), .A2(n6374), .B1(n6456), .B2(n5609), .ZN(n5599)
         );
  AOI21_X1 U5437 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6368), .A(n5599), .ZN(
        n4936) );
  AOI21_X1 U5438 ( .B1(n5429), .B2(n5597), .A(n4936), .ZN(n4423) );
  OAI22_X1 U5439 ( .A1(n4424), .A2(n4936), .B1(n4423), .B2(n3090), .ZN(U3461)
         );
  INV_X1 U5440 ( .A(n4931), .ZN(n6366) );
  INV_X1 U5441 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4915) );
  AOI22_X1 U5442 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4915), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4109), .ZN(n4929) );
  NOR2_X1 U5443 ( .A1(n6376), .A2(n4930), .ZN(n4432) );
  INV_X1 U5444 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4920) );
  NOR3_X1 U5445 ( .A1(n4429), .A2(n4427), .A3(n4428), .ZN(n4430) );
  AOI21_X1 U5446 ( .B1(n5429), .B2(n4920), .A(n4430), .ZN(n4431) );
  OAI21_X1 U5447 ( .B1(n5396), .B2(n4928), .A(n4431), .ZN(n6336) );
  AOI222_X1 U5448 ( .A1(n6366), .A2(n4433), .B1(n4929), .B2(n4432), .C1(n6336), 
        .C2(n5597), .ZN(n4436) );
  AOI22_X1 U5449 ( .A1(n4434), .A2(n6366), .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n4936), .ZN(n4435) );
  OAI21_X1 U5450 ( .B1(n4436), .B2(n4936), .A(n4435), .ZN(U3460) );
  XNOR2_X1 U5451 ( .A(n4438), .B(n4437), .ZN(n4509) );
  OR2_X1 U5452 ( .A1(n4387), .A2(n4439), .ZN(n4440) );
  NAND2_X1 U5453 ( .A1(n4396), .A2(n4440), .ZN(n5748) );
  INV_X1 U5454 ( .A(n5748), .ZN(n4443) );
  INV_X1 U5455 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6406) );
  NOR2_X1 U5456 ( .A1(n6684), .A2(n6406), .ZN(n4506) );
  AOI21_X1 U5457 ( .B1(n5919), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4506), 
        .ZN(n4441) );
  OAI21_X1 U5458 ( .B1(n5741), .B2(n5914), .A(n4441), .ZN(n4442) );
  AOI21_X1 U5459 ( .B1(n5909), .B2(n4443), .A(n4442), .ZN(n4444) );
  OAI21_X1 U5460 ( .B1(n4509), .B2(n3056), .A(n4444), .ZN(U2983) );
  NAND2_X1 U5461 ( .A1(n4395), .A2(n4445), .ZN(n4446) );
  NAND2_X1 U5462 ( .A1(n4589), .A2(n4446), .ZN(n4511) );
  AOI21_X1 U5463 ( .B1(n4448), .B2(n4399), .A(n4447), .ZN(n5710) );
  INV_X1 U5464 ( .A(n5710), .ZN(n4449) );
  OAI222_X1 U5465 ( .A1(n5126), .A2(n4511), .B1(n5776), .B2(n5713), .C1(n5122), 
        .C2(n4449), .ZN(U2854) );
  INV_X1 U5466 ( .A(n6101), .ZN(n6051) );
  XNOR2_X1 U5467 ( .A(n4451), .B(n3104), .ZN(n4455) );
  INV_X1 U5468 ( .A(n4923), .ZN(n4454) );
  INV_X1 U5469 ( .A(n4452), .ZN(n4453) );
  OAI211_X1 U5470 ( .C1(n4427), .C2(n3104), .A(n3189), .B(n4453), .ZN(n4464)
         );
  AOI22_X1 U5471 ( .A1(n5429), .A2(n4455), .B1(n4454), .B2(n4464), .ZN(n4463)
         );
  NAND2_X1 U5472 ( .A1(n4457), .A2(n4456), .ZN(n4926) );
  INV_X1 U5473 ( .A(n4458), .ZN(n4459) );
  MUX2_X1 U5474 ( .A(n4459), .B(n3104), .S(n4427), .Z(n4460) );
  NAND3_X1 U5475 ( .A1(n4926), .A2(n4461), .A3(n4460), .ZN(n4462) );
  OAI211_X1 U5476 ( .C1(n6051), .C2(n4928), .A(n4463), .B(n4462), .ZN(n5400)
         );
  AOI22_X1 U5477 ( .A1(n5400), .A2(n5597), .B1(n4464), .B2(n6366), .ZN(n4465)
         );
  INV_X1 U5478 ( .A(n4936), .ZN(n5601) );
  MUX2_X1 U5479 ( .A(n3104), .B(n4465), .S(n5601), .Z(n4466) );
  INV_X1 U5480 ( .A(n4466), .ZN(U3456) );
  XNOR2_X1 U5481 ( .A(n4468), .B(n3058), .ZN(n4516) );
  OAI21_X1 U5482 ( .B1(n5343), .B2(n4498), .A(n5955), .ZN(n4499) );
  NOR2_X1 U5483 ( .A1(n5948), .A2(n4469), .ZN(n4496) );
  INV_X1 U5484 ( .A(n4496), .ZN(n4472) );
  OAI211_X1 U5485 ( .C1(n4520), .C2(n4472), .A(n4471), .B(n4470), .ZN(n4473)
         );
  NAND2_X1 U5486 ( .A1(n4499), .A2(n4473), .ZN(n4475) );
  AND2_X1 U5487 ( .A1(n5917), .A2(REIP_REG_5__SCAN_IN), .ZN(n4512) );
  AOI21_X1 U5488 ( .B1(n5944), .B2(n5710), .A(n4512), .ZN(n4474) );
  OAI211_X1 U5489 ( .C1(n4516), .C2(n5394), .A(n4475), .B(n4474), .ZN(U3013)
         );
  INV_X1 U5490 ( .A(DATAI_5_), .ZN(n5872) );
  OAI222_X1 U5491 ( .A1(n4511), .A2(n5507), .B1(n5152), .B2(n5872), .C1(n5151), 
        .C2(n3622), .ZN(U2886) );
  INV_X1 U5492 ( .A(DATAI_3_), .ZN(n5868) );
  INV_X1 U5493 ( .A(EAX_REG_3__SCAN_IN), .ZN(n5830) );
  OAI222_X1 U5494 ( .A1(n5748), .A2(n5507), .B1(n5152), .B2(n5868), .C1(n5151), 
        .C2(n5830), .ZN(U2888) );
  OAI222_X1 U5495 ( .A1(n4477), .A2(n5126), .B1(n5776), .B2(n4736), .C1(n5122), 
        .C2(n4476), .ZN(U2858) );
  AOI22_X1 U5496 ( .A1(n4194), .A2(n3016), .B1(EBX_REG_3__SCAN_IN), .B2(n5103), 
        .ZN(n4480) );
  OAI21_X1 U5497 ( .B1(n5748), .B2(n5126), .A(n4480), .ZN(U2856) );
  INV_X1 U5498 ( .A(n4481), .ZN(n4484) );
  INV_X1 U5499 ( .A(n4482), .ZN(n4483) );
  AOI21_X1 U5500 ( .B1(n4484), .B2(n4930), .A(n4483), .ZN(n5915) );
  AOI21_X1 U5501 ( .B1(n5371), .B2(n4485), .A(n4930), .ZN(n4492) );
  INV_X1 U5502 ( .A(REIP_REG_0__SCAN_IN), .ZN(n4490) );
  AOI21_X1 U5503 ( .B1(n4487), .B2(n4930), .A(n4486), .ZN(n5757) );
  NAND2_X1 U5504 ( .A1(n5944), .A2(n5757), .ZN(n4489) );
  OAI211_X1 U5505 ( .C1(n6684), .C2(n4490), .A(n4489), .B(n4488), .ZN(n4491)
         );
  AOI211_X1 U5506 ( .C1(n5951), .C2(n5915), .A(n4492), .B(n4491), .ZN(n4493)
         );
  INV_X1 U5507 ( .A(n4493), .ZN(U3018) );
  XNOR2_X1 U5508 ( .A(n4494), .B(n4495), .ZN(n4596) );
  NOR2_X1 U5509 ( .A1(n5342), .A2(n4496), .ZN(n4503) );
  NOR2_X1 U5510 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4503), .ZN(n4497)
         );
  AOI22_X1 U5511 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4499), .B1(n4498), 
        .B2(n4497), .ZN(n4502) );
  XOR2_X1 U5512 ( .A(n4447), .B(n4500), .Z(n5771) );
  AND2_X1 U5513 ( .A1(n5917), .A2(REIP_REG_6__SCAN_IN), .ZN(n4592) );
  AOI21_X1 U5514 ( .B1(n5944), .B2(n5771), .A(n4592), .ZN(n4501) );
  OAI211_X1 U5515 ( .C1(n5394), .C2(n4596), .A(n4502), .B(n4501), .ZN(U3012)
         );
  OAI21_X1 U5516 ( .B1(n5940), .B2(n5942), .A(n5955), .ZN(n4519) );
  NOR2_X1 U5517 ( .A1(n4504), .A2(n4503), .ZN(n4750) );
  AOI22_X1 U5518 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4519), .B1(n4750), 
        .B2(n4505), .ZN(n4508) );
  AOI21_X1 U5519 ( .B1(n5944), .B2(n3016), .A(n4506), .ZN(n4507) );
  OAI211_X1 U5520 ( .C1(n4509), .C2(n5394), .A(n4508), .B(n4507), .ZN(U3015)
         );
  INV_X1 U5521 ( .A(n5757), .ZN(n4510) );
  OAI222_X1 U5522 ( .A1(n5126), .A2(n5922), .B1(n5776), .B2(n5760), .C1(n5122), 
        .C2(n4510), .ZN(U2859) );
  INV_X1 U5523 ( .A(n4511), .ZN(n5716) );
  AOI21_X1 U5524 ( .B1(n5919), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4512), 
        .ZN(n4513) );
  OAI21_X1 U5525 ( .B1(n5721), .B2(n5914), .A(n4513), .ZN(n4514) );
  AOI21_X1 U5526 ( .B1(n5716), .B2(n5909), .A(n4514), .ZN(n4515) );
  OAI21_X1 U5527 ( .B1(n4516), .B2(n3056), .A(n4515), .ZN(U2981) );
  OAI22_X1 U5528 ( .A1(n6688), .A2(n5729), .B1(n6505), .B2(n6684), .ZN(n4518)
         );
  AOI21_X1 U5529 ( .B1(n4519), .B2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4518), 
        .ZN(n4522) );
  OAI211_X1 U5530 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n4750), .B(n4520), .ZN(n4521) );
  OAI211_X1 U5531 ( .C1(n5394), .C2(n4559), .A(n4522), .B(n4521), .ZN(U3014)
         );
  NOR2_X2 U5532 ( .A1(n4740), .A2(n4101), .ZN(n6294) );
  INV_X1 U5533 ( .A(n6294), .ZN(n4629) );
  NAND3_X1 U5534 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6231), .A3(n6337), .ZN(n4696) );
  NOR2_X1 U5535 ( .A1(n6468), .A2(n4696), .ZN(n4530) );
  INV_X1 U5536 ( .A(n4530), .ZN(n4747) );
  INV_X1 U5537 ( .A(n6191), .ZN(n6281) );
  INV_X1 U5538 ( .A(n4608), .ZN(n4524) );
  INV_X1 U5539 ( .A(n5424), .ZN(n4528) );
  NOR2_X1 U5540 ( .A1(n4526), .A2(n6224), .ZN(n4527) );
  AOI21_X1 U5541 ( .B1(n4528), .B2(n4527), .A(n6271), .ZN(n4532) );
  INV_X1 U5542 ( .A(n5420), .ZN(n4802) );
  NAND2_X1 U5543 ( .A1(n4802), .A2(n5396), .ZN(n6187) );
  NOR2_X1 U5544 ( .A1(n6187), .A2(n4679), .ZN(n4698) );
  AOI21_X1 U5545 ( .B1(n4698), .B2(n6461), .A(n4530), .ZN(n4534) );
  AOI22_X1 U5546 ( .A1(n4532), .A2(n4534), .B1(n6271), .B2(n4696), .ZN(n4531)
         );
  NAND2_X1 U5547 ( .A1(n6281), .A2(n4531), .ZN(n4742) );
  NOR2_X2 U5548 ( .A1(n5866), .A2(n5416), .ZN(n6293) );
  INV_X1 U5549 ( .A(n4532), .ZN(n4533) );
  OAI22_X1 U5550 ( .A1(n4534), .A2(n4533), .B1(n6367), .B2(n4696), .ZN(n4741)
         );
  AOI22_X1 U5551 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n4742), .B1(n6293), 
        .B2(n4741), .ZN(n4540) );
  INV_X1 U5552 ( .A(DATAI_26_), .ZN(n4535) );
  NOR2_X1 U5553 ( .A1(n5213), .A2(n4535), .ZN(n6241) );
  NOR2_X2 U5554 ( .A1(n4537), .A2(n6465), .ZN(n4792) );
  INV_X1 U5555 ( .A(DATAI_18_), .ZN(n4538) );
  NOR2_X1 U5556 ( .A1(n6275), .A2(n4538), .ZN(n6295) );
  AOI22_X1 U5557 ( .A1(n6241), .A2(n4792), .B1(n4801), .B2(n6295), .ZN(n4539)
         );
  OAI211_X1 U5558 ( .C1(n4629), .C2(n4747), .A(n4540), .B(n4539), .ZN(U3062)
         );
  NOR2_X2 U5559 ( .A1(n4740), .A2(n5127), .ZN(n6326) );
  INV_X1 U5560 ( .A(n6326), .ZN(n4632) );
  INV_X1 U5561 ( .A(DATAI_7_), .ZN(n5876) );
  NOR2_X2 U5562 ( .A1(n5876), .A2(n5416), .ZN(n6324) );
  AOI22_X1 U5563 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n4742), .B1(n6324), 
        .B2(n4741), .ZN(n4544) );
  INV_X1 U5564 ( .A(DATAI_31_), .ZN(n4541) );
  NOR2_X1 U5565 ( .A1(n5213), .A2(n4541), .ZN(n6264) );
  INV_X1 U5566 ( .A(DATAI_23_), .ZN(n4542) );
  NOR2_X1 U5567 ( .A1(n5213), .A2(n4542), .ZN(n6328) );
  AOI22_X1 U5568 ( .A1(n6264), .A2(n4792), .B1(n4801), .B2(n6328), .ZN(n4543)
         );
  OAI211_X1 U5569 ( .C1(n4632), .C2(n4747), .A(n4544), .B(n4543), .ZN(U3067)
         );
  INV_X1 U5570 ( .A(n3573), .ZN(n4545) );
  NOR2_X2 U5571 ( .A1(n4740), .A2(n4545), .ZN(n6318) );
  INV_X1 U5572 ( .A(n6318), .ZN(n4635) );
  INV_X1 U5573 ( .A(DATAI_6_), .ZN(n5874) );
  NOR2_X2 U5574 ( .A1(n5874), .A2(n5416), .ZN(n6317) );
  AOI22_X1 U5575 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n4742), .B1(n6317), 
        .B2(n4741), .ZN(n4549) );
  INV_X1 U5576 ( .A(DATAI_30_), .ZN(n4546) );
  NOR2_X1 U5577 ( .A1(n5213), .A2(n4546), .ZN(n6257) );
  INV_X1 U5578 ( .A(DATAI_22_), .ZN(n4547) );
  NOR2_X2 U5579 ( .A1(n5213), .A2(n4547), .ZN(n6319) );
  AOI22_X1 U5580 ( .A1(n6257), .A2(n4792), .B1(n4801), .B2(n6319), .ZN(n4548)
         );
  OAI211_X1 U5581 ( .C1(n4635), .C2(n4747), .A(n4549), .B(n4548), .ZN(U3066)
         );
  NOR2_X2 U5582 ( .A1(n4740), .A2(n4550), .ZN(n6288) );
  INV_X1 U5583 ( .A(n6288), .ZN(n4620) );
  NOR2_X2 U5584 ( .A1(n5864), .A2(n5416), .ZN(n6287) );
  AOI22_X1 U5585 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n4742), .B1(n6287), 
        .B2(n4741), .ZN(n4554) );
  INV_X1 U5586 ( .A(DATAI_25_), .ZN(n4551) );
  NOR2_X1 U5587 ( .A1(n5213), .A2(n4551), .ZN(n6237) );
  INV_X1 U5588 ( .A(DATAI_17_), .ZN(n4552) );
  NOR2_X1 U5589 ( .A1(n6275), .A2(n4552), .ZN(n6289) );
  AOI22_X1 U5590 ( .A1(n6237), .A2(n4792), .B1(n4801), .B2(n6289), .ZN(n4553)
         );
  OAI211_X1 U5591 ( .C1(n4620), .C2(n4747), .A(n4554), .B(n4553), .ZN(U3061)
         );
  OAI22_X1 U5592 ( .A1(n5553), .A2(n4555), .B1(n6684), .B2(n6505), .ZN(n4557)
         );
  NOR2_X1 U5593 ( .A1(n5733), .A2(n6275), .ZN(n4556) );
  AOI211_X1 U5594 ( .C1(n5897), .C2(n5722), .A(n4557), .B(n4556), .ZN(n4558)
         );
  OAI21_X1 U5595 ( .B1(n3056), .B2(n4559), .A(n4558), .ZN(U2982) );
  XOR2_X1 U5596 ( .A(n4561), .B(n4560), .Z(n5943) );
  INV_X1 U5597 ( .A(n5943), .ZN(n4786) );
  INV_X1 U5598 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4562) );
  OAI222_X1 U5599 ( .A1(n4786), .A2(n5122), .B1(n4562), .B2(n5776), .C1(n5903), 
        .C2(n5126), .ZN(U2857) );
  OAI21_X1 U5600 ( .B1(n3067), .B2(n4563), .A(n4346), .ZN(n5696) );
  AOI21_X1 U5601 ( .B1(n4566), .B2(n4565), .A(n4564), .ZN(n5931) );
  AOI22_X1 U5602 ( .A1(n5931), .A2(n4194), .B1(EBX_REG_7__SCAN_IN), .B2(n5103), 
        .ZN(n4567) );
  OAI21_X1 U5603 ( .B1(n5696), .B2(n5126), .A(n4567), .ZN(U2852) );
  NAND2_X1 U5604 ( .A1(n4526), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5423) );
  NOR2_X1 U5605 ( .A1(n5423), .A2(n3074), .ZN(n5419) );
  NAND2_X1 U5606 ( .A1(n5419), .A2(n5957), .ZN(n4568) );
  NAND2_X1 U5607 ( .A1(n4568), .A2(n6464), .ZN(n4574) );
  AND2_X1 U5608 ( .A1(n5420), .A2(n4426), .ZN(n6024) );
  NAND2_X1 U5609 ( .A1(n6024), .A2(n6101), .ZN(n6140) );
  NOR2_X1 U5610 ( .A1(n6231), .A2(n4606), .ZN(n6169) );
  INV_X1 U5611 ( .A(n6169), .ZN(n4569) );
  OAI21_X1 U5612 ( .B1(n6140), .B2(n3582), .A(n4569), .ZN(n4572) );
  NAND2_X1 U5613 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4611), .ZN(n6132) );
  INV_X1 U5614 ( .A(n6132), .ZN(n4575) );
  OAI22_X1 U5615 ( .A1(n4574), .A2(n4572), .B1(n6464), .B2(n4575), .ZN(n4570)
         );
  NAND2_X1 U5616 ( .A1(n6288), .A2(n6169), .ZN(n4580) );
  NAND2_X1 U5617 ( .A1(n4526), .A2(n3581), .ZN(n6218) );
  INV_X1 U5618 ( .A(n4617), .ZN(n4571) );
  NAND2_X1 U5619 ( .A1(n4526), .A2(n6465), .ZN(n5960) );
  NOR2_X1 U5620 ( .A1(n5960), .A2(n3074), .ZN(n4616) );
  AOI22_X1 U5621 ( .A1(n6237), .A2(n6156), .B1(n6181), .B2(n6289), .ZN(n4579)
         );
  INV_X1 U5622 ( .A(n4572), .ZN(n4573) );
  OR2_X1 U5623 ( .A1(n4574), .A2(n4573), .ZN(n4577) );
  NAND2_X1 U5624 ( .A1(n4575), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4576) );
  NAND2_X1 U5625 ( .A1(n4577), .A2(n4576), .ZN(n6170) );
  NAND2_X1 U5626 ( .A1(n6170), .A2(n6287), .ZN(n4578) );
  NAND3_X1 U5627 ( .A1(n4580), .A2(n4579), .A3(n4578), .ZN(n4581) );
  AOI21_X1 U5628 ( .B1(n6171), .B2(INSTQUEUE_REG_11__1__SCAN_IN), .A(n4581), 
        .ZN(n4582) );
  INV_X1 U5629 ( .A(n4582), .ZN(U3109) );
  NAND2_X1 U5630 ( .A1(n6318), .A2(n6169), .ZN(n4585) );
  AOI22_X1 U5631 ( .A1(n6257), .A2(n6156), .B1(n6181), .B2(n6319), .ZN(n4584)
         );
  NAND2_X1 U5632 ( .A1(n6170), .A2(n6317), .ZN(n4583) );
  NAND3_X1 U5633 ( .A1(n4585), .A2(n4584), .A3(n4583), .ZN(n4586) );
  AOI21_X1 U5634 ( .B1(n6171), .B2(INSTQUEUE_REG_11__6__SCAN_IN), .A(n4586), 
        .ZN(n4587) );
  INV_X1 U5635 ( .A(n4587), .ZN(U3114) );
  AOI21_X1 U5636 ( .B1(n4590), .B2(n4589), .A(n3067), .ZN(n5773) );
  INV_X1 U5637 ( .A(n5773), .ZN(n4591) );
  OAI222_X1 U5638 ( .A1(n4591), .A2(n5507), .B1(n5152), .B2(n5874), .C1(n5151), 
        .C2(n3630), .ZN(U2885) );
  AOI21_X1 U5639 ( .B1(n5919), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n4592), 
        .ZN(n4593) );
  OAI21_X1 U5640 ( .B1(n5705), .B2(n5914), .A(n4593), .ZN(n4594) );
  AOI21_X1 U5641 ( .B1(n5773), .B2(n5909), .A(n4594), .ZN(n4595) );
  OAI21_X1 U5642 ( .B1(n3056), .B2(n4596), .A(n4595), .ZN(U2980) );
  OAI222_X1 U5643 ( .A1(n5696), .A2(n5507), .B1(n5152), .B2(n5876), .C1(n5151), 
        .C2(n3638), .ZN(U2884) );
  NOR2_X2 U5644 ( .A1(n4740), .A2(n4597), .ZN(n6312) );
  INV_X1 U5645 ( .A(n6312), .ZN(n4626) );
  NOR2_X2 U5646 ( .A1(n5872), .A2(n5416), .ZN(n6311) );
  AOI22_X1 U5647 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n4742), .B1(n6311), 
        .B2(n4741), .ZN(n4601) );
  INV_X1 U5648 ( .A(DATAI_29_), .ZN(n4598) );
  NOR2_X1 U5649 ( .A1(n5213), .A2(n4598), .ZN(n6253) );
  INV_X1 U5650 ( .A(DATAI_21_), .ZN(n4599) );
  NOR2_X2 U5651 ( .A1(n5213), .A2(n4599), .ZN(n6313) );
  AOI22_X1 U5652 ( .A1(n6253), .A2(n4792), .B1(n4801), .B2(n6313), .ZN(n4600)
         );
  OAI211_X1 U5653 ( .C1(n4626), .C2(n4747), .A(n4601), .B(n4600), .ZN(U3065)
         );
  NOR2_X2 U5654 ( .A1(n4740), .A2(n4602), .ZN(n6300) );
  INV_X1 U5655 ( .A(n6300), .ZN(n4623) );
  NOR2_X2 U5656 ( .A1(n5868), .A2(n5416), .ZN(n6299) );
  AOI22_X1 U5657 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n4742), .B1(n6299), 
        .B2(n4741), .ZN(n4605) );
  NAND2_X1 U5658 ( .A1(n5909), .A2(DATAI_27_), .ZN(n6304) );
  INV_X1 U5659 ( .A(n6304), .ZN(n6245) );
  INV_X1 U5660 ( .A(DATAI_19_), .ZN(n4603) );
  NOR2_X2 U5661 ( .A1(n5213), .A2(n4603), .ZN(n6301) );
  AOI22_X1 U5662 ( .A1(n6245), .A2(n4792), .B1(n4801), .B2(n6301), .ZN(n4604)
         );
  OAI211_X1 U5663 ( .C1(n4623), .C2(n4747), .A(n4605), .B(n4604), .ZN(U3063)
         );
  OR2_X1 U5664 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4606), .ZN(n4764)
         );
  NAND3_X1 U5665 ( .A1(n6051), .A2(n6461), .A3(n6024), .ZN(n4607) );
  AND2_X1 U5666 ( .A1(n4607), .A2(n4764), .ZN(n4615) );
  INV_X1 U5667 ( .A(n4615), .ZN(n4613) );
  INV_X1 U5668 ( .A(n5957), .ZN(n5427) );
  NAND2_X1 U5669 ( .A1(n6185), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6186) );
  OAI21_X1 U5670 ( .B1(n5427), .B2(n3074), .A(n6186), .ZN(n5425) );
  INV_X1 U5671 ( .A(n5419), .ZN(n4610) );
  OAI21_X1 U5672 ( .B1(n5425), .B2(n4610), .A(n6464), .ZN(n4614) );
  NAND2_X1 U5673 ( .A1(n4611), .A2(n6231), .ZN(n6018) );
  AOI21_X1 U5674 ( .B1(n6271), .B2(n6018), .A(n6191), .ZN(n4612) );
  OAI21_X1 U5675 ( .B1(n4613), .B2(n4614), .A(n4612), .ZN(n4760) );
  OAI22_X1 U5676 ( .A1(n4615), .A2(n4614), .B1(n6367), .B2(n6018), .ZN(n4759)
         );
  AOI22_X1 U5677 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n4760), .B1(n6287), 
        .B2(n4759), .ZN(n4619) );
  NAND2_X1 U5678 ( .A1(n4616), .A2(n5427), .ZN(n4714) );
  NOR2_X2 U5679 ( .A1(n4617), .A2(n5957), .ZN(n6045) );
  AOI22_X1 U5680 ( .A1(n4793), .A2(n6289), .B1(n6045), .B2(n6237), .ZN(n4618)
         );
  OAI211_X1 U5681 ( .C1(n4764), .C2(n4620), .A(n4619), .B(n4618), .ZN(U3045)
         );
  AOI22_X1 U5682 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n4760), .B1(n6299), 
        .B2(n4759), .ZN(n4622) );
  AOI22_X1 U5683 ( .A1(n4793), .A2(n6301), .B1(n6045), .B2(n6245), .ZN(n4621)
         );
  OAI211_X1 U5684 ( .C1(n4764), .C2(n4623), .A(n4622), .B(n4621), .ZN(U3047)
         );
  AOI22_X1 U5685 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n4760), .B1(n6311), 
        .B2(n4759), .ZN(n4625) );
  AOI22_X1 U5686 ( .A1(n4793), .A2(n6313), .B1(n6045), .B2(n6253), .ZN(n4624)
         );
  OAI211_X1 U5687 ( .C1(n4764), .C2(n4626), .A(n4625), .B(n4624), .ZN(U3049)
         );
  AOI22_X1 U5688 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n4760), .B1(n6293), 
        .B2(n4759), .ZN(n4628) );
  AOI22_X1 U5689 ( .A1(n4793), .A2(n6295), .B1(n6045), .B2(n6241), .ZN(n4627)
         );
  OAI211_X1 U5690 ( .C1(n4764), .C2(n4629), .A(n4628), .B(n4627), .ZN(U3046)
         );
  AOI22_X1 U5691 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n4760), .B1(n6324), 
        .B2(n4759), .ZN(n4631) );
  AOI22_X1 U5692 ( .A1(n4793), .A2(n6328), .B1(n6045), .B2(n6264), .ZN(n4630)
         );
  OAI211_X1 U5693 ( .C1(n4764), .C2(n4632), .A(n4631), .B(n4630), .ZN(U3051)
         );
  AOI22_X1 U5694 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n4760), .B1(n6317), 
        .B2(n4759), .ZN(n4634) );
  AOI22_X1 U5695 ( .A1(n4793), .A2(n6319), .B1(n6045), .B2(n6257), .ZN(n4633)
         );
  OAI211_X1 U5696 ( .C1(n4764), .C2(n4635), .A(n4634), .B(n4633), .ZN(U3050)
         );
  NOR2_X2 U5697 ( .A1(n4740), .A2(n5787), .ZN(n6273) );
  INV_X1 U5698 ( .A(n6273), .ZN(n4671) );
  NOR2_X2 U5699 ( .A1(n6603), .A2(n5416), .ZN(n6272) );
  AOI22_X1 U5700 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n4742), .B1(n6272), 
        .B2(n4741), .ZN(n4639) );
  INV_X1 U5701 ( .A(DATAI_24_), .ZN(n4636) );
  NOR2_X1 U5702 ( .A1(n5213), .A2(n4636), .ZN(n6233) );
  INV_X1 U5703 ( .A(DATAI_16_), .ZN(n4637) );
  AOI22_X1 U5704 ( .A1(n6233), .A2(n4792), .B1(n4801), .B2(n6283), .ZN(n4638)
         );
  OAI211_X1 U5705 ( .C1(n4671), .C2(n4747), .A(n4639), .B(n4638), .ZN(U3060)
         );
  INV_X1 U5706 ( .A(n4641), .ZN(n4642) );
  XNOR2_X1 U5707 ( .A(n4640), .B(n4642), .ZN(n5932) );
  NAND2_X1 U5708 ( .A1(n5932), .A2(n5916), .ZN(n4645) );
  AND2_X1 U5709 ( .A1(n5917), .A2(REIP_REG_7__SCAN_IN), .ZN(n5930) );
  NOR2_X1 U5710 ( .A1(n5914), .A2(n5694), .ZN(n4643) );
  AOI211_X1 U5711 ( .C1(n5919), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5930), 
        .B(n4643), .ZN(n4644) );
  OAI211_X1 U5712 ( .C1(n5213), .C2(n5696), .A(n4645), .B(n4644), .ZN(U2979)
         );
  NAND2_X1 U5713 ( .A1(n6312), .A2(n6169), .ZN(n4648) );
  AOI22_X1 U5714 ( .A1(n6253), .A2(n6156), .B1(n6181), .B2(n6313), .ZN(n4647)
         );
  NAND2_X1 U5715 ( .A1(n6170), .A2(n6311), .ZN(n4646) );
  NAND3_X1 U5716 ( .A1(n4648), .A2(n4647), .A3(n4646), .ZN(n4649) );
  AOI21_X1 U5717 ( .B1(n6171), .B2(INSTQUEUE_REG_11__5__SCAN_IN), .A(n4649), 
        .ZN(n4650) );
  INV_X1 U5718 ( .A(n4650), .ZN(U3113) );
  OR2_X1 U5719 ( .A1(n6101), .A2(n6271), .ZN(n6021) );
  NAND2_X1 U5720 ( .A1(n5396), .A2(n5420), .ZN(n5959) );
  NAND2_X1 U5721 ( .A1(n5959), .A2(n6464), .ZN(n4652) );
  NOR2_X2 U5722 ( .A1(n5424), .A2(n5960), .ZN(n6097) );
  INV_X1 U5723 ( .A(n5956), .ZN(n4651) );
  INV_X1 U5724 ( .A(n6125), .ZN(n6126) );
  AOI211_X1 U5725 ( .C1(n6021), .C2(n4652), .A(n6097), .B(n6126), .ZN(n4656)
         );
  NAND3_X1 U5726 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6344), .A3(n6337), .ZN(n6107) );
  NOR2_X1 U5727 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6107), .ZN(n6096)
         );
  AND2_X1 U5728 ( .A1(n4657), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6027) );
  INV_X1 U5729 ( .A(n6027), .ZN(n6221) );
  INV_X1 U5730 ( .A(n4700), .ZN(n4653) );
  OR2_X1 U5731 ( .A1(n4653), .A2(n6138), .ZN(n4683) );
  AOI21_X1 U5732 ( .B1(n4683), .B2(STATE2_REG_2__SCAN_IN), .A(n5416), .ZN(
        n4677) );
  OAI211_X1 U5733 ( .C1(n6458), .C2(n6096), .A(n6221), .B(n4677), .ZN(n4655)
         );
  INV_X1 U5734 ( .A(n5959), .ZN(n6102) );
  NAND2_X1 U5735 ( .A1(n6464), .A2(n6224), .ZN(n6022) );
  NOR2_X1 U5736 ( .A1(n6102), .A2(n6022), .ZN(n4654) );
  INV_X1 U5737 ( .A(n6098), .ZN(n4769) );
  INV_X1 U5738 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4664) );
  INV_X1 U5739 ( .A(n6313), .ZN(n6256) );
  NAND2_X1 U5740 ( .A1(n6101), .A2(n6464), .ZN(n6223) );
  OR2_X1 U5741 ( .A1(n6223), .A2(n5959), .ZN(n4660) );
  NOR2_X1 U5742 ( .A1(n4657), .A2(n6367), .ZN(n6230) );
  INV_X1 U5743 ( .A(n4683), .ZN(n4658) );
  NAND2_X1 U5744 ( .A1(n6230), .A2(n4658), .ZN(n4659) );
  NAND2_X1 U5745 ( .A1(n4660), .A2(n4659), .ZN(n6095) );
  AOI22_X1 U5746 ( .A1(n6097), .A2(n6253), .B1(n6311), .B2(n6095), .ZN(n4661)
         );
  OAI21_X1 U5747 ( .B1(n6125), .B2(n6256), .A(n4661), .ZN(n4662) );
  AOI21_X1 U5748 ( .B1(n6312), .B2(n6096), .A(n4662), .ZN(n4663) );
  OAI21_X1 U5749 ( .B1(n4769), .B2(n4664), .A(n4663), .ZN(U3089) );
  INV_X1 U5750 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4668) );
  INV_X1 U5751 ( .A(n6301), .ZN(n6248) );
  AOI22_X1 U5752 ( .A1(n6097), .A2(n6245), .B1(n6299), .B2(n6095), .ZN(n4665)
         );
  OAI21_X1 U5753 ( .B1(n6125), .B2(n6248), .A(n4665), .ZN(n4666) );
  AOI21_X1 U5754 ( .B1(n6300), .B2(n6096), .A(n4666), .ZN(n4667) );
  OAI21_X1 U5755 ( .B1(n4769), .B2(n4668), .A(n4667), .ZN(U3087) );
  AOI22_X1 U5756 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n4760), .B1(n6272), 
        .B2(n4759), .ZN(n4670) );
  AOI22_X1 U5757 ( .A1(n4793), .A2(n6283), .B1(n6045), .B2(n6233), .ZN(n4669)
         );
  OAI211_X1 U5758 ( .C1(n4764), .C2(n4671), .A(n4670), .B(n4669), .ZN(U3044)
         );
  NAND2_X1 U5759 ( .A1(n6273), .A2(n6169), .ZN(n4674) );
  AOI22_X1 U5760 ( .A1(n6233), .A2(n6156), .B1(n6181), .B2(n6283), .ZN(n4673)
         );
  NAND2_X1 U5761 ( .A1(n6170), .A2(n6272), .ZN(n4672) );
  NAND3_X1 U5762 ( .A1(n4674), .A2(n4673), .A3(n4672), .ZN(n4675) );
  AOI21_X1 U5763 ( .B1(n6171), .B2(INSTQUEUE_REG_11__0__SCAN_IN), .A(n4675), 
        .ZN(n4676) );
  INV_X1 U5764 ( .A(n4676), .ZN(U3108) );
  NAND3_X1 U5765 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6337), .ZN(n6194) );
  NOR2_X1 U5766 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6194), .ZN(n6180)
         );
  INV_X1 U5767 ( .A(n6230), .ZN(n6139) );
  OAI211_X1 U5768 ( .C1(n6458), .C2(n6180), .A(n6139), .B(n4677), .ZN(n4678)
         );
  INV_X1 U5769 ( .A(n4678), .ZN(n4682) );
  INV_X1 U5770 ( .A(n4679), .ZN(n5405) );
  NAND2_X1 U5771 ( .A1(n6185), .A2(n3581), .ZN(n6211) );
  OAI21_X1 U5772 ( .B1(n6212), .B2(n6181), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4680) );
  OAI211_X1 U5773 ( .C1(n5405), .C2(n6187), .A(n4680), .B(n6464), .ZN(n4681)
         );
  NAND2_X1 U5774 ( .A1(n4682), .A2(n4681), .ZN(n6182) );
  INV_X1 U5775 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4686) );
  OAI22_X1 U5776 ( .A1(n6223), .A2(n6187), .B1(n6221), .B2(n4683), .ZN(n6179)
         );
  AOI22_X1 U5777 ( .A1(n6181), .A2(n6245), .B1(n6299), .B2(n6179), .ZN(n4685)
         );
  AOI22_X1 U5778 ( .A1(n6300), .A2(n6180), .B1(n6301), .B2(n6212), .ZN(n4684)
         );
  OAI211_X1 U5779 ( .C1(n4773), .C2(n4686), .A(n4685), .B(n4684), .ZN(U3119)
         );
  INV_X1 U5780 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4689) );
  AOI22_X1 U5781 ( .A1(n6181), .A2(n6264), .B1(n6324), .B2(n6179), .ZN(n4688)
         );
  AOI22_X1 U5782 ( .A1(n6326), .A2(n6180), .B1(n6328), .B2(n6212), .ZN(n4687)
         );
  OAI211_X1 U5783 ( .C1(n4773), .C2(n4689), .A(n4688), .B(n4687), .ZN(U3123)
         );
  INV_X1 U5784 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4692) );
  AOI22_X1 U5785 ( .A1(n6181), .A2(n6253), .B1(n6311), .B2(n6179), .ZN(n4691)
         );
  AOI22_X1 U5786 ( .A1(n6312), .A2(n6180), .B1(n6313), .B2(n6212), .ZN(n4690)
         );
  OAI211_X1 U5787 ( .C1(n4773), .C2(n4692), .A(n4691), .B(n4690), .ZN(U3121)
         );
  INV_X1 U5788 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4695) );
  AOI22_X1 U5789 ( .A1(n6181), .A2(n6257), .B1(n6317), .B2(n6179), .ZN(n4694)
         );
  AOI22_X1 U5790 ( .A1(n6318), .A2(n6180), .B1(n6319), .B2(n6212), .ZN(n4693)
         );
  OAI211_X1 U5791 ( .C1(n4773), .C2(n4695), .A(n4694), .B(n4693), .ZN(U3122)
         );
  NOR2_X1 U5792 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4696), .ZN(n4794)
         );
  INV_X1 U5793 ( .A(n4792), .ZN(n4697) );
  AOI21_X1 U5794 ( .B1(n4697), .B2(n4714), .A(n6224), .ZN(n4699) );
  NOR2_X1 U5795 ( .A1(n4699), .A2(n4698), .ZN(n4702) );
  OR2_X1 U5796 ( .A1(n6138), .A2(n4700), .ZN(n5958) );
  INV_X1 U5797 ( .A(n5958), .ZN(n4701) );
  OAI21_X1 U5798 ( .B1(n4701), .B2(n6367), .A(n4803), .ZN(n5963) );
  AOI211_X1 U5799 ( .C1(n6464), .C2(n4702), .A(n6230), .B(n5963), .ZN(n4703)
         );
  OAI21_X1 U5800 ( .B1(n4794), .B2(n6458), .A(n4703), .ZN(n4704) );
  INV_X1 U5801 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4708) );
  INV_X1 U5802 ( .A(n6237), .ZN(n6292) );
  OAI22_X1 U5803 ( .A1(n6021), .A2(n6187), .B1(n6221), .B2(n5958), .ZN(n4791)
         );
  AOI22_X1 U5804 ( .A1(n4792), .A2(n6289), .B1(n6287), .B2(n4791), .ZN(n4705)
         );
  OAI21_X1 U5805 ( .B1(n4714), .B2(n6292), .A(n4705), .ZN(n4706) );
  AOI21_X1 U5806 ( .B1(n6288), .B2(n4794), .A(n4706), .ZN(n4707) );
  OAI21_X1 U5807 ( .B1(n4798), .B2(n4708), .A(n4707), .ZN(U3053) );
  INV_X1 U5808 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4712) );
  INV_X1 U5809 ( .A(n6233), .ZN(n6286) );
  AOI22_X1 U5810 ( .A1(n4792), .A2(n6283), .B1(n6272), .B2(n4791), .ZN(n4709)
         );
  OAI21_X1 U5811 ( .B1(n6286), .B2(n4714), .A(n4709), .ZN(n4710) );
  AOI21_X1 U5812 ( .B1(n6273), .B2(n4794), .A(n4710), .ZN(n4711) );
  OAI21_X1 U5813 ( .B1(n4798), .B2(n4712), .A(n4711), .ZN(U3052) );
  INV_X1 U5814 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4717) );
  AOI22_X1 U5815 ( .A1(n4792), .A2(n6301), .B1(n6299), .B2(n4791), .ZN(n4713)
         );
  OAI21_X1 U5816 ( .B1(n4714), .B2(n6304), .A(n4713), .ZN(n4715) );
  AOI21_X1 U5817 ( .B1(n6300), .B2(n4794), .A(n4715), .ZN(n4716) );
  OAI21_X1 U5818 ( .B1(n4798), .B2(n4717), .A(n4716), .ZN(U3055) );
  INV_X1 U5819 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4720) );
  AOI22_X1 U5820 ( .A1(n4792), .A2(n6328), .B1(n6324), .B2(n4791), .ZN(n4719)
         );
  AOI22_X1 U5821 ( .A1(n6326), .A2(n4794), .B1(n4793), .B2(n6264), .ZN(n4718)
         );
  OAI211_X1 U5822 ( .C1(n4798), .C2(n4720), .A(n4719), .B(n4718), .ZN(U3059)
         );
  INV_X1 U5823 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4723) );
  AOI22_X1 U5824 ( .A1(n4792), .A2(n6313), .B1(n6311), .B2(n4791), .ZN(n4722)
         );
  AOI22_X1 U5825 ( .A1(n6312), .A2(n4794), .B1(n4793), .B2(n6253), .ZN(n4721)
         );
  OAI211_X1 U5826 ( .C1(n4798), .C2(n4723), .A(n4722), .B(n4721), .ZN(U3057)
         );
  INV_X1 U5827 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4726) );
  AOI22_X1 U5828 ( .A1(n4792), .A2(n6319), .B1(n6317), .B2(n4791), .ZN(n4725)
         );
  AOI22_X1 U5829 ( .A1(n6318), .A2(n4794), .B1(n4793), .B2(n6257), .ZN(n4724)
         );
  OAI211_X1 U5830 ( .C1(n4798), .C2(n4726), .A(n4725), .B(n4724), .ZN(U3058)
         );
  INV_X1 U5831 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4729) );
  AOI22_X1 U5832 ( .A1(n4792), .A2(n6295), .B1(n6293), .B2(n4791), .ZN(n4728)
         );
  AOI22_X1 U5833 ( .A1(n6294), .A2(n4794), .B1(n4793), .B2(n6241), .ZN(n4727)
         );
  OAI211_X1 U5834 ( .C1(n4798), .C2(n4729), .A(n4728), .B(n4727), .ZN(U3054)
         );
  INV_X1 U5835 ( .A(DATAI_8_), .ZN(n5878) );
  INV_X1 U5836 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6620) );
  OAI222_X1 U5837 ( .A1(n4845), .A2(n5507), .B1(n5152), .B2(n5878), .C1(n5151), 
        .C2(n6620), .ZN(U2883) );
  INV_X1 U5838 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4730) );
  OAI222_X1 U5839 ( .A1(n4845), .A2(n5126), .B1(n5776), .B2(n4730), .C1(n5122), 
        .C2(n4778), .ZN(U2851) );
  NAND2_X1 U5840 ( .A1(n4974), .A2(n4731), .ZN(n4732) );
  INV_X1 U5841 ( .A(n5767), .ZN(n5715) );
  NAND2_X1 U5842 ( .A1(n5715), .A2(n5272), .ZN(n4734) );
  AOI22_X1 U5843 ( .A1(n5764), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n5723), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4733) );
  OAI211_X1 U5844 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n5738), .A(n4734), 
        .B(n4733), .ZN(n4739) );
  OAI22_X1 U5845 ( .A1(n4332), .A2(n5671), .B1(n5754), .B2(REIP_REG_1__SCAN_IN), .ZN(n4738) );
  NAND2_X1 U5846 ( .A1(n4974), .A2(n4735), .ZN(n5759) );
  OAI22_X1 U5847 ( .A1(n5761), .A2(n4736), .B1(n5396), .B2(n5759), .ZN(n4737)
         );
  OR3_X1 U5848 ( .A1(n4739), .A2(n4738), .A3(n4737), .ZN(U2826) );
  NOR2_X2 U5849 ( .A1(n4740), .A2(n3306), .ZN(n6306) );
  INV_X1 U5850 ( .A(n6306), .ZN(n4763) );
  NOR2_X2 U5851 ( .A1(n5870), .A2(n5416), .ZN(n6305) );
  AOI22_X1 U5852 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4742), .B1(n6305), 
        .B2(n4741), .ZN(n4746) );
  INV_X1 U5853 ( .A(DATAI_28_), .ZN(n4743) );
  NOR2_X1 U5854 ( .A1(n5213), .A2(n4743), .ZN(n6249) );
  INV_X1 U5855 ( .A(DATAI_20_), .ZN(n4744) );
  NOR2_X2 U5856 ( .A1(n5213), .A2(n4744), .ZN(n6307) );
  AOI22_X1 U5857 ( .A1(n6249), .A2(n4792), .B1(n4801), .B2(n6307), .ZN(n4745)
         );
  OAI211_X1 U5858 ( .C1(n4763), .C2(n4747), .A(n4746), .B(n4745), .ZN(U3064)
         );
  XNOR2_X1 U5859 ( .A(n3071), .B(n4749), .ZN(n4856) );
  INV_X1 U5860 ( .A(n4752), .ZN(n4779) );
  OAI21_X1 U5861 ( .B1(n5343), .B2(n4779), .A(n2998), .ZN(n4870) );
  NAND2_X1 U5862 ( .A1(n4751), .A2(n4750), .ZN(n5935) );
  NOR2_X1 U5863 ( .A1(n4752), .A2(n5935), .ZN(n4868) );
  AOI22_X1 U5864 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n4870), .B1(n4868), 
        .B2(n4753), .ZN(n4758) );
  AOI21_X1 U5865 ( .B1(n4756), .B2(n4755), .A(n4754), .ZN(n5686) );
  AND2_X1 U5866 ( .A1(n5917), .A2(REIP_REG_9__SCAN_IN), .ZN(n4852) );
  AOI21_X1 U5867 ( .B1(n5686), .B2(n5944), .A(n4852), .ZN(n4757) );
  OAI211_X1 U5868 ( .C1(n4856), .C2(n5394), .A(n4758), .B(n4757), .ZN(U3009)
         );
  AOI22_X1 U5869 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n4760), .B1(n6305), 
        .B2(n4759), .ZN(n4762) );
  AOI22_X1 U5870 ( .A1(n4793), .A2(n6307), .B1(n6045), .B2(n6249), .ZN(n4761)
         );
  OAI211_X1 U5871 ( .C1(n4764), .C2(n4763), .A(n4762), .B(n4761), .ZN(U3048)
         );
  INV_X1 U5872 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4768) );
  INV_X1 U5873 ( .A(n6307), .ZN(n6252) );
  AOI22_X1 U5874 ( .A1(n6097), .A2(n6249), .B1(n6305), .B2(n6095), .ZN(n4765)
         );
  OAI21_X1 U5875 ( .B1(n6125), .B2(n6252), .A(n4765), .ZN(n4766) );
  AOI21_X1 U5876 ( .B1(n6306), .B2(n6096), .A(n4766), .ZN(n4767) );
  OAI21_X1 U5877 ( .B1(n4769), .B2(n4768), .A(n4767), .ZN(U3088) );
  INV_X1 U5878 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4772) );
  AOI22_X1 U5879 ( .A1(n6181), .A2(n6249), .B1(n6305), .B2(n6179), .ZN(n4771)
         );
  AOI22_X1 U5880 ( .A1(n6306), .A2(n6180), .B1(n6307), .B2(n6212), .ZN(n4770)
         );
  OAI211_X1 U5881 ( .C1(n4773), .C2(n4772), .A(n4771), .B(n4770), .ZN(U3120)
         );
  XOR2_X1 U5882 ( .A(n3070), .B(n4775), .Z(n4844) );
  INV_X1 U5883 ( .A(n2998), .ZN(n4776) );
  AOI22_X1 U5884 ( .A1(n5917), .A2(REIP_REG_8__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n4776), .ZN(n4777) );
  OAI21_X1 U5885 ( .B1(n6688), .B2(n4778), .A(n4777), .ZN(n4782) );
  AOI211_X1 U5886 ( .C1(n4780), .C2(n5938), .A(n4779), .B(n5935), .ZN(n4781)
         );
  AOI211_X1 U5887 ( .C1(n4844), .C2(n5951), .A(n4782), .B(n4781), .ZN(n4783)
         );
  INV_X1 U5888 ( .A(n4783), .ZN(U3010) );
  NOR2_X1 U5889 ( .A1(n5759), .A2(n5420), .ZN(n4788) );
  INV_X1 U5890 ( .A(n5913), .ZN(n4784) );
  AOI22_X1 U5891 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n5764), .B1(n5763), 
        .B2(n4784), .ZN(n4785) );
  OAI21_X1 U5892 ( .B1(n5671), .B2(n4786), .A(n4785), .ZN(n4787) );
  AOI211_X1 U5893 ( .C1(n5743), .C2(EBX_REG_2__SCAN_IN), .A(n4788), .B(n4787), 
        .ZN(n4790) );
  OAI211_X1 U5894 ( .C1(REIP_REG_1__SCAN_IN), .C2(n5754), .A(
        REIP_REG_2__SCAN_IN), .B(n5755), .ZN(n5752) );
  OAI221_X1 U5895 ( .B1(REIP_REG_2__SCAN_IN), .B2(REIP_REG_1__SCAN_IN), .C1(
        REIP_REG_2__SCAN_IN), .C2(n5724), .A(n5752), .ZN(n4789) );
  OAI211_X1 U5896 ( .C1(n5767), .C2(n5903), .A(n4790), .B(n4789), .ZN(U2825)
         );
  INV_X1 U5897 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4797) );
  AOI22_X1 U5898 ( .A1(n4792), .A2(n6307), .B1(n6305), .B2(n4791), .ZN(n4796)
         );
  AOI22_X1 U5899 ( .A1(n6306), .A2(n4794), .B1(n4793), .B2(n6249), .ZN(n4795)
         );
  OAI211_X1 U5900 ( .C1(n4798), .C2(n4797), .A(n4796), .B(n4795), .ZN(U3056)
         );
  XOR2_X1 U5901 ( .A(n4799), .B(n4348), .Z(n5689) );
  INV_X1 U5902 ( .A(n5689), .ZN(n4857) );
  AOI22_X1 U5903 ( .A1(n5686), .A2(n4194), .B1(EBX_REG_9__SCAN_IN), .B2(n5103), 
        .ZN(n4800) );
  OAI21_X1 U5904 ( .B1(n4857), .B2(n5126), .A(n4800), .ZN(U2850) );
  OR2_X1 U5905 ( .A1(n5424), .A2(n6218), .ZN(n4808) );
  AOI21_X1 U5906 ( .B1(n4838), .B2(n4808), .A(n6224), .ZN(n4805) );
  NAND2_X1 U5907 ( .A1(n4802), .A2(n4426), .ZN(n6222) );
  NAND2_X1 U5908 ( .A1(n6222), .A2(n6464), .ZN(n6227) );
  NAND2_X1 U5909 ( .A1(n6468), .A2(n6058), .ZN(n4807) );
  OAI21_X1 U5910 ( .B1(n6138), .B2(n6367), .A(n4803), .ZN(n6228) );
  AOI211_X1 U5911 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4807), .A(n6230), .B(
        n6228), .ZN(n4804) );
  OAI211_X1 U5912 ( .C1(n4805), .C2(n6227), .A(n4804), .B(n6231), .ZN(n4806)
         );
  INV_X1 U5913 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4812) );
  INV_X1 U5914 ( .A(n4807), .ZN(n4840) );
  INV_X1 U5915 ( .A(n6241), .ZN(n6298) );
  NAND2_X1 U5916 ( .A1(n6138), .A2(n6231), .ZN(n6019) );
  OAI22_X1 U5917 ( .A1(n6021), .A2(n6222), .B1(n6221), .B2(n6019), .ZN(n4836)
         );
  AOI22_X1 U5918 ( .A1(n6080), .A2(n6295), .B1(n6293), .B2(n4836), .ZN(n4809)
         );
  OAI21_X1 U5919 ( .B1(n4838), .B2(n6298), .A(n4809), .ZN(n4810) );
  AOI21_X1 U5920 ( .B1(n6294), .B2(n4840), .A(n4810), .ZN(n4811) );
  OAI21_X1 U5921 ( .B1(n4843), .B2(n4812), .A(n4811), .ZN(U3070) );
  INV_X1 U5922 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n6653) );
  INV_X1 U5923 ( .A(n6253), .ZN(n6316) );
  AOI22_X1 U5924 ( .A1(n6080), .A2(n6313), .B1(n6311), .B2(n4836), .ZN(n4813)
         );
  OAI21_X1 U5925 ( .B1(n4838), .B2(n6316), .A(n4813), .ZN(n4814) );
  AOI21_X1 U5926 ( .B1(n6312), .B2(n4840), .A(n4814), .ZN(n4815) );
  OAI21_X1 U5927 ( .B1(n4843), .B2(n6653), .A(n4815), .ZN(U3073) );
  INV_X1 U5928 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4819) );
  AOI22_X1 U5929 ( .A1(n6080), .A2(n6283), .B1(n6272), .B2(n4836), .ZN(n4816)
         );
  OAI21_X1 U5930 ( .B1(n4838), .B2(n6286), .A(n4816), .ZN(n4817) );
  AOI21_X1 U5931 ( .B1(n6273), .B2(n4840), .A(n4817), .ZN(n4818) );
  OAI21_X1 U5932 ( .B1(n4843), .B2(n4819), .A(n4818), .ZN(U3068) );
  INV_X1 U5933 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4823) );
  INV_X1 U5934 ( .A(n6257), .ZN(n6322) );
  AOI22_X1 U5935 ( .A1(n6080), .A2(n6319), .B1(n6317), .B2(n4836), .ZN(n4820)
         );
  OAI21_X1 U5936 ( .B1(n4838), .B2(n6322), .A(n4820), .ZN(n4821) );
  AOI21_X1 U5937 ( .B1(n6318), .B2(n4840), .A(n4821), .ZN(n4822) );
  OAI21_X1 U5938 ( .B1(n4843), .B2(n4823), .A(n4822), .ZN(U3074) );
  INV_X1 U5939 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4827) );
  AOI22_X1 U5940 ( .A1(n6080), .A2(n6301), .B1(n6299), .B2(n4836), .ZN(n4824)
         );
  OAI21_X1 U5941 ( .B1(n4838), .B2(n6304), .A(n4824), .ZN(n4825) );
  AOI21_X1 U5942 ( .B1(n6300), .B2(n4840), .A(n4825), .ZN(n4826) );
  OAI21_X1 U5943 ( .B1(n4843), .B2(n4827), .A(n4826), .ZN(U3071) );
  INV_X1 U5944 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4831) );
  INV_X1 U5945 ( .A(n6264), .ZN(n6333) );
  AOI22_X1 U5946 ( .A1(n6080), .A2(n6328), .B1(n6324), .B2(n4836), .ZN(n4828)
         );
  OAI21_X1 U5947 ( .B1(n4838), .B2(n6333), .A(n4828), .ZN(n4829) );
  AOI21_X1 U5948 ( .B1(n6326), .B2(n4840), .A(n4829), .ZN(n4830) );
  OAI21_X1 U5949 ( .B1(n4843), .B2(n4831), .A(n4830), .ZN(U3075) );
  INV_X1 U5950 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4835) );
  INV_X1 U5951 ( .A(n6249), .ZN(n6310) );
  AOI22_X1 U5952 ( .A1(n6080), .A2(n6307), .B1(n6305), .B2(n4836), .ZN(n4832)
         );
  OAI21_X1 U5953 ( .B1(n4838), .B2(n6310), .A(n4832), .ZN(n4833) );
  AOI21_X1 U5954 ( .B1(n6306), .B2(n4840), .A(n4833), .ZN(n4834) );
  OAI21_X1 U5955 ( .B1(n4843), .B2(n4835), .A(n4834), .ZN(U3072) );
  INV_X1 U5956 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4842) );
  AOI22_X1 U5957 ( .A1(n6080), .A2(n6289), .B1(n6287), .B2(n4836), .ZN(n4837)
         );
  OAI21_X1 U5958 ( .B1(n4838), .B2(n6292), .A(n4837), .ZN(n4839) );
  AOI21_X1 U5959 ( .B1(n6288), .B2(n4840), .A(n4839), .ZN(n4841) );
  OAI21_X1 U5960 ( .B1(n4843), .B2(n4842), .A(n4841), .ZN(U3069) );
  INV_X1 U5961 ( .A(n4844), .ZN(n4851) );
  INV_X1 U5962 ( .A(n4845), .ZN(n4849) );
  AOI22_X1 U5963 ( .A1(n5919), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n5917), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n4846) );
  OAI21_X1 U5964 ( .B1(n5914), .B2(n4847), .A(n4846), .ZN(n4848) );
  AOI21_X1 U5965 ( .B1(n4849), .B2(n5909), .A(n4848), .ZN(n4850) );
  OAI21_X1 U5966 ( .B1(n4851), .B2(n3056), .A(n4850), .ZN(U2978) );
  AOI21_X1 U5967 ( .B1(n5919), .B2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n4852), 
        .ZN(n4853) );
  OAI21_X1 U5968 ( .B1(n5687), .B2(n5914), .A(n4853), .ZN(n4854) );
  AOI21_X1 U5969 ( .B1(n5689), .B2(n5909), .A(n4854), .ZN(n4855) );
  OAI21_X1 U5970 ( .B1(n4856), .B2(n3056), .A(n4855), .ZN(U2977) );
  INV_X1 U5971 ( .A(DATAI_9_), .ZN(n5880) );
  INV_X1 U5972 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6670) );
  OAI222_X1 U5973 ( .A1(n5507), .A2(n4857), .B1(n5152), .B2(n5880), .C1(n5151), 
        .C2(n6670), .ZN(U2882) );
  NOR2_X1 U5974 ( .A1(n4860), .A2(n4859), .ZN(n4861) );
  OR2_X1 U5975 ( .A1(n4858), .A2(n4861), .ZN(n5673) );
  INV_X1 U5976 ( .A(DATAI_10_), .ZN(n5882) );
  INV_X1 U5977 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5819) );
  OAI222_X1 U5978 ( .A1(n5673), .A2(n5507), .B1(n5152), .B2(n5882), .C1(n5151), 
        .C2(n5819), .ZN(U2881) );
  OAI21_X1 U5979 ( .B1(n4754), .B2(n4862), .A(n4876), .ZN(n5670) );
  OAI222_X1 U5980 ( .A1(n5673), .A2(n5126), .B1(n5776), .B2(n4863), .C1(n5122), 
        .C2(n5670), .ZN(U2849) );
  NAND2_X1 U5981 ( .A1(n5254), .A2(n4864), .ZN(n4866) );
  XOR2_X1 U5982 ( .A(n4866), .B(n4865), .Z(n5269) );
  OAI211_X1 U5983 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A(n4868), .B(n4867), .ZN(n4872) );
  INV_X1 U5984 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6417) );
  OAI22_X1 U5985 ( .A1(n5670), .A2(n6688), .B1(n6417), .B2(n6684), .ZN(n4869)
         );
  AOI21_X1 U5986 ( .B1(n4870), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n4869), 
        .ZN(n4871) );
  OAI211_X1 U5987 ( .C1(n5269), .C2(n5394), .A(n4872), .B(n4871), .ZN(U3008)
         );
  NOR2_X1 U5988 ( .A1(n4858), .A2(n4873), .ZN(n4874) );
  OR2_X1 U5989 ( .A1(n4890), .A2(n4874), .ZN(n5264) );
  AOI21_X1 U5990 ( .B1(n4877), .B2(n4876), .A(n4875), .ZN(n5924) );
  AOI22_X1 U5991 ( .A1(n5924), .A2(n4194), .B1(EBX_REG_11__SCAN_IN), .B2(n5103), .ZN(n4878) );
  OAI21_X1 U5992 ( .B1(n5264), .B2(n5126), .A(n4878), .ZN(U2848) );
  AOI22_X1 U5993 ( .A1(n5148), .A2(DATAI_11_), .B1(n5783), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n4879) );
  OAI21_X1 U5994 ( .B1(n5264), .B2(n5507), .A(n4879), .ZN(U2880) );
  INV_X1 U5995 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6416) );
  NAND2_X1 U5996 ( .A1(n5724), .A2(n4880), .ZN(n5676) );
  NOR2_X1 U5997 ( .A1(n6416), .A2(n5676), .ZN(n5668) );
  INV_X1 U5998 ( .A(n4881), .ZN(n4882) );
  OAI21_X1 U5999 ( .B1(n4882), .B2(n5754), .A(n5755), .ZN(n5659) );
  OAI221_X1 U6000 ( .B1(REIP_REG_11__SCAN_IN), .B2(REIP_REG_10__SCAN_IN), .C1(
        REIP_REG_11__SCAN_IN), .C2(n5668), .A(n5659), .ZN(n4887) );
  INV_X1 U6001 ( .A(n5260), .ZN(n4885) );
  AOI22_X1 U6002 ( .A1(EBX_REG_11__SCAN_IN), .A2(n5743), .B1(n5758), .B2(n5924), .ZN(n4883) );
  OAI211_X1 U6003 ( .C1(n5683), .C2(n3692), .A(n4883), .B(n5712), .ZN(n4884)
         );
  AOI21_X1 U6004 ( .B1(n5763), .B2(n4885), .A(n4884), .ZN(n4886) );
  OAI211_X1 U6005 ( .C1(n5264), .C2(n5695), .A(n4887), .B(n4886), .ZN(U2816)
         );
  OAI21_X1 U6006 ( .B1(n4890), .B2(n4889), .A(n4888), .ZN(n5665) );
  OAI21_X1 U6007 ( .B1(n4875), .B2(n4891), .A(n5042), .ZN(n5658) );
  OAI222_X1 U6008 ( .A1(n5665), .A2(n5126), .B1(n5776), .B2(n5661), .C1(n5122), 
        .C2(n5658), .ZN(U2847) );
  INV_X1 U6009 ( .A(DATAI_12_), .ZN(n4892) );
  OAI222_X1 U6010 ( .A1(n5665), .A2(n5507), .B1(n5151), .B2(n4893), .C1(n5152), 
        .C2(n4892), .ZN(U2879) );
  AOI22_X1 U6011 ( .A1(n4897), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n4896), .B2(EBX_REG_31__SCAN_IN), .ZN(n4898) );
  INV_X1 U6012 ( .A(n4983), .ZN(n5053) );
  NOR2_X1 U6013 ( .A1(n4941), .A2(n5281), .ZN(n4903) );
  NOR3_X1 U6014 ( .A1(n4901), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4902) );
  AOI22_X1 U6015 ( .A1(n4939), .A2(n4903), .B1(n5524), .B2(n4902), .ZN(n4904)
         );
  XNOR2_X1 U6016 ( .A(n4904), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4961)
         );
  NAND2_X1 U6017 ( .A1(n4961), .A2(n5951), .ZN(n4919) );
  INV_X1 U6018 ( .A(n4914), .ZN(n4908) );
  NAND2_X1 U6019 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5306) );
  INV_X1 U6020 ( .A(n5948), .ZN(n4905) );
  NOR2_X1 U6021 ( .A1(n4905), .A2(n5342), .ZN(n5386) );
  OAI21_X1 U6022 ( .B1(n4907), .B2(n5386), .A(n4906), .ZN(n5558) );
  OAI21_X1 U6023 ( .B1(n4908), .B2(n5343), .A(n5300), .ZN(n4943) );
  OAI21_X1 U6024 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5343), .A(n5282), 
        .ZN(n4917) );
  INV_X1 U6025 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6450) );
  NOR2_X1 U6026 ( .A1(n6684), .A2(n6450), .ZN(n4957) );
  INV_X1 U6027 ( .A(n4909), .ZN(n4910) );
  NAND2_X1 U6028 ( .A1(n4911), .A2(n4910), .ZN(n6686) );
  NOR2_X1 U6029 ( .A1(n6686), .A2(n4912), .ZN(n5560) );
  INV_X1 U6030 ( .A(n5306), .ZN(n4913) );
  NAND2_X1 U6031 ( .A1(n5560), .A2(n4913), .ZN(n5289) );
  NOR2_X1 U6032 ( .A1(n5289), .A2(n4914), .ZN(n5278) );
  AND4_X1 U6033 ( .A1(n5278), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n4915), .ZN(n4916) );
  AOI211_X1 U6034 ( .C1(n4917), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n4957), .B(n4916), .ZN(n4918) );
  OAI211_X1 U6035 ( .C1(n5053), .C2(n6688), .A(n4919), .B(n4918), .ZN(U2987)
         );
  XNOR2_X1 U6036 ( .A(n4427), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4925)
         );
  XNOR2_X1 U6037 ( .A(n4920), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4921)
         );
  NAND2_X1 U6038 ( .A1(n5429), .A2(n4921), .ZN(n4922) );
  OAI21_X1 U6039 ( .B1(n4925), .B2(n4923), .A(n4922), .ZN(n4924) );
  AOI21_X1 U6040 ( .B1(n4926), .B2(n4925), .A(n4924), .ZN(n4927) );
  OAI21_X1 U6041 ( .B1(n5420), .B2(n4928), .A(n4927), .ZN(n5397) );
  NOR3_X1 U6042 ( .A1(n6376), .A2(n4930), .A3(n4929), .ZN(n4933) );
  INV_X1 U6043 ( .A(n4427), .ZN(n4934) );
  NOR3_X1 U6044 ( .A1(n4934), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n4931), 
        .ZN(n4932) );
  AOI211_X1 U6045 ( .C1(n5397), .C2(n5597), .A(n4933), .B(n4932), .ZN(n4937)
         );
  AOI21_X1 U6046 ( .B1(n4934), .B2(n6366), .A(n4936), .ZN(n4935) );
  OAI22_X1 U6047 ( .A1(n4937), .A2(n4936), .B1(n4935), .B2(n3321), .ZN(U3459)
         );
  OAI222_X1 U6048 ( .A1(n5133), .A2(n5126), .B1(n4938), .B2(n5776), .C1(n4946), 
        .C2(n5122), .ZN(U2830) );
  NOR2_X1 U6049 ( .A1(n4939), .A2(n4940), .ZN(n4942) );
  XNOR2_X1 U6050 ( .A(n4942), .B(n4941), .ZN(n5159) );
  INV_X1 U6051 ( .A(n4943), .ZN(n4948) );
  INV_X1 U6052 ( .A(n5278), .ZN(n4944) );
  NAND2_X1 U6053 ( .A1(n5917), .A2(REIP_REG_29__SCAN_IN), .ZN(n5154) );
  OAI21_X1 U6054 ( .B1(n4944), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5154), 
        .ZN(n4945) );
  INV_X1 U6055 ( .A(n4945), .ZN(n4947) );
  INV_X1 U6056 ( .A(n4949), .ZN(n4950) );
  OAI21_X1 U6057 ( .B1(n5159), .B2(n5394), .A(n4950), .ZN(U2989) );
  NAND2_X1 U6058 ( .A1(n4952), .A2(n4951), .ZN(n4956) );
  AOI22_X1 U6059 ( .A1(n4954), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n4953), .ZN(n4955) );
  XNOR2_X1 U6060 ( .A(n4956), .B(n4955), .ZN(n5130) );
  AOI21_X1 U6061 ( .B1(n5919), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n4957), 
        .ZN(n4958) );
  OAI21_X1 U6062 ( .B1(n5914), .B2(n4959), .A(n4958), .ZN(n4960) );
  AOI21_X1 U6063 ( .B1(n4961), .B2(n5916), .A(n4960), .ZN(n4962) );
  OAI21_X1 U6064 ( .B1(n5130), .B2(n6275), .A(n4962), .ZN(U2955) );
  INV_X1 U6065 ( .A(n4977), .ZN(n4963) );
  NAND2_X1 U6066 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .ZN(
        n4976) );
  AOI21_X1 U6067 ( .B1(n4963), .B2(n4976), .A(n4994), .ZN(n4981) );
  AOI21_X1 U6068 ( .B1(n4963), .B2(REIP_REG_29__SCAN_IN), .A(
        REIP_REG_30__SCAN_IN), .ZN(n4967) );
  AOI22_X1 U6069 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n5764), .B1(n5763), 
        .B2(n4964), .ZN(n4966) );
  NAND2_X1 U6070 ( .A1(n5743), .A2(EBX_REG_30__SCAN_IN), .ZN(n4965) );
  OAI211_X1 U6071 ( .C1(n4981), .C2(n4967), .A(n4966), .B(n4965), .ZN(n4968)
         );
  AOI21_X1 U6072 ( .B1(n3086), .B2(n5758), .A(n4968), .ZN(n4969) );
  OAI21_X1 U6073 ( .B1(n3069), .B2(n5695), .A(n4969), .ZN(U2797) );
  AOI22_X1 U6074 ( .A1(n5780), .A2(DATAI_30_), .B1(n5783), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n4973) );
  NOR3_X1 U6075 ( .A1(n5783), .A2(n5127), .A3(n4970), .ZN(n4971) );
  NAND2_X1 U6076 ( .A1(n5784), .A2(DATAI_14_), .ZN(n4972) );
  OAI211_X1 U6077 ( .C1(n3069), .C2(n5507), .A(n4973), .B(n4972), .ZN(U2861)
         );
  INV_X1 U6078 ( .A(n4974), .ZN(n4975) );
  NOR4_X1 U6079 ( .A1(n4975), .A2(n6363), .A3(n6485), .A4(n5052), .ZN(n4979)
         );
  NOR3_X1 U6080 ( .A1(n4977), .A2(REIP_REG_31__SCAN_IN), .A3(n4976), .ZN(n4978) );
  AOI211_X1 U6081 ( .C1(PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n5764), .A(n4979), 
        .B(n4978), .ZN(n4980) );
  OAI21_X1 U6082 ( .B1(n4981), .B2(n6450), .A(n4980), .ZN(n4982) );
  AOI21_X1 U6083 ( .B1(n4983), .B2(n5758), .A(n4982), .ZN(n4984) );
  INV_X1 U6084 ( .A(n4986), .ZN(n4987) );
  AOI21_X1 U6085 ( .B1(n4988), .B2(n5058), .A(n4987), .ZN(n5167) );
  INV_X1 U6086 ( .A(n5167), .ZN(n5136) );
  NAND3_X1 U6087 ( .A1(n5438), .A2(REIP_REG_27__SCAN_IN), .A3(n6514), .ZN(
        n4990) );
  AOI22_X1 U6088 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n5764), .B1(n5763), 
        .B2(n5164), .ZN(n4989) );
  OAI211_X1 U6089 ( .C1(n5054), .C2(n5761), .A(n4990), .B(n4989), .ZN(n4993)
         );
  OAI21_X1 U6090 ( .B1(n5061), .B2(n4991), .A(n4216), .ZN(n5286) );
  NOR2_X1 U6091 ( .A1(n5286), .A2(n5671), .ZN(n4992) );
  AOI211_X1 U6092 ( .C1(REIP_REG_28__SCAN_IN), .C2(n4994), .A(n4993), .B(n4992), .ZN(n4995) );
  OAI21_X1 U6093 ( .B1(n5136), .B2(n5695), .A(n4995), .ZN(U2799) );
  NAND2_X1 U6094 ( .A1(n4997), .A2(n4998), .ZN(n5098) );
  XNOR2_X1 U6095 ( .A(n5098), .B(n4999), .ZN(n5517) );
  INV_X1 U6096 ( .A(n5000), .ZN(n5002) );
  AOI22_X1 U6097 ( .A1(n5002), .A2(n5001), .B1(n4117), .B2(n5000), .ZN(n5003)
         );
  XNOR2_X1 U6098 ( .A(n5004), .B(n5003), .ZN(n5094) );
  AOI21_X1 U6099 ( .B1(n5724), .B2(n5005), .A(REIP_REG_20__SCAN_IN), .ZN(n5006) );
  AOI21_X1 U6100 ( .B1(n5724), .B2(n5488), .A(n5723), .ZN(n5489) );
  OAI22_X1 U6101 ( .A1(n5006), .A2(n5489), .B1(n4156), .B2(n5761), .ZN(n5009)
         );
  INV_X1 U6102 ( .A(n5210), .ZN(n5007) );
  INV_X1 U6103 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5208) );
  OAI22_X1 U6104 ( .A1(n5007), .A2(n5738), .B1(n5683), .B2(n5208), .ZN(n5008)
         );
  AOI211_X1 U6105 ( .C1(n5094), .C2(n5758), .A(n5009), .B(n5008), .ZN(n5010)
         );
  OAI21_X1 U6106 ( .B1(n5517), .B2(n5695), .A(n5010), .ZN(U2807) );
  NAND2_X1 U6107 ( .A1(n4997), .A2(n5011), .ZN(n5545) );
  INV_X1 U6108 ( .A(n5545), .ZN(n5014) );
  NAND2_X1 U6109 ( .A1(n4997), .A2(n5012), .ZN(n5096) );
  INV_X1 U6110 ( .A(n5357), .ZN(n5021) );
  OAI21_X1 U6111 ( .B1(n5018), .B2(n4117), .A(n5016), .ZN(n5020) );
  OAI211_X1 U6112 ( .C1(n5018), .C2(n4117), .A(n5357), .B(n5016), .ZN(n5099)
         );
  INV_X1 U6113 ( .A(n5099), .ZN(n5019) );
  AOI21_X1 U6114 ( .B1(n5021), .B2(n5020), .A(n5019), .ZN(n5566) );
  AOI21_X1 U6115 ( .B1(n5724), .B2(n5022), .A(n5723), .ZN(n5628) );
  INV_X1 U6116 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6429) );
  NOR2_X1 U6117 ( .A1(n5754), .A2(n5022), .ZN(n5498) );
  AOI22_X1 U6118 ( .A1(EBX_REG_18__SCAN_IN), .A2(n5743), .B1(n5498), .B2(n6429), .ZN(n5023) );
  OAI21_X1 U6119 ( .B1(n5628), .B2(n6429), .A(n5023), .ZN(n5026) );
  NAND2_X1 U6120 ( .A1(n5763), .A2(n5219), .ZN(n5024) );
  OAI211_X1 U6121 ( .C1(n5683), .C2(n3745), .A(n5712), .B(n5024), .ZN(n5025)
         );
  AOI211_X1 U6122 ( .C1(n5566), .C2(n5758), .A(n5026), .B(n5025), .ZN(n5027)
         );
  OAI21_X1 U6123 ( .B1(n5222), .B2(n5695), .A(n5027), .ZN(U2809) );
  NAND2_X1 U6124 ( .A1(n4997), .A2(n5114), .ZN(n5118) );
  XNOR2_X1 U6125 ( .A(n5118), .B(n5106), .ZN(n5237) );
  OAI21_X1 U6126 ( .B1(n5646), .B2(n5754), .A(n5755), .ZN(n5647) );
  AOI22_X1 U6127 ( .A1(EBX_REG_15__SCAN_IN), .A2(n5743), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5647), .ZN(n5028) );
  OAI211_X1 U6128 ( .C1(n5683), .C2(n5029), .A(n5028), .B(n5712), .ZN(n5032)
         );
  NAND2_X1 U6129 ( .A1(n5724), .A2(n5646), .ZN(n5625) );
  NOR2_X1 U6130 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5625), .ZN(n5634) );
  AND2_X1 U6131 ( .A1(n5763), .A2(n5234), .ZN(n5030) );
  OR2_X1 U6132 ( .A1(n5634), .A2(n5030), .ZN(n5031) );
  NOR2_X1 U6133 ( .A1(n5032), .A2(n5031), .ZN(n5035) );
  AOI21_X1 U6134 ( .B1(n5033), .B2(n5119), .A(n5111), .ZN(n5581) );
  NAND2_X1 U6135 ( .A1(n5581), .A2(n5758), .ZN(n5034) );
  OAI211_X1 U6136 ( .C1(n5237), .C2(n5695), .A(n5035), .B(n5034), .ZN(U2812)
         );
  OAI21_X1 U6137 ( .B1(n3064), .B2(n5037), .A(n5036), .ZN(n5252) );
  INV_X1 U6138 ( .A(n5252), .ZN(n5039) );
  NAND2_X1 U6139 ( .A1(n5039), .A2(n2999), .ZN(n5051) );
  NAND3_X1 U6140 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .ZN(n5040) );
  NOR3_X1 U6141 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5040), .A3(n5676), .ZN(n5663) );
  OAI21_X1 U6142 ( .B1(n5663), .B2(n5659), .A(REIP_REG_13__SCAN_IN), .ZN(n5050) );
  INV_X1 U6143 ( .A(n5041), .ZN(n5249) );
  AOI21_X1 U6144 ( .B1(n5043), .B2(n5042), .A(n5121), .ZN(n5593) );
  INV_X1 U6145 ( .A(n5593), .ZN(n5124) );
  OAI22_X1 U6146 ( .A1(n5125), .A2(n5761), .B1(n5671), .B2(n5124), .ZN(n5044)
         );
  AOI21_X1 U6147 ( .B1(n5763), .B2(n5249), .A(n5044), .ZN(n5049) );
  INV_X1 U6148 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6633) );
  NAND3_X1 U6149 ( .A1(n5724), .A2(n5045), .A3(n6633), .ZN(n5046) );
  OAI211_X1 U6150 ( .C1(n5683), .C2(n5247), .A(n5712), .B(n5046), .ZN(n5047)
         );
  INV_X1 U6151 ( .A(n5047), .ZN(n5048) );
  NAND4_X1 U6152 ( .A1(n5051), .A2(n5050), .A3(n5049), .A4(n5048), .ZN(U2814)
         );
  OAI22_X1 U6153 ( .A1(n5053), .A2(n5122), .B1(n5776), .B2(n5052), .ZN(U2828)
         );
  OAI222_X1 U6154 ( .A1(n5136), .A2(n5126), .B1(n5054), .B2(n5776), .C1(n5286), 
        .C2(n5122), .ZN(U2831) );
  NAND2_X1 U6155 ( .A1(n5055), .A2(n5056), .ZN(n5057) );
  NAND2_X1 U6156 ( .A1(n5058), .A2(n5057), .ZN(n5435) );
  NOR2_X1 U6157 ( .A1(n5066), .A2(n5059), .ZN(n5060) );
  OR2_X1 U6158 ( .A1(n5061), .A2(n5060), .ZN(n5296) );
  OAI222_X1 U6159 ( .A1(n5435), .A2(n5126), .B1(n5062), .B2(n5776), .C1(n5122), 
        .C2(n5296), .ZN(U2832) );
  OAI21_X1 U6160 ( .B1(n5076), .B2(n5064), .A(n5055), .ZN(n5445) );
  AND2_X1 U6161 ( .A1(n5072), .A2(n5065), .ZN(n5067) );
  OR2_X1 U6162 ( .A1(n5067), .A2(n5066), .ZN(n5444) );
  OAI222_X1 U6163 ( .A1(n5445), .A2(n5126), .B1(n5776), .B2(n5068), .C1(n5444), 
        .C2(n5122), .ZN(U2833) );
  NAND2_X1 U6164 ( .A1(n5069), .A2(n5070), .ZN(n5071) );
  NAND2_X1 U6165 ( .A1(n5072), .A2(n5071), .ZN(n5554) );
  INV_X1 U6166 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5077) );
  NOR2_X1 U6167 ( .A1(n5073), .A2(n5074), .ZN(n5075) );
  OR2_X1 U6168 ( .A1(n5076), .A2(n5075), .ZN(n5523) );
  OAI222_X1 U6169 ( .A1(n5554), .A2(n5122), .B1(n5077), .B2(n5776), .C1(n5523), 
        .C2(n5126), .ZN(U2834) );
  AND2_X1 U6170 ( .A1(n5079), .A2(n5078), .ZN(n5080) );
  OR2_X1 U6171 ( .A1(n5080), .A2(n5073), .ZN(n5187) );
  OAI21_X1 U6172 ( .B1(n4322), .B2(n5081), .A(n5069), .ZN(n5467) );
  OAI222_X1 U6173 ( .A1(n5187), .A2(n5126), .B1(n5460), .B2(n5776), .C1(n5467), 
        .C2(n5122), .ZN(U2835) );
  AND2_X1 U6174 ( .A1(n5083), .A2(n5082), .ZN(n5084) );
  OR2_X1 U6175 ( .A1(n5084), .A2(n4323), .ZN(n5486) );
  OR2_X1 U6176 ( .A1(n5085), .A2(n5086), .ZN(n5087) );
  NAND2_X1 U6177 ( .A1(n4262), .A2(n5087), .ZN(n5482) );
  OAI222_X1 U6178 ( .A1(n5486), .A2(n5122), .B1(n5478), .B2(n5776), .C1(n5482), 
        .C2(n5126), .ZN(U2837) );
  NOR2_X1 U6179 ( .A1(n5089), .A2(n5088), .ZN(n5090) );
  OR2_X1 U6180 ( .A1(n5085), .A2(n5090), .ZN(n5200) );
  XOR2_X1 U6181 ( .A(n5092), .B(n5091), .Z(n5492) );
  INV_X1 U6182 ( .A(n5492), .ZN(n5093) );
  OAI222_X1 U6183 ( .A1(n5200), .A2(n5126), .B1(n5496), .B2(n5776), .C1(n5093), 
        .C2(n5122), .ZN(U2838) );
  INV_X1 U6184 ( .A(n5094), .ZN(n5349) );
  OAI222_X1 U6185 ( .A1(n5349), .A2(n5122), .B1(n5776), .B2(n4156), .C1(n5517), 
        .C2(n5126), .ZN(U2839) );
  NAND2_X1 U6186 ( .A1(n5096), .A2(n5095), .ZN(n5097) );
  INV_X1 U6187 ( .A(n5534), .ZN(n5102) );
  INV_X1 U6188 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5101) );
  XOR2_X1 U6189 ( .A(n5100), .B(n5099), .Z(n6689) );
  OAI222_X1 U6190 ( .A1(n5126), .A2(n5102), .B1(n5101), .B2(n5776), .C1(n5122), 
        .C2(n6689), .ZN(U2840) );
  AOI22_X1 U6191 ( .A1(n5566), .A2(n4194), .B1(EBX_REG_18__SCAN_IN), .B2(n5103), .ZN(n5104) );
  OAI21_X1 U6192 ( .B1(n5222), .B2(n5126), .A(n5104), .ZN(U2841) );
  AND2_X1 U6193 ( .A1(n4997), .A2(n5105), .ZN(n5543) );
  OR2_X1 U6194 ( .A1(n5118), .A2(n5106), .ZN(n5108) );
  AND2_X1 U6195 ( .A1(n5108), .A2(n5107), .ZN(n5109) );
  INV_X1 U6196 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5112) );
  OAI21_X1 U6197 ( .B1(n5111), .B2(n5110), .A(n3010), .ZN(n5645) );
  OAI222_X1 U6198 ( .A1(n5641), .A2(n5126), .B1(n5776), .B2(n5112), .C1(n5122), 
        .C2(n5645), .ZN(U2843) );
  INV_X1 U6199 ( .A(n5581), .ZN(n5113) );
  OAI222_X1 U6200 ( .A1(n5122), .A2(n5113), .B1(n5126), .B2(n5237), .C1(n6671), 
        .C2(n5776), .ZN(U2844) );
  INV_X1 U6201 ( .A(n5114), .ZN(n5116) );
  NAND3_X1 U6202 ( .A1(n5036), .A2(n5116), .A3(n5115), .ZN(n5117) );
  INV_X1 U6203 ( .A(n5654), .ZN(n5150) );
  INV_X1 U6204 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5123) );
  OAI21_X1 U6205 ( .B1(n5121), .B2(n5120), .A(n5119), .ZN(n5657) );
  OAI222_X1 U6206 ( .A1(n5126), .A2(n5150), .B1(n5776), .B2(n5123), .C1(n5122), 
        .C2(n5657), .ZN(U2845) );
  OAI222_X1 U6207 ( .A1(n5126), .A2(n5252), .B1(n5776), .B2(n5125), .C1(n5122), 
        .C2(n5124), .ZN(U2846) );
  NAND2_X1 U6208 ( .A1(n5151), .A2(n5127), .ZN(n5129) );
  AOI22_X1 U6209 ( .A1(n5780), .A2(DATAI_31_), .B1(n5783), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5128) );
  OAI21_X1 U6210 ( .B1(n5130), .B2(n5129), .A(n5128), .ZN(U2860) );
  AOI22_X1 U6211 ( .A1(n5780), .A2(DATAI_29_), .B1(n5783), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5132) );
  NAND2_X1 U6212 ( .A1(n5784), .A2(DATAI_13_), .ZN(n5131) );
  OAI211_X1 U6213 ( .C1(n5133), .C2(n5507), .A(n5132), .B(n5131), .ZN(U2862)
         );
  AOI22_X1 U6214 ( .A1(n5780), .A2(DATAI_28_), .B1(n5783), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5135) );
  NAND2_X1 U6215 ( .A1(n5784), .A2(DATAI_12_), .ZN(n5134) );
  OAI211_X1 U6216 ( .C1(n5136), .C2(n5507), .A(n5135), .B(n5134), .ZN(U2863)
         );
  AOI22_X1 U6217 ( .A1(n5784), .A2(DATAI_11_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n5783), .ZN(n5138) );
  NAND2_X1 U6218 ( .A1(n5780), .A2(DATAI_27_), .ZN(n5137) );
  OAI211_X1 U6219 ( .C1(n5435), .C2(n5507), .A(n5138), .B(n5137), .ZN(U2864)
         );
  AOI22_X1 U6220 ( .A1(n5784), .A2(DATAI_10_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n5783), .ZN(n5140) );
  NAND2_X1 U6221 ( .A1(n5780), .A2(DATAI_26_), .ZN(n5139) );
  OAI211_X1 U6222 ( .C1(n5445), .C2(n5507), .A(n5140), .B(n5139), .ZN(U2865)
         );
  AOI22_X1 U6223 ( .A1(n5784), .A2(DATAI_9_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n5783), .ZN(n5142) );
  NAND2_X1 U6224 ( .A1(n5780), .A2(DATAI_25_), .ZN(n5141) );
  OAI211_X1 U6225 ( .C1(n5523), .C2(n5507), .A(n5142), .B(n5141), .ZN(U2866)
         );
  AOI22_X1 U6226 ( .A1(n5784), .A2(DATAI_8_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n5783), .ZN(n5144) );
  NAND2_X1 U6227 ( .A1(n5780), .A2(DATAI_24_), .ZN(n5143) );
  OAI211_X1 U6228 ( .C1(n5187), .C2(n5507), .A(n5144), .B(n5143), .ZN(U2867)
         );
  AOI22_X1 U6229 ( .A1(n5780), .A2(DATAI_18_), .B1(n5783), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U6230 ( .A1(n5784), .A2(DATAI_2_), .ZN(n5145) );
  OAI211_X1 U6231 ( .C1(n5222), .C2(n5507), .A(n5146), .B(n5145), .ZN(U2873)
         );
  AOI22_X1 U6232 ( .A1(n5148), .A2(DATAI_15_), .B1(n5783), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5147) );
  OAI21_X1 U6233 ( .B1(n5237), .B2(n5507), .A(n5147), .ZN(U2876) );
  AOI22_X1 U6234 ( .A1(n5148), .A2(DATAI_14_), .B1(n5783), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5149) );
  OAI21_X1 U6235 ( .B1(n5150), .B2(n5507), .A(n5149), .ZN(U2877) );
  INV_X1 U6236 ( .A(DATAI_13_), .ZN(n5889) );
  INV_X1 U6237 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5813) );
  OAI222_X1 U6238 ( .A1(n5252), .A2(n5507), .B1(n5152), .B2(n5889), .C1(n5813), 
        .C2(n5151), .ZN(U2878) );
  NAND2_X1 U6239 ( .A1(n5919), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5153)
         );
  OAI211_X1 U6240 ( .C1(n5914), .C2(n5155), .A(n5154), .B(n5153), .ZN(n5156)
         );
  AOI21_X1 U6241 ( .B1(n5157), .B2(n5909), .A(n5156), .ZN(n5158) );
  OAI21_X1 U6242 ( .B1(n5159), .B2(n3056), .A(n5158), .ZN(U2957) );
  NAND3_X1 U6243 ( .A1(n3514), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5228), .ZN(n5162) );
  AND2_X1 U6244 ( .A1(n5177), .A2(n5559), .ZN(n5160) );
  NAND2_X1 U6245 ( .A1(n5161), .A2(n5160), .ZN(n5169) );
  INV_X1 U6246 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5309) );
  AOI22_X1 U6247 ( .A1(n5162), .A2(n5169), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5309), .ZN(n5163) );
  XNOR2_X1 U6248 ( .A(n5163), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5295)
         );
  NAND2_X1 U6249 ( .A1(n5897), .A2(n5164), .ZN(n5165) );
  NAND2_X1 U6250 ( .A1(n5917), .A2(REIP_REG_28__SCAN_IN), .ZN(n5287) );
  OAI211_X1 U6251 ( .C1(n5553), .C2(n6650), .A(n5165), .B(n5287), .ZN(n5166)
         );
  AOI21_X1 U6252 ( .B1(n5167), .B2(n5909), .A(n5166), .ZN(n5168) );
  OAI21_X1 U6253 ( .B1(n3056), .B2(n5295), .A(n5168), .ZN(U2958) );
  NAND2_X1 U6254 ( .A1(n5170), .A2(n5169), .ZN(n5171) );
  XNOR2_X1 U6255 ( .A(n5171), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5303)
         );
  INV_X1 U6256 ( .A(n5435), .ZN(n5174) );
  NAND2_X1 U6257 ( .A1(n5917), .A2(REIP_REG_27__SCAN_IN), .ZN(n5297) );
  NAND2_X1 U6258 ( .A1(n5919), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5172)
         );
  OAI211_X1 U6259 ( .C1(n5914), .C2(n5442), .A(n5297), .B(n5172), .ZN(n5173)
         );
  AOI21_X1 U6260 ( .B1(n5174), .B2(n5909), .A(n5173), .ZN(n5175) );
  OAI21_X1 U6261 ( .B1(n5303), .B2(n3056), .A(n5175), .ZN(U2959) );
  NOR2_X1 U6262 ( .A1(n5177), .A2(n5176), .ZN(n5178) );
  XOR2_X1 U6263 ( .A(n5178), .B(n3514), .Z(n5314) );
  NAND2_X1 U6264 ( .A1(n5917), .A2(REIP_REG_26__SCAN_IN), .ZN(n5308) );
  OAI21_X1 U6265 ( .B1(n5553), .B2(n5179), .A(n5308), .ZN(n5181) );
  NOR2_X1 U6266 ( .A1(n5445), .A2(n6275), .ZN(n5180) );
  AOI211_X1 U6267 ( .C1(n5897), .C2(n5447), .A(n5181), .B(n5180), .ZN(n5182)
         );
  OAI21_X1 U6268 ( .B1(n5314), .B2(n3056), .A(n5182), .ZN(U2960) );
  INV_X1 U6269 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6662) );
  NOR3_X1 U6270 ( .A1(n3075), .A2(n6662), .A3(n5315), .ZN(n5184) );
  OAI22_X1 U6271 ( .A1(n5193), .A2(n5315), .B1(n5185), .B2(n5184), .ZN(n5186)
         );
  XNOR2_X1 U6272 ( .A(n5186), .B(n6606), .ZN(n5321) );
  INV_X1 U6273 ( .A(n5187), .ZN(n5464) );
  INV_X1 U6274 ( .A(n5463), .ZN(n5189) );
  NAND2_X1 U6275 ( .A1(n5917), .A2(REIP_REG_24__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6276 ( .A1(n5919), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5188)
         );
  OAI211_X1 U6277 ( .C1(n5914), .C2(n5189), .A(n5317), .B(n5188), .ZN(n5190)
         );
  AOI21_X1 U6278 ( .B1(n5464), .B2(n5909), .A(n5190), .ZN(n5191) );
  OAI21_X1 U6279 ( .B1(n5321), .B2(n3056), .A(n5191), .ZN(U2962) );
  XNOR2_X1 U6280 ( .A(n3497), .B(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5192)
         );
  XNOR2_X1 U6281 ( .A(n5193), .B(n5192), .ZN(n5331) );
  NAND2_X1 U6282 ( .A1(n5917), .A2(REIP_REG_22__SCAN_IN), .ZN(n5322) );
  OAI21_X1 U6283 ( .B1(n5553), .B2(n5477), .A(n5322), .ZN(n5195) );
  NOR2_X1 U6284 ( .A1(n5482), .A2(n6275), .ZN(n5194) );
  AOI211_X1 U6285 ( .C1(n5897), .C2(n5483), .A(n5195), .B(n5194), .ZN(n5196)
         );
  OAI21_X1 U6286 ( .B1(n5331), .B2(n3056), .A(n5196), .ZN(U2964) );
  AOI21_X1 U6287 ( .B1(n5199), .B2(n5198), .A(n5197), .ZN(n5338) );
  NAND2_X1 U6288 ( .A1(n5917), .A2(REIP_REG_21__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6289 ( .A1(n5919), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5201)
         );
  OAI211_X1 U6290 ( .C1(n5914), .C2(n5491), .A(n5333), .B(n5201), .ZN(n5202)
         );
  AOI21_X1 U6291 ( .B1(n5514), .B2(n5909), .A(n5202), .ZN(n5203) );
  OAI21_X1 U6292 ( .B1(n5338), .B2(n3056), .A(n5203), .ZN(U2965) );
  INV_X1 U6293 ( .A(n5204), .ZN(n5205) );
  AOI21_X1 U6294 ( .B1(n5207), .B2(n5206), .A(n5205), .ZN(n5339) );
  NAND2_X1 U6295 ( .A1(n5339), .A2(n5916), .ZN(n5212) );
  NAND2_X1 U6296 ( .A1(n5917), .A2(REIP_REG_20__SCAN_IN), .ZN(n5348) );
  OAI21_X1 U6297 ( .B1(n5553), .B2(n5208), .A(n5348), .ZN(n5209) );
  AOI21_X1 U6298 ( .B1(n5897), .B2(n5210), .A(n5209), .ZN(n5211) );
  OAI211_X1 U6299 ( .C1(n5213), .C2(n5517), .A(n5212), .B(n5211), .ZN(U2966)
         );
  OR2_X1 U6300 ( .A1(n5214), .A2(n5564), .ZN(n5216) );
  MUX2_X1 U6301 ( .A(n5216), .B(n5215), .S(n3075), .Z(n5217) );
  XNOR2_X1 U6302 ( .A(n5217), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5567)
         );
  NAND2_X1 U6303 ( .A1(n5567), .A2(n5916), .ZN(n5221) );
  OAI22_X1 U6304 ( .A1(n5553), .A2(n3745), .B1(n6684), .B2(n6429), .ZN(n5218)
         );
  AOI21_X1 U6305 ( .B1(n5897), .B2(n5219), .A(n5218), .ZN(n5220) );
  OAI211_X1 U6306 ( .C1(n6275), .C2(n5222), .A(n5221), .B(n5220), .ZN(U2968)
         );
  XNOR2_X1 U6307 ( .A(n3497), .B(n5574), .ZN(n5223) );
  XNOR2_X1 U6308 ( .A(n4255), .B(n5223), .ZN(n5575) );
  INV_X1 U6309 ( .A(n5641), .ZN(n5782) );
  AOI22_X1 U6310 ( .A1(n5919), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n5917), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5224) );
  OAI21_X1 U6311 ( .B1(n5640), .B2(n5914), .A(n5224), .ZN(n5225) );
  AOI21_X1 U6312 ( .B1(n5782), .B2(n5909), .A(n5225), .ZN(n5226) );
  OAI21_X1 U6313 ( .B1(n3056), .B2(n5575), .A(n5226), .ZN(U2970) );
  NAND2_X1 U6314 ( .A1(n5228), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5230) );
  NAND3_X1 U6315 ( .A1(n5240), .A2(n3075), .A3(n5238), .ZN(n5229) );
  OAI21_X1 U6316 ( .B1(n5240), .B2(n5230), .A(n5229), .ZN(n5231) );
  XNOR2_X1 U6317 ( .A(n5231), .B(n4305), .ZN(n5582) );
  NAND2_X1 U6318 ( .A1(n5582), .A2(n5916), .ZN(n5236) );
  INV_X1 U6319 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5232) );
  OAI22_X1 U6320 ( .A1(n5553), .A2(n5029), .B1(n6684), .B2(n5232), .ZN(n5233)
         );
  AOI21_X1 U6321 ( .B1(n5897), .B2(n5234), .A(n5233), .ZN(n5235) );
  OAI211_X1 U6322 ( .C1(n5237), .C2(n6275), .A(n5236), .B(n5235), .ZN(U2971)
         );
  XNOR2_X1 U6323 ( .A(n3497), .B(n5238), .ZN(n5239) );
  XNOR2_X1 U6324 ( .A(n5240), .B(n5239), .ZN(n5363) );
  NOR2_X1 U6325 ( .A1(n5914), .A2(n5652), .ZN(n5243) );
  INV_X1 U6326 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5241) );
  OAI22_X1 U6327 ( .A1(n5553), .A2(n5241), .B1(n6684), .B2(n6424), .ZN(n5242)
         );
  AOI211_X1 U6328 ( .C1(n5654), .C2(n5909), .A(n5243), .B(n5242), .ZN(n5244)
         );
  OAI21_X1 U6329 ( .B1(n3056), .B2(n5363), .A(n5244), .ZN(U2972) );
  XNOR2_X1 U6330 ( .A(n5246), .B(n5245), .ZN(n5588) );
  NAND2_X1 U6331 ( .A1(n5588), .A2(n5916), .ZN(n5251) );
  OAI22_X1 U6332 ( .A1(n5553), .A2(n5247), .B1(n6684), .B2(n6633), .ZN(n5248)
         );
  AOI21_X1 U6333 ( .B1(n5897), .B2(n5249), .A(n5248), .ZN(n5250) );
  OAI211_X1 U6334 ( .C1(n5252), .C2(n6275), .A(n5251), .B(n5250), .ZN(U2973)
         );
  NAND2_X1 U6335 ( .A1(n5253), .A2(n5254), .ZN(n5258) );
  INV_X1 U6336 ( .A(n5381), .ZN(n5256) );
  NOR2_X1 U6337 ( .A1(n5256), .A2(n5255), .ZN(n5257) );
  NAND2_X1 U6338 ( .A1(n5258), .A2(n5257), .ZN(n5382) );
  OAI21_X1 U6339 ( .B1(n5258), .B2(n5257), .A(n5382), .ZN(n5259) );
  INV_X1 U6340 ( .A(n5259), .ZN(n5926) );
  NAND2_X1 U6341 ( .A1(n5926), .A2(n5916), .ZN(n5263) );
  AND2_X1 U6342 ( .A1(n5917), .A2(REIP_REG_11__SCAN_IN), .ZN(n5923) );
  NOR2_X1 U6343 ( .A1(n5914), .A2(n5260), .ZN(n5261) );
  AOI211_X1 U6344 ( .C1(n5919), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n5923), 
        .B(n5261), .ZN(n5262) );
  OAI211_X1 U6345 ( .C1(n6275), .C2(n5264), .A(n5263), .B(n5262), .ZN(U2975)
         );
  INV_X1 U6346 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5265) );
  OAI22_X1 U6347 ( .A1(n5553), .A2(n5265), .B1(n6684), .B2(n6417), .ZN(n5267)
         );
  NOR2_X1 U6348 ( .A1(n5673), .A2(n6275), .ZN(n5266) );
  AOI211_X1 U6349 ( .C1(n5897), .C2(n5674), .A(n5267), .B(n5266), .ZN(n5268)
         );
  OAI21_X1 U6350 ( .B1(n5269), .B2(n3056), .A(n5268), .ZN(U2976) );
  INV_X1 U6351 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U6352 ( .A1(n5897), .A2(n5270), .ZN(n5277) );
  INV_X1 U6353 ( .A(n5271), .ZN(n5273) );
  AOI22_X1 U6354 ( .A1(n5273), .A2(n5916), .B1(n5909), .B2(n5272), .ZN(n5276)
         );
  NAND2_X1 U6355 ( .A1(n5919), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5274)
         );
  NAND4_X1 U6356 ( .A1(n5277), .A2(n5276), .A3(n5275), .A4(n5274), .ZN(U2985)
         );
  NAND3_X1 U6357 ( .A1(n5278), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5281), .ZN(n5279) );
  OAI211_X1 U6358 ( .C1(n5282), .C2(n5281), .A(n5280), .B(n5279), .ZN(n5283)
         );
  AOI21_X1 U6359 ( .B1(n3086), .B2(n5944), .A(n5283), .ZN(n5284) );
  OAI21_X1 U6360 ( .B1(n5285), .B2(n5394), .A(n5284), .ZN(U2988) );
  INV_X1 U6361 ( .A(n5286), .ZN(n5293) );
  INV_X1 U6362 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U6363 ( .A1(n5290), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5288) );
  OAI21_X1 U6364 ( .B1(n5289), .B2(n5288), .A(n5287), .ZN(n5292) );
  OR2_X1 U6365 ( .A1(n5289), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5298)
         );
  AOI21_X1 U6366 ( .B1(n5300), .B2(n5298), .A(n5290), .ZN(n5291) );
  AOI211_X1 U6367 ( .C1(n5293), .C2(n5944), .A(n5292), .B(n5291), .ZN(n5294)
         );
  OAI21_X1 U6368 ( .B1(n5295), .B2(n5394), .A(n5294), .ZN(U2990) );
  INV_X1 U6369 ( .A(n5296), .ZN(n5439) );
  OAI211_X1 U6370 ( .C1(n5300), .C2(n5299), .A(n5298), .B(n5297), .ZN(n5301)
         );
  AOI21_X1 U6371 ( .B1(n5944), .B2(n5439), .A(n5301), .ZN(n5302) );
  OAI21_X1 U6372 ( .B1(n5303), .B2(n5394), .A(n5302), .ZN(U2991) );
  INV_X1 U6373 ( .A(n5444), .ZN(n5312) );
  INV_X1 U6374 ( .A(n5558), .ZN(n5310) );
  INV_X1 U6375 ( .A(n5560), .ZN(n5304) );
  AOI21_X1 U6376 ( .B1(n5309), .B2(n5559), .A(n5304), .ZN(n5305) );
  NAND2_X1 U6377 ( .A1(n5306), .A2(n5305), .ZN(n5307) );
  OAI211_X1 U6378 ( .C1(n5310), .C2(n5309), .A(n5308), .B(n5307), .ZN(n5311)
         );
  AOI21_X1 U6379 ( .B1(n5944), .B2(n5312), .A(n5311), .ZN(n5313) );
  OAI21_X1 U6380 ( .B1(n5314), .B2(n5394), .A(n5313), .ZN(U2992) );
  NOR3_X1 U6381 ( .A1(n5335), .A2(n5323), .A3(n5315), .ZN(n5316) );
  OAI21_X1 U6382 ( .B1(INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n5316), .A(n5558), 
        .ZN(n5318) );
  OAI211_X1 U6383 ( .C1(n5467), .C2(n6688), .A(n5318), .B(n5317), .ZN(n5319)
         );
  INV_X1 U6384 ( .A(n5319), .ZN(n5320) );
  OAI21_X1 U6385 ( .B1(n5321), .B2(n5394), .A(n5320), .ZN(U2994) );
  INV_X1 U6386 ( .A(n5322), .ZN(n5327) );
  INV_X1 U6387 ( .A(n5323), .ZN(n5324) );
  NOR3_X1 U6388 ( .A1(n5335), .A2(n5325), .A3(n5324), .ZN(n5326) );
  AOI211_X1 U6389 ( .C1(n5332), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5327), .B(n5326), .ZN(n5330) );
  INV_X1 U6390 ( .A(n5486), .ZN(n5328) );
  NAND2_X1 U6391 ( .A1(n5328), .A2(n5944), .ZN(n5329) );
  OAI211_X1 U6392 ( .C1(n5331), .C2(n5394), .A(n5330), .B(n5329), .ZN(U2996)
         );
  NAND2_X1 U6393 ( .A1(n5332), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5334) );
  OAI211_X1 U6394 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5335), .A(n5334), .B(n5333), .ZN(n5336) );
  AOI21_X1 U6395 ( .B1(n5944), .B2(n5492), .A(n5336), .ZN(n5337) );
  OAI21_X1 U6396 ( .B1(n5338), .B2(n5394), .A(n5337), .ZN(U2997) );
  INV_X1 U6397 ( .A(n5339), .ZN(n5352) );
  AOI221_X1 U6398 ( .B1(n5342), .B2(n5564), .C1(n5341), .C2(n5564), .A(n5340), 
        .ZN(n5570) );
  OAI21_X1 U6399 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5343), .A(n5570), 
        .ZN(n6693) );
  NOR2_X1 U6400 ( .A1(n5344), .A2(n6686), .ZN(n5345) );
  NAND2_X1 U6401 ( .A1(n5346), .A2(n5345), .ZN(n5347) );
  OAI211_X1 U6402 ( .C1(n5349), .C2(n6688), .A(n5348), .B(n5347), .ZN(n5350)
         );
  AOI21_X1 U6403 ( .B1(n6693), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5350), 
        .ZN(n5351) );
  OAI21_X1 U6404 ( .B1(n5352), .B2(n5394), .A(n5351), .ZN(U2998) );
  OR3_X1 U6405 ( .A1(n4255), .A2(n3075), .A3(n5574), .ZN(n5355) );
  NOR2_X1 U6406 ( .A1(n5228), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5353)
         );
  NAND2_X1 U6407 ( .A1(n4255), .A2(n5353), .ZN(n5354) );
  NAND2_X1 U6408 ( .A1(n5355), .A2(n5354), .ZN(n5356) );
  XNOR2_X1 U6409 ( .A(n5356), .B(n5564), .ZN(n5546) );
  NAND2_X1 U6410 ( .A1(n5546), .A2(n5951), .ZN(n5361) );
  AOI21_X1 U6411 ( .B1(n5358), .B2(n3010), .A(n5357), .ZN(n5768) );
  NAND2_X1 U6412 ( .A1(n5917), .A2(REIP_REG_17__SCAN_IN), .ZN(n5551) );
  OAI21_X1 U6413 ( .B1(n5563), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5551), 
        .ZN(n5359) );
  AOI21_X1 U6414 ( .B1(n5768), .B2(n5944), .A(n5359), .ZN(n5360) );
  OAI211_X1 U6415 ( .C1(n5362), .C2(n5564), .A(n5361), .B(n5360), .ZN(U3001)
         );
  NOR2_X1 U6416 ( .A1(n5363), .A2(n5394), .ZN(n5380) );
  INV_X1 U6417 ( .A(n5374), .ZN(n5364) );
  NOR4_X1 U6418 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5929), .A3(n5373), 
        .A4(n5364), .ZN(n5379) );
  NOR2_X1 U6419 ( .A1(n5366), .A2(n5365), .ZN(n5367) );
  OAI21_X1 U6420 ( .B1(n5368), .B2(n5367), .A(n5374), .ZN(n5369) );
  NOR2_X1 U6421 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5369), .ZN(n5591)
         );
  NAND2_X1 U6422 ( .A1(n5374), .A2(n5370), .ZN(n5590) );
  INV_X1 U6423 ( .A(n5371), .ZN(n5372) );
  OAI21_X1 U6424 ( .B1(n5373), .B2(n5590), .A(n5372), .ZN(n5589) );
  OAI211_X1 U6425 ( .C1(n5375), .C2(n5374), .A(n5589), .B(n5385), .ZN(n5587)
         );
  OAI21_X1 U6426 ( .B1(n5591), .B2(n5587), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5377) );
  NAND2_X1 U6427 ( .A1(n5917), .A2(REIP_REG_14__SCAN_IN), .ZN(n5376) );
  OAI211_X1 U6428 ( .C1(n5657), .C2(n6688), .A(n5377), .B(n5376), .ZN(n5378)
         );
  OR3_X1 U6429 ( .A1(n5380), .A2(n5379), .A3(n5378), .ZN(U3004) );
  NAND2_X1 U6430 ( .A1(n5382), .A2(n5381), .ZN(n5384) );
  XNOR2_X1 U6431 ( .A(n3497), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5383)
         );
  XNOR2_X1 U6432 ( .A(n5384), .B(n5383), .ZN(n5902) );
  OAI21_X1 U6433 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n5386), .A(n5385), 
        .ZN(n5389) );
  NOR2_X1 U6434 ( .A1(n5929), .A2(n5387), .ZN(n5388) );
  AOI22_X1 U6435 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n5389), .B1(n5388), .B2(n3500), .ZN(n5391) );
  NAND2_X1 U6436 ( .A1(n5917), .A2(REIP_REG_12__SCAN_IN), .ZN(n5390) );
  OAI211_X1 U6437 ( .C1(n5658), .C2(n6688), .A(n5391), .B(n5390), .ZN(n5392)
         );
  INV_X1 U6438 ( .A(n5392), .ZN(n5393) );
  OAI21_X1 U6439 ( .B1(n5902), .B2(n5394), .A(n5393), .ZN(U3006) );
  NOR2_X1 U6440 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6376), .ZN(n6459) );
  OAI211_X1 U6441 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4526), .A(n5423), .B(
        n6464), .ZN(n5395) );
  OAI21_X1 U6442 ( .B1(n5396), .B2(n6459), .A(n5395), .ZN(n5418) );
  OR2_X1 U6443 ( .A1(n6341), .A2(n5397), .ZN(n5399) );
  NAND2_X1 U6444 ( .A1(n6341), .A2(n3321), .ZN(n5398) );
  MUX2_X1 U6445 ( .A(n5400), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6341), 
        .Z(n6345) );
  NAND3_X1 U6446 ( .A1(n6343), .A2(n6345), .A3(n6376), .ZN(n5403) );
  NAND2_X1 U6447 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5609), .ZN(n5411) );
  INV_X1 U6448 ( .A(n5411), .ZN(n5401) );
  NAND2_X1 U6449 ( .A1(n5403), .A2(n5402), .ZN(n6348) );
  INV_X1 U6450 ( .A(n4428), .ZN(n5404) );
  NAND2_X1 U6451 ( .A1(n6348), .A2(n5404), .ZN(n5415) );
  NAND2_X1 U6452 ( .A1(n6341), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5410) );
  OR2_X1 U6453 ( .A1(n5406), .A2(n5405), .ZN(n5407) );
  XNOR2_X1 U6454 ( .A(n5407), .B(n3522), .ZN(n5725) );
  OR2_X1 U6455 ( .A1(n5725), .A2(n5408), .ZN(n5409) );
  AOI21_X1 U6456 ( .B1(n5410), .B2(n5409), .A(STATE2_REG_1__SCAN_IN), .ZN(
        n5413) );
  NOR2_X1 U6457 ( .A1(n3522), .A2(n5411), .ZN(n5412) );
  INV_X1 U6458 ( .A(n6356), .ZN(n5414) );
  NAND2_X1 U6459 ( .A1(n5415), .A2(n5414), .ZN(n6358) );
  INV_X1 U6460 ( .A(n6456), .ZN(n6360) );
  OAI21_X1 U6461 ( .B1(n6358), .B2(FLUSH_REG_SCAN_IN), .A(n6360), .ZN(n5417)
         );
  NAND2_X1 U6462 ( .A1(n5417), .A2(n5416), .ZN(n6466) );
  MUX2_X1 U6463 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5418), .S(n6466), 
        .Z(U3464) );
  AOI21_X1 U6464 ( .B1(n3074), .B2(n5423), .A(n5419), .ZN(n5421) );
  OAI22_X1 U6465 ( .A1(n5421), .A2(n6271), .B1(n5420), .B2(n6459), .ZN(n5422)
         );
  MUX2_X1 U6466 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5422), .S(n6466), 
        .Z(U3463) );
  NOR2_X1 U6467 ( .A1(n5424), .A2(n5423), .ZN(n6050) );
  NOR2_X1 U6468 ( .A1(n5425), .A2(n6050), .ZN(n5426) );
  OAI222_X1 U6469 ( .A1(n6022), .A2(n5427), .B1(n6271), .B2(n5426), .C1(n6459), 
        .C2(n6051), .ZN(n5428) );
  MUX2_X1 U6470 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5428), .S(n6466), 
        .Z(U3462) );
  NAND2_X1 U6471 ( .A1(n6462), .A2(n6368), .ZN(n5825) );
  INV_X2 U6472 ( .A(n5825), .ZN(n5816) );
  INV_X1 U6473 ( .A(n5429), .ZN(n6335) );
  AOI21_X1 U6474 ( .B1(n6335), .B2(n5839), .A(n6391), .ZN(n5430) );
  INV_X2 U6475 ( .A(n5824), .ZN(n5835) );
  AND2_X1 U6476 ( .A1(n5835), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI21_X1 U6477 ( .B1(n5432), .B2(MEMORYFETCH_REG_SCAN_IN), .A(n5431), .ZN(
        n5433) );
  INV_X1 U6478 ( .A(n5433), .ZN(U2788) );
  INV_X1 U6479 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6440) );
  AOI22_X1 U6480 ( .A1(EBX_REG_27__SCAN_IN), .A2(n5743), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n5764), .ZN(n5434) );
  OAI21_X1 U6481 ( .B1(n5451), .B2(n6440), .A(n5434), .ZN(n5437) );
  NOR2_X1 U6482 ( .A1(n5435), .A2(n5695), .ZN(n5436) );
  AOI211_X1 U6483 ( .C1(n5438), .C2(n6440), .A(n5437), .B(n5436), .ZN(n5441)
         );
  NAND2_X1 U6484 ( .A1(n5439), .A2(n5758), .ZN(n5440) );
  OAI211_X1 U6485 ( .C1(n5738), .C2(n5442), .A(n5441), .B(n5440), .ZN(U2800)
         );
  NOR2_X1 U6486 ( .A1(REIP_REG_26__SCAN_IN), .A2(n5443), .ZN(n5450) );
  AOI22_X1 U6487 ( .A1(EBX_REG_26__SCAN_IN), .A2(n5743), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n5764), .ZN(n5449) );
  OAI22_X1 U6488 ( .A1(n5445), .A2(n5695), .B1(n5671), .B2(n5444), .ZN(n5446)
         );
  AOI21_X1 U6489 ( .B1(n5447), .B2(n5763), .A(n5446), .ZN(n5448) );
  OAI211_X1 U6490 ( .C1(n5451), .C2(n5450), .A(n5449), .B(n5448), .ZN(U2801)
         );
  INV_X1 U6491 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6436) );
  NAND2_X1 U6492 ( .A1(n5452), .A2(n6436), .ZN(n5459) );
  AOI21_X1 U6493 ( .B1(n5470), .B2(n5459), .A(n6438), .ZN(n5455) );
  OAI22_X1 U6494 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5453), .B1(n3950), .B2(
        n5683), .ZN(n5454) );
  AOI211_X1 U6495 ( .C1(n5743), .C2(EBX_REG_25__SCAN_IN), .A(n5455), .B(n5454), 
        .ZN(n5458) );
  OAI22_X1 U6496 ( .A1(n5523), .A2(n5695), .B1(n5671), .B2(n5554), .ZN(n5456)
         );
  INV_X1 U6497 ( .A(n5456), .ZN(n5457) );
  OAI211_X1 U6498 ( .C1(n5531), .C2(n5738), .A(n5458), .B(n5457), .ZN(U2802)
         );
  INV_X1 U6499 ( .A(n5459), .ZN(n5462) );
  OAI22_X1 U6500 ( .A1(n5470), .A2(n6436), .B1(n5460), .B2(n5761), .ZN(n5461)
         );
  AOI211_X1 U6501 ( .C1(n5764), .C2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5462), 
        .B(n5461), .ZN(n5466) );
  AOI22_X1 U6502 ( .A1(n5464), .A2(n2999), .B1(n5463), .B2(n5763), .ZN(n5465)
         );
  OAI211_X1 U6503 ( .C1(n5467), .C2(n5671), .A(n5466), .B(n5465), .ZN(U2803)
         );
  AND2_X1 U6504 ( .A1(n5724), .A2(n5468), .ZN(n5481) );
  AOI21_X1 U6505 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5481), .A(
        REIP_REG_23__SCAN_IN), .ZN(n5469) );
  INV_X1 U6506 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6525) );
  OAI22_X1 U6507 ( .A1(n5470), .A2(n5469), .B1(n6525), .B2(n5683), .ZN(n5471)
         );
  AOI21_X1 U6508 ( .B1(EBX_REG_23__SCAN_IN), .B2(n5743), .A(n5471), .ZN(n5475)
         );
  INV_X1 U6509 ( .A(n5472), .ZN(n5508) );
  INV_X1 U6510 ( .A(n5473), .ZN(n5504) );
  AOI22_X1 U6511 ( .A1(n5508), .A2(n2999), .B1(n5758), .B2(n5504), .ZN(n5474)
         );
  OAI211_X1 U6512 ( .C1(n5476), .C2(n5738), .A(n5475), .B(n5474), .ZN(U2804)
         );
  INV_X1 U6513 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6434) );
  OAI21_X1 U6514 ( .B1(REIP_REG_21__SCAN_IN), .B2(n5754), .A(n5489), .ZN(n5480) );
  OAI22_X1 U6515 ( .A1(n5478), .A2(n5761), .B1(n5477), .B2(n5683), .ZN(n5479)
         );
  AOI221_X1 U6516 ( .B1(n5481), .B2(n6434), .C1(n5480), .C2(
        REIP_REG_22__SCAN_IN), .A(n5479), .ZN(n5485) );
  INV_X1 U6517 ( .A(n5482), .ZN(n5511) );
  AOI22_X1 U6518 ( .A1(n5511), .A2(n2999), .B1(n5483), .B2(n5763), .ZN(n5484)
         );
  OAI211_X1 U6519 ( .C1(n5486), .C2(n5671), .A(n5485), .B(n5484), .ZN(U2805)
         );
  NAND2_X1 U6520 ( .A1(n5724), .A2(n6433), .ZN(n5487) );
  OAI22_X1 U6521 ( .A1(n6433), .A2(n5489), .B1(n5488), .B2(n5487), .ZN(n5490)
         );
  AOI21_X1 U6522 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n5764), .A(n5490), 
        .ZN(n5495) );
  INV_X1 U6523 ( .A(n5491), .ZN(n5493) );
  AOI222_X1 U6524 ( .A1(n5514), .A2(n2999), .B1(n5493), .B2(n5763), .C1(n5758), 
        .C2(n5492), .ZN(n5494) );
  OAI211_X1 U6525 ( .C1(n5496), .C2(n5761), .A(n5495), .B(n5494), .ZN(U2806)
         );
  INV_X1 U6526 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6685) );
  INV_X1 U6527 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5541) );
  OAI211_X1 U6528 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n5498), .B(n5497), .ZN(n5499) );
  OAI211_X1 U6529 ( .C1(n5683), .C2(n5541), .A(n5499), .B(n5712), .ZN(n5500)
         );
  AOI21_X1 U6530 ( .B1(EBX_REG_19__SCAN_IN), .B2(n5743), .A(n5500), .ZN(n5503)
         );
  OAI22_X1 U6531 ( .A1(n6689), .A2(n5671), .B1(n5537), .B2(n5738), .ZN(n5501)
         );
  AOI21_X1 U6532 ( .B1(n5534), .B2(n2999), .A(n5501), .ZN(n5502) );
  OAI211_X1 U6533 ( .C1(n5628), .C2(n6685), .A(n5503), .B(n5502), .ZN(U2808)
         );
  AOI22_X1 U6534 ( .A1(n5508), .A2(n5772), .B1(n4194), .B2(n5504), .ZN(n5505)
         );
  OAI21_X1 U6535 ( .B1(n5776), .B2(n5506), .A(n5505), .ZN(U2836) );
  AOI22_X1 U6536 ( .A1(n5508), .A2(n5781), .B1(n5780), .B2(DATAI_23_), .ZN(
        n5510) );
  AOI22_X1 U6537 ( .A1(n5784), .A2(DATAI_7_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n5783), .ZN(n5509) );
  NAND2_X1 U6538 ( .A1(n5510), .A2(n5509), .ZN(U2868) );
  AOI22_X1 U6539 ( .A1(n5511), .A2(n5781), .B1(n5780), .B2(DATAI_22_), .ZN(
        n5513) );
  AOI22_X1 U6540 ( .A1(n5784), .A2(DATAI_6_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n5783), .ZN(n5512) );
  NAND2_X1 U6541 ( .A1(n5513), .A2(n5512), .ZN(U2869) );
  AOI22_X1 U6542 ( .A1(n5514), .A2(n5781), .B1(n5780), .B2(DATAI_21_), .ZN(
        n5516) );
  AOI22_X1 U6543 ( .A1(n5784), .A2(DATAI_5_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n5783), .ZN(n5515) );
  NAND2_X1 U6544 ( .A1(n5516), .A2(n5515), .ZN(U2870) );
  INV_X1 U6545 ( .A(n5517), .ZN(n5518) );
  AOI22_X1 U6546 ( .A1(n5518), .A2(n5781), .B1(n5780), .B2(DATAI_20_), .ZN(
        n5520) );
  AOI22_X1 U6547 ( .A1(n5784), .A2(DATAI_4_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n5783), .ZN(n5519) );
  NAND2_X1 U6548 ( .A1(n5520), .A2(n5519), .ZN(U2871) );
  AOI22_X1 U6549 ( .A1(n5534), .A2(n5781), .B1(n5780), .B2(DATAI_19_), .ZN(
        n5522) );
  AOI22_X1 U6550 ( .A1(n5784), .A2(DATAI_3_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n5783), .ZN(n5521) );
  NAND2_X1 U6551 ( .A1(n5522), .A2(n5521), .ZN(U2872) );
  AOI22_X1 U6552 ( .A1(n5917), .A2(REIP_REG_25__SCAN_IN), .B1(n5919), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5530) );
  INV_X1 U6553 ( .A(n5523), .ZN(n5528) );
  AOI21_X1 U6554 ( .B1(n5526), .B2(n5525), .A(n5524), .ZN(n5527) );
  INV_X1 U6555 ( .A(n5527), .ZN(n5556) );
  AOI22_X1 U6556 ( .A1(n5528), .A2(n5909), .B1(n5916), .B2(n5556), .ZN(n5529)
         );
  OAI211_X1 U6557 ( .C1(n5914), .C2(n5531), .A(n5530), .B(n5529), .ZN(U2961)
         );
  XNOR2_X1 U6558 ( .A(n5533), .B(n5532), .ZN(n6687) );
  NAND2_X1 U6559 ( .A1(n6687), .A2(n5916), .ZN(n5536) );
  NAND2_X1 U6560 ( .A1(n5534), .A2(n5909), .ZN(n5535) );
  OAI211_X1 U6561 ( .C1(n5914), .C2(n5537), .A(n5536), .B(n5535), .ZN(n5538)
         );
  INV_X1 U6562 ( .A(n5538), .ZN(n5540) );
  NAND2_X1 U6563 ( .A1(n5917), .A2(REIP_REG_19__SCAN_IN), .ZN(n5539) );
  OAI211_X1 U6564 ( .C1(n5541), .C2(n5553), .A(n5540), .B(n5539), .ZN(U2967)
         );
  INV_X1 U6565 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5626) );
  OR2_X1 U6566 ( .A1(n5543), .A2(n5542), .ZN(n5544) );
  NAND2_X1 U6567 ( .A1(n5545), .A2(n5544), .ZN(n5630) );
  NAND2_X1 U6568 ( .A1(n5546), .A2(n5916), .ZN(n5549) );
  INV_X1 U6569 ( .A(n5633), .ZN(n5547) );
  NAND2_X1 U6570 ( .A1(n5897), .A2(n5547), .ZN(n5548) );
  OAI211_X1 U6571 ( .C1(n6275), .C2(n5630), .A(n5549), .B(n5548), .ZN(n5550)
         );
  INV_X1 U6572 ( .A(n5550), .ZN(n5552) );
  OAI211_X1 U6573 ( .C1(n5626), .C2(n5553), .A(n5552), .B(n5551), .ZN(U2969)
         );
  INV_X1 U6574 ( .A(n5554), .ZN(n5555) );
  AOI22_X1 U6575 ( .A1(n5556), .A2(n5951), .B1(n5944), .B2(n5555), .ZN(n5562)
         );
  NOR2_X1 U6576 ( .A1(n6684), .A2(n6438), .ZN(n5557) );
  AOI221_X1 U6577 ( .B1(n5560), .B2(n5559), .C1(n5558), .C2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5557), .ZN(n5561) );
  NAND2_X1 U6578 ( .A1(n5562), .A2(n5561), .ZN(U2993) );
  NOR3_X1 U6579 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5564), .A3(n5563), 
        .ZN(n5565) );
  AOI21_X1 U6580 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5917), .A(n5565), .ZN(n5569) );
  AOI22_X1 U6581 ( .A1(n5567), .A2(n5951), .B1(n5944), .B2(n5566), .ZN(n5568)
         );
  OAI211_X1 U6582 ( .C1(n5570), .C2(n6626), .A(n5569), .B(n5568), .ZN(U3000)
         );
  NAND2_X1 U6583 ( .A1(n5571), .A2(n5574), .ZN(n5579) );
  NOR3_X1 U6584 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n5929), .A3(n5573), 
        .ZN(n5580) );
  AOI211_X1 U6585 ( .C1(n5573), .C2(n5572), .A(n5580), .B(n5925), .ZN(n5586)
         );
  OAI222_X1 U6586 ( .A1(n5575), .A2(n5394), .B1(n6688), .B2(n5645), .C1(n5574), 
        .C2(n5586), .ZN(n5576) );
  INV_X1 U6587 ( .A(n5576), .ZN(n5578) );
  NAND2_X1 U6588 ( .A1(n5917), .A2(REIP_REG_16__SCAN_IN), .ZN(n5577) );
  OAI211_X1 U6589 ( .C1(n5929), .C2(n5579), .A(n5578), .B(n5577), .ZN(U3002)
         );
  NOR2_X1 U6590 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n5580), .ZN(n5585)
         );
  AOI22_X1 U6591 ( .A1(n5582), .A2(n5951), .B1(n5944), .B2(n5581), .ZN(n5584)
         );
  NAND2_X1 U6592 ( .A1(n5917), .A2(REIP_REG_15__SCAN_IN), .ZN(n5583) );
  OAI211_X1 U6593 ( .C1(n5586), .C2(n5585), .A(n5584), .B(n5583), .ZN(U3003)
         );
  AOI22_X1 U6594 ( .A1(n5588), .A2(n5951), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5587), .ZN(n5595) );
  OAI22_X1 U6595 ( .A1(n5590), .A2(n5589), .B1(n6633), .B2(n6684), .ZN(n5592)
         );
  AOI211_X1 U6596 ( .C1(n5944), .C2(n5593), .A(n5592), .B(n5591), .ZN(n5594)
         );
  NAND2_X1 U6597 ( .A1(n5595), .A2(n5594), .ZN(U3005) );
  INV_X1 U6598 ( .A(n5725), .ZN(n5596) );
  NAND4_X1 U6599 ( .A1(n5599), .A2(n5598), .A3(n5597), .A4(n5596), .ZN(n5600)
         );
  OAI21_X1 U6600 ( .B1(n5601), .B2(n3522), .A(n5600), .ZN(U3455) );
  AOI21_X1 U6601 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6529), .A(n6393), .ZN(n5607) );
  INV_X1 U6602 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5602) );
  NOR2_X2 U6603 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6392), .ZN(n6491) );
  AOI21_X1 U6604 ( .B1(n5607), .B2(n5602), .A(n6491), .ZN(U2789) );
  NAND2_X1 U6605 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6486), .ZN(n5605) );
  OAI21_X1 U6606 ( .B1(n5603), .B2(n6374), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5604) );
  OAI21_X1 U6607 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5605), .A(n5604), .ZN(
        U2790) );
  NOR2_X1 U6608 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5608) );
  OAI21_X1 U6609 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5608), .A(n6480), .ZN(n5606)
         );
  OAI21_X1 U6610 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6480), .A(n5606), .ZN(
        U2791) );
  NOR2_X1 U6611 ( .A1(n6491), .A2(n5607), .ZN(n6455) );
  OAI21_X1 U6612 ( .B1(BS16_N), .B2(n5608), .A(n6455), .ZN(n6453) );
  OAI21_X1 U6613 ( .B1(n6455), .B2(n6224), .A(n6453), .ZN(U2792) );
  OAI21_X1 U6614 ( .B1(n5610), .B2(n5609), .A(n3056), .ZN(U2793) );
  NOR4_X1 U6615 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n5614) );
  NOR4_X1 U6616 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n5613) );
  NOR4_X1 U6617 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5612) );
  NOR4_X1 U6618 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n5611) );
  NAND4_X1 U6619 ( .A1(n5614), .A2(n5613), .A3(n5612), .A4(n5611), .ZN(n5620)
         );
  NOR4_X1 U6620 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n5618) );
  AOI211_X1 U6621 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_8__SCAN_IN), .B(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5617) );
  NOR4_X1 U6622 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n5616) );
  NOR4_X1 U6623 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n5615) );
  NAND4_X1 U6624 ( .A1(n5618), .A2(n5617), .A3(n5616), .A4(n5615), .ZN(n5619)
         );
  NOR2_X1 U6625 ( .A1(n5620), .A2(n5619), .ZN(n6478) );
  INV_X1 U6626 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5622) );
  NOR3_X1 U6627 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_1__SCAN_IN), .ZN(n5623) );
  OAI21_X1 U6628 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5623), .A(n6478), .ZN(n5621)
         );
  OAI21_X1 U6629 ( .B1(n6478), .B2(n5622), .A(n5621), .ZN(U2794) );
  INV_X1 U6630 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6656) );
  NOR2_X1 U6631 ( .A1(REIP_REG_1__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .ZN(n6472) );
  OAI21_X1 U6632 ( .B1(n5623), .B2(n6472), .A(n6478), .ZN(n5624) );
  OAI21_X1 U6633 ( .B1(n6478), .B2(n6656), .A(n5624), .ZN(U2795) );
  INV_X1 U6634 ( .A(n5712), .ZN(n5727) );
  NOR2_X1 U6635 ( .A1(n5232), .A2(n5625), .ZN(n5635) );
  AOI21_X1 U6636 ( .B1(REIP_REG_16__SCAN_IN), .B2(n5635), .A(
        REIP_REG_17__SCAN_IN), .ZN(n5627) );
  OAI22_X1 U6637 ( .A1(n5628), .A2(n5627), .B1(n5626), .B2(n5683), .ZN(n5629)
         );
  AOI211_X1 U6638 ( .C1(n5743), .C2(EBX_REG_17__SCAN_IN), .A(n5727), .B(n5629), 
        .ZN(n5632) );
  AOI22_X1 U6639 ( .A1(n5777), .A2(n2999), .B1(n5758), .B2(n5768), .ZN(n5631)
         );
  OAI211_X1 U6640 ( .C1(n5633), .C2(n5738), .A(n5632), .B(n5631), .ZN(U2810)
         );
  INV_X1 U6642 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6427) );
  OAI33_X1 U6643 ( .A1(1'b0), .A2(n5635), .A3(REIP_REG_16__SCAN_IN), .B1(n6427), .B2(n5634), .B3(n5647), .ZN(n5637) );
  OAI211_X1 U6644 ( .C1(n5683), .C2(n5638), .A(n5637), .B(n5712), .ZN(n5639)
         );
  AOI21_X1 U6645 ( .B1(EBX_REG_16__SCAN_IN), .B2(n5743), .A(n5639), .ZN(n5644)
         );
  OAI22_X1 U6646 ( .A1(n5641), .A2(n5695), .B1(n5640), .B2(n5738), .ZN(n5642)
         );
  INV_X1 U6647 ( .A(n5642), .ZN(n5643) );
  OAI211_X1 U6648 ( .C1(n5671), .C2(n5645), .A(n5644), .B(n5643), .ZN(U2811)
         );
  OR2_X1 U6649 ( .A1(n5754), .A2(n5646), .ZN(n5649) );
  AOI22_X1 U6650 ( .A1(EBX_REG_14__SCAN_IN), .A2(n5743), .B1(
        REIP_REG_14__SCAN_IN), .B2(n5647), .ZN(n5648) );
  OAI21_X1 U6651 ( .B1(n5650), .B2(n5649), .A(n5648), .ZN(n5651) );
  AOI211_X1 U6652 ( .C1(n5764), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5727), 
        .B(n5651), .ZN(n5656) );
  INV_X1 U6653 ( .A(n5652), .ZN(n5653) );
  AOI22_X1 U6654 ( .A1(n5654), .A2(n2999), .B1(n5653), .B2(n5763), .ZN(n5655)
         );
  OAI211_X1 U6655 ( .C1(n5671), .C2(n5657), .A(n5656), .B(n5655), .ZN(U2813)
         );
  INV_X1 U6656 ( .A(n5658), .ZN(n5664) );
  AOI22_X1 U6657 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n5764), .B1(
        REIP_REG_12__SCAN_IN), .B2(n5659), .ZN(n5660) );
  OAI211_X1 U6658 ( .C1(n5761), .C2(n5661), .A(n5660), .B(n5712), .ZN(n5662)
         );
  AOI211_X1 U6659 ( .C1(n5664), .C2(n5758), .A(n5663), .B(n5662), .ZN(n5667)
         );
  INV_X1 U6660 ( .A(n5665), .ZN(n5899) );
  AOI22_X1 U6661 ( .A1(n5899), .A2(n2999), .B1(n5898), .B2(n5763), .ZN(n5666)
         );
  NAND2_X1 U6662 ( .A1(n5667), .A2(n5666), .ZN(U2815) );
  AOI22_X1 U6663 ( .A1(EBX_REG_10__SCAN_IN), .A2(n5743), .B1(n5668), .B2(n6417), .ZN(n5669) );
  OAI21_X1 U6664 ( .B1(n5671), .B2(n5670), .A(n5669), .ZN(n5672) );
  AOI211_X1 U6665 ( .C1(n5764), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5727), 
        .B(n5672), .ZN(n5679) );
  INV_X1 U6666 ( .A(n5673), .ZN(n5675) );
  AOI22_X1 U6667 ( .A1(n5675), .A2(n2999), .B1(n5763), .B2(n5674), .ZN(n5678)
         );
  NOR2_X1 U6668 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5676), .ZN(n5685) );
  OAI21_X1 U6669 ( .B1(n5685), .B2(n5680), .A(REIP_REG_10__SCAN_IN), .ZN(n5677) );
  NAND3_X1 U6670 ( .A1(n5679), .A2(n5678), .A3(n5677), .ZN(U2817) );
  AOI22_X1 U6671 ( .A1(EBX_REG_9__SCAN_IN), .A2(n5743), .B1(
        REIP_REG_9__SCAN_IN), .B2(n5680), .ZN(n5681) );
  OAI211_X1 U6672 ( .C1(n5683), .C2(n5682), .A(n5681), .B(n5712), .ZN(n5684)
         );
  AOI211_X1 U6673 ( .C1(n5686), .C2(n5758), .A(n5685), .B(n5684), .ZN(n5691)
         );
  INV_X1 U6674 ( .A(n5687), .ZN(n5688) );
  AOI22_X1 U6675 ( .A1(n5689), .A2(n2999), .B1(n5763), .B2(n5688), .ZN(n5690)
         );
  NAND2_X1 U6676 ( .A1(n5691), .A2(n5690), .ZN(U2818) );
  AOI21_X1 U6677 ( .B1(n5764), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5727), 
        .ZN(n5702) );
  AOI22_X1 U6678 ( .A1(EBX_REG_7__SCAN_IN), .A2(n5743), .B1(n5758), .B2(n5931), 
        .ZN(n5701) );
  INV_X1 U6679 ( .A(n5693), .ZN(n5692) );
  OAI21_X1 U6680 ( .B1(n5692), .B2(n5754), .A(n5755), .ZN(n5717) );
  NOR3_X1 U6681 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5754), .A3(n5693), .ZN(n5704)
         );
  OAI22_X1 U6682 ( .A1(n5696), .A2(n5695), .B1(n5694), .B2(n5738), .ZN(n5697)
         );
  AOI221_X1 U6683 ( .B1(n5717), .B2(REIP_REG_7__SCAN_IN), .C1(n5704), .C2(
        REIP_REG_7__SCAN_IN), .A(n5697), .ZN(n5700) );
  INV_X1 U6684 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6413) );
  NAND3_X1 U6685 ( .A1(n5724), .A2(n5698), .A3(n6413), .ZN(n5699) );
  NAND4_X1 U6686 ( .A1(n5702), .A2(n5701), .A3(n5700), .A4(n5699), .ZN(U2820)
         );
  AOI22_X1 U6687 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n5764), .B1(n5758), 
        .B2(n5771), .ZN(n5709) );
  NOR2_X1 U6688 ( .A1(n5775), .A2(n5761), .ZN(n5703) );
  AOI211_X1 U6689 ( .C1(n5717), .C2(REIP_REG_6__SCAN_IN), .A(n5704), .B(n5703), 
        .ZN(n5708) );
  INV_X1 U6690 ( .A(n5705), .ZN(n5706) );
  AOI22_X1 U6691 ( .A1(n5773), .A2(n2999), .B1(n5706), .B2(n5763), .ZN(n5707)
         );
  NAND4_X1 U6692 ( .A1(n5709), .A2(n5708), .A3(n5707), .A4(n5712), .ZN(U2821)
         );
  AOI22_X1 U6693 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n5764), .B1(n5758), 
        .B2(n5710), .ZN(n5711) );
  OAI211_X1 U6694 ( .C1(n5761), .C2(n5713), .A(n5712), .B(n5711), .ZN(n5714)
         );
  AOI21_X1 U6695 ( .B1(n5716), .B2(n5715), .A(n5714), .ZN(n5720) );
  OAI221_X1 U6696 ( .B1(REIP_REG_5__SCAN_IN), .B2(n5724), .C1(
        REIP_REG_5__SCAN_IN), .C2(n5718), .A(n5717), .ZN(n5719) );
  OAI211_X1 U6697 ( .C1(n5738), .C2(n5721), .A(n5720), .B(n5719), .ZN(U2822)
         );
  INV_X1 U6698 ( .A(n5722), .ZN(n5739) );
  AOI21_X1 U6699 ( .B1(n5724), .B2(n5728), .A(n5723), .ZN(n5753) );
  OAI22_X1 U6700 ( .A1(n5753), .A2(n6505), .B1(n5725), .B2(n5759), .ZN(n5726)
         );
  AOI211_X1 U6701 ( .C1(n5764), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5727), 
        .B(n5726), .ZN(n5737) );
  NOR3_X1 U6702 ( .A1(REIP_REG_4__SCAN_IN), .A2(n5754), .A3(n5728), .ZN(n5735)
         );
  NAND2_X1 U6703 ( .A1(n5743), .A2(EBX_REG_4__SCAN_IN), .ZN(n5732) );
  INV_X1 U6704 ( .A(n5729), .ZN(n5730) );
  NAND2_X1 U6705 ( .A1(n5758), .A2(n5730), .ZN(n5731) );
  OAI211_X1 U6706 ( .C1(n5767), .C2(n5733), .A(n5732), .B(n5731), .ZN(n5734)
         );
  NOR2_X1 U6707 ( .A1(n5735), .A2(n5734), .ZN(n5736) );
  OAI211_X1 U6708 ( .C1(n5739), .C2(n5738), .A(n5737), .B(n5736), .ZN(U2823)
         );
  INV_X1 U6709 ( .A(n5759), .ZN(n5740) );
  NAND2_X1 U6710 ( .A1(n5740), .A2(n6101), .ZN(n5747) );
  INV_X1 U6711 ( .A(n5741), .ZN(n5742) );
  AOI22_X1 U6712 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n5764), .B1(n5763), 
        .B2(n5742), .ZN(n5746) );
  NAND2_X1 U6713 ( .A1(n5743), .A2(EBX_REG_3__SCAN_IN), .ZN(n5745) );
  NAND2_X1 U6714 ( .A1(n5758), .A2(n3016), .ZN(n5744) );
  NAND4_X1 U6715 ( .A1(n5747), .A2(n5746), .A3(n5745), .A4(n5744), .ZN(n5750)
         );
  NOR2_X1 U6716 ( .A1(n5767), .A2(n5748), .ZN(n5749) );
  NOR2_X1 U6717 ( .A1(n5750), .A2(n5749), .ZN(n5751) );
  OAI221_X1 U6718 ( .B1(n5753), .B2(n6406), .C1(n5753), .C2(n5752), .A(n5751), 
        .ZN(U2824) );
  NAND2_X1 U6719 ( .A1(n5755), .A2(n5754), .ZN(n5756) );
  AOI22_X1 U6720 ( .A1(n5758), .A2(n5757), .B1(REIP_REG_0__SCAN_IN), .B2(n5756), .ZN(n5766) );
  OAI22_X1 U6721 ( .A1(n5761), .A2(n5760), .B1(n3582), .B2(n5759), .ZN(n5762)
         );
  AOI221_X1 U6722 ( .B1(n5764), .B2(PHYADDRPOINTER_REG_0__SCAN_IN), .C1(n5763), 
        .C2(PHYADDRPOINTER_REG_0__SCAN_IN), .A(n5762), .ZN(n5765) );
  OAI211_X1 U6723 ( .C1(n5767), .C2(n5922), .A(n5766), .B(n5765), .ZN(U2827)
         );
  AOI22_X1 U6724 ( .A1(n5777), .A2(n5772), .B1(n4194), .B2(n5768), .ZN(n5769)
         );
  OAI21_X1 U6725 ( .B1(n5776), .B2(n5770), .A(n5769), .ZN(U2842) );
  AOI22_X1 U6726 ( .A1(n5773), .A2(n5772), .B1(n4194), .B2(n5771), .ZN(n5774)
         );
  OAI21_X1 U6727 ( .B1(n5776), .B2(n5775), .A(n5774), .ZN(U2853) );
  AOI22_X1 U6728 ( .A1(n5777), .A2(n5781), .B1(n5780), .B2(DATAI_17_), .ZN(
        n5779) );
  AOI22_X1 U6729 ( .A1(n5784), .A2(DATAI_1_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n5783), .ZN(n5778) );
  NAND2_X1 U6730 ( .A1(n5779), .A2(n5778), .ZN(U2874) );
  AOI22_X1 U6731 ( .A1(n5782), .A2(n5781), .B1(n5780), .B2(DATAI_16_), .ZN(
        n5786) );
  AOI22_X1 U6732 ( .A1(n5784), .A2(DATAI_0_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n5783), .ZN(n5785) );
  NAND2_X1 U6733 ( .A1(n5786), .A2(n5785), .ZN(U2875) );
  INV_X1 U6734 ( .A(UWORD_REG_14__SCAN_IN), .ZN(n6601) );
  AOI22_X1 U6735 ( .A1(EAX_REG_30__SCAN_IN), .A2(n5805), .B1(n5835), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n5788) );
  OAI21_X1 U6736 ( .B1(n6601), .B2(n5825), .A(n5788), .ZN(U2893) );
  INV_X1 U6737 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n6515) );
  AOI22_X1 U6738 ( .A1(EAX_REG_29__SCAN_IN), .A2(n5805), .B1(n5816), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n5789) );
  OAI21_X1 U6739 ( .B1(n6515), .B2(n5824), .A(n5789), .ZN(U2894) );
  INV_X1 U6740 ( .A(EAX_REG_28__SCAN_IN), .ZN(n5858) );
  AOI22_X1 U6741 ( .A1(n5816), .A2(UWORD_REG_12__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n5790) );
  OAI21_X1 U6742 ( .B1(n5858), .B2(n5809), .A(n5790), .ZN(U2895) );
  INV_X1 U6743 ( .A(EAX_REG_27__SCAN_IN), .ZN(n5856) );
  AOI22_X1 U6744 ( .A1(n5816), .A2(UWORD_REG_11__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n5791) );
  OAI21_X1 U6745 ( .B1(n5856), .B2(n5809), .A(n5791), .ZN(U2896) );
  INV_X1 U6746 ( .A(EAX_REG_26__SCAN_IN), .ZN(n5793) );
  AOI22_X1 U6747 ( .A1(n5816), .A2(UWORD_REG_10__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n5792) );
  OAI21_X1 U6748 ( .B1(n5793), .B2(n5809), .A(n5792), .ZN(U2897) );
  INV_X1 U6749 ( .A(EAX_REG_25__SCAN_IN), .ZN(n5795) );
  AOI22_X1 U6750 ( .A1(n5816), .A2(UWORD_REG_9__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n5794) );
  OAI21_X1 U6751 ( .B1(n5795), .B2(n5809), .A(n5794), .ZN(U2898) );
  INV_X1 U6752 ( .A(EAX_REG_24__SCAN_IN), .ZN(n5797) );
  AOI22_X1 U6753 ( .A1(n5816), .A2(UWORD_REG_8__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n5796) );
  OAI21_X1 U6754 ( .B1(n5797), .B2(n5809), .A(n5796), .ZN(U2899) );
  INV_X1 U6755 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6623) );
  AOI22_X1 U6756 ( .A1(n5816), .A2(UWORD_REG_7__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n5798) );
  OAI21_X1 U6757 ( .B1(n6623), .B2(n5809), .A(n5798), .ZN(U2900) );
  INV_X1 U6758 ( .A(EAX_REG_22__SCAN_IN), .ZN(n5800) );
  AOI22_X1 U6759 ( .A1(n5816), .A2(UWORD_REG_6__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n5799) );
  OAI21_X1 U6760 ( .B1(n5800), .B2(n5809), .A(n5799), .ZN(U2901) );
  INV_X1 U6761 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n6504) );
  AOI22_X1 U6762 ( .A1(EAX_REG_21__SCAN_IN), .A2(n5805), .B1(n5816), .B2(
        UWORD_REG_5__SCAN_IN), .ZN(n5801) );
  OAI21_X1 U6763 ( .B1(n6504), .B2(n5824), .A(n5801), .ZN(U2902) );
  INV_X1 U6764 ( .A(EAX_REG_20__SCAN_IN), .ZN(n5803) );
  AOI22_X1 U6765 ( .A1(n5816), .A2(UWORD_REG_4__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n5802) );
  OAI21_X1 U6766 ( .B1(n5803), .B2(n5809), .A(n5802), .ZN(U2903) );
  INV_X1 U6767 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6636) );
  AOI22_X1 U6768 ( .A1(DATAO_REG_19__SCAN_IN), .A2(n5835), .B1(n5816), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n5804) );
  OAI21_X1 U6769 ( .B1(n6636), .B2(n5809), .A(n5804), .ZN(U2904) );
  INV_X1 U6770 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n6666) );
  AOI22_X1 U6771 ( .A1(EAX_REG_18__SCAN_IN), .A2(n5805), .B1(n5816), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n5806) );
  OAI21_X1 U6772 ( .B1(n6666), .B2(n5824), .A(n5806), .ZN(U2905) );
  INV_X1 U6773 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6648) );
  AOI22_X1 U6774 ( .A1(n5816), .A2(UWORD_REG_1__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5807) );
  OAI21_X1 U6775 ( .B1(n6648), .B2(n5809), .A(n5807), .ZN(U2906) );
  INV_X1 U6776 ( .A(EAX_REG_16__SCAN_IN), .ZN(n5844) );
  AOI22_X1 U6777 ( .A1(n5816), .A2(UWORD_REG_0__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5808) );
  OAI21_X1 U6778 ( .B1(n5844), .B2(n5809), .A(n5808), .ZN(U2907) );
  INV_X1 U6779 ( .A(EAX_REG_15__SCAN_IN), .ZN(n5896) );
  AOI22_X1 U6780 ( .A1(n5816), .A2(LWORD_REG_15__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5810) );
  OAI21_X1 U6781 ( .B1(n5896), .B2(n5837), .A(n5810), .ZN(U2908) );
  AOI22_X1 U6782 ( .A1(n5816), .A2(LWORD_REG_14__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5811) );
  OAI21_X1 U6783 ( .B1(n3846), .B2(n5837), .A(n5811), .ZN(U2909) );
  AOI22_X1 U6784 ( .A1(n5816), .A2(LWORD_REG_13__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n5812) );
  OAI21_X1 U6785 ( .B1(n5813), .B2(n5837), .A(n5812), .ZN(U2910) );
  INV_X1 U6786 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n6625) );
  AOI22_X1 U6787 ( .A1(EAX_REG_12__SCAN_IN), .A2(n5814), .B1(n5816), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n5815) );
  OAI21_X1 U6788 ( .B1(n6625), .B2(n5824), .A(n5815), .ZN(U2911) );
  INV_X1 U6789 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5884) );
  AOI22_X1 U6790 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n5816), .B1(n5835), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5817) );
  OAI21_X1 U6791 ( .B1(n5884), .B2(n5837), .A(n5817), .ZN(U2912) );
  AOI22_X1 U6792 ( .A1(n5816), .A2(LWORD_REG_10__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5818) );
  OAI21_X1 U6793 ( .B1(n5819), .B2(n5837), .A(n5818), .ZN(U2913) );
  AOI22_X1 U6794 ( .A1(n5816), .A2(LWORD_REG_9__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5820) );
  OAI21_X1 U6795 ( .B1(n6670), .B2(n5837), .A(n5820), .ZN(U2914) );
  AOI22_X1 U6796 ( .A1(n5816), .A2(LWORD_REG_8__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5821) );
  OAI21_X1 U6797 ( .B1(n6620), .B2(n5837), .A(n5821), .ZN(U2915) );
  AOI22_X1 U6798 ( .A1(n5816), .A2(LWORD_REG_7__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5822) );
  OAI21_X1 U6799 ( .B1(n3638), .B2(n5837), .A(n5822), .ZN(U2916) );
  AOI22_X1 U6800 ( .A1(n5816), .A2(LWORD_REG_6__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5823) );
  OAI21_X1 U6801 ( .B1(n3630), .B2(n5837), .A(n5823), .ZN(U2917) );
  INV_X1 U6802 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n5826) );
  INV_X1 U6803 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n6640) );
  OAI222_X1 U6804 ( .A1(n5826), .A2(n5825), .B1(n5837), .B2(n3622), .C1(n5824), 
        .C2(n6640), .ZN(U2918) );
  AOI22_X1 U6805 ( .A1(n5816), .A2(LWORD_REG_4__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5827) );
  OAI21_X1 U6806 ( .B1(n5828), .B2(n5837), .A(n5827), .ZN(U2919) );
  AOI22_X1 U6807 ( .A1(n5816), .A2(LWORD_REG_3__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5829) );
  OAI21_X1 U6808 ( .B1(n5830), .B2(n5837), .A(n5829), .ZN(U2920) );
  AOI22_X1 U6809 ( .A1(n5816), .A2(LWORD_REG_2__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5831) );
  OAI21_X1 U6810 ( .B1(n5832), .B2(n5837), .A(n5831), .ZN(U2921) );
  AOI22_X1 U6811 ( .A1(n5816), .A2(LWORD_REG_1__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n5833) );
  OAI21_X1 U6812 ( .B1(n5834), .B2(n5837), .A(n5833), .ZN(U2922) );
  AOI22_X1 U6813 ( .A1(n5816), .A2(LWORD_REG_0__SCAN_IN), .B1(n5835), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5836) );
  OAI21_X1 U6814 ( .B1(n5838), .B2(n5837), .A(n5836), .ZN(U2923) );
  INV_X1 U6815 ( .A(n5839), .ZN(n6364) );
  AND2_X2 U6816 ( .A1(n5840), .A2(n6364), .ZN(n5887) );
  AND2_X1 U6817 ( .A1(n6485), .A2(READY_N), .ZN(n5841) );
  OR2_X2 U6818 ( .A1(n5842), .A2(n5841), .ZN(n5892) );
  AOI22_X1 U6819 ( .A1(n5893), .A2(DATAI_0_), .B1(UWORD_REG_0__SCAN_IN), .B2(
        n5892), .ZN(n5843) );
  OAI21_X1 U6820 ( .B1(n5844), .B2(n5895), .A(n5843), .ZN(U2924) );
  AOI22_X1 U6821 ( .A1(n5893), .A2(DATAI_1_), .B1(UWORD_REG_1__SCAN_IN), .B2(
        n5892), .ZN(n5845) );
  OAI21_X1 U6822 ( .B1(n6648), .B2(n5895), .A(n5845), .ZN(U2925) );
  AOI22_X1 U6823 ( .A1(EAX_REG_18__SCAN_IN), .A2(n5887), .B1(
        UWORD_REG_2__SCAN_IN), .B2(n5892), .ZN(n5846) );
  OAI21_X1 U6824 ( .B1(n5890), .B2(n5866), .A(n5846), .ZN(U2926) );
  AOI22_X1 U6825 ( .A1(EAX_REG_19__SCAN_IN), .A2(n5887), .B1(
        UWORD_REG_3__SCAN_IN), .B2(n5892), .ZN(n5847) );
  OAI21_X1 U6826 ( .B1(n5890), .B2(n5868), .A(n5847), .ZN(U2927) );
  AOI22_X1 U6827 ( .A1(EAX_REG_20__SCAN_IN), .A2(n5887), .B1(
        UWORD_REG_4__SCAN_IN), .B2(n5892), .ZN(n5848) );
  OAI21_X1 U6828 ( .B1(n5890), .B2(n5870), .A(n5848), .ZN(U2928) );
  AOI22_X1 U6829 ( .A1(EAX_REG_21__SCAN_IN), .A2(n5887), .B1(
        UWORD_REG_5__SCAN_IN), .B2(n5892), .ZN(n5849) );
  OAI21_X1 U6830 ( .B1(n5890), .B2(n5872), .A(n5849), .ZN(U2929) );
  AOI22_X1 U6831 ( .A1(EAX_REG_22__SCAN_IN), .A2(n5887), .B1(
        UWORD_REG_6__SCAN_IN), .B2(n5892), .ZN(n5850) );
  OAI21_X1 U6832 ( .B1(n5890), .B2(n5874), .A(n5850), .ZN(U2930) );
  AOI22_X1 U6833 ( .A1(EAX_REG_23__SCAN_IN), .A2(n5887), .B1(
        UWORD_REG_7__SCAN_IN), .B2(n5892), .ZN(n5851) );
  OAI21_X1 U6834 ( .B1(n5890), .B2(n5876), .A(n5851), .ZN(U2931) );
  AOI22_X1 U6835 ( .A1(EAX_REG_24__SCAN_IN), .A2(n5887), .B1(
        UWORD_REG_8__SCAN_IN), .B2(n5892), .ZN(n5852) );
  OAI21_X1 U6836 ( .B1(n5890), .B2(n5878), .A(n5852), .ZN(U2932) );
  AOI22_X1 U6837 ( .A1(EAX_REG_25__SCAN_IN), .A2(n5887), .B1(
        UWORD_REG_9__SCAN_IN), .B2(n5892), .ZN(n5853) );
  OAI21_X1 U6838 ( .B1(n5890), .B2(n5880), .A(n5853), .ZN(U2933) );
  AOI22_X1 U6839 ( .A1(EAX_REG_26__SCAN_IN), .A2(n5887), .B1(
        UWORD_REG_10__SCAN_IN), .B2(n5892), .ZN(n5854) );
  OAI21_X1 U6840 ( .B1(n5890), .B2(n5882), .A(n5854), .ZN(U2934) );
  AOI22_X1 U6841 ( .A1(n5893), .A2(DATAI_11_), .B1(UWORD_REG_11__SCAN_IN), 
        .B2(n5892), .ZN(n5855) );
  OAI21_X1 U6842 ( .B1(n5856), .B2(n5895), .A(n5855), .ZN(U2935) );
  AOI22_X1 U6843 ( .A1(n5893), .A2(DATAI_12_), .B1(UWORD_REG_12__SCAN_IN), 
        .B2(n5892), .ZN(n5857) );
  OAI21_X1 U6844 ( .B1(n5858), .B2(n5895), .A(n5857), .ZN(U2936) );
  AOI22_X1 U6845 ( .A1(EAX_REG_29__SCAN_IN), .A2(n5887), .B1(
        UWORD_REG_13__SCAN_IN), .B2(n5892), .ZN(n5859) );
  OAI21_X1 U6846 ( .B1(n5890), .B2(n5889), .A(n5859), .ZN(U2937) );
  INV_X1 U6847 ( .A(n5892), .ZN(n5861) );
  AOI22_X1 U6848 ( .A1(EAX_REG_30__SCAN_IN), .A2(n5887), .B1(n5893), .B2(
        DATAI_14_), .ZN(n5860) );
  OAI21_X1 U6849 ( .B1(n5861), .B2(n6601), .A(n5860), .ZN(U2938) );
  AOI22_X1 U6850 ( .A1(EAX_REG_0__SCAN_IN), .A2(n5887), .B1(
        LWORD_REG_0__SCAN_IN), .B2(n5892), .ZN(n5862) );
  OAI21_X1 U6851 ( .B1(n5890), .B2(n6603), .A(n5862), .ZN(U2939) );
  AOI22_X1 U6852 ( .A1(EAX_REG_1__SCAN_IN), .A2(n5887), .B1(
        LWORD_REG_1__SCAN_IN), .B2(n5892), .ZN(n5863) );
  OAI21_X1 U6853 ( .B1(n5890), .B2(n5864), .A(n5863), .ZN(U2940) );
  AOI22_X1 U6854 ( .A1(EAX_REG_2__SCAN_IN), .A2(n5887), .B1(
        LWORD_REG_2__SCAN_IN), .B2(n5892), .ZN(n5865) );
  OAI21_X1 U6855 ( .B1(n5890), .B2(n5866), .A(n5865), .ZN(U2941) );
  AOI22_X1 U6856 ( .A1(EAX_REG_3__SCAN_IN), .A2(n5887), .B1(
        LWORD_REG_3__SCAN_IN), .B2(n5892), .ZN(n5867) );
  OAI21_X1 U6857 ( .B1(n5890), .B2(n5868), .A(n5867), .ZN(U2942) );
  AOI22_X1 U6858 ( .A1(EAX_REG_4__SCAN_IN), .A2(n5887), .B1(
        LWORD_REG_4__SCAN_IN), .B2(n5892), .ZN(n5869) );
  OAI21_X1 U6859 ( .B1(n5890), .B2(n5870), .A(n5869), .ZN(U2943) );
  AOI22_X1 U6860 ( .A1(EAX_REG_5__SCAN_IN), .A2(n5887), .B1(
        LWORD_REG_5__SCAN_IN), .B2(n5892), .ZN(n5871) );
  OAI21_X1 U6861 ( .B1(n5890), .B2(n5872), .A(n5871), .ZN(U2944) );
  AOI22_X1 U6862 ( .A1(EAX_REG_6__SCAN_IN), .A2(n5887), .B1(
        LWORD_REG_6__SCAN_IN), .B2(n5892), .ZN(n5873) );
  OAI21_X1 U6863 ( .B1(n5890), .B2(n5874), .A(n5873), .ZN(U2945) );
  AOI22_X1 U6864 ( .A1(EAX_REG_7__SCAN_IN), .A2(n5887), .B1(
        LWORD_REG_7__SCAN_IN), .B2(n5892), .ZN(n5875) );
  OAI21_X1 U6865 ( .B1(n5890), .B2(n5876), .A(n5875), .ZN(U2946) );
  AOI22_X1 U6866 ( .A1(EAX_REG_8__SCAN_IN), .A2(n5887), .B1(
        LWORD_REG_8__SCAN_IN), .B2(n5892), .ZN(n5877) );
  OAI21_X1 U6867 ( .B1(n5890), .B2(n5878), .A(n5877), .ZN(U2947) );
  AOI22_X1 U6868 ( .A1(EAX_REG_9__SCAN_IN), .A2(n5887), .B1(
        LWORD_REG_9__SCAN_IN), .B2(n5892), .ZN(n5879) );
  OAI21_X1 U6869 ( .B1(n5890), .B2(n5880), .A(n5879), .ZN(U2948) );
  AOI22_X1 U6870 ( .A1(EAX_REG_10__SCAN_IN), .A2(n5887), .B1(
        LWORD_REG_10__SCAN_IN), .B2(n5892), .ZN(n5881) );
  OAI21_X1 U6871 ( .B1(n5890), .B2(n5882), .A(n5881), .ZN(U2949) );
  AOI22_X1 U6872 ( .A1(n5893), .A2(DATAI_11_), .B1(LWORD_REG_11__SCAN_IN), 
        .B2(n5892), .ZN(n5883) );
  OAI21_X1 U6873 ( .B1(n5884), .B2(n5895), .A(n5883), .ZN(U2950) );
  AOI22_X1 U6874 ( .A1(EAX_REG_12__SCAN_IN), .A2(n5887), .B1(
        LWORD_REG_12__SCAN_IN), .B2(n5892), .ZN(n5886) );
  NAND2_X1 U6875 ( .A1(n5893), .A2(DATAI_12_), .ZN(n5885) );
  NAND2_X1 U6876 ( .A1(n5886), .A2(n5885), .ZN(U2951) );
  AOI22_X1 U6877 ( .A1(EAX_REG_13__SCAN_IN), .A2(n5887), .B1(
        LWORD_REG_13__SCAN_IN), .B2(n5892), .ZN(n5888) );
  OAI21_X1 U6878 ( .B1(n5890), .B2(n5889), .A(n5888), .ZN(U2952) );
  AOI22_X1 U6879 ( .A1(n5893), .A2(DATAI_14_), .B1(LWORD_REG_14__SCAN_IN), 
        .B2(n5892), .ZN(n5891) );
  OAI21_X1 U6880 ( .B1(n3846), .B2(n5895), .A(n5891), .ZN(U2953) );
  AOI22_X1 U6881 ( .A1(n5893), .A2(DATAI_15_), .B1(LWORD_REG_15__SCAN_IN), 
        .B2(n5892), .ZN(n5894) );
  OAI21_X1 U6882 ( .B1(n5896), .B2(n5895), .A(n5894), .ZN(U2954) );
  AOI22_X1 U6883 ( .A1(n5917), .A2(REIP_REG_12__SCAN_IN), .B1(n5919), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5901) );
  AOI22_X1 U6884 ( .A1(n5899), .A2(n5909), .B1(n5898), .B2(n5897), .ZN(n5900)
         );
  OAI211_X1 U6885 ( .C1(n5902), .C2(n3056), .A(n5901), .B(n5900), .ZN(U2974)
         );
  AOI22_X1 U6886 ( .A1(n5917), .A2(REIP_REG_2__SCAN_IN), .B1(n5919), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5912) );
  INV_X1 U6887 ( .A(n5903), .ZN(n5910) );
  INV_X1 U6888 ( .A(n5904), .ZN(n5906) );
  NAND2_X1 U6889 ( .A1(n5906), .A2(n5905), .ZN(n5907) );
  XNOR2_X1 U6890 ( .A(n5908), .B(n5907), .ZN(n5950) );
  AOI22_X1 U6891 ( .A1(n5910), .A2(n5909), .B1(n5950), .B2(n5916), .ZN(n5911)
         );
  OAI211_X1 U6892 ( .C1(n5914), .C2(n5913), .A(n5912), .B(n5911), .ZN(U2984)
         );
  AOI22_X1 U6893 ( .A1(n5917), .A2(REIP_REG_0__SCAN_IN), .B1(n5916), .B2(n5915), .ZN(n5921) );
  OAI21_X1 U6894 ( .B1(n5919), .B2(n5918), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5920) );
  OAI211_X1 U6895 ( .C1(n5922), .C2(n6275), .A(n5921), .B(n5920), .ZN(U2986)
         );
  AOI21_X1 U6896 ( .B1(n5924), .B2(n5944), .A(n5923), .ZN(n5928) );
  AOI22_X1 U6897 ( .A1(n5926), .A2(n5951), .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n5925), .ZN(n5927) );
  OAI211_X1 U6898 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n5929), .A(n5928), .B(n5927), .ZN(U3007) );
  AOI21_X1 U6899 ( .B1(n5944), .B2(n5931), .A(n5930), .ZN(n5934) );
  NAND2_X1 U6900 ( .A1(n5932), .A2(n5951), .ZN(n5933) );
  OAI211_X1 U6901 ( .C1(n5935), .C2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n5934), 
        .B(n5933), .ZN(n5936) );
  INV_X1 U6902 ( .A(n5936), .ZN(n5937) );
  OAI21_X1 U6903 ( .B1(n2998), .B2(n5938), .A(n5937), .ZN(U3011) );
  AOI221_X1 U6904 ( .B1(n5954), .B2(n5942), .C1(n5941), .C2(n5942), .A(n5940), 
        .ZN(n5947) );
  INV_X1 U6905 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6404) );
  NAND2_X1 U6906 ( .A1(n5944), .A2(n5943), .ZN(n5945) );
  OAI21_X1 U6907 ( .B1(n6404), .B2(n6684), .A(n5945), .ZN(n5946) );
  NOR2_X1 U6908 ( .A1(n5947), .A2(n5946), .ZN(n5953) );
  NOR2_X1 U6909 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n5948), .ZN(n5949)
         );
  AOI22_X1 U6910 ( .A1(n5951), .A2(n5950), .B1(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .B2(n5949), .ZN(n5952) );
  OAI211_X1 U6911 ( .C1(n5955), .C2(n5954), .A(n5953), .B(n5952), .ZN(U3016)
         );
  NOR2_X1 U6912 ( .A1(n3525), .A2(n6466), .ZN(U3019) );
  INV_X1 U6913 ( .A(n6283), .ZN(n6236) );
  OAI22_X1 U6914 ( .A1(n6021), .A2(n5959), .B1(n5958), .B2(n6139), .ZN(n5982)
         );
  NAND3_X1 U6915 ( .A1(n6231), .A2(n6344), .A3(n6337), .ZN(n5994) );
  NOR2_X1 U6916 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5994), .ZN(n5983)
         );
  AOI22_X1 U6917 ( .A1(n6272), .A2(n5982), .B1(n6273), .B2(n5983), .ZN(n5968)
         );
  NOR2_X1 U6918 ( .A1(n5959), .A2(n6101), .ZN(n5989) );
  INV_X1 U6919 ( .A(n5960), .ZN(n5961) );
  NOR3_X1 U6920 ( .A1(n6001), .A2(n6327), .A3(n6271), .ZN(n5962) );
  INV_X1 U6921 ( .A(n6022), .ZN(n6278) );
  NOR2_X1 U6922 ( .A1(n5962), .A2(n6278), .ZN(n5966) );
  INV_X1 U6923 ( .A(n5983), .ZN(n5964) );
  AOI211_X1 U6924 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5964), .A(n6027), .B(
        n5963), .ZN(n5965) );
  AOI22_X1 U6925 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n5984), .B1(n6233), 
        .B2(n6327), .ZN(n5967) );
  OAI211_X1 U6926 ( .C1(n6236), .C2(n6017), .A(n5968), .B(n5967), .ZN(U3020)
         );
  AOI22_X1 U6927 ( .A1(n6287), .A2(n5982), .B1(n6288), .B2(n5983), .ZN(n5970)
         );
  AOI22_X1 U6928 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n5984), .B1(n6289), 
        .B2(n6001), .ZN(n5969) );
  OAI211_X1 U6929 ( .C1(n6292), .C2(n5979), .A(n5970), .B(n5969), .ZN(U3021)
         );
  AOI22_X1 U6930 ( .A1(n6294), .A2(n5983), .B1(n6293), .B2(n5982), .ZN(n5972)
         );
  AOI22_X1 U6931 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(n5984), .B1(n6295), 
        .B2(n6001), .ZN(n5971) );
  OAI211_X1 U6932 ( .C1(n6298), .C2(n5979), .A(n5972), .B(n5971), .ZN(U3022)
         );
  AOI22_X1 U6933 ( .A1(n6299), .A2(n5982), .B1(n6300), .B2(n5983), .ZN(n5974)
         );
  AOI22_X1 U6934 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n5984), .B1(n6301), 
        .B2(n6001), .ZN(n5973) );
  OAI211_X1 U6935 ( .C1(n6304), .C2(n5979), .A(n5974), .B(n5973), .ZN(U3023)
         );
  AOI22_X1 U6936 ( .A1(n6306), .A2(n5983), .B1(n6305), .B2(n5982), .ZN(n5976)
         );
  AOI22_X1 U6937 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n5984), .B1(n6307), 
        .B2(n6001), .ZN(n5975) );
  OAI211_X1 U6938 ( .C1(n6310), .C2(n5979), .A(n5976), .B(n5975), .ZN(U3024)
         );
  AOI22_X1 U6939 ( .A1(n6312), .A2(n5983), .B1(n6311), .B2(n5982), .ZN(n5978)
         );
  AOI22_X1 U6940 ( .A1(INSTQUEUE_REG_0__5__SCAN_IN), .A2(n5984), .B1(n6313), 
        .B2(n6001), .ZN(n5977) );
  OAI211_X1 U6941 ( .C1(n6316), .C2(n5979), .A(n5978), .B(n5977), .ZN(U3025)
         );
  INV_X1 U6942 ( .A(n6319), .ZN(n6260) );
  AOI22_X1 U6943 ( .A1(n6318), .A2(n5983), .B1(n6317), .B2(n5982), .ZN(n5981)
         );
  AOI22_X1 U6944 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(n5984), .B1(n6257), 
        .B2(n6327), .ZN(n5980) );
  OAI211_X1 U6945 ( .C1(n6260), .C2(n6017), .A(n5981), .B(n5980), .ZN(U3026)
         );
  INV_X1 U6946 ( .A(n6328), .ZN(n6268) );
  AOI22_X1 U6947 ( .A1(n6326), .A2(n5983), .B1(n6324), .B2(n5982), .ZN(n5986)
         );
  AOI22_X1 U6948 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n5984), .B1(n6264), 
        .B2(n6327), .ZN(n5985) );
  OAI211_X1 U6949 ( .C1(n6268), .C2(n6017), .A(n5986), .B(n5985), .ZN(U3027)
         );
  NOR2_X1 U6950 ( .A1(n6468), .A2(n5994), .ZN(n6012) );
  AOI22_X1 U6951 ( .A1(n6233), .A2(n6001), .B1(n6273), .B2(n6012), .ZN(n5998)
         );
  INV_X1 U6952 ( .A(n5987), .ZN(n5988) );
  OAI21_X1 U6953 ( .B1(n5988), .B2(n6224), .A(n6464), .ZN(n5995) );
  NAND2_X1 U6954 ( .A1(n5989), .A2(n6461), .ZN(n5991) );
  INV_X1 U6955 ( .A(n6012), .ZN(n5990) );
  AND2_X1 U6956 ( .A1(n5991), .A2(n5990), .ZN(n5996) );
  INV_X1 U6957 ( .A(n5996), .ZN(n5993) );
  AOI21_X1 U6958 ( .B1(n6271), .B2(n5994), .A(n6191), .ZN(n5992) );
  OAI21_X1 U6959 ( .B1(n5995), .B2(n5993), .A(n5992), .ZN(n6014) );
  OAI22_X1 U6960 ( .A1(n5996), .A2(n5995), .B1(n6367), .B2(n5994), .ZN(n6013)
         );
  AOI22_X1 U6961 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n6014), .B1(n6272), 
        .B2(n6013), .ZN(n5997) );
  OAI211_X1 U6962 ( .C1(n6049), .C2(n6236), .A(n5998), .B(n5997), .ZN(U3028)
         );
  INV_X1 U6963 ( .A(n6289), .ZN(n6240) );
  AOI22_X1 U6964 ( .A1(n6237), .A2(n6001), .B1(n6288), .B2(n6012), .ZN(n6000)
         );
  AOI22_X1 U6965 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n6014), .B1(n6287), 
        .B2(n6013), .ZN(n5999) );
  OAI211_X1 U6966 ( .C1(n6049), .C2(n6240), .A(n6000), .B(n5999), .ZN(U3029)
         );
  INV_X1 U6967 ( .A(n6295), .ZN(n6244) );
  AOI22_X1 U6968 ( .A1(n6294), .A2(n6012), .B1(n6001), .B2(n6241), .ZN(n6003)
         );
  AOI22_X1 U6969 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n6014), .B1(n6293), 
        .B2(n6013), .ZN(n6002) );
  OAI211_X1 U6970 ( .C1(n6049), .C2(n6244), .A(n6003), .B(n6002), .ZN(U3030)
         );
  AOI22_X1 U6971 ( .A1(n6023), .A2(n6301), .B1(n6300), .B2(n6012), .ZN(n6005)
         );
  AOI22_X1 U6972 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n6014), .B1(n6299), 
        .B2(n6013), .ZN(n6004) );
  OAI211_X1 U6973 ( .C1(n6304), .C2(n6017), .A(n6005), .B(n6004), .ZN(U3031)
         );
  AOI22_X1 U6974 ( .A1(n6306), .A2(n6012), .B1(n6023), .B2(n6307), .ZN(n6007)
         );
  AOI22_X1 U6975 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n6014), .B1(n6305), 
        .B2(n6013), .ZN(n6006) );
  OAI211_X1 U6976 ( .C1(n6310), .C2(n6017), .A(n6007), .B(n6006), .ZN(U3032)
         );
  AOI22_X1 U6977 ( .A1(n6312), .A2(n6012), .B1(n6023), .B2(n6313), .ZN(n6009)
         );
  AOI22_X1 U6978 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n6014), .B1(n6311), 
        .B2(n6013), .ZN(n6008) );
  OAI211_X1 U6979 ( .C1(n6316), .C2(n6017), .A(n6009), .B(n6008), .ZN(U3033)
         );
  AOI22_X1 U6980 ( .A1(n6318), .A2(n6012), .B1(n6023), .B2(n6319), .ZN(n6011)
         );
  AOI22_X1 U6981 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n6014), .B1(n6317), 
        .B2(n6013), .ZN(n6010) );
  OAI211_X1 U6982 ( .C1(n6322), .C2(n6017), .A(n6011), .B(n6010), .ZN(U3034)
         );
  AOI22_X1 U6983 ( .A1(n6326), .A2(n6012), .B1(n6023), .B2(n6328), .ZN(n6016)
         );
  AOI22_X1 U6984 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n6014), .B1(n6324), 
        .B2(n6013), .ZN(n6015) );
  OAI211_X1 U6985 ( .C1(n6333), .C2(n6017), .A(n6016), .B(n6015), .ZN(U3035)
         );
  NOR2_X1 U6986 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6018), .ZN(n6044)
         );
  INV_X1 U6987 ( .A(n6024), .ZN(n6020) );
  OAI22_X1 U6988 ( .A1(n6021), .A2(n6020), .B1(n6019), .B2(n6139), .ZN(n6043)
         );
  AOI22_X1 U6989 ( .A1(n6044), .A2(n6273), .B1(n6272), .B2(n6043), .ZN(n6030)
         );
  OAI21_X1 U6990 ( .B1(n6023), .B2(n6045), .A(n6022), .ZN(n6026) );
  NAND2_X1 U6991 ( .A1(n6051), .A2(n6024), .ZN(n6025) );
  AOI21_X1 U6992 ( .B1(n6026), .B2(n6025), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n6028) );
  NOR2_X1 U6993 ( .A1(n6027), .A2(n6228), .ZN(n6136) );
  AOI22_X1 U6994 ( .A1(n6046), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n6045), 
        .B2(n6283), .ZN(n6029) );
  OAI211_X1 U6995 ( .C1(n6286), .C2(n6049), .A(n6030), .B(n6029), .ZN(U3036)
         );
  AOI22_X1 U6996 ( .A1(n6044), .A2(n6288), .B1(n6287), .B2(n6043), .ZN(n6032)
         );
  AOI22_X1 U6997 ( .A1(n6046), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n6045), 
        .B2(n6289), .ZN(n6031) );
  OAI211_X1 U6998 ( .C1(n6049), .C2(n6292), .A(n6032), .B(n6031), .ZN(U3037)
         );
  AOI22_X1 U6999 ( .A1(n6294), .A2(n6044), .B1(n6293), .B2(n6043), .ZN(n6034)
         );
  AOI22_X1 U7000 ( .A1(n6046), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n6045), 
        .B2(n6295), .ZN(n6033) );
  OAI211_X1 U7001 ( .C1(n6049), .C2(n6298), .A(n6034), .B(n6033), .ZN(U3038)
         );
  AOI22_X1 U7002 ( .A1(n6044), .A2(n6300), .B1(n6299), .B2(n6043), .ZN(n6036)
         );
  AOI22_X1 U7003 ( .A1(n6046), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n6045), 
        .B2(n6301), .ZN(n6035) );
  OAI211_X1 U7004 ( .C1(n6049), .C2(n6304), .A(n6036), .B(n6035), .ZN(U3039)
         );
  AOI22_X1 U7005 ( .A1(n6306), .A2(n6044), .B1(n6305), .B2(n6043), .ZN(n6038)
         );
  AOI22_X1 U7006 ( .A1(n6046), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n6045), 
        .B2(n6307), .ZN(n6037) );
  OAI211_X1 U7007 ( .C1(n6049), .C2(n6310), .A(n6038), .B(n6037), .ZN(U3040)
         );
  AOI22_X1 U7008 ( .A1(n6312), .A2(n6044), .B1(n6311), .B2(n6043), .ZN(n6040)
         );
  AOI22_X1 U7009 ( .A1(n6046), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n6045), 
        .B2(n6313), .ZN(n6039) );
  OAI211_X1 U7010 ( .C1(n6049), .C2(n6316), .A(n6040), .B(n6039), .ZN(U3041)
         );
  AOI22_X1 U7011 ( .A1(n6318), .A2(n6044), .B1(n6317), .B2(n6043), .ZN(n6042)
         );
  AOI22_X1 U7012 ( .A1(n6046), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n6045), 
        .B2(n6319), .ZN(n6041) );
  OAI211_X1 U7013 ( .C1(n6049), .C2(n6322), .A(n6042), .B(n6041), .ZN(U3042)
         );
  AOI22_X1 U7014 ( .A1(n6326), .A2(n6044), .B1(n6324), .B2(n6043), .ZN(n6048)
         );
  AOI22_X1 U7015 ( .A1(n6046), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n6045), 
        .B2(n6328), .ZN(n6047) );
  OAI211_X1 U7016 ( .C1(n6049), .C2(n6333), .A(n6048), .B(n6047), .ZN(U3043)
         );
  NOR2_X1 U7017 ( .A1(n6050), .A2(n6271), .ZN(n6056) );
  INV_X1 U7018 ( .A(n6222), .ZN(n6270) );
  NAND3_X1 U7019 ( .A1(n6270), .A2(n6051), .A3(n6461), .ZN(n6052) );
  NAND2_X1 U7020 ( .A1(n6052), .A2(n6053), .ZN(n6054) );
  AOI22_X1 U7021 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6058), .B1(n6056), .B2(
        n6054), .ZN(n6086) );
  INV_X1 U7022 ( .A(n6272), .ZN(n6061) );
  INV_X1 U7023 ( .A(n6053), .ZN(n6081) );
  AOI22_X1 U7024 ( .A1(n6273), .A2(n6081), .B1(n6283), .B2(n6097), .ZN(n6060)
         );
  INV_X1 U7025 ( .A(n6054), .ZN(n6055) );
  NAND2_X1 U7026 ( .A1(n6056), .A2(n6055), .ZN(n6057) );
  OAI211_X1 U7027 ( .C1(n6464), .C2(n6058), .A(n6057), .B(n6281), .ZN(n6082)
         );
  AOI22_X1 U7028 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6082), .B1(n6233), 
        .B2(n6080), .ZN(n6059) );
  OAI211_X1 U7029 ( .C1(n6086), .C2(n6061), .A(n6060), .B(n6059), .ZN(U3076)
         );
  INV_X1 U7030 ( .A(n6287), .ZN(n6064) );
  AOI22_X1 U7031 ( .A1(n6288), .A2(n6081), .B1(n6289), .B2(n6097), .ZN(n6063)
         );
  AOI22_X1 U7032 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6082), .B1(n6237), 
        .B2(n6080), .ZN(n6062) );
  OAI211_X1 U7033 ( .C1(n6086), .C2(n6064), .A(n6063), .B(n6062), .ZN(U3077)
         );
  INV_X1 U7034 ( .A(n6293), .ZN(n6067) );
  AOI22_X1 U7035 ( .A1(n6294), .A2(n6081), .B1(n6295), .B2(n6097), .ZN(n6066)
         );
  AOI22_X1 U7036 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6082), .B1(n6241), 
        .B2(n6080), .ZN(n6065) );
  OAI211_X1 U7037 ( .C1(n6086), .C2(n6067), .A(n6066), .B(n6065), .ZN(U3078)
         );
  INV_X1 U7038 ( .A(n6299), .ZN(n6070) );
  AOI22_X1 U7039 ( .A1(n6081), .A2(n6300), .B1(n6245), .B2(n6080), .ZN(n6069)
         );
  AOI22_X1 U7040 ( .A1(n6082), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n6301), 
        .B2(n6097), .ZN(n6068) );
  OAI211_X1 U7041 ( .C1(n6086), .C2(n6070), .A(n6069), .B(n6068), .ZN(U3079)
         );
  INV_X1 U7042 ( .A(n6305), .ZN(n6073) );
  AOI22_X1 U7043 ( .A1(n6306), .A2(n6081), .B1(n6249), .B2(n6080), .ZN(n6072)
         );
  AOI22_X1 U7044 ( .A1(n6082), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n6307), 
        .B2(n6097), .ZN(n6071) );
  OAI211_X1 U7045 ( .C1(n6086), .C2(n6073), .A(n6072), .B(n6071), .ZN(U3080)
         );
  INV_X1 U7046 ( .A(n6311), .ZN(n6076) );
  AOI22_X1 U7047 ( .A1(n6312), .A2(n6081), .B1(n6313), .B2(n6097), .ZN(n6075)
         );
  AOI22_X1 U7048 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6082), .B1(n6253), 
        .B2(n6080), .ZN(n6074) );
  OAI211_X1 U7049 ( .C1(n6086), .C2(n6076), .A(n6075), .B(n6074), .ZN(U3081)
         );
  INV_X1 U7050 ( .A(n6317), .ZN(n6079) );
  AOI22_X1 U7051 ( .A1(n6318), .A2(n6081), .B1(n6319), .B2(n6097), .ZN(n6078)
         );
  AOI22_X1 U7052 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6082), .B1(n6257), 
        .B2(n6080), .ZN(n6077) );
  OAI211_X1 U7053 ( .C1(n6086), .C2(n6079), .A(n6078), .B(n6077), .ZN(U3082)
         );
  INV_X1 U7054 ( .A(n6324), .ZN(n6085) );
  AOI22_X1 U7055 ( .A1(n6326), .A2(n6081), .B1(n6264), .B2(n6080), .ZN(n6084)
         );
  AOI22_X1 U7056 ( .A1(n6082), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n6328), 
        .B2(n6097), .ZN(n6083) );
  OAI211_X1 U7057 ( .C1(n6086), .C2(n6085), .A(n6084), .B(n6083), .ZN(U3083)
         );
  AOI22_X1 U7058 ( .A1(n6272), .A2(n6095), .B1(n6273), .B2(n6096), .ZN(n6088)
         );
  AOI22_X1 U7059 ( .A1(n6098), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6233), 
        .B2(n6097), .ZN(n6087) );
  OAI211_X1 U7060 ( .C1(n6236), .C2(n6125), .A(n6088), .B(n6087), .ZN(U3084)
         );
  AOI22_X1 U7061 ( .A1(n6287), .A2(n6095), .B1(n6288), .B2(n6096), .ZN(n6090)
         );
  AOI22_X1 U7062 ( .A1(n6098), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6237), 
        .B2(n6097), .ZN(n6089) );
  OAI211_X1 U7063 ( .C1(n6240), .C2(n6125), .A(n6090), .B(n6089), .ZN(U3085)
         );
  AOI22_X1 U7064 ( .A1(n6294), .A2(n6096), .B1(n6293), .B2(n6095), .ZN(n6092)
         );
  AOI22_X1 U7065 ( .A1(n6098), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6241), 
        .B2(n6097), .ZN(n6091) );
  OAI211_X1 U7066 ( .C1(n6244), .C2(n6125), .A(n6092), .B(n6091), .ZN(U3086)
         );
  AOI22_X1 U7067 ( .A1(n6318), .A2(n6096), .B1(n6317), .B2(n6095), .ZN(n6094)
         );
  AOI22_X1 U7068 ( .A1(n6098), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6257), 
        .B2(n6097), .ZN(n6093) );
  OAI211_X1 U7069 ( .C1(n6260), .C2(n6125), .A(n6094), .B(n6093), .ZN(U3090)
         );
  AOI22_X1 U7070 ( .A1(n6326), .A2(n6096), .B1(n6324), .B2(n6095), .ZN(n6100)
         );
  AOI22_X1 U7071 ( .A1(n6098), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6264), 
        .B2(n6097), .ZN(n6099) );
  OAI211_X1 U7072 ( .C1(n6268), .C2(n6125), .A(n6100), .B(n6099), .ZN(U3091)
         );
  INV_X1 U7073 ( .A(n6162), .ZN(n6122) );
  NOR2_X1 U7074 ( .A1(n6468), .A2(n6107), .ZN(n6127) );
  AOI22_X1 U7075 ( .A1(n6283), .A2(n6122), .B1(n6273), .B2(n6127), .ZN(n6111)
         );
  AND2_X1 U7076 ( .A1(n6101), .A2(n6461), .ZN(n6269) );
  AOI21_X1 U7077 ( .B1(n6269), .B2(n6102), .A(n6127), .ZN(n6109) );
  INV_X1 U7078 ( .A(n6109), .ZN(n6106) );
  INV_X1 U7079 ( .A(n6103), .ZN(n6104) );
  OAI21_X1 U7080 ( .B1(n6104), .B2(n6224), .A(n6464), .ZN(n6108) );
  AOI21_X1 U7081 ( .B1(n6271), .B2(n6107), .A(n6191), .ZN(n6105) );
  OAI21_X1 U7082 ( .B1(n6106), .B2(n6108), .A(n6105), .ZN(n6129) );
  OAI22_X1 U7083 ( .A1(n6109), .A2(n6108), .B1(n6367), .B2(n6107), .ZN(n6128)
         );
  AOI22_X1 U7084 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n6129), .B1(n6272), 
        .B2(n6128), .ZN(n6110) );
  OAI211_X1 U7085 ( .C1(n6286), .C2(n6125), .A(n6111), .B(n6110), .ZN(U3092)
         );
  AOI22_X1 U7086 ( .A1(n6237), .A2(n6126), .B1(n6288), .B2(n6127), .ZN(n6113)
         );
  AOI22_X1 U7087 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n6129), .B1(n6287), 
        .B2(n6128), .ZN(n6112) );
  OAI211_X1 U7088 ( .C1(n6240), .C2(n6162), .A(n6113), .B(n6112), .ZN(U3093)
         );
  AOI22_X1 U7089 ( .A1(n6294), .A2(n6127), .B1(n6122), .B2(n6295), .ZN(n6115)
         );
  AOI22_X1 U7090 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n6129), .B1(n6293), 
        .B2(n6128), .ZN(n6114) );
  OAI211_X1 U7091 ( .C1(n6298), .C2(n6125), .A(n6115), .B(n6114), .ZN(U3094)
         );
  AOI22_X1 U7092 ( .A1(n6301), .A2(n6122), .B1(n6300), .B2(n6127), .ZN(n6117)
         );
  AOI22_X1 U7093 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n6129), .B1(n6299), 
        .B2(n6128), .ZN(n6116) );
  OAI211_X1 U7094 ( .C1(n6304), .C2(n6125), .A(n6117), .B(n6116), .ZN(U3095)
         );
  AOI22_X1 U7095 ( .A1(n6306), .A2(n6127), .B1(n6126), .B2(n6249), .ZN(n6119)
         );
  AOI22_X1 U7096 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n6129), .B1(n6305), 
        .B2(n6128), .ZN(n6118) );
  OAI211_X1 U7097 ( .C1(n6252), .C2(n6162), .A(n6119), .B(n6118), .ZN(U3096)
         );
  AOI22_X1 U7098 ( .A1(n6312), .A2(n6127), .B1(n6122), .B2(n6313), .ZN(n6121)
         );
  AOI22_X1 U7099 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n6129), .B1(n6311), 
        .B2(n6128), .ZN(n6120) );
  OAI211_X1 U7100 ( .C1(n6316), .C2(n6125), .A(n6121), .B(n6120), .ZN(U3097)
         );
  AOI22_X1 U7101 ( .A1(n6318), .A2(n6127), .B1(n6122), .B2(n6319), .ZN(n6124)
         );
  AOI22_X1 U7102 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n6129), .B1(n6317), 
        .B2(n6128), .ZN(n6123) );
  OAI211_X1 U7103 ( .C1(n6322), .C2(n6125), .A(n6124), .B(n6123), .ZN(U3098)
         );
  AOI22_X1 U7104 ( .A1(n6326), .A2(n6127), .B1(n6126), .B2(n6264), .ZN(n6131)
         );
  AOI22_X1 U7105 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n6129), .B1(n6324), 
        .B2(n6128), .ZN(n6130) );
  OAI211_X1 U7106 ( .C1(n6268), .C2(n6162), .A(n6131), .B(n6130), .ZN(U3099)
         );
  NOR2_X1 U7107 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6132), .ZN(n6157)
         );
  AOI22_X1 U7108 ( .A1(n6283), .A2(n6156), .B1(n6273), .B2(n6157), .ZN(n6143)
         );
  NAND2_X1 U7109 ( .A1(n6174), .A2(n6162), .ZN(n6133) );
  AOI21_X1 U7110 ( .B1(n6133), .B2(STATEBS16_REG_SCAN_IN), .A(n6271), .ZN(
        n6137) );
  INV_X1 U7111 ( .A(n6157), .ZN(n6134) );
  AOI22_X1 U7112 ( .A1(n6137), .A2(n6140), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n6134), .ZN(n6135) );
  OAI211_X1 U7113 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6367), .A(n6136), .B(n6135), .ZN(n6159) );
  INV_X1 U7114 ( .A(n6137), .ZN(n6141) );
  NAND2_X1 U7115 ( .A1(n6138), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6220) );
  OAI22_X1 U7116 ( .A1(n6141), .A2(n6140), .B1(n6139), .B2(n6220), .ZN(n6158)
         );
  AOI22_X1 U7117 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n6159), .B1(n6272), 
        .B2(n6158), .ZN(n6142) );
  OAI211_X1 U7118 ( .C1(n6286), .C2(n6162), .A(n6143), .B(n6142), .ZN(U3100)
         );
  AOI22_X1 U7119 ( .A1(n6289), .A2(n6156), .B1(n6288), .B2(n6157), .ZN(n6145)
         );
  AOI22_X1 U7120 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n6159), .B1(n6287), 
        .B2(n6158), .ZN(n6144) );
  OAI211_X1 U7121 ( .C1(n6292), .C2(n6162), .A(n6145), .B(n6144), .ZN(U3101)
         );
  AOI22_X1 U7122 ( .A1(n6294), .A2(n6157), .B1(n6295), .B2(n6156), .ZN(n6147)
         );
  AOI22_X1 U7123 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(n6159), .B1(n6293), 
        .B2(n6158), .ZN(n6146) );
  OAI211_X1 U7124 ( .C1(n6298), .C2(n6162), .A(n6147), .B(n6146), .ZN(U3102)
         );
  AOI22_X1 U7125 ( .A1(n6301), .A2(n6156), .B1(n6300), .B2(n6157), .ZN(n6149)
         );
  AOI22_X1 U7126 ( .A1(INSTQUEUE_REG_10__3__SCAN_IN), .A2(n6159), .B1(n6299), 
        .B2(n6158), .ZN(n6148) );
  OAI211_X1 U7127 ( .C1(n6304), .C2(n6162), .A(n6149), .B(n6148), .ZN(U3103)
         );
  AOI22_X1 U7128 ( .A1(n6306), .A2(n6157), .B1(n6307), .B2(n6156), .ZN(n6151)
         );
  AOI22_X1 U7129 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n6159), .B1(n6305), 
        .B2(n6158), .ZN(n6150) );
  OAI211_X1 U7130 ( .C1(n6310), .C2(n6162), .A(n6151), .B(n6150), .ZN(U3104)
         );
  AOI22_X1 U7131 ( .A1(n6312), .A2(n6157), .B1(n6313), .B2(n6156), .ZN(n6153)
         );
  AOI22_X1 U7132 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n6159), .B1(n6311), 
        .B2(n6158), .ZN(n6152) );
  OAI211_X1 U7133 ( .C1(n6316), .C2(n6162), .A(n6153), .B(n6152), .ZN(U3105)
         );
  AOI22_X1 U7134 ( .A1(n6318), .A2(n6157), .B1(n6319), .B2(n6156), .ZN(n6155)
         );
  AOI22_X1 U7135 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n6159), .B1(n6317), 
        .B2(n6158), .ZN(n6154) );
  OAI211_X1 U7136 ( .C1(n6322), .C2(n6162), .A(n6155), .B(n6154), .ZN(U3106)
         );
  AOI22_X1 U7137 ( .A1(n6326), .A2(n6157), .B1(n6328), .B2(n6156), .ZN(n6161)
         );
  AOI22_X1 U7138 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n6159), .B1(n6324), 
        .B2(n6158), .ZN(n6160) );
  OAI211_X1 U7139 ( .C1(n6333), .C2(n6162), .A(n6161), .B(n6160), .ZN(U3107)
         );
  AOI22_X1 U7140 ( .A1(n6294), .A2(n6169), .B1(n6295), .B2(n6181), .ZN(n6164)
         );
  AOI22_X1 U7141 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6171), .B1(n6293), 
        .B2(n6170), .ZN(n6163) );
  OAI211_X1 U7142 ( .C1(n6298), .C2(n6174), .A(n6164), .B(n6163), .ZN(U3110)
         );
  AOI22_X1 U7143 ( .A1(n6300), .A2(n6169), .B1(n6301), .B2(n6181), .ZN(n6166)
         );
  AOI22_X1 U7144 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6171), .B1(n6299), 
        .B2(n6170), .ZN(n6165) );
  OAI211_X1 U7145 ( .C1(n6304), .C2(n6174), .A(n6166), .B(n6165), .ZN(U3111)
         );
  AOI22_X1 U7146 ( .A1(n6306), .A2(n6169), .B1(n6307), .B2(n6181), .ZN(n6168)
         );
  AOI22_X1 U7147 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6171), .B1(n6305), 
        .B2(n6170), .ZN(n6167) );
  OAI211_X1 U7148 ( .C1(n6310), .C2(n6174), .A(n6168), .B(n6167), .ZN(U3112)
         );
  AOI22_X1 U7149 ( .A1(n6326), .A2(n6169), .B1(n6328), .B2(n6181), .ZN(n6173)
         );
  AOI22_X1 U7150 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6171), .B1(n6324), 
        .B2(n6170), .ZN(n6172) );
  OAI211_X1 U7151 ( .C1(n6333), .C2(n6174), .A(n6173), .B(n6172), .ZN(U3115)
         );
  AOI22_X1 U7152 ( .A1(n6272), .A2(n6179), .B1(n6273), .B2(n6180), .ZN(n6176)
         );
  AOI22_X1 U7153 ( .A1(n6182), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n6233), 
        .B2(n6181), .ZN(n6175) );
  OAI211_X1 U7154 ( .C1(n6236), .C2(n6211), .A(n6176), .B(n6175), .ZN(U3116)
         );
  AOI22_X1 U7155 ( .A1(n6287), .A2(n6179), .B1(n6288), .B2(n6180), .ZN(n6178)
         );
  AOI22_X1 U7156 ( .A1(n6182), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n6237), 
        .B2(n6181), .ZN(n6177) );
  OAI211_X1 U7157 ( .C1(n6240), .C2(n6211), .A(n6178), .B(n6177), .ZN(U3117)
         );
  AOI22_X1 U7158 ( .A1(n6294), .A2(n6180), .B1(n6293), .B2(n6179), .ZN(n6184)
         );
  AOI22_X1 U7159 ( .A1(n6182), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n6241), 
        .B2(n6181), .ZN(n6183) );
  OAI211_X1 U7160 ( .C1(n6244), .C2(n6211), .A(n6184), .B(n6183), .ZN(U3118)
         );
  NOR2_X1 U7161 ( .A1(n6468), .A2(n6194), .ZN(n6213) );
  AOI22_X1 U7162 ( .A1(n6283), .A2(n6263), .B1(n6273), .B2(n6213), .ZN(n6198)
         );
  NAND2_X1 U7163 ( .A1(n6464), .A2(n6186), .ZN(n6195) );
  INV_X1 U7164 ( .A(n6187), .ZN(n6188) );
  NAND2_X1 U7165 ( .A1(n6188), .A2(n6269), .ZN(n6190) );
  INV_X1 U7166 ( .A(n6213), .ZN(n6189) );
  AND2_X1 U7167 ( .A1(n6190), .A2(n6189), .ZN(n6196) );
  INV_X1 U7168 ( .A(n6196), .ZN(n6193) );
  AOI21_X1 U7169 ( .B1(n6271), .B2(n6194), .A(n6191), .ZN(n6192) );
  OAI21_X1 U7170 ( .B1(n6195), .B2(n6193), .A(n6192), .ZN(n6215) );
  OAI22_X1 U7171 ( .A1(n6196), .A2(n6195), .B1(n6367), .B2(n6194), .ZN(n6214)
         );
  AOI22_X1 U7172 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n6215), .B1(n6272), 
        .B2(n6214), .ZN(n6197) );
  OAI211_X1 U7173 ( .C1(n6286), .C2(n6211), .A(n6198), .B(n6197), .ZN(U3124)
         );
  AOI22_X1 U7174 ( .A1(n6237), .A2(n6212), .B1(n6288), .B2(n6213), .ZN(n6200)
         );
  AOI22_X1 U7175 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n6215), .B1(n6287), 
        .B2(n6214), .ZN(n6199) );
  OAI211_X1 U7176 ( .C1(n6240), .C2(n6225), .A(n6200), .B(n6199), .ZN(U3125)
         );
  AOI22_X1 U7177 ( .A1(n6294), .A2(n6213), .B1(n6241), .B2(n6212), .ZN(n6202)
         );
  AOI22_X1 U7178 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n6215), .B1(n6293), 
        .B2(n6214), .ZN(n6201) );
  OAI211_X1 U7179 ( .C1(n6244), .C2(n6225), .A(n6202), .B(n6201), .ZN(U3126)
         );
  AOI22_X1 U7180 ( .A1(n6245), .A2(n6212), .B1(n6300), .B2(n6213), .ZN(n6204)
         );
  AOI22_X1 U7181 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n6215), .B1(n6299), 
        .B2(n6214), .ZN(n6203) );
  OAI211_X1 U7182 ( .C1(n6248), .C2(n6225), .A(n6204), .B(n6203), .ZN(U3127)
         );
  AOI22_X1 U7183 ( .A1(n6306), .A2(n6213), .B1(n6249), .B2(n6212), .ZN(n6206)
         );
  AOI22_X1 U7184 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n6215), .B1(n6305), 
        .B2(n6214), .ZN(n6205) );
  OAI211_X1 U7185 ( .C1(n6252), .C2(n6225), .A(n6206), .B(n6205), .ZN(U3128)
         );
  AOI22_X1 U7186 ( .A1(n6312), .A2(n6213), .B1(n6253), .B2(n6212), .ZN(n6208)
         );
  AOI22_X1 U7187 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n6215), .B1(n6311), 
        .B2(n6214), .ZN(n6207) );
  OAI211_X1 U7188 ( .C1(n6256), .C2(n6225), .A(n6208), .B(n6207), .ZN(U3129)
         );
  AOI22_X1 U7189 ( .A1(n6318), .A2(n6213), .B1(n6319), .B2(n6263), .ZN(n6210)
         );
  AOI22_X1 U7190 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n6215), .B1(n6317), 
        .B2(n6214), .ZN(n6209) );
  OAI211_X1 U7191 ( .C1(n6322), .C2(n6211), .A(n6210), .B(n6209), .ZN(U3130)
         );
  AOI22_X1 U7192 ( .A1(n6326), .A2(n6213), .B1(n6264), .B2(n6212), .ZN(n6217)
         );
  AOI22_X1 U7193 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n6215), .B1(n6324), 
        .B2(n6214), .ZN(n6216) );
  OAI211_X1 U7194 ( .C1(n6268), .C2(n6225), .A(n6217), .B(n6216), .ZN(U3131)
         );
  INV_X1 U7195 ( .A(n6218), .ZN(n6219) );
  OAI22_X1 U7196 ( .A1(n6223), .A2(n6222), .B1(n6221), .B2(n6220), .ZN(n6261)
         );
  NOR2_X1 U7197 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6274), .ZN(n6262)
         );
  AOI22_X1 U7198 ( .A1(n6272), .A2(n6261), .B1(n6273), .B2(n6262), .ZN(n6235)
         );
  INV_X1 U7199 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6231) );
  AOI21_X1 U7200 ( .B1(n6225), .B2(n6332), .A(n6224), .ZN(n6226) );
  NOR2_X1 U7201 ( .A1(n6227), .A2(n6226), .ZN(n6229) );
  NOR4_X1 U7202 ( .A1(n6231), .A2(n6230), .A3(n6229), .A4(n6228), .ZN(n6232)
         );
  AOI22_X1 U7203 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n6265), .B1(n6233), 
        .B2(n6263), .ZN(n6234) );
  OAI211_X1 U7204 ( .C1(n6236), .C2(n6332), .A(n6235), .B(n6234), .ZN(U3132)
         );
  AOI22_X1 U7205 ( .A1(n6287), .A2(n6261), .B1(n6288), .B2(n6262), .ZN(n6239)
         );
  AOI22_X1 U7206 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n6265), .B1(n6237), 
        .B2(n6263), .ZN(n6238) );
  OAI211_X1 U7207 ( .C1(n6240), .C2(n6332), .A(n6239), .B(n6238), .ZN(U3133)
         );
  AOI22_X1 U7208 ( .A1(n6294), .A2(n6262), .B1(n6293), .B2(n6261), .ZN(n6243)
         );
  AOI22_X1 U7209 ( .A1(INSTQUEUE_REG_14__2__SCAN_IN), .A2(n6265), .B1(n6241), 
        .B2(n6263), .ZN(n6242) );
  OAI211_X1 U7210 ( .C1(n6244), .C2(n6332), .A(n6243), .B(n6242), .ZN(U3134)
         );
  AOI22_X1 U7211 ( .A1(n6299), .A2(n6261), .B1(n6300), .B2(n6262), .ZN(n6247)
         );
  AOI22_X1 U7212 ( .A1(INSTQUEUE_REG_14__3__SCAN_IN), .A2(n6265), .B1(n6245), 
        .B2(n6263), .ZN(n6246) );
  OAI211_X1 U7213 ( .C1(n6248), .C2(n6332), .A(n6247), .B(n6246), .ZN(U3135)
         );
  AOI22_X1 U7214 ( .A1(n6306), .A2(n6262), .B1(n6305), .B2(n6261), .ZN(n6251)
         );
  AOI22_X1 U7215 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n6265), .B1(n6249), 
        .B2(n6263), .ZN(n6250) );
  OAI211_X1 U7216 ( .C1(n6252), .C2(n6332), .A(n6251), .B(n6250), .ZN(U3136)
         );
  AOI22_X1 U7217 ( .A1(n6312), .A2(n6262), .B1(n6311), .B2(n6261), .ZN(n6255)
         );
  AOI22_X1 U7218 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n6265), .B1(n6253), 
        .B2(n6263), .ZN(n6254) );
  OAI211_X1 U7219 ( .C1(n6256), .C2(n6332), .A(n6255), .B(n6254), .ZN(U3137)
         );
  AOI22_X1 U7220 ( .A1(n6318), .A2(n6262), .B1(n6317), .B2(n6261), .ZN(n6259)
         );
  AOI22_X1 U7221 ( .A1(INSTQUEUE_REG_14__6__SCAN_IN), .A2(n6265), .B1(n6257), 
        .B2(n6263), .ZN(n6258) );
  OAI211_X1 U7222 ( .C1(n6260), .C2(n6332), .A(n6259), .B(n6258), .ZN(U3138)
         );
  AOI22_X1 U7223 ( .A1(n6326), .A2(n6262), .B1(n6324), .B2(n6261), .ZN(n6267)
         );
  AOI22_X1 U7224 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n6265), .B1(n6264), 
        .B2(n6263), .ZN(n6266) );
  OAI211_X1 U7225 ( .C1(n6268), .C2(n6332), .A(n6267), .B(n6266), .ZN(U3139)
         );
  AOI21_X1 U7226 ( .B1(n6270), .B2(n6269), .A(n6325), .ZN(n6277) );
  OAI22_X1 U7227 ( .A1(n6277), .A2(n6271), .B1(n6274), .B2(n6367), .ZN(n6323)
         );
  AOI22_X1 U7228 ( .A1(n6325), .A2(n6273), .B1(n6272), .B2(n6323), .ZN(n6285)
         );
  INV_X1 U7229 ( .A(n6274), .ZN(n6282) );
  AOI21_X1 U7230 ( .B1(n6276), .B2(n4526), .A(n6275), .ZN(n6279) );
  OAI21_X1 U7231 ( .B1(n6279), .B2(n6278), .A(n6277), .ZN(n6280) );
  OAI211_X1 U7232 ( .C1(n6282), .C2(n6464), .A(n6281), .B(n6280), .ZN(n6329)
         );
  AOI22_X1 U7233 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6329), .B1(n6283), 
        .B2(n6327), .ZN(n6284) );
  OAI211_X1 U7234 ( .C1(n6286), .C2(n6332), .A(n6285), .B(n6284), .ZN(U3140)
         );
  AOI22_X1 U7235 ( .A1(n6325), .A2(n6288), .B1(n6287), .B2(n6323), .ZN(n6291)
         );
  AOI22_X1 U7236 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n6329), .B1(n6289), 
        .B2(n6327), .ZN(n6290) );
  OAI211_X1 U7237 ( .C1(n6292), .C2(n6332), .A(n6291), .B(n6290), .ZN(U3141)
         );
  AOI22_X1 U7238 ( .A1(n6294), .A2(n6325), .B1(n6293), .B2(n6323), .ZN(n6297)
         );
  AOI22_X1 U7239 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n6329), .B1(n6295), 
        .B2(n6327), .ZN(n6296) );
  OAI211_X1 U7240 ( .C1(n6298), .C2(n6332), .A(n6297), .B(n6296), .ZN(U3142)
         );
  AOI22_X1 U7241 ( .A1(n6325), .A2(n6300), .B1(n6299), .B2(n6323), .ZN(n6303)
         );
  AOI22_X1 U7242 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n6329), .B1(n6301), 
        .B2(n6327), .ZN(n6302) );
  OAI211_X1 U7243 ( .C1(n6304), .C2(n6332), .A(n6303), .B(n6302), .ZN(U3143)
         );
  AOI22_X1 U7244 ( .A1(n6306), .A2(n6325), .B1(n6305), .B2(n6323), .ZN(n6309)
         );
  AOI22_X1 U7245 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n6329), .B1(n6307), 
        .B2(n6327), .ZN(n6308) );
  OAI211_X1 U7246 ( .C1(n6310), .C2(n6332), .A(n6309), .B(n6308), .ZN(U3144)
         );
  AOI22_X1 U7247 ( .A1(n6312), .A2(n6325), .B1(n6311), .B2(n6323), .ZN(n6315)
         );
  AOI22_X1 U7248 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6329), .B1(n6313), 
        .B2(n6327), .ZN(n6314) );
  OAI211_X1 U7249 ( .C1(n6316), .C2(n6332), .A(n6315), .B(n6314), .ZN(U3145)
         );
  AOI22_X1 U7250 ( .A1(n6318), .A2(n6325), .B1(n6317), .B2(n6323), .ZN(n6321)
         );
  AOI22_X1 U7251 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n6329), .B1(n6319), 
        .B2(n6327), .ZN(n6320) );
  OAI211_X1 U7252 ( .C1(n6322), .C2(n6332), .A(n6321), .B(n6320), .ZN(U3146)
         );
  AOI22_X1 U7253 ( .A1(n6326), .A2(n6325), .B1(n6324), .B2(n6323), .ZN(n6331)
         );
  AOI22_X1 U7254 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6329), .B1(n6328), 
        .B2(n6327), .ZN(n6330) );
  OAI211_X1 U7255 ( .C1(n6333), .C2(n6332), .A(n6331), .B(n6330), .ZN(U3147)
         );
  OAI211_X1 U7256 ( .C1(n3090), .C2(n6335), .A(n6334), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6338) );
  OAI21_X1 U7257 ( .B1(n6337), .B2(n6338), .A(n6336), .ZN(n6340) );
  NAND2_X1 U7258 ( .A1(n6338), .A2(n6337), .ZN(n6339) );
  OAI21_X1 U7259 ( .B1(n6341), .B2(n6340), .A(n6339), .ZN(n6342) );
  AOI222_X1 U7260 ( .A1(n6344), .A2(n6343), .B1(n6344), .B2(n6342), .C1(n6343), 
        .C2(n6342), .ZN(n6347) );
  INV_X1 U7261 ( .A(n6345), .ZN(n6346) );
  AOI222_X1 U7262 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6347), .B1(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6346), .C1(n6347), .C2(n6346), 
        .ZN(n6357) );
  INV_X1 U7263 ( .A(n6348), .ZN(n6354) );
  INV_X1 U7264 ( .A(n6349), .ZN(n6353) );
  OAI21_X1 U7265 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6350), 
        .ZN(n6351) );
  NAND4_X1 U7266 ( .A1(n6354), .A2(n6353), .A3(n6352), .A4(n6351), .ZN(n6355)
         );
  AOI211_X1 U7267 ( .C1(n6357), .C2(n3525), .A(n6356), .B(n6355), .ZN(n6373)
         );
  INV_X1 U7268 ( .A(n6358), .ZN(n6463) );
  AOI21_X1 U7269 ( .B1(n6463), .B2(n6360), .A(n6359), .ZN(n6372) );
  AOI22_X1 U7270 ( .A1(n6373), .A2(n6361), .B1(READY_N), .B2(n5816), .ZN(n6362) );
  AOI21_X1 U7271 ( .B1(n6364), .B2(n6363), .A(n6362), .ZN(n6365) );
  AOI21_X1 U7272 ( .B1(n6486), .B2(n6366), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n6370) );
  NAND2_X1 U7273 ( .A1(READY_N), .A2(n6367), .ZN(n6381) );
  AOI21_X1 U7274 ( .B1(n6381), .B2(n6457), .A(n6368), .ZN(n6369) );
  AOI21_X1 U7275 ( .B1(n6457), .B2(n6370), .A(n6369), .ZN(n6371) );
  OAI211_X1 U7276 ( .C1(n6373), .C2(n6374), .A(n6372), .B(n6371), .ZN(U3148)
         );
  OAI21_X1 U7277 ( .B1(READY_N), .B2(n6375), .A(n6374), .ZN(n6379) );
  AOI211_X1 U7278 ( .C1(n6457), .C2(n6381), .A(n6385), .B(n6376), .ZN(n6377)
         );
  AOI211_X1 U7279 ( .C1(n6457), .C2(n6379), .A(n6378), .B(n6377), .ZN(n6380)
         );
  INV_X1 U7280 ( .A(n6380), .ZN(U3149) );
  NAND3_X1 U7281 ( .A1(n6382), .A2(n6381), .A3(n6456), .ZN(n6384) );
  OAI21_X1 U7282 ( .B1(n6385), .B2(n6384), .A(n6383), .ZN(U3150) );
  AND2_X1 U7283 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6452), .ZN(U3151) );
  AND2_X1 U7284 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6452), .ZN(U3152) );
  AND2_X1 U7285 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6452), .ZN(U3153) );
  AND2_X1 U7286 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6452), .ZN(U3154) );
  INV_X1 U7287 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6635) );
  NOR2_X1 U7288 ( .A1(n6455), .A2(n6635), .ZN(U3155) );
  AND2_X1 U7289 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6452), .ZN(U3156) );
  INV_X1 U7290 ( .A(DATAWIDTH_REG_25__SCAN_IN), .ZN(n6618) );
  NOR2_X1 U7291 ( .A1(n6455), .A2(n6618), .ZN(U3157) );
  AND2_X1 U7292 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6452), .ZN(U3158) );
  AND2_X1 U7293 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6452), .ZN(U3159) );
  AND2_X1 U7294 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6452), .ZN(U3160) );
  AND2_X1 U7295 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6452), .ZN(U3161) );
  INV_X1 U7296 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6638) );
  NOR2_X1 U7297 ( .A1(n6455), .A2(n6638), .ZN(U3162) );
  AND2_X1 U7298 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6452), .ZN(U3163) );
  AND2_X1 U7299 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6452), .ZN(U3164) );
  AND2_X1 U7300 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6452), .ZN(U3165) );
  AND2_X1 U7301 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6452), .ZN(U3166) );
  INV_X1 U7302 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6668) );
  NOR2_X1 U7303 ( .A1(n6455), .A2(n6668), .ZN(U3167) );
  AND2_X1 U7304 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6452), .ZN(U3168) );
  AND2_X1 U7305 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6452), .ZN(U3169) );
  AND2_X1 U7306 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6452), .ZN(U3170) );
  AND2_X1 U7307 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6452), .ZN(U3171) );
  AND2_X1 U7308 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6452), .ZN(U3172) );
  AND2_X1 U7309 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6452), .ZN(U3173) );
  AND2_X1 U7310 ( .A1(n6452), .A2(DATAWIDTH_REG_8__SCAN_IN), .ZN(U3174) );
  AND2_X1 U7311 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6452), .ZN(U3175) );
  AND2_X1 U7312 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6452), .ZN(U3176) );
  AND2_X1 U7313 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6452), .ZN(U3177) );
  AND2_X1 U7314 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6452), .ZN(U3178) );
  AND2_X1 U7315 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6452), .ZN(U3179) );
  AND2_X1 U7316 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6452), .ZN(U3180) );
  AOI22_X1 U7317 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .B1(
        STATE_REG_1__SCAN_IN), .B2(READY_N), .ZN(n6399) );
  AND2_X1 U7318 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6389) );
  INV_X1 U7319 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6387) );
  INV_X1 U7320 ( .A(NA_N), .ZN(n6396) );
  AOI211_X1 U7321 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6396), .A(
        STATE_REG_0__SCAN_IN), .B(n6395), .ZN(n6401) );
  AOI221_X1 U7322 ( .B1(n6389), .B2(n6480), .C1(n6387), .C2(n6480), .A(n6401), 
        .ZN(n6386) );
  OAI21_X1 U7323 ( .B1(n6395), .B2(n6399), .A(n6386), .ZN(U3181) );
  NOR2_X1 U7324 ( .A1(n6393), .A2(n6387), .ZN(n6397) );
  NAND2_X1 U7325 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6388) );
  OAI21_X1 U7326 ( .B1(n6397), .B2(n6389), .A(n6388), .ZN(n6390) );
  OAI211_X1 U7327 ( .C1(n6392), .C2(n6483), .A(n6391), .B(n6390), .ZN(U3182)
         );
  AOI221_X1 U7328 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6483), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6394) );
  AOI221_X1 U7329 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6394), .C2(HOLD), .A(n6393), .ZN(n6400) );
  AOI21_X1 U7330 ( .B1(n6397), .B2(n6396), .A(n6395), .ZN(n6398) );
  OAI22_X1 U7331 ( .A1(n6401), .A2(n6400), .B1(n6399), .B2(n6398), .ZN(U3183)
         );
  NAND2_X1 U7332 ( .A1(n6491), .A2(n6529), .ZN(n6449) );
  INV_X1 U7333 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6622) );
  INV_X1 U7334 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U7335 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6491), .ZN(n6445) );
  OAI222_X1 U7336 ( .A1(n6449), .A2(n6404), .B1(n6622), .B2(n6491), .C1(n6402), 
        .C2(n6445), .ZN(U3184) );
  AOI22_X1 U7337 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6443), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6480), .ZN(n6403) );
  OAI21_X1 U7338 ( .B1(n6404), .B2(n6445), .A(n6403), .ZN(U3185) );
  AOI22_X1 U7339 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6443), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6480), .ZN(n6405) );
  OAI21_X1 U7340 ( .B1(n6406), .B2(n6445), .A(n6405), .ZN(U3186) );
  AOI22_X1 U7341 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6443), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6480), .ZN(n6407) );
  OAI21_X1 U7342 ( .B1(n6505), .B2(n6445), .A(n6407), .ZN(U3187) );
  INV_X1 U7343 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6409) );
  AOI22_X1 U7344 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6443), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6480), .ZN(n6408) );
  OAI21_X1 U7345 ( .B1(n6409), .B2(n6445), .A(n6408), .ZN(U3188) );
  AOI22_X1 U7346 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6443), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6480), .ZN(n6410) );
  OAI21_X1 U7347 ( .B1(n6411), .B2(n6445), .A(n6410), .ZN(U3189) );
  AOI22_X1 U7348 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6443), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6480), .ZN(n6412) );
  OAI21_X1 U7349 ( .B1(n6413), .B2(n6445), .A(n6412), .ZN(U3190) );
  AOI22_X1 U7350 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6443), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6480), .ZN(n6414) );
  OAI21_X1 U7351 ( .B1(n6415), .B2(n6445), .A(n6414), .ZN(U3191) );
  INV_X1 U7352 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6652) );
  OAI222_X1 U7353 ( .A1(n6445), .A2(n6416), .B1(n6652), .B2(n6491), .C1(n6417), 
        .C2(n6449), .ZN(U3192) );
  INV_X1 U7354 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n6665) );
  INV_X1 U7355 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6419) );
  OAI222_X1 U7356 ( .A1(n6445), .A2(n6417), .B1(n6665), .B2(n6491), .C1(n6419), 
        .C2(n6449), .ZN(U3193) );
  AOI22_X1 U7357 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6443), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6480), .ZN(n6418) );
  OAI21_X1 U7358 ( .B1(n6419), .B2(n6445), .A(n6418), .ZN(U3194) );
  AOI22_X1 U7359 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6443), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6480), .ZN(n6420) );
  OAI21_X1 U7360 ( .B1(n6421), .B2(n6445), .A(n6420), .ZN(U3195) );
  AOI22_X1 U7361 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6443), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6480), .ZN(n6422) );
  OAI21_X1 U7362 ( .B1(n6633), .B2(n6445), .A(n6422), .ZN(U3196) );
  AOI22_X1 U7363 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6443), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6480), .ZN(n6423) );
  OAI21_X1 U7364 ( .B1(n6424), .B2(n6445), .A(n6423), .ZN(U3197) );
  AOI22_X1 U7365 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6443), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6480), .ZN(n6425) );
  OAI21_X1 U7366 ( .B1(n5232), .B2(n6445), .A(n6425), .ZN(U3198) );
  AOI22_X1 U7367 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6443), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6480), .ZN(n6426) );
  OAI21_X1 U7368 ( .B1(n6427), .B2(n6445), .A(n6426), .ZN(U3199) );
  INV_X1 U7369 ( .A(n6445), .ZN(n6447) );
  AOI22_X1 U7370 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6447), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6480), .ZN(n6428) );
  OAI21_X1 U7371 ( .B1(n6429), .B2(n6449), .A(n6428), .ZN(U3200) );
  AOI22_X1 U7372 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6447), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6480), .ZN(n6430) );
  OAI21_X1 U7373 ( .B1(n6685), .B2(n6449), .A(n6430), .ZN(U3201) );
  AOI22_X1 U7374 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6443), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6480), .ZN(n6431) );
  OAI21_X1 U7375 ( .B1(n6685), .B2(n6445), .A(n6431), .ZN(U3202) );
  AOI22_X1 U7376 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6447), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6480), .ZN(n6432) );
  OAI21_X1 U7377 ( .B1(n6433), .B2(n6449), .A(n6432), .ZN(U3203) );
  INV_X1 U7378 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6604) );
  OAI222_X1 U7379 ( .A1(n6445), .A2(n6433), .B1(n6604), .B2(n6491), .C1(n6434), 
        .C2(n6449), .ZN(U3204) );
  INV_X1 U7380 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6641) );
  OAI222_X1 U7381 ( .A1(n6445), .A2(n6434), .B1(n6641), .B2(n6491), .C1(n4265), 
        .C2(n6449), .ZN(U3205) );
  AOI22_X1 U7382 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6447), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6480), .ZN(n6435) );
  OAI21_X1 U7383 ( .B1(n6436), .B2(n6449), .A(n6435), .ZN(U3206) );
  INV_X1 U7384 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6632) );
  OAI222_X1 U7385 ( .A1(n6449), .A2(n6438), .B1(n6632), .B2(n6491), .C1(n6436), 
        .C2(n6445), .ZN(U3207) );
  AOI22_X1 U7386 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6443), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6480), .ZN(n6437) );
  OAI21_X1 U7387 ( .B1(n6438), .B2(n6445), .A(n6437), .ZN(U3208) );
  AOI22_X1 U7388 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6447), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6480), .ZN(n6439) );
  OAI21_X1 U7389 ( .B1(n6440), .B2(n6449), .A(n6439), .ZN(U3209) );
  INV_X1 U7390 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6514) );
  AOI22_X1 U7391 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6447), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6480), .ZN(n6441) );
  OAI21_X1 U7392 ( .B1(n6514), .B2(n6449), .A(n6441), .ZN(U3210) );
  AOI22_X1 U7393 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6443), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6480), .ZN(n6442) );
  OAI21_X1 U7394 ( .B1(n6514), .B2(n6445), .A(n6442), .ZN(U3211) );
  INV_X1 U7395 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6446) );
  AOI22_X1 U7396 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6443), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6480), .ZN(n6444) );
  OAI21_X1 U7397 ( .B1(n6446), .B2(n6445), .A(n6444), .ZN(U3212) );
  AOI22_X1 U7398 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6447), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6480), .ZN(n6448) );
  OAI21_X1 U7399 ( .B1(n6450), .B2(n6449), .A(n6448), .ZN(U3213) );
  MUX2_X1 U7400 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6491), .Z(U3445) );
  MUX2_X1 U7401 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6491), .Z(U3446) );
  MUX2_X1 U7402 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6491), .Z(U3447) );
  MUX2_X1 U7403 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6491), .Z(U3448) );
  INV_X1 U7404 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6471) );
  INV_X1 U7405 ( .A(n6453), .ZN(n6451) );
  AOI21_X1 U7406 ( .B1(n6471), .B2(n6452), .A(n6451), .ZN(U3451) );
  INV_X1 U7407 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6454) );
  OAI21_X1 U7408 ( .B1(n6455), .B2(n6454), .A(n6453), .ZN(U3452) );
  OAI221_X1 U7409 ( .B1(n6458), .B2(STATE2_REG_0__SCAN_IN), .C1(n6458), .C2(
        n6457), .A(n6456), .ZN(U3453) );
  INV_X1 U7410 ( .A(n6466), .ZN(n6469) );
  INV_X1 U7411 ( .A(n6459), .ZN(n6460) );
  AOI222_X1 U7412 ( .A1(n6465), .A2(n6464), .B1(n6463), .B2(n6462), .C1(n6461), 
        .C2(n6460), .ZN(n6467) );
  AOI22_X1 U7413 ( .A1(n6469), .A2(n6468), .B1(n6467), .B2(n6466), .ZN(U3465)
         );
  NOR3_X1 U7414 ( .A1(n6471), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_0__SCAN_IN), .ZN(n6470) );
  AOI221_X1 U7415 ( .B1(n6472), .B2(n6471), .C1(REIP_REG_0__SCAN_IN), .C2(
        REIP_REG_1__SCAN_IN), .A(n6470), .ZN(n6474) );
  INV_X1 U7416 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6473) );
  INV_X1 U7417 ( .A(n6478), .ZN(n6475) );
  AOI22_X1 U7418 ( .A1(n6478), .A2(n6474), .B1(n6473), .B2(n6475), .ZN(U3468)
         );
  NOR2_X1 U7419 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6477) );
  INV_X1 U7420 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6476) );
  AOI22_X1 U7421 ( .A1(n6478), .A2(n6477), .B1(n6476), .B2(n6475), .ZN(U3469)
         );
  NAND2_X1 U7422 ( .A1(n6480), .A2(W_R_N_REG_SCAN_IN), .ZN(n6479) );
  OAI21_X1 U7423 ( .B1(n6480), .B2(READREQUEST_REG_SCAN_IN), .A(n6479), .ZN(
        U3470) );
  AOI211_X1 U7424 ( .C1(n6483), .C2(n5816), .A(n6482), .B(n6481), .ZN(n6490)
         );
  OAI211_X1 U7425 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6485), .A(
        STATE2_REG_2__SCAN_IN), .B(n6484), .ZN(n6487) );
  AOI21_X1 U7426 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6487), .A(n6486), .ZN(
        n6489) );
  NAND2_X1 U7427 ( .A1(n6490), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6488) );
  OAI21_X1 U7428 ( .B1(n6490), .B2(n6489), .A(n6488), .ZN(U3472) );
  MUX2_X1 U7429 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6491), .Z(U3473) );
  INV_X1 U7430 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n6617) );
  INV_X1 U7431 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n6607) );
  AOI22_X1 U7432 ( .A1(n6617), .A2(keyinput100), .B1(keyinput114), .B2(n6607), 
        .ZN(n6492) );
  OAI221_X1 U7433 ( .B1(n6617), .B2(keyinput100), .C1(n6607), .C2(keyinput114), 
        .A(n6492), .ZN(n6500) );
  AOI22_X1 U7434 ( .A1(n6640), .A2(keyinput96), .B1(n6626), .B2(keyinput109), 
        .ZN(n6493) );
  OAI221_X1 U7435 ( .B1(n6640), .B2(keyinput96), .C1(n6626), .C2(keyinput109), 
        .A(n6493), .ZN(n6499) );
  INV_X1 U7436 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n6495) );
  AOI22_X1 U7437 ( .A1(n4729), .A2(keyinput72), .B1(keyinput90), .B2(n6495), 
        .ZN(n6494) );
  OAI221_X1 U7438 ( .B1(n4729), .B2(keyinput72), .C1(n6495), .C2(keyinput90), 
        .A(n6494), .ZN(n6498) );
  AOI22_X1 U7439 ( .A1(n6662), .A2(keyinput71), .B1(n6653), .B2(keyinput94), 
        .ZN(n6496) );
  OAI221_X1 U7440 ( .B1(n6662), .B2(keyinput71), .C1(n6653), .C2(keyinput94), 
        .A(n6496), .ZN(n6497) );
  NOR4_X1 U7441 ( .A1(n6500), .A2(n6499), .A3(n6498), .A4(n6497), .ZN(n6537)
         );
  AOI22_X1 U7442 ( .A1(ADDRESS_REG_21__SCAN_IN), .A2(keyinput118), .B1(
        EBX_REG_20__SCAN_IN), .B2(keyinput81), .ZN(n6501) );
  OAI221_X1 U7443 ( .B1(ADDRESS_REG_21__SCAN_IN), .B2(keyinput118), .C1(
        EBX_REG_20__SCAN_IN), .C2(keyinput81), .A(n6501), .ZN(n6510) );
  AOI22_X1 U7444 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(keyinput99), .B1(
        DATAO_REG_19__SCAN_IN), .B2(keyinput74), .ZN(n6502) );
  OAI221_X1 U7445 ( .B1(DATAWIDTH_REG_25__SCAN_IN), .B2(keyinput99), .C1(
        DATAO_REG_19__SCAN_IN), .C2(keyinput74), .A(n6502), .ZN(n6509) );
  AOI22_X1 U7446 ( .A1(n6505), .A2(keyinput105), .B1(keyinput85), .B2(n6504), 
        .ZN(n6503) );
  OAI221_X1 U7447 ( .B1(n6505), .B2(keyinput105), .C1(n6504), .C2(keyinput85), 
        .A(n6503), .ZN(n6508) );
  AOI22_X1 U7448 ( .A1(n6666), .A2(keyinput77), .B1(n6636), .B2(keyinput119), 
        .ZN(n6506) );
  OAI221_X1 U7449 ( .B1(n6666), .B2(keyinput77), .C1(n6636), .C2(keyinput119), 
        .A(n6506), .ZN(n6507) );
  NOR4_X1 U7450 ( .A1(n6510), .A2(n6509), .A3(n6508), .A4(n6507), .ZN(n6536)
         );
  INV_X1 U7451 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6512) );
  AOI22_X1 U7452 ( .A1(n6512), .A2(keyinput124), .B1(keyinput91), .B2(n6668), 
        .ZN(n6511) );
  OAI221_X1 U7453 ( .B1(n6512), .B2(keyinput124), .C1(n6668), .C2(keyinput91), 
        .A(n6511), .ZN(n6522) );
  AOI22_X1 U7454 ( .A1(n6515), .A2(keyinput70), .B1(n6514), .B2(keyinput107), 
        .ZN(n6513) );
  OAI221_X1 U7455 ( .B1(n6515), .B2(keyinput70), .C1(n6514), .C2(keyinput107), 
        .A(n6513), .ZN(n6521) );
  AOI22_X1 U7456 ( .A1(n6517), .A2(keyinput66), .B1(keyinput84), .B2(n6603), 
        .ZN(n6516) );
  OAI221_X1 U7457 ( .B1(n6517), .B2(keyinput66), .C1(n6603), .C2(keyinput84), 
        .A(n6516), .ZN(n6520) );
  AOI22_X1 U7458 ( .A1(n3522), .A2(keyinput65), .B1(keyinput117), .B2(n6633), 
        .ZN(n6518) );
  OAI221_X1 U7459 ( .B1(n3522), .B2(keyinput65), .C1(n6633), .C2(keyinput117), 
        .A(n6518), .ZN(n6519) );
  NOR4_X1 U7460 ( .A1(n6522), .A2(n6521), .A3(n6520), .A4(n6519), .ZN(n6535)
         );
  AOI22_X1 U7461 ( .A1(n6665), .A2(keyinput86), .B1(keyinput79), .B2(n6656), 
        .ZN(n6523) );
  OAI221_X1 U7462 ( .B1(n6665), .B2(keyinput86), .C1(n6656), .C2(keyinput79), 
        .A(n6523), .ZN(n6533) );
  AOI22_X1 U7463 ( .A1(n6525), .A2(keyinput101), .B1(keyinput68), .B2(n6601), 
        .ZN(n6524) );
  OAI221_X1 U7464 ( .B1(n6525), .B2(keyinput101), .C1(n6601), .C2(keyinput68), 
        .A(n6524), .ZN(n6532) );
  INV_X1 U7465 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n6527) );
  AOI22_X1 U7466 ( .A1(n6652), .A2(keyinput127), .B1(n6527), .B2(keyinput126), 
        .ZN(n6526) );
  OAI221_X1 U7467 ( .B1(n6652), .B2(keyinput127), .C1(n6527), .C2(keyinput126), 
        .A(n6526), .ZN(n6531) );
  AOI22_X1 U7468 ( .A1(n6529), .A2(keyinput102), .B1(keyinput108), .B2(n6685), 
        .ZN(n6528) );
  OAI221_X1 U7469 ( .B1(n6529), .B2(keyinput102), .C1(n6685), .C2(keyinput108), 
        .A(n6528), .ZN(n6530) );
  NOR4_X1 U7470 ( .A1(n6533), .A2(n6532), .A3(n6531), .A4(n6530), .ZN(n6534)
         );
  AND4_X1 U7471 ( .A1(n6537), .A2(n6536), .A3(n6535), .A4(n6534), .ZN(n6683)
         );
  OAI22_X1 U7472 ( .A1(INSTQUEUE_REG_8__3__SCAN_IN), .A2(keyinput88), .B1(
        keyinput104), .B2(DATAI_7_), .ZN(n6538) );
  AOI221_X1 U7473 ( .B1(INSTQUEUE_REG_8__3__SCAN_IN), .B2(keyinput88), .C1(
        DATAI_7_), .C2(keyinput104), .A(n6538), .ZN(n6545) );
  OAI22_X1 U7474 ( .A1(EBX_REG_15__SCAN_IN), .A2(keyinput64), .B1(
        DATAO_REG_12__SCAN_IN), .B2(keyinput67), .ZN(n6539) );
  AOI221_X1 U7475 ( .B1(EBX_REG_15__SCAN_IN), .B2(keyinput64), .C1(keyinput67), 
        .C2(DATAO_REG_12__SCAN_IN), .A(n6539), .ZN(n6544) );
  OAI22_X1 U7476 ( .A1(EBX_REG_30__SCAN_IN), .A2(keyinput112), .B1(
        DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput73), .ZN(n6540) );
  AOI221_X1 U7477 ( .B1(EBX_REG_30__SCAN_IN), .B2(keyinput112), .C1(keyinput73), .C2(DATAWIDTH_REG_20__SCAN_IN), .A(n6540), .ZN(n6543) );
  OAI22_X1 U7478 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(keyinput113), .B1(
        keyinput98), .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n6541) );
  AOI221_X1 U7479 ( .B1(INSTQUEUE_REG_6__1__SCAN_IN), .B2(keyinput113), .C1(
        INSTQUEUE_REG_13__6__SCAN_IN), .C2(keyinput98), .A(n6541), .ZN(n6542)
         );
  NAND4_X1 U7480 ( .A1(n6545), .A2(n6544), .A3(n6543), .A4(n6542), .ZN(n6573)
         );
  OAI22_X1 U7481 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(keyinput69), .B1(
        keyinput116), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6546) );
  AOI221_X1 U7482 ( .B1(INSTQUEUE_REG_9__4__SCAN_IN), .B2(keyinput69), .C1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .C2(keyinput116), .A(n6546), .ZN(
        n6553) );
  OAI22_X1 U7483 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(keyinput111), 
        .B1(keyinput92), .B2(ADDRESS_REG_0__SCAN_IN), .ZN(n6547) );
  AOI221_X1 U7484 ( .B1(INSTADDRPOINTER_REG_24__SCAN_IN), .B2(keyinput111), 
        .C1(ADDRESS_REG_0__SCAN_IN), .C2(keyinput92), .A(n6547), .ZN(n6552) );
  OAI22_X1 U7485 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(keyinput83), .B1(
        keyinput80), .B2(ADDRESS_REG_20__SCAN_IN), .ZN(n6548) );
  AOI221_X1 U7486 ( .B1(INSTQUEUE_REG_7__5__SCAN_IN), .B2(keyinput83), .C1(
        ADDRESS_REG_20__SCAN_IN), .C2(keyinput80), .A(n6548), .ZN(n6551) );
  OAI22_X1 U7487 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(keyinput106), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(keyinput93), .ZN(n6549) );
  AOI221_X1 U7488 ( .B1(INSTQUEUE_REG_7__3__SCAN_IN), .B2(keyinput106), .C1(
        keyinput93), .C2(ADDRESS_REG_23__SCAN_IN), .A(n6549), .ZN(n6550) );
  NAND4_X1 U7489 ( .A1(n6553), .A2(n6552), .A3(n6551), .A4(n6550), .ZN(n6572)
         );
  OAI22_X1 U7490 ( .A1(EAX_REG_8__SCAN_IN), .A2(keyinput97), .B1(
        LWORD_REG_11__SCAN_IN), .B2(keyinput75), .ZN(n6554) );
  AOI221_X1 U7491 ( .B1(EAX_REG_8__SCAN_IN), .B2(keyinput97), .C1(keyinput75), 
        .C2(LWORD_REG_11__SCAN_IN), .A(n6554), .ZN(n6561) );
  OAI22_X1 U7492 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(keyinput122), .B1(
        DATAWIDTH_REG_27__SCAN_IN), .B2(keyinput110), .ZN(n6555) );
  AOI221_X1 U7493 ( .B1(INSTQUEUE_REG_15__0__SCAN_IN), .B2(keyinput122), .C1(
        keyinput110), .C2(DATAWIDTH_REG_27__SCAN_IN), .A(n6555), .ZN(n6560) );
  OAI22_X1 U7494 ( .A1(EAX_REG_23__SCAN_IN), .A2(keyinput78), .B1(
        DATAWIDTH_REG_8__SCAN_IN), .B2(keyinput125), .ZN(n6556) );
  AOI221_X1 U7495 ( .B1(EAX_REG_23__SCAN_IN), .B2(keyinput78), .C1(keyinput125), .C2(DATAWIDTH_REG_8__SCAN_IN), .A(n6556), .ZN(n6559) );
  OAI22_X1 U7496 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(keyinput120), .B1(
        keyinput121), .B2(EAX_REG_10__SCAN_IN), .ZN(n6557) );
  AOI221_X1 U7497 ( .B1(INSTQUEUE_REG_14__4__SCAN_IN), .B2(keyinput120), .C1(
        EAX_REG_10__SCAN_IN), .C2(keyinput121), .A(n6557), .ZN(n6558) );
  NAND4_X1 U7498 ( .A1(n6561), .A2(n6560), .A3(n6559), .A4(n6558), .ZN(n6571)
         );
  OAI22_X1 U7499 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(keyinput123), .B1(
        keyinput89), .B2(EAX_REG_17__SCAN_IN), .ZN(n6562) );
  AOI221_X1 U7500 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput123), 
        .C1(EAX_REG_17__SCAN_IN), .C2(keyinput89), .A(n6562), .ZN(n6569) );
  OAI22_X1 U7501 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(keyinput87), .B1(
        keyinput103), .B2(DATAI_27_), .ZN(n6563) );
  AOI221_X1 U7502 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(keyinput87), .C1(
        DATAI_27_), .C2(keyinput103), .A(n6563), .ZN(n6568) );
  OAI22_X1 U7503 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(keyinput76), .B1(
        DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput82), .ZN(n6564) );
  AOI221_X1 U7504 ( .B1(INSTQUEUE_REG_7__6__SCAN_IN), .B2(keyinput76), .C1(
        keyinput82), .C2(DATAWIDTH_REG_0__SCAN_IN), .A(n6564), .ZN(n6567) );
  OAI22_X1 U7505 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(keyinput95), .B1(
        keyinput115), .B2(EAX_REG_9__SCAN_IN), .ZN(n6565) );
  AOI221_X1 U7506 ( .B1(INSTQUEUE_REG_6__0__SCAN_IN), .B2(keyinput95), .C1(
        EAX_REG_9__SCAN_IN), .C2(keyinput115), .A(n6565), .ZN(n6566) );
  NAND4_X1 U7507 ( .A1(n6569), .A2(n6568), .A3(n6567), .A4(n6566), .ZN(n6570)
         );
  NOR4_X1 U7508 ( .A1(n6573), .A2(n6572), .A3(n6571), .A4(n6570), .ZN(n6682)
         );
  AOI22_X1 U7509 ( .A1(DATAO_REG_19__SCAN_IN), .A2(keyinput10), .B1(
        INSTQUEUE_REG_0__3__SCAN_IN), .B2(keyinput62), .ZN(n6574) );
  OAI221_X1 U7510 ( .B1(DATAO_REG_19__SCAN_IN), .B2(keyinput10), .C1(
        INSTQUEUE_REG_0__3__SCAN_IN), .C2(keyinput62), .A(n6574), .ZN(n6581)
         );
  AOI22_X1 U7511 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(keyinput18), .B1(
        REIP_REG_28__SCAN_IN), .B2(keyinput43), .ZN(n6575) );
  OAI221_X1 U7512 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput18), .C1(
        REIP_REG_28__SCAN_IN), .C2(keyinput43), .A(n6575), .ZN(n6580) );
  AOI22_X1 U7513 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(keyinput5), .B1(
        INSTQUEUE_REG_3__5__SCAN_IN), .B2(keyinput2), .ZN(n6576) );
  OAI221_X1 U7514 ( .B1(INSTQUEUE_REG_9__4__SCAN_IN), .B2(keyinput5), .C1(
        INSTQUEUE_REG_3__5__SCAN_IN), .C2(keyinput2), .A(n6576), .ZN(n6579) );
  AOI22_X1 U7515 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(keyinput23), .B1(
        STATE_REG_2__SCAN_IN), .B2(keyinput38), .ZN(n6577) );
  OAI221_X1 U7516 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(keyinput23), .C1(
        STATE_REG_2__SCAN_IN), .C2(keyinput38), .A(n6577), .ZN(n6578) );
  NOR4_X1 U7517 ( .A1(n6581), .A2(n6580), .A3(n6579), .A4(n6578), .ZN(n6615)
         );
  AOI22_X1 U7518 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(keyinput37), .B1(
        INSTQUEUE_REG_7__6__SCAN_IN), .B2(keyinput12), .ZN(n6582) );
  OAI221_X1 U7519 ( .B1(PHYADDRPOINTER_REG_23__SCAN_IN), .B2(keyinput37), .C1(
        INSTQUEUE_REG_7__6__SCAN_IN), .C2(keyinput12), .A(n6582), .ZN(n6589)
         );
  AOI22_X1 U7520 ( .A1(DATAI_7_), .A2(keyinput40), .B1(
        INSTQUEUE_REG_5__1__SCAN_IN), .B2(keyinput60), .ZN(n6583) );
  OAI221_X1 U7521 ( .B1(DATAI_7_), .B2(keyinput40), .C1(
        INSTQUEUE_REG_5__1__SCAN_IN), .C2(keyinput60), .A(n6583), .ZN(n6588)
         );
  AOI22_X1 U7522 ( .A1(LWORD_REG_11__SCAN_IN), .A2(keyinput11), .B1(
        INSTQUEUE_REG_15__0__SCAN_IN), .B2(keyinput58), .ZN(n6584) );
  OAI221_X1 U7523 ( .B1(LWORD_REG_11__SCAN_IN), .B2(keyinput11), .C1(
        INSTQUEUE_REG_15__0__SCAN_IN), .C2(keyinput58), .A(n6584), .ZN(n6587)
         );
  AOI22_X1 U7524 ( .A1(DATAO_REG_21__SCAN_IN), .A2(keyinput21), .B1(
        INSTQUEUE_REG_8__6__SCAN_IN), .B2(keyinput26), .ZN(n6585) );
  OAI221_X1 U7525 ( .B1(DATAO_REG_21__SCAN_IN), .B2(keyinput21), .C1(
        INSTQUEUE_REG_8__6__SCAN_IN), .C2(keyinput26), .A(n6585), .ZN(n6586)
         );
  NOR4_X1 U7526 ( .A1(n6589), .A2(n6588), .A3(n6587), .A4(n6586), .ZN(n6614)
         );
  AOI22_X1 U7527 ( .A1(DATAO_REG_29__SCAN_IN), .A2(keyinput6), .B1(
        INSTQUEUE_REG_13__6__SCAN_IN), .B2(keyinput34), .ZN(n6590) );
  OAI221_X1 U7528 ( .B1(DATAO_REG_29__SCAN_IN), .B2(keyinput6), .C1(
        INSTQUEUE_REG_13__6__SCAN_IN), .C2(keyinput34), .A(n6590), .ZN(n6597)
         );
  AOI22_X1 U7529 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(keyinput61), .B1(
        REIP_REG_19__SCAN_IN), .B2(keyinput44), .ZN(n6591) );
  OAI221_X1 U7530 ( .B1(DATAWIDTH_REG_8__SCAN_IN), .B2(keyinput61), .C1(
        REIP_REG_19__SCAN_IN), .C2(keyinput44), .A(n6591), .ZN(n6596) );
  AOI22_X1 U7531 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(keyinput52), .B1(
        INSTQUEUE_REG_7__5__SCAN_IN), .B2(keyinput19), .ZN(n6592) );
  OAI221_X1 U7532 ( .B1(PHYADDRPOINTER_REG_25__SCAN_IN), .B2(keyinput52), .C1(
        INSTQUEUE_REG_7__5__SCAN_IN), .C2(keyinput19), .A(n6592), .ZN(n6595)
         );
  AOI22_X1 U7533 ( .A1(EAX_REG_10__SCAN_IN), .A2(keyinput57), .B1(
        INSTQUEUE_REG_6__1__SCAN_IN), .B2(keyinput49), .ZN(n6593) );
  OAI221_X1 U7534 ( .B1(EAX_REG_10__SCAN_IN), .B2(keyinput57), .C1(
        INSTQUEUE_REG_6__1__SCAN_IN), .C2(keyinput49), .A(n6593), .ZN(n6594)
         );
  NOR4_X1 U7535 ( .A1(n6597), .A2(n6596), .A3(n6595), .A4(n6594), .ZN(n6613)
         );
  INV_X1 U7536 ( .A(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n6599) );
  AOI22_X1 U7537 ( .A1(REIP_REG_4__SCAN_IN), .A2(keyinput41), .B1(n6599), .B2(
        keyinput42), .ZN(n6598) );
  OAI221_X1 U7538 ( .B1(REIP_REG_4__SCAN_IN), .B2(keyinput41), .C1(n6599), 
        .C2(keyinput42), .A(n6598), .ZN(n6611) );
  AOI22_X1 U7539 ( .A1(n4729), .A2(keyinput8), .B1(keyinput4), .B2(n6601), 
        .ZN(n6600) );
  OAI221_X1 U7540 ( .B1(n4729), .B2(keyinput8), .C1(n6601), .C2(keyinput4), 
        .A(n6600), .ZN(n6610) );
  AOI22_X1 U7541 ( .A1(n6604), .A2(keyinput16), .B1(keyinput20), .B2(n6603), 
        .ZN(n6602) );
  OAI221_X1 U7542 ( .B1(n6604), .B2(keyinput16), .C1(n6603), .C2(keyinput20), 
        .A(n6602), .ZN(n6609) );
  AOI22_X1 U7543 ( .A1(n6607), .A2(keyinput50), .B1(keyinput47), .B2(n6606), 
        .ZN(n6605) );
  OAI221_X1 U7544 ( .B1(n6607), .B2(keyinput50), .C1(n6606), .C2(keyinput47), 
        .A(n6605), .ZN(n6608) );
  NOR4_X1 U7545 ( .A1(n6611), .A2(n6610), .A3(n6609), .A4(n6608), .ZN(n6612)
         );
  NAND4_X1 U7546 ( .A1(n6615), .A2(n6614), .A3(n6613), .A4(n6612), .ZN(n6681)
         );
  AOI22_X1 U7547 ( .A1(n6618), .A2(keyinput35), .B1(n6617), .B2(keyinput36), 
        .ZN(n6616) );
  OAI221_X1 U7548 ( .B1(n6618), .B2(keyinput35), .C1(n6617), .C2(keyinput36), 
        .A(n6616), .ZN(n6630) );
  AOI22_X1 U7549 ( .A1(n4819), .A2(keyinput31), .B1(keyinput33), .B2(n6620), 
        .ZN(n6619) );
  OAI221_X1 U7550 ( .B1(n4819), .B2(keyinput31), .C1(n6620), .C2(keyinput33), 
        .A(n6619), .ZN(n6629) );
  AOI22_X1 U7551 ( .A1(n6623), .A2(keyinput14), .B1(keyinput28), .B2(n6622), 
        .ZN(n6621) );
  OAI221_X1 U7552 ( .B1(n6623), .B2(keyinput14), .C1(n6622), .C2(keyinput28), 
        .A(n6621), .ZN(n6628) );
  AOI22_X1 U7553 ( .A1(n6626), .A2(keyinput45), .B1(keyinput3), .B2(n6625), 
        .ZN(n6624) );
  OAI221_X1 U7554 ( .B1(n6626), .B2(keyinput45), .C1(n6625), .C2(keyinput3), 
        .A(n6624), .ZN(n6627) );
  NOR4_X1 U7555 ( .A1(n6630), .A2(n6629), .A3(n6628), .A4(n6627), .ZN(n6679)
         );
  AOI22_X1 U7556 ( .A1(n6633), .A2(keyinput53), .B1(keyinput29), .B2(n6632), 
        .ZN(n6631) );
  OAI221_X1 U7557 ( .B1(n6633), .B2(keyinput53), .C1(n6632), .C2(keyinput29), 
        .A(n6631), .ZN(n6645) );
  AOI22_X1 U7558 ( .A1(n6636), .A2(keyinput55), .B1(keyinput46), .B2(n6635), 
        .ZN(n6634) );
  OAI221_X1 U7559 ( .B1(n6636), .B2(keyinput55), .C1(n6635), .C2(keyinput46), 
        .A(n6634), .ZN(n6644) );
  AOI22_X1 U7560 ( .A1(n6638), .A2(keyinput9), .B1(n3522), .B2(keyinput1), 
        .ZN(n6637) );
  OAI221_X1 U7561 ( .B1(n6638), .B2(keyinput9), .C1(n3522), .C2(keyinput1), 
        .A(n6637), .ZN(n6643) );
  AOI22_X1 U7562 ( .A1(n6641), .A2(keyinput54), .B1(keyinput32), .B2(n6640), 
        .ZN(n6639) );
  OAI221_X1 U7563 ( .B1(n6641), .B2(keyinput54), .C1(n6640), .C2(keyinput32), 
        .A(n6639), .ZN(n6642) );
  NOR4_X1 U7564 ( .A1(n6645), .A2(n6644), .A3(n6643), .A4(n6642), .ZN(n6678)
         );
  AOI22_X1 U7565 ( .A1(n6648), .A2(keyinput25), .B1(n6647), .B2(keyinput48), 
        .ZN(n6646) );
  OAI221_X1 U7566 ( .B1(n6648), .B2(keyinput25), .C1(n6647), .C2(keyinput48), 
        .A(n6646), .ZN(n6660) );
  AOI22_X1 U7567 ( .A1(n6650), .A2(keyinput59), .B1(n4668), .B2(keyinput24), 
        .ZN(n6649) );
  OAI221_X1 U7568 ( .B1(n6650), .B2(keyinput59), .C1(n4668), .C2(keyinput24), 
        .A(n6649), .ZN(n6659) );
  AOI22_X1 U7569 ( .A1(n6653), .A2(keyinput30), .B1(keyinput63), .B2(n6652), 
        .ZN(n6651) );
  OAI221_X1 U7570 ( .B1(n6653), .B2(keyinput30), .C1(n6652), .C2(keyinput63), 
        .A(n6651), .ZN(n6658) );
  INV_X1 U7571 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n6655) );
  AOI22_X1 U7572 ( .A1(n6656), .A2(keyinput15), .B1(n6655), .B2(keyinput56), 
        .ZN(n6654) );
  OAI221_X1 U7573 ( .B1(n6656), .B2(keyinput15), .C1(n6655), .C2(keyinput56), 
        .A(n6654), .ZN(n6657) );
  NOR4_X1 U7574 ( .A1(n6660), .A2(n6659), .A3(n6658), .A4(n6657), .ZN(n6677)
         );
  INV_X1 U7575 ( .A(DATAI_27_), .ZN(n6663) );
  AOI22_X1 U7576 ( .A1(n6663), .A2(keyinput39), .B1(n6662), .B2(keyinput7), 
        .ZN(n6661) );
  OAI221_X1 U7577 ( .B1(n6663), .B2(keyinput39), .C1(n6662), .C2(keyinput7), 
        .A(n6661), .ZN(n6675) );
  AOI22_X1 U7578 ( .A1(n6666), .A2(keyinput13), .B1(keyinput22), .B2(n6665), 
        .ZN(n6664) );
  OAI221_X1 U7579 ( .B1(n6666), .B2(keyinput13), .C1(n6665), .C2(keyinput22), 
        .A(n6664), .ZN(n6674) );
  AOI22_X1 U7580 ( .A1(n4156), .A2(keyinput17), .B1(keyinput27), .B2(n6668), 
        .ZN(n6667) );
  OAI221_X1 U7581 ( .B1(n4156), .B2(keyinput17), .C1(n6668), .C2(keyinput27), 
        .A(n6667), .ZN(n6673) );
  AOI22_X1 U7582 ( .A1(n6671), .A2(keyinput0), .B1(keyinput51), .B2(n6670), 
        .ZN(n6669) );
  OAI221_X1 U7583 ( .B1(n6671), .B2(keyinput0), .C1(n6670), .C2(keyinput51), 
        .A(n6669), .ZN(n6672) );
  NOR4_X1 U7584 ( .A1(n6675), .A2(n6674), .A3(n6673), .A4(n6672), .ZN(n6676)
         );
  NAND4_X1 U7585 ( .A1(n6679), .A2(n6678), .A3(n6677), .A4(n6676), .ZN(n6680)
         );
  AOI211_X1 U7586 ( .C1(n6683), .C2(n6682), .A(n6681), .B(n6680), .ZN(n6695)
         );
  OAI22_X1 U7587 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n6686), .B1(n6685), .B2(n6684), .ZN(n6692) );
  INV_X1 U7588 ( .A(n6687), .ZN(n6690) );
  OAI22_X1 U7589 ( .A1(n6690), .A2(n5394), .B1(n6689), .B2(n6688), .ZN(n6691)
         );
  AOI211_X1 U7590 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n6693), .A(n6692), .B(n6691), .ZN(n6694) );
  XNOR2_X1 U7591 ( .A(n6695), .B(n6694), .ZN(U2999) );
  CLKBUF_X1 U34680 ( .A(n4120), .Z(n4291) );
  CLKBUF_X1 U3484 ( .A(n4123), .Z(n4178) );
  CLKBUF_X1 U3487 ( .A(n4102), .Z(n4550) );
  NAND2_X1 U3741 ( .A1(n4890), .A2(n4889), .ZN(n4888) );
  CLKBUF_X1 U3974 ( .A(n5939), .Z(n2998) );
endmodule

