

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9560, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9571,
         n9572, n9573, n9574, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932;

  INV_X2 U11004 ( .A(n19155), .ZN(n16264) );
  INV_X1 U11005 ( .A(n15965), .ZN(n16013) );
  NOR2_X2 U11006 ( .A1(n13016), .A2(n18858), .ZN(n18855) );
  AND2_X1 U11007 ( .A1(n11703), .A2(n11719), .ZN(n9676) );
  CLKBUF_X1 U11008 ( .A(n10412), .Z(n13740) );
  XNOR2_X1 U11009 ( .A(n11383), .B(n11382), .ZN(n11541) );
  AND2_X1 U11010 ( .A1(n10298), .A2(n10290), .ZN(n10412) );
  NOR2_X1 U11011 ( .A1(n10286), .A2(n9829), .ZN(n10403) );
  OAI22_X1 U11012 ( .A1(n13571), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11545), 
        .B2(n11522), .ZN(n11383) );
  CLKBUF_X2 U11013 ( .A(n10277), .Z(n10274) );
  AND2_X1 U11014 ( .A1(n19023), .A2(n10264), .ZN(n10299) );
  CLKBUF_X3 U11015 ( .A(n12691), .Z(n9568) );
  AND2_X1 U11017 ( .A1(n12420), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12383) );
  AND2_X1 U11018 ( .A1(n13936), .A2(n12401), .ZN(n11072) );
  CLKBUF_X2 U11019 ( .A(n11251), .Z(n12155) );
  CLKBUF_X1 U11020 ( .A(n12675), .Z(n17100) );
  CLKBUF_X2 U11021 ( .A(n11419), .Z(n12013) );
  NAND4_X1 U11022 ( .A1(n18783), .A2(n18777), .A3(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A4(n18769), .ZN(n17090) );
  INV_X1 U11023 ( .A(n14276), .ZN(n14290) );
  INV_X1 U11024 ( .A(n9618), .ZN(n17142) );
  INV_X1 U11025 ( .A(n9564), .ZN(n17141) );
  NAND2_X1 U11026 ( .A1(n9573), .A2(n10874), .ZN(n10879) );
  AND4_X1 U11027 ( .A1(n11246), .A2(n11245), .A3(n11244), .A4(n11243), .ZN(
        n11247) );
  AND2_X1 U11028 ( .A1(n10889), .A2(n10874), .ZN(n9593) );
  AND4_X1 U11029 ( .A1(n11189), .A2(n11188), .A3(n11187), .A4(n11186), .ZN(
        n11210) );
  AND2_X1 U11030 ( .A1(n11196), .A2(n13345), .ZN(n11467) );
  CLKBUF_X2 U11031 ( .A(n10191), .Z(n9584) );
  CLKBUF_X1 U11032 ( .A(n18579), .Z(n9560) );
  NOR2_X1 U11033 ( .A1(n18386), .A2(n18477), .ZN(n18579) );
  INV_X1 U11035 ( .A(n20930), .ZN(n9562) );
  CLKBUF_X3 U11036 ( .A(n11266), .Z(n12014) );
  NAND2_X1 U11037 ( .A1(n11386), .A2(n11333), .ZN(n11454) );
  INV_X1 U11038 ( .A(n9567), .ZN(n12364) );
  AOI21_X1 U11040 ( .B1(n11454), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11361), .ZN(n11366) );
  NAND2_X1 U11041 ( .A1(n11447), .A2(n20676), .ZN(n11450) );
  CLKBUF_X3 U11042 ( .A(n10239), .Z(n10862) );
  AND2_X1 U11043 ( .A1(n12575), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10331) );
  AND2_X1 U11044 ( .A1(n12575), .A2(n10115), .ZN(n10376) );
  INV_X1 U11045 ( .A(n13035), .ZN(n10701) );
  NAND2_X1 U11046 ( .A1(n10298), .A2(n10059), .ZN(n19500) );
  NOR2_X1 U11047 ( .A1(n9874), .A2(n14276), .ZN(n14168) );
  NAND4_X2 U11048 ( .A1(n11314), .A2(n11313), .A3(n11312), .A4(n11311), .ZN(
        n11328) );
  INV_X1 U11049 ( .A(n11764), .ZN(n12201) );
  CLKBUF_X3 U11050 ( .A(n10239), .Z(n14242) );
  CLKBUF_X2 U11051 ( .A(n9569), .Z(n10771) );
  AND2_X1 U11052 ( .A1(n9830), .A2(n14011), .ZN(n19323) );
  INV_X1 U11053 ( .A(n9805), .ZN(n15798) );
  AND2_X2 U11055 ( .A1(n14399), .A2(n9975), .ZN(n14316) );
  BUF_X1 U11057 ( .A(n9916), .Z(n14236) );
  AND2_X1 U11058 ( .A1(n9712), .A2(n9648), .ZN(n15330) );
  AND2_X1 U11059 ( .A1(n9572), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10389) );
  NOR2_X1 U11060 ( .A1(n17785), .A2(n17784), .ZN(n17783) );
  INV_X1 U11061 ( .A(n17199), .ZN(n18187) );
  NOR3_X1 U11062 ( .A1(n14392), .A2(n9673), .A3(n9875), .ZN(n14306) );
  NAND2_X1 U11063 ( .A1(n13512), .A2(n11719), .ZN(n13527) );
  NAND2_X1 U11064 ( .A1(n13892), .A2(n13918), .ZN(n13917) );
  INV_X2 U11065 ( .A(n12700), .ZN(n17137) );
  INV_X1 U11066 ( .A(n17666), .ZN(n17682) );
  NOR2_X1 U11067 ( .A1(n18804), .A2(n9617), .ZN(n17816) );
  INV_X1 U11068 ( .A(n13675), .ZN(n13674) );
  INV_X1 U11069 ( .A(n17819), .ZN(n17811) );
  XNOR2_X1 U11070 ( .A(n11541), .B(n11540), .ZN(n11696) );
  XOR2_X1 U11071 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11637), .Z(
        n9563) );
  OR2_X1 U11072 ( .A1(n12648), .A2(n12647), .ZN(n9564) );
  INV_X2 U11073 ( .A(n17113), .ZN(n17149) );
  NAND2_X1 U11074 ( .A1(n12640), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15478) );
  NAND2_X2 U11075 ( .A1(n15599), .A2(n12629), .ZN(n12265) );
  AND2_X4 U11076 ( .A1(n11202), .A2(n11190), .ZN(n11462) );
  OR2_X1 U11077 ( .A1(n10274), .A2(n9692), .ZN(n9694) );
  NOR2_X2 U11078 ( .A1(n9691), .A2(n10274), .ZN(n19294) );
  NAND2_X2 U11079 ( .A1(n10178), .A2(n10115), .ZN(n10179) );
  OR2_X1 U11081 ( .A1(n18769), .A2(n18617), .ZN(n12685) );
  NOR3_X4 U11082 ( .A1(n9877), .A2(n9876), .A3(n9670), .ZN(n14304) );
  NAND2_X2 U11083 ( .A1(n13101), .A2(n11325), .ZN(n11348) );
  AND2_X2 U11084 ( .A1(n13332), .A2(n12217), .ZN(n13101) );
  NAND2_X1 U11085 ( .A1(n14002), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9566) );
  NOR3_X1 U11086 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n10317), .ZN(n10318) );
  NOR2_X2 U11087 ( .A1(n13642), .A2(n13641), .ZN(n13656) );
  NAND2_X2 U11088 ( .A1(n9776), .A2(n9774), .ZN(n15197) );
  INV_X2 U11090 ( .A(n15727), .ZN(n18181) );
  NAND2_X2 U11091 ( .A1(n14973), .A2(n12473), .ZN(n12493) );
  NAND3_X2 U11092 ( .A1(n10481), .A2(n11148), .A3(n13887), .ZN(n13888) );
  NAND2_X2 U11095 ( .A1(n10154), .A2(n10153), .ZN(n10718) );
  INV_X2 U11096 ( .A(n13870), .ZN(n11447) );
  OAI222_X1 U11097 ( .A1(n14455), .A2(n14575), .B1(n14191), .B2(n19994), .C1(
        n14184), .C2(n14457), .ZN(P1_U2844) );
  NAND2_X4 U11098 ( .A1(n12650), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n17113) );
  AND2_X2 U11099 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n12643), .ZN(
        n12650) );
  NAND2_X2 U11100 ( .A1(n10128), .A2(n10127), .ZN(n10183) );
  AOI21_X2 U11101 ( .B1(n15162), .B2(n15158), .A(n15160), .ZN(n12623) );
  INV_X4 U11103 ( .A(n13017), .ZN(n13016) );
  XOR2_X2 U11104 ( .A(n18771), .B(n17347), .Z(n17818) );
  AND3_X2 U11105 ( .A1(n12684), .A2(n9938), .A3(n9935), .ZN(n17347) );
  BUF_X2 U11106 ( .A(n10309), .Z(n9571) );
  BUF_X8 U11107 ( .A(n10309), .Z(n9572) );
  AND2_X2 U11108 ( .A1(n10316), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10309) );
  AOI211_X1 U11109 ( .C1(n16248), .C2(n15266), .A(n15118), .B(n15117), .ZN(
        n15119) );
  NAND2_X1 U11110 ( .A1(n9770), .A2(n15442), .ZN(n15217) );
  NAND2_X1 U11111 ( .A1(n9772), .A2(n9771), .ZN(n15445) );
  OR2_X1 U11112 ( .A1(n15490), .A2(n9595), .ZN(n9841) );
  NAND2_X1 U11113 ( .A1(n15227), .A2(n10567), .ZN(n15490) );
  NAND2_X1 U11114 ( .A1(n15237), .A2(n15235), .ZN(n15227) );
  XNOR2_X1 U11115 ( .A(n14247), .B(n14246), .ZN(n14262) );
  NAND2_X1 U11116 ( .A1(n9728), .A2(n16024), .ZN(n11613) );
  AND2_X1 U11117 ( .A1(n12771), .A2(n12770), .ZN(n17493) );
  NAND2_X1 U11118 ( .A1(n11555), .A2(n11563), .ZN(n11720) );
  OR2_X1 U11119 ( .A1(n12915), .A2(n12759), .ZN(n17611) );
  NOR3_X1 U11121 ( .A1(n14800), .A2(n14079), .A3(n9663), .ZN(n9884) );
  NAND2_X1 U11122 ( .A1(n19994), .A2(n20134), .ZN(n14455) );
  CLKBUF_X2 U11123 ( .A(n18048), .Z(n9586) );
  NOR2_X1 U11125 ( .A1(n10489), .A2(n10483), .ZN(n10482) );
  CLKBUF_X2 U11126 ( .A(n10239), .Z(n10858) );
  AND3_X2 U11127 ( .A1(n9828), .A2(n9593), .A3(n10194), .ZN(n10744) );
  AOI211_X1 U11128 ( .C1(n9574), .C2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n12732), .B(n12731), .ZN(n17316) );
  INV_X1 U11129 ( .A(n10889), .ZN(n9573) );
  CLKBUF_X2 U11130 ( .A(n10212), .Z(n13035) );
  BUF_X2 U11131 ( .A(n13661), .Z(n9581) );
  INV_X2 U11132 ( .A(n19196), .ZN(n12416) );
  BUF_X2 U11133 ( .A(n11328), .Z(n20102) );
  INV_X2 U11134 ( .A(n10718), .ZN(n10874) );
  CLKBUF_X2 U11135 ( .A(n11420), .Z(n12173) );
  CLKBUF_X2 U11136 ( .A(n11819), .Z(n11835) );
  CLKBUF_X2 U11137 ( .A(n11273), .Z(n12183) );
  CLKBUF_X2 U11138 ( .A(n11422), .Z(n11423) );
  CLKBUF_X2 U11139 ( .A(n11461), .Z(n12182) );
  BUF_X2 U11140 ( .A(n11467), .Z(n9576) );
  CLKBUF_X2 U11141 ( .A(n10311), .Z(n12571) );
  BUF_X1 U11142 ( .A(n12829), .Z(n9579) );
  CLKBUF_X2 U11143 ( .A(n10307), .Z(n12570) );
  INV_X4 U11144 ( .A(n10053), .ZN(n16899) );
  INV_X1 U11145 ( .A(n12829), .ZN(n12721) );
  INV_X1 U11146 ( .A(n12367), .ZN(n12375) );
  CLKBUF_X2 U11147 ( .A(n11372), .Z(n12015) );
  INV_X4 U11148 ( .A(n17090), .ZN(n12701) );
  INV_X4 U11149 ( .A(n17108), .ZN(n17131) );
  NOR3_X1 U11150 ( .A1(n18769), .A2(n18777), .A3(n16867), .ZN(n12829) );
  AND2_X1 U11151 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13346) );
  INV_X4 U11152 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n20806) );
  INV_X1 U11153 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20676) );
  OR2_X1 U11154 ( .A1(n9926), .A2(n9769), .ZN(n9768) );
  NOR2_X1 U11155 ( .A1(n15274), .A2(n10045), .ZN(n10044) );
  AOI21_X1 U11156 ( .B1(n15107), .B2(n9624), .A(n9709), .ZN(n9708) );
  OAI21_X1 U11157 ( .B1(n15418), .B2(n9607), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9889) );
  NAND2_X1 U11158 ( .A1(n9898), .A2(n9613), .ZN(n16198) );
  XNOR2_X1 U11159 ( .A(n12204), .B(n12203), .ZN(n14281) );
  OR2_X1 U11160 ( .A1(n15478), .A2(n15449), .ZN(n15448) );
  XNOR2_X1 U11161 ( .A(n9987), .B(n14287), .ZN(n14554) );
  NAND2_X1 U11162 ( .A1(n9841), .A2(n9839), .ZN(n12612) );
  AND2_X1 U11163 ( .A1(n14400), .A2(n14409), .ZN(n15848) );
  NAND2_X1 U11164 ( .A1(n11172), .A2(n11171), .ZN(n15501) );
  NAND2_X1 U11165 ( .A1(n11165), .A2(n11164), .ZN(n15225) );
  NAND2_X1 U11166 ( .A1(n12472), .A2(n12471), .ZN(n12473) );
  NAND2_X1 U11167 ( .A1(n10866), .A2(n10865), .ZN(n14247) );
  NOR2_X1 U11168 ( .A1(n10034), .A2(n11161), .ZN(n10033) );
  AND2_X1 U11169 ( .A1(n14869), .A2(n14858), .ZN(n10866) );
  NAND2_X1 U11170 ( .A1(n11158), .A2(n20886), .ZN(n9894) );
  NOR2_X1 U11171 ( .A1(n14899), .A2(n14212), .ZN(n14965) );
  NAND2_X1 U11172 ( .A1(n14922), .A2(n10048), .ZN(n14899) );
  INV_X1 U11173 ( .A(n15106), .ZN(n9706) );
  OR2_X1 U11174 ( .A1(n9958), .A2(n9955), .ZN(n9954) );
  NOR2_X2 U11175 ( .A1(n15013), .A2(n14921), .ZN(n14922) );
  AND2_X1 U11176 ( .A1(n10683), .A2(n10684), .ZN(n9707) );
  AND2_X1 U11177 ( .A1(n11612), .A2(n9634), .ZN(n9958) );
  AND2_X1 U11178 ( .A1(n10439), .A2(n10438), .ZN(n10508) );
  AND2_X1 U11179 ( .A1(n10553), .A2(n10552), .ZN(n11167) );
  AND2_X1 U11180 ( .A1(n15150), .A2(n9868), .ZN(n9867) );
  XNOR2_X1 U11181 ( .A(n11600), .B(n11599), .ZN(n11766) );
  NAND2_X1 U11182 ( .A1(n13527), .A2(n13526), .ZN(n13525) );
  AND2_X1 U11183 ( .A1(n10517), .A2(n10516), .ZN(n10535) );
  OR2_X1 U11184 ( .A1(n19328), .A2(n10544), .ZN(n10517) );
  OR2_X1 U11185 ( .A1(n10649), .A2(n10593), .ZN(n18860) );
  OAI21_X1 U11186 ( .B1(n10399), .B2(n10365), .A(n9695), .ZN(n10366) );
  OR2_X1 U11187 ( .A1(n10654), .A2(n10655), .ZN(n10661) );
  AND2_X1 U11188 ( .A1(n10300), .A2(n10299), .ZN(n10511) );
  AND2_X1 U11189 ( .A1(n10300), .A2(n10290), .ZN(n10359) );
  AND2_X1 U11190 ( .A1(n10300), .A2(n10059), .ZN(n19614) );
  INV_X1 U11191 ( .A(n10278), .ZN(n10298) );
  OR2_X1 U11192 ( .A1(n10281), .A2(n10280), .ZN(n19555) );
  OAI21_X2 U11193 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18811), .A(n9617), 
        .ZN(n17827) );
  NAND2_X1 U11194 ( .A1(n11476), .A2(n14825), .ZN(n11563) );
  NAND2_X1 U11195 ( .A1(n10651), .A2(n10670), .ZN(n10649) );
  OR2_X1 U11196 ( .A1(n12253), .A2(n12252), .ZN(n13322) );
  AND2_X1 U11197 ( .A1(n13237), .A2(n12260), .ZN(n13325) );
  OR2_X1 U11198 ( .A1(n18606), .A2(n18657), .ZN(n9617) );
  CLKBUF_X1 U11199 ( .A(n12246), .Z(n14011) );
  NOR2_X1 U11200 ( .A1(n10269), .A2(n12246), .ZN(n9698) );
  NAND2_X1 U11201 ( .A1(n10267), .A2(n10266), .ZN(n15568) );
  NOR2_X1 U11202 ( .A1(n13804), .A2(n13803), .ZN(n19923) );
  NAND2_X1 U11203 ( .A1(n11475), .A2(n11474), .ZN(n14825) );
  NAND2_X1 U11204 ( .A1(n12255), .A2(n12254), .ZN(n15584) );
  AND2_X1 U11205 ( .A1(n10270), .A2(n19023), .ZN(n10290) );
  AND2_X1 U11206 ( .A1(n10767), .A2(n10256), .ZN(n10769) );
  NAND2_X1 U11207 ( .A1(n9918), .A2(n9917), .ZN(n10246) );
  XNOR2_X1 U11208 ( .A(n11453), .B(n20250), .ZN(n13328) );
  INV_X2 U11209 ( .A(n13414), .ZN(n20052) );
  AOI21_X1 U11210 ( .B1(n13082), .B2(n13081), .A(n19873), .ZN(n13107) );
  OR2_X1 U11211 ( .A1(n10255), .A2(n10254), .ZN(n10767) );
  XNOR2_X1 U11212 ( .A(n11528), .B(n11527), .ZN(n20171) );
  NAND2_X1 U11213 ( .A1(n11363), .A2(n11362), .ZN(n11453) );
  NOR2_X1 U11214 ( .A1(n10258), .A2(n10257), .ZN(n10259) );
  NAND2_X1 U11215 ( .A1(n11451), .A2(n11441), .ZN(n11704) );
  NAND2_X1 U11216 ( .A1(n11526), .A2(n11418), .ZN(n11451) );
  INV_X2 U11217 ( .A(n17357), .ZN(n17392) );
  NAND2_X1 U11218 ( .A1(n11459), .A2(n11458), .ZN(n20250) );
  AND2_X1 U11219 ( .A1(n13051), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13049) );
  OR2_X1 U11220 ( .A1(n13536), .A2(n13535), .ZN(n13627) );
  AND2_X1 U11221 ( .A1(n13934), .A2(n10892), .ZN(n14003) );
  NAND2_X1 U11222 ( .A1(n12994), .A2(n9606), .ZN(n13052) );
  OAI211_X1 U11223 ( .C1(n10233), .C2(n10231), .A(n10209), .B(n10208), .ZN(
        n10222) );
  AOI21_X1 U11224 ( .B1(n10862), .B2(P2_REIP_REG_1__SCAN_IN), .A(n9833), .ZN(
        n9832) );
  NAND2_X1 U11225 ( .A1(n10204), .A2(n10057), .ZN(n10233) );
  AND2_X1 U11226 ( .A1(n11522), .A2(n11417), .ZN(n11418) );
  AND2_X1 U11227 ( .A1(n10203), .A2(n10202), .ZN(n10057) );
  AND2_X1 U11228 ( .A1(n10192), .A2(n16348), .ZN(n11115) );
  AND2_X1 U11229 ( .A1(n9950), .A2(n11344), .ZN(n9949) );
  INV_X1 U11230 ( .A(n18151), .ZN(n16820) );
  NAND2_X1 U11231 ( .A1(n10892), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10231) );
  AND2_X1 U11232 ( .A1(n10881), .A2(n10213), .ZN(n14002) );
  AND2_X1 U11233 ( .A1(n12587), .A2(n10198), .ZN(n10204) );
  NAND2_X1 U11234 ( .A1(n11319), .A2(n10073), .ZN(n11334) );
  OAI211_X1 U11235 ( .C1(n11523), .C2(n13242), .A(n11437), .B(n11436), .ZN(
        n11527) );
  AOI211_X1 U11236 ( .C1(n17137), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n12720), .B(n12719), .ZN(n17323) );
  INV_X1 U11237 ( .A(n10487), .ZN(n10491) );
  AND2_X1 U11238 ( .A1(n11315), .A2(n11336), .ZN(n11319) );
  NAND2_X1 U11239 ( .A1(n9593), .A2(n10190), .ZN(n16321) );
  INV_X1 U11240 ( .A(n18163), .ZN(n15724) );
  AND3_X1 U11241 ( .A1(n11340), .A2(n13213), .A3(n9725), .ZN(n13104) );
  AND2_X1 U11242 ( .A1(n12854), .A2(n9743), .ZN(n18163) );
  AND3_X1 U11243 ( .A1(n9633), .A2(n12696), .A3(n9940), .ZN(n17336) );
  OAI211_X2 U11244 ( .C1(n12700), .C2(n18244), .A(n12876), .B(n12875), .ZN(
        n17240) );
  AND3_X1 U11245 ( .A1(n10372), .A2(n10375), .A3(n9902), .ZN(n10926) );
  NAND2_X1 U11246 ( .A1(n9916), .A2(n9915), .ZN(n10199) );
  AND2_X2 U11247 ( .A1(n9916), .A2(n9584), .ZN(n10194) );
  AND2_X1 U11248 ( .A1(n13413), .A2(n20084), .ZN(n13213) );
  INV_X1 U11249 ( .A(n20084), .ZN(n13242) );
  INV_X2 U11250 ( .A(U212), .ZN(n16458) );
  BUF_X1 U11251 ( .A(n10191), .Z(n9582) );
  INV_X1 U11252 ( .A(n11324), .ZN(n13359) );
  OR2_X1 U11253 ( .A1(n10353), .A2(n10352), .ZN(n10468) );
  NOR2_X2 U11254 ( .A1(n20084), .A2(n11328), .ZN(n13410) );
  OR2_X1 U11255 ( .A1(n11261), .A2(n11260), .ZN(n11324) );
  OR2_X1 U11256 ( .A1(n11434), .A2(n11433), .ZN(n11542) );
  AND4_X1 U11257 ( .A1(n11282), .A2(n11281), .A3(n11280), .A4(n11279), .ZN(
        n11293) );
  AND4_X1 U11258 ( .A1(n11286), .A2(n11285), .A3(n11284), .A4(n11283), .ZN(
        n11292) );
  AND3_X1 U11259 ( .A1(n9714), .A2(n11217), .A3(n11211), .ZN(n9589) );
  AND4_X1 U11260 ( .A1(n11265), .A2(n11264), .A3(n11263), .A4(n11262), .ZN(
        n10072) );
  AND4_X1 U11261 ( .A1(n10139), .A2(n10138), .A3(n10137), .A4(n10136), .ZN(
        n10140) );
  AND4_X1 U11262 ( .A1(n11238), .A2(n11237), .A3(n11236), .A4(n11235), .ZN(
        n11249) );
  AND4_X1 U11263 ( .A1(n11278), .A2(n11277), .A3(n11276), .A4(n11275), .ZN(
        n11294) );
  AND4_X1 U11264 ( .A1(n11206), .A2(n11205), .A3(n11204), .A4(n11203), .ZN(
        n11207) );
  AND4_X1 U11265 ( .A1(n11194), .A2(n11193), .A3(n11192), .A4(n11191), .ZN(
        n11209) );
  NAND2_X2 U11266 ( .A1(n18800), .A2(n18685), .ZN(n18743) );
  BUF_X2 U11267 ( .A(n12675), .Z(n17143) );
  INV_X2 U11268 ( .A(n12721), .ZN(n17148) );
  BUF_X4 U11269 ( .A(n12690), .Z(n9574) );
  AND4_X1 U11270 ( .A1(n11242), .A2(n11241), .A3(n11240), .A4(n11239), .ZN(
        n11248) );
  AND4_X1 U11271 ( .A1(n11302), .A2(n11301), .A3(n11300), .A4(n11299), .ZN(
        n11313) );
  AND4_X1 U11272 ( .A1(n11306), .A2(n11305), .A3(n11304), .A4(n11303), .ZN(
        n11312) );
  CLKBUF_X2 U11273 ( .A(n11478), .Z(n12184) );
  NOR2_X2 U11274 ( .A1(n18634), .A2(n18433), .ZN(n18526) );
  BUF_X2 U11275 ( .A(n10306), .Z(n12569) );
  AND2_X2 U11276 ( .A1(n9572), .A2(n10115), .ZN(n12393) );
  NAND2_X2 U11277 ( .A1(n19868), .A2(n19739), .ZN(n19792) );
  AND2_X1 U11278 ( .A1(n10131), .A2(n10115), .ZN(n10132) );
  INV_X1 U11279 ( .A(n17088), .ZN(n17140) );
  NAND2_X1 U11280 ( .A1(n18769), .A2(n12650), .ZN(n17004) );
  INV_X2 U11281 ( .A(n16490), .ZN(U215) );
  NAND2_X1 U11282 ( .A1(n9822), .A2(n9821), .ZN(n12700) );
  AND2_X2 U11283 ( .A1(n11197), .A2(n13340), .ZN(n11421) );
  CLKBUF_X1 U11284 ( .A(n12156), .Z(n12176) );
  INV_X2 U11285 ( .A(n18817), .ZN(n18800) );
  INV_X2 U11286 ( .A(n18137), .ZN(n9577) );
  INV_X2 U11287 ( .A(n16492), .ZN(n16494) );
  OR2_X1 U11288 ( .A1(n16868), .A2(n12649), .ZN(n9616) );
  AND2_X2 U11289 ( .A1(n13936), .A2(n10458), .ZN(n10306) );
  AND2_X1 U11290 ( .A1(n11184), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11195) );
  OR3_X2 U11291 ( .A1(n16867), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10053) );
  NAND4_X1 U11292 ( .A1(n18777), .A2(n18783), .A3(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17108) );
  AND3_X2 U11293 ( .A1(n10078), .A2(n10077), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12575) );
  NAND2_X1 U11294 ( .A1(n20806), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12648) );
  AND2_X2 U11295 ( .A1(n9761), .A2(n10458), .ZN(n10307) );
  AND2_X1 U11296 ( .A1(n10083), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13936) );
  NAND2_X1 U11297 ( .A1(n18777), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12649) );
  NAND2_X1 U11298 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16868) );
  INV_X1 U11299 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15577) );
  NOR2_X1 U11300 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14004) );
  OR2_X1 U11301 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16867) );
  NOR2_X2 U11302 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14830) );
  AND2_X1 U11304 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13340) );
  OR2_X1 U11305 ( .A1(n12613), .A2(n9777), .ZN(n9776) );
  NAND2_X1 U11306 ( .A1(n14141), .A2(n14142), .ZN(n14301) );
  OR2_X4 U11307 ( .A1(n14219), .A2(n11179), .ZN(n15134) );
  AND2_X4 U11308 ( .A1(n14830), .A2(n13346), .ZN(n11230) );
  OAI211_X1 U11309 ( .C1(n10233), .C2(n10231), .A(n10209), .B(n10208), .ZN(
        n9578) );
  NOR3_X2 U11310 ( .A1(n17275), .A2(n17241), .A3(n17198), .ZN(n17236) );
  OAI21_X2 U11311 ( .B1(n10110), .B2(n10109), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9765) );
  OR2_X1 U11312 ( .A1(n11563), .A2(n11562), .ZN(n11577) );
  NAND2_X2 U11313 ( .A1(n10193), .A2(n10228), .ZN(n10237) );
  INV_X1 U11314 ( .A(n10770), .ZN(n9580) );
  NAND2_X1 U11315 ( .A1(n14002), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10241) );
  AND2_X2 U11316 ( .A1(n10749), .A2(n9584), .ZN(n10185) );
  OR2_X1 U11317 ( .A1(n12261), .A2(n10291), .ZN(n19357) );
  OR3_X1 U11318 ( .A1(n12261), .A2(n12246), .A3(n10271), .ZN(n10399) );
  NOR2_X4 U11319 ( .A1(n15116), .A2(n15099), .ZN(n15098) );
  OR2_X1 U11320 ( .A1(n20112), .A2(n20084), .ZN(n13661) );
  BUF_X2 U11321 ( .A(n12261), .Z(n15599) );
  BUF_X2 U11322 ( .A(n11160), .Z(n11162) );
  INV_X2 U11323 ( .A(n12521), .ZN(n10017) );
  INV_X2 U11324 ( .A(n19852), .ZN(n16322) );
  NAND2_X1 U11326 ( .A1(n10104), .A2(n10103), .ZN(n10191) );
  BUF_X1 U11327 ( .A(n17192), .Z(n9585) );
  NAND2_X2 U11328 ( .A1(n14352), .A2(n9979), .ZN(n14407) );
  XNOR2_X2 U11329 ( .A(n14995), .B(n12440), .ZN(n14988) );
  NOR2_X2 U11330 ( .A1(n14979), .A2(n12444), .ZN(n12469) );
  NOR2_X4 U11331 ( .A1(n14407), .A2(n14408), .ZN(n14399) );
  AND2_X4 U11332 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10739) );
  AND2_X2 U11333 ( .A1(n13758), .A2(n13893), .ZN(n13892) );
  NOR2_X2 U11334 ( .A1(n13719), .A2(n13759), .ZN(n13758) );
  NOR2_X2 U11335 ( .A1(n13647), .A2(n13646), .ZN(n13648) );
  OAI21_X2 U11336 ( .B1(n14141), .B2(n14142), .A(n14301), .ZN(n14575) );
  AND2_X4 U11337 ( .A1(n14316), .A2(n12125), .ZN(n14141) );
  AOI21_X1 U11338 ( .B1(n9864), .B2(n9862), .A(n15140), .ZN(n9861) );
  NOR2_X1 U11339 ( .A1(n9866), .A2(n10658), .ZN(n9862) );
  NAND2_X1 U11340 ( .A1(n20084), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11460) );
  AOI21_X1 U11341 ( .B1(n9864), .B2(n9859), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n9858) );
  INV_X1 U11342 ( .A(n9866), .ZN(n9859) );
  NAND2_X1 U11343 ( .A1(n11326), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11522) );
  AND2_X1 U11344 ( .A1(n11379), .A2(n13242), .ZN(n11683) );
  NOR2_X1 U11345 ( .A1(n11326), .A2(n20676), .ZN(n11379) );
  AND4_X1 U11346 ( .A1(n10443), .A2(n10442), .A3(n10441), .A4(n10440), .ZN(
        n10457) );
  AND3_X1 U11347 ( .A1(n10448), .A2(n10447), .A3(n10446), .ZN(n10456) );
  INV_X1 U11348 ( .A(n10559), .ZN(n11175) );
  CLKBUF_X1 U11349 ( .A(n10559), .Z(n14239) );
  AOI21_X1 U11350 ( .B1(n15197), .B2(n9933), .A(n9931), .ZN(n9926) );
  NAND2_X1 U11351 ( .A1(n12773), .A2(n17632), .ZN(n12774) );
  NAND2_X1 U11352 ( .A1(n12772), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12773) );
  OAI21_X1 U11353 ( .B1(n19357), .B2(n11036), .A(n9693), .ZN(n10401) );
  INV_X1 U11354 ( .A(n10197), .ZN(n10198) );
  NAND2_X1 U11355 ( .A1(n10463), .A2(n10462), .ZN(n10474) );
  OR2_X1 U11357 ( .A1(n10397), .A2(n10396), .ZN(n10931) );
  INV_X1 U11358 ( .A(n9864), .ZN(n9860) );
  NAND2_X1 U11359 ( .A1(n9856), .A2(n9855), .ZN(n9854) );
  INV_X1 U11360 ( .A(n9858), .ZN(n9856) );
  INV_X1 U11361 ( .A(n9861), .ZN(n9855) );
  NAND2_X1 U11362 ( .A1(n9861), .A2(n9863), .ZN(n9853) );
  NAND2_X1 U11363 ( .A1(n9864), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9863) );
  NAND2_X1 U11364 ( .A1(n10469), .A2(n10183), .ZN(n10184) );
  AND2_X1 U11365 ( .A1(n14426), .A2(n9981), .ZN(n9980) );
  AND2_X1 U11366 ( .A1(n14430), .A2(n11939), .ZN(n9981) );
  OAI21_X1 U11367 ( .B1(n11613), .B2(n9956), .A(n9952), .ZN(n11622) );
  NAND2_X1 U11368 ( .A1(n9957), .A2(n11615), .ZN(n9956) );
  INV_X1 U11369 ( .A(n9953), .ZN(n9952) );
  INV_X1 U11370 ( .A(n11619), .ZN(n9957) );
  INV_X1 U11371 ( .A(n11586), .ZN(n11518) );
  INV_X1 U11372 ( .A(n14273), .ZN(n14176) );
  AND2_X2 U11373 ( .A1(n11326), .A2(n20122), .ZN(n11320) );
  NOR3_X1 U11374 ( .A1(n10625), .A2(n10591), .A3(P2_EBX_REG_20__SCAN_IN), .ZN(
        n10629) );
  OR2_X1 U11375 ( .A1(n10625), .A2(n10591), .ZN(n10630) );
  INV_X1 U11376 ( .A(n10469), .ZN(n9916) );
  NAND2_X1 U11377 ( .A1(n13028), .A2(n10657), .ZN(n9869) );
  NOR2_X1 U11378 ( .A1(n12612), .A2(n10635), .ZN(n10647) );
  NOR2_X1 U11379 ( .A1(n15160), .A2(n12620), .ZN(n10646) );
  NAND2_X1 U11380 ( .A1(n9996), .A2(n15078), .ZN(n9995) );
  INV_X1 U11381 ( .A(n14017), .ZN(n9996) );
  OAI21_X1 U11382 ( .B1(n15188), .B2(n9932), .A(n12619), .ZN(n9931) );
  NAND2_X1 U11383 ( .A1(n15196), .A2(n12617), .ZN(n9932) );
  NOR2_X1 U11384 ( .A1(n15188), .A2(n9934), .ZN(n9933) );
  INV_X1 U11385 ( .A(n12617), .ZN(n9934) );
  NAND2_X1 U11386 ( .A1(n9701), .A2(n19196), .ZN(n9700) );
  INV_X1 U11387 ( .A(n10926), .ZN(n10472) );
  AND2_X1 U11388 ( .A1(n10902), .A2(n10470), .ZN(n10904) );
  INV_X1 U11389 ( .A(n10904), .ZN(n11063) );
  AND2_X1 U11390 ( .A1(n19206), .A2(n9582), .ZN(n10130) );
  INV_X1 U11391 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10078) );
  INV_X1 U11392 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10077) );
  INV_X1 U11393 ( .A(n16980), .ZN(n12675) );
  OR2_X1 U11394 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15717), .ZN(
        n12670) );
  INV_X1 U11395 ( .A(n17004), .ZN(n12690) );
  NOR2_X1 U11396 ( .A1(n12760), .A2(n9944), .ZN(n9943) );
  OAI21_X1 U11397 ( .B1(n12762), .B2(n12761), .A(n17734), .ZN(n12765) );
  INV_X1 U11398 ( .A(n17347), .ZN(n12932) );
  CLKBUF_X1 U11399 ( .A(n11323), .Z(n13384) );
  NAND2_X1 U11400 ( .A1(n11695), .A2(n20134), .ZN(n13385) );
  AND2_X1 U11401 ( .A1(n9977), .A2(n9976), .ZN(n9975) );
  INV_X1 U11402 ( .A(n14330), .ZN(n9976) );
  AND2_X1 U11403 ( .A1(n11991), .A2(n11990), .ZN(n14416) );
  OAI21_X1 U11404 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n16150), .A(n11686), 
        .ZN(n11687) );
  AND2_X1 U11405 ( .A1(n14965), .A2(n9678), .ZN(n14869) );
  INV_X1 U11406 ( .A(n14871), .ZN(n10037) );
  NOR2_X1 U11407 ( .A1(n11113), .A2(n11114), .ZN(n14251) );
  INV_X1 U11408 ( .A(n15094), .ZN(n14231) );
  NOR3_X1 U11409 ( .A1(n14932), .A2(n9997), .A3(n14017), .ZN(n15079) );
  OR2_X1 U11410 ( .A1(n14935), .A2(n10644), .ZN(n15178) );
  AND2_X1 U11411 ( .A1(n9775), .A2(n15206), .ZN(n9774) );
  OR3_X1 U11412 ( .A1(n12615), .A2(n9779), .A3(n9778), .ZN(n9775) );
  AND2_X1 U11413 ( .A1(n10766), .A2(n13167), .ZN(n11181) );
  NAND2_X1 U11414 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17039), .ZN(n17022) );
  NOR2_X1 U11415 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9821) );
  INV_X1 U11416 ( .A(n12648), .ZN(n9822) );
  NAND2_X1 U11417 ( .A1(n17509), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12771) );
  AOI21_X1 U11418 ( .B1(n17855), .B2(n17632), .A(n17508), .ZN(n12770) );
  NAND2_X1 U11419 ( .A1(n17553), .A2(n17906), .ZN(n17539) );
  AND2_X1 U11420 ( .A1(n12765), .A2(n12763), .ZN(n9810) );
  NAND2_X1 U11421 ( .A1(n17632), .A2(n17952), .ZN(n12763) );
  AND2_X1 U11422 ( .A1(n12809), .A2(n12808), .ZN(n18157) );
  NOR3_X1 U11423 ( .A1(n12807), .A2(n12806), .A3(n12805), .ZN(n12808) );
  AND2_X1 U11424 ( .A1(n16039), .A2(n20057), .ZN(n16007) );
  INV_X1 U11425 ( .A(n20060), .ZN(n19879) );
  OR2_X1 U11426 ( .A1(n14202), .A2(n15022), .ZN(n12961) );
  NAND2_X1 U11427 ( .A1(n20371), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11643) );
  NOR2_X1 U11428 ( .A1(n10416), .A2(n10415), .ZN(n10421) );
  NAND2_X1 U11429 ( .A1(n11640), .A2(n11639), .ZN(n11666) );
  OR2_X1 U11430 ( .A1(n11648), .A2(n11650), .ZN(n11640) );
  INV_X1 U11431 ( .A(n10199), .ZN(n10200) );
  NAND2_X1 U11432 ( .A1(n10211), .A2(n9573), .ZN(n10186) );
  INV_X1 U11433 ( .A(n17336), .ZN(n12918) );
  AOI21_X1 U11434 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n18640), .A(
        n12784), .ZN(n12785) );
  NAND2_X1 U11435 ( .A1(n13359), .A2(n20112), .ZN(n11531) );
  CLKBUF_X1 U11436 ( .A(n11478), .Z(n12059) );
  CLKBUF_X1 U11437 ( .A(n11230), .Z(n12106) );
  AND2_X1 U11438 ( .A1(n11517), .A2(n11516), .ZN(n11586) );
  OR2_X1 U11439 ( .A1(n11668), .A2(n11505), .ZN(n11517) );
  NOR2_X1 U11440 ( .A1(n14276), .A2(n13381), .ZN(n13501) );
  INV_X1 U11441 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n9872) );
  OR2_X1 U11442 ( .A1(n11414), .A2(n11413), .ZN(n11543) );
  NAND2_X1 U11443 ( .A1(n20122), .A2(n11710), .ZN(n13068) );
  NAND2_X1 U11444 ( .A1(n11316), .A2(n13359), .ZN(n11317) );
  NOR2_X1 U11445 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n11185), .ZN(
        n11196) );
  AOI21_X1 U11446 ( .B1(n13212), .B2(n13075), .A(n13104), .ZN(n11325) );
  INV_X1 U11447 ( .A(n10591), .ZN(n9912) );
  NOR2_X1 U11448 ( .A1(P2_EBX_REG_21__SCAN_IN), .A2(P2_EBX_REG_20__SCAN_IN), 
        .ZN(n9911) );
  NAND2_X1 U11449 ( .A1(n9704), .A2(n10238), .ZN(n9705) );
  NAND2_X1 U11450 ( .A1(n10003), .A2(n15422), .ZN(n10002) );
  INV_X1 U11451 ( .A(n15436), .ZN(n10003) );
  NAND2_X1 U11452 ( .A1(n9845), .A2(n9843), .ZN(n9842) );
  INV_X1 U11453 ( .A(n10579), .ZN(n9844) );
  XNOR2_X1 U11454 ( .A(n11166), .B(n11167), .ZN(n11160) );
  NOR2_X1 U11455 ( .A1(n10383), .A2(n9903), .ZN(n9902) );
  NAND2_X1 U11456 ( .A1(n14242), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10227) );
  OAI21_X1 U11457 ( .B1(n10241), .B2(n10485), .A(n10224), .ZN(n10225) );
  NAND2_X1 U11458 ( .A1(n10311), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10080) );
  AOI21_X1 U11459 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n16335), .A(
        n10465), .ZN(n10697) );
  NOR2_X1 U11460 ( .A1(n10464), .A2(n10473), .ZN(n10465) );
  OR2_X1 U11461 ( .A1(n12747), .A2(n17331), .ZN(n12734) );
  NOR2_X1 U11462 ( .A1(n20806), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12906) );
  INV_X1 U11463 ( .A(n20122), .ZN(n11323) );
  AND2_X1 U11464 ( .A1(n9978), .A2(n14389), .ZN(n9977) );
  AND2_X1 U11465 ( .A1(n14344), .A2(n12040), .ZN(n9978) );
  NAND2_X1 U11466 ( .A1(n14832), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12167) );
  INV_X1 U11467 ( .A(n14041), .ZN(n9982) );
  NAND2_X1 U11468 ( .A1(n11818), .A2(n11817), .ZN(n14047) );
  INV_X1 U11469 ( .A(n11713), .ZN(n11764) );
  NAND2_X1 U11470 ( .A1(n14598), .A2(n9690), .ZN(n11635) );
  NOR2_X1 U11471 ( .A1(n14736), .A2(n14698), .ZN(n9959) );
  NOR2_X1 U11472 ( .A1(n13903), .A2(n13902), .ZN(n13925) );
  AND2_X1 U11473 ( .A1(n13530), .A2(n14276), .ZN(n14273) );
  NAND2_X1 U11474 ( .A1(n11553), .A2(n11552), .ZN(n11560) );
  NOR2_X1 U11475 ( .A1(n13364), .A2(n13067), .ZN(n13357) );
  INV_X1 U11476 ( .A(n11683), .ZN(n11668) );
  INV_X1 U11477 ( .A(n11543), .ZN(n11448) );
  NAND2_X1 U11478 ( .A1(n11356), .A2(n20210), .ZN(n11446) );
  NAND2_X1 U11479 ( .A1(n13328), .A2(n20676), .ZN(n11475) );
  NAND2_X1 U11480 ( .A1(n10585), .A2(n18944), .ZN(n10581) );
  NAND2_X1 U11481 ( .A1(n10581), .A2(n10670), .ZN(n10589) );
  NAND2_X1 U11482 ( .A1(n14236), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10476) );
  NAND2_X1 U11483 ( .A1(n10724), .A2(n10470), .ZN(n10477) );
  INV_X1 U11484 ( .A(n14969), .ZN(n10021) );
  NAND2_X1 U11485 ( .A1(n9591), .A2(n10027), .ZN(n10026) );
  INV_X1 U11486 ( .A(n9686), .ZN(n10027) );
  NOR2_X1 U11487 ( .A1(n16234), .A2(n9974), .ZN(n9973) );
  INV_X1 U11488 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n9974) );
  NAND2_X1 U11489 ( .A1(n10257), .A2(n10258), .ZN(n9885) );
  NAND2_X1 U11490 ( .A1(n9832), .A2(n9835), .ZN(n10215) );
  NAND2_X1 U11491 ( .A1(n9838), .A2(n9836), .ZN(n10216) );
  AND2_X1 U11492 ( .A1(n12416), .A2(n10900), .ZN(n10902) );
  INV_X1 U11493 ( .A(n13060), .ZN(n10005) );
  NAND2_X1 U11494 ( .A1(n10674), .A2(n10673), .ZN(n10675) );
  INV_X1 U11495 ( .A(n15131), .ZN(n10674) );
  AND2_X1 U11496 ( .A1(n10052), .A2(n10051), .ZN(n10050) );
  AND2_X1 U11497 ( .A1(n12634), .A2(n14992), .ZN(n10052) );
  NAND2_X1 U11498 ( .A1(n9929), .A2(n15205), .ZN(n9925) );
  INV_X1 U11499 ( .A(n9928), .ZN(n9927) );
  AOI21_X1 U11500 ( .B1(n9931), .B2(n12622), .A(n10066), .ZN(n9928) );
  NOR2_X1 U11501 ( .A1(n12620), .A2(n9930), .ZN(n9929) );
  INV_X1 U11502 ( .A(n9933), .ZN(n9930) );
  NAND2_X1 U11503 ( .A1(n11168), .A2(n11167), .ZN(n11176) );
  NOR2_X1 U11504 ( .A1(n13604), .A2(n10042), .ZN(n10041) );
  INV_X1 U11505 ( .A(n13597), .ZN(n10042) );
  INV_X1 U11507 ( .A(n13825), .ZN(n9993) );
  NAND2_X1 U11508 ( .A1(n11151), .A2(n11150), .ZN(n11153) );
  NOR2_X1 U11509 ( .A1(n10918), .A2(n10917), .ZN(n10924) );
  NAND2_X1 U11510 ( .A1(n10014), .A2(n12266), .ZN(n12268) );
  NAND2_X1 U11511 ( .A1(n10116), .A2(n10115), .ZN(n9764) );
  NOR2_X1 U11512 ( .A1(n16820), .A2(n18157), .ZN(n12883) );
  NOR2_X1 U11513 ( .A1(n14122), .A2(n14121), .ZN(n15714) );
  NOR2_X1 U11514 ( .A1(n17577), .A2(n9747), .ZN(n9746) );
  NAND2_X1 U11515 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n9747) );
  NAND2_X1 U11516 ( .A1(n9684), .A2(n17648), .ZN(n12984) );
  NAND2_X1 U11517 ( .A1(n9941), .A2(n17632), .ZN(n9942) );
  NOR2_X1 U11518 ( .A1(n17744), .A2(n17745), .ZN(n12942) );
  NAND2_X1 U11519 ( .A1(n12915), .A2(n12759), .ZN(n12762) );
  NOR2_X1 U11520 ( .A1(n17327), .A2(n12734), .ZN(n12754) );
  XNOR2_X1 U11521 ( .A(n17347), .B(n17336), .ZN(n12745) );
  NOR2_X1 U11522 ( .A1(n18181), .A2(n18187), .ZN(n12890) );
  OAI21_X1 U11523 ( .B1(n12794), .B2(n12793), .A(n12904), .ZN(n12973) );
  AOI211_X1 U11524 ( .C1(n17156), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n12864), .B(n12863), .ZN(n12865) );
  NOR2_X1 U11525 ( .A1(n9791), .A2(n9784), .ZN(n9783) );
  INV_X1 U11526 ( .A(n12811), .ZN(n9791) );
  NAND2_X1 U11527 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n9785) );
  NAND2_X1 U11528 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n9745) );
  NAND2_X1 U11529 ( .A1(n20760), .A2(n13791), .ZN(n19898) );
  NAND2_X1 U11530 ( .A1(n14303), .A2(n14331), .ZN(n9875) );
  INV_X2 U11531 ( .A(n11328), .ZN(n13413) );
  NOR2_X1 U11532 ( .A1(n9986), .A2(n14302), .ZN(n9985) );
  INV_X1 U11533 ( .A(n14142), .ZN(n9986) );
  AND2_X1 U11534 ( .A1(n14549), .A2(n12142), .ZN(n12197) );
  OR2_X1 U11535 ( .A1(n12121), .A2(n14322), .ZN(n12146) );
  AND2_X1 U11536 ( .A1(n14626), .A2(n9687), .ZN(n9960) );
  AND2_X1 U11537 ( .A1(n9980), .A2(n14416), .ZN(n9979) );
  NOR2_X1 U11538 ( .A1(n11954), .A2(n14360), .ZN(n11955) );
  NAND2_X1 U11539 ( .A1(n11955), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11988) );
  AND2_X1 U11540 ( .A1(n14088), .A2(n14089), .ZN(n14090) );
  NAND2_X1 U11541 ( .A1(n11754), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11758) );
  NAND2_X1 U11542 ( .A1(n11729), .A2(n11728), .ZN(n13526) );
  AND2_X1 U11543 ( .A1(n14753), .A2(n14694), .ZN(n14740) );
  NOR3_X1 U11544 ( .A1(n14800), .A2(n14079), .A3(n9883), .ZN(n14450) );
  NOR2_X1 U11545 ( .A1(n14800), .A2(n14079), .ZN(n14106) );
  NOR2_X1 U11546 ( .A1(n14642), .A2(n14636), .ZN(n14781) );
  NOR2_X1 U11547 ( .A1(n9626), .A2(n9729), .ZN(n9728) );
  INV_X1 U11548 ( .A(n11607), .ZN(n9729) );
  NAND2_X1 U11549 ( .A1(n9881), .A2(n9880), .ZN(n13903) );
  INV_X1 U11550 ( .A(n13765), .ZN(n9880) );
  XNOR2_X1 U11551 ( .A(n11560), .B(n13775), .ZN(n13610) );
  INV_X1 U11552 ( .A(n13381), .ZN(n13530) );
  NAND2_X1 U11553 ( .A1(n11720), .A2(n20082), .ZN(n20214) );
  NOR2_X1 U11554 ( .A1(n11720), .A2(n9587), .ZN(n20483) );
  OR2_X1 U11555 ( .A1(n10691), .A2(n10690), .ZN(n14235) );
  OR2_X1 U11556 ( .A1(n10680), .A2(n10679), .ZN(n10691) );
  AND2_X1 U11557 ( .A1(n10633), .A2(n10632), .ZN(n14927) );
  AND2_X1 U11558 ( .A1(n13039), .A2(n14903), .ZN(n14905) );
  NAND2_X1 U11559 ( .A1(n15554), .A2(n10939), .ZN(n15533) );
  NOR2_X2 U11560 ( .A1(n13052), .A2(n14893), .ZN(n13051) );
  NAND2_X1 U11561 ( .A1(n12994), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12993) );
  OR2_X1 U11562 ( .A1(n15011), .A2(n15010), .ZN(n15013) );
  NAND2_X1 U11563 ( .A1(n13012), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13014) );
  AND2_X1 U11564 ( .A1(n13656), .A2(n9649), .ZN(n13833) );
  INV_X1 U11565 ( .A(n13754), .ZN(n10030) );
  NAND2_X1 U11566 ( .A1(n13007), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13006) );
  INV_X1 U11567 ( .A(n9885), .ZN(n10265) );
  AND2_X1 U11568 ( .A1(n9869), .A2(n15326), .ZN(n9866) );
  INV_X1 U11569 ( .A(n9869), .ZN(n9865) );
  NAND2_X1 U11570 ( .A1(n15328), .A2(n15326), .ZN(n9868) );
  AND2_X1 U11571 ( .A1(n12640), .A2(n9612), .ZN(n15152) );
  NAND2_X1 U11572 ( .A1(n12640), .A2(n9610), .ZN(n15331) );
  OAI21_X1 U11573 ( .B1(n9772), .B2(n9713), .A(n10647), .ZN(n9712) );
  NAND2_X1 U11574 ( .A1(n12640), .A2(n11178), .ZN(n15333) );
  AND2_X1 U11575 ( .A1(n11092), .A2(n11091), .ZN(n14017) );
  OR2_X1 U11576 ( .A1(n13965), .A2(n14934), .ZN(n14932) );
  NAND2_X1 U11577 ( .A1(n9773), .A2(n16199), .ZN(n15207) );
  NAND2_X1 U11578 ( .A1(n12613), .A2(n9779), .ZN(n9773) );
  INV_X1 U11579 ( .A(n12612), .ZN(n9771) );
  AND2_X1 U11580 ( .A1(n15517), .A2(n10010), .ZN(n15455) );
  AND2_X1 U11581 ( .A1(n9655), .A2(n10011), .ZN(n10010) );
  INV_X1 U11582 ( .A(n15467), .ZN(n10011) );
  NAND2_X1 U11583 ( .A1(n15517), .A2(n9655), .ZN(n15479) );
  AND2_X1 U11584 ( .A1(n15517), .A2(n10012), .ZN(n15481) );
  INV_X1 U11585 ( .A(n10480), .ZN(n9760) );
  INV_X1 U11586 ( .A(n10479), .ZN(n9759) );
  NOR2_X1 U11587 ( .A1(n10324), .A2(n10323), .ZN(n13400) );
  AND2_X1 U11588 ( .A1(n13257), .A2(n13258), .ZN(n13256) );
  AND2_X1 U11589 ( .A1(n18828), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12629) );
  NAND2_X1 U11590 ( .A1(n15601), .A2(n12636), .ZN(n12637) );
  OAI21_X1 U11591 ( .B1(n10097), .B2(n10096), .A(n10115), .ZN(n10104) );
  NAND2_X1 U11592 ( .A1(n10102), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10103) );
  INV_X1 U11593 ( .A(n10095), .ZN(n10096) );
  NOR2_X1 U11594 ( .A1(n12898), .A2(n18163), .ZN(n16496) );
  NOR2_X1 U11595 ( .A1(n18151), .A2(n15706), .ZN(n17408) );
  NAND2_X1 U11596 ( .A1(n9749), .A2(n9748), .ZN(n16597) );
  NAND2_X1 U11597 ( .A1(n9590), .A2(n12981), .ZN(n9748) );
  OR2_X1 U11598 ( .A1(n16613), .A2(n9665), .ZN(n9749) );
  OR2_X1 U11599 ( .A1(n16613), .A2(n17545), .ZN(n9750) );
  INV_X1 U11600 ( .A(n16838), .ZN(n9590) );
  NAND2_X1 U11601 ( .A1(n17121), .A2(n9736), .ZN(n9737) );
  NOR2_X1 U11602 ( .A1(n14125), .A2(n16745), .ZN(n9736) );
  NOR2_X1 U11603 ( .A1(n17159), .A2(n17163), .ZN(n9738) );
  INV_X1 U11604 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n20864) );
  NAND2_X1 U11605 ( .A1(n12644), .A2(n18623), .ZN(n16980) );
  NOR2_X1 U11606 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12644) );
  INV_X1 U11607 ( .A(n9622), .ZN(n17056) );
  INV_X1 U11608 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n20809) );
  AOI21_X1 U11609 ( .B1(n17131), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n12692), .ZN(n12697) );
  NOR2_X1 U11610 ( .A1(n12661), .A2(n20864), .ZN(n12692) );
  INV_X1 U11611 ( .A(n12671), .ZN(n9937) );
  NAND2_X1 U11612 ( .A1(n12674), .A2(n12673), .ZN(n9936) );
  NAND2_X1 U11613 ( .A1(n12681), .A2(n12680), .ZN(n12682) );
  AOI21_X1 U11614 ( .B1(n17137), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n12679), .ZN(n12680) );
  NOR2_X1 U11615 ( .A1(n10053), .A2(n17128), .ZN(n12679) );
  AND2_X1 U11616 ( .A1(n12740), .A2(n9824), .ZN(n9823) );
  NOR2_X1 U11617 ( .A1(n9826), .A2(n9825), .ZN(n9824) );
  OAI22_X1 U11618 ( .A1(n17088), .A2(n17024), .B1(n17090), .B2(n20773), .ZN(
        n9825) );
  NOR2_X1 U11619 ( .A1(n9565), .A2(n18154), .ZN(n12737) );
  NOR2_X1 U11620 ( .A1(n17501), .A2(n17502), .ZN(n17486) );
  AND2_X1 U11621 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n9755) );
  NOR2_X1 U11622 ( .A1(n16374), .A2(n16362), .ZN(n16359) );
  NOR2_X1 U11623 ( .A1(n9608), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9947) );
  NAND2_X1 U11624 ( .A1(n17475), .A2(n9806), .ZN(n15742) );
  AND2_X1 U11625 ( .A1(n17632), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9806) );
  NOR2_X2 U11626 ( .A1(n12775), .A2(n17484), .ZN(n17475) );
  NAND2_X1 U11627 ( .A1(n17493), .A2(n17843), .ZN(n17492) );
  INV_X1 U11628 ( .A(n17851), .ZN(n9801) );
  INV_X1 U11629 ( .A(n17595), .ZN(n9802) );
  OAI21_X1 U11630 ( .B1(n17612), .B2(n17506), .A(n12767), .ZN(n12768) );
  OR3_X1 U11631 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17539), .ZN(n12767) );
  NAND3_X1 U11632 ( .A1(n12768), .A2(n17525), .A3(n17878), .ZN(n17520) );
  NOR2_X1 U11633 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n12766), .ZN(
        n17553) );
  NAND4_X1 U11634 ( .A1(n9808), .A2(n17943), .A3(n9810), .A4(n9621), .ZN(
        n17604) );
  NAND2_X1 U11635 ( .A1(n9941), .A2(n9807), .ZN(n9808) );
  AND2_X1 U11636 ( .A1(n17632), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9807) );
  AND2_X1 U11637 ( .A1(n12765), .A2(n12764), .ZN(n17612) );
  NOR2_X1 U11638 ( .A1(n12880), .A2(n15724), .ZN(n18611) );
  INV_X1 U11639 ( .A(n17316), .ZN(n16403) );
  NOR2_X1 U11640 ( .A1(n9816), .A2(n9819), .ZN(n9813) );
  INV_X1 U11641 ( .A(n9818), .ZN(n9816) );
  NAND2_X1 U11642 ( .A1(n9814), .A2(n9812), .ZN(n9921) );
  NOR2_X1 U11643 ( .A1(n9813), .A2(n17756), .ZN(n9812) );
  OR2_X1 U11644 ( .A1(n9817), .A2(n17783), .ZN(n9814) );
  NOR2_X1 U11645 ( .A1(n9818), .A2(n9625), .ZN(n9817) );
  AND2_X1 U11646 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12751), .ZN(
        n12752) );
  INV_X1 U11647 ( .A(n17783), .ZN(n9815) );
  NOR2_X1 U11648 ( .A1(n12750), .A2(n17797), .ZN(n17785) );
  XNOR2_X1 U11649 ( .A(n9914), .B(n9913), .ZN(n17798) );
  INV_X1 U11650 ( .A(n12748), .ZN(n9913) );
  NOR2_X1 U11651 ( .A1(n17817), .A2(n12744), .ZN(n17806) );
  INV_X1 U11652 ( .A(n16868), .ZN(n18623) );
  AND2_X1 U11653 ( .A1(n13412), .A2(n13156), .ZN(n20760) );
  AND2_X1 U11654 ( .A1(n14540), .A2(n13386), .ZN(n15961) );
  AND2_X1 U11655 ( .A1(n14540), .A2(n13391), .ZN(n15959) );
  INV_X1 U11656 ( .A(n14540), .ZN(n15957) );
  NAND2_X1 U11657 ( .A1(n19879), .A2(n12207), .ZN(n16039) );
  AND2_X1 U11658 ( .A1(n12206), .A2(n12205), .ZN(n16031) );
  AND2_X1 U11659 ( .A1(n13364), .A2(n11694), .ZN(n20060) );
  NOR2_X1 U11660 ( .A1(n16318), .A2(n19714), .ZN(n18829) );
  NOR2_X1 U11661 ( .A1(n14864), .A2(n13016), .ZN(n14197) );
  OR2_X1 U11662 ( .A1(n14197), .A2(n15087), .ZN(n14857) );
  NOR2_X1 U11663 ( .A1(n14865), .A2(n15102), .ZN(n14864) );
  INV_X2 U11664 ( .A(n15027), .ZN(n15022) );
  AND2_X1 U11665 ( .A1(n15027), .A2(n9584), .ZN(n15018) );
  NAND2_X1 U11666 ( .A1(n14247), .A2(n10867), .ZN(n14202) );
  NAND2_X1 U11667 ( .A1(n18832), .A2(n12628), .ZN(n16259) );
  AND2_X1 U11668 ( .A1(n16259), .A2(n13407), .ZN(n19175) );
  NAND3_X1 U11669 ( .A1(n19802), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19656), 
        .ZN(n19179) );
  INV_X1 U11670 ( .A(n19169), .ZN(n16245) );
  XNOR2_X1 U11671 ( .A(n14251), .B(n14250), .ZN(n19045) );
  INV_X1 U11672 ( .A(n10008), .ZN(n10007) );
  OAI21_X1 U11673 ( .B1(n14259), .B2(n16295), .A(n14258), .ZN(n10008) );
  XNOR2_X1 U11674 ( .A(n9847), .B(n9620), .ZN(n14270) );
  NAND2_X1 U11675 ( .A1(n9848), .A2(n9641), .ZN(n9847) );
  NAND2_X1 U11676 ( .A1(n15116), .A2(n10047), .ZN(n15273) );
  NAND2_X1 U11677 ( .A1(n15275), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10046) );
  XNOR2_X1 U11678 ( .A(n9766), .B(n9656), .ZN(n15374) );
  NAND2_X1 U11679 ( .A1(n9768), .A2(n9767), .ZN(n9766) );
  INV_X1 U11680 ( .A(n16294), .ZN(n16280) );
  NAND2_X1 U11681 ( .A1(n15400), .A2(n13277), .ZN(n16297) );
  AND2_X1 U11682 ( .A1(n11181), .A2(n19842), .ZN(n16301) );
  INV_X1 U11683 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19837) );
  OR2_X1 U11684 ( .A1(n15584), .A2(n13231), .ZN(n19830) );
  INV_X1 U11685 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19828) );
  INV_X1 U11686 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n18828) );
  INV_X1 U11687 ( .A(n18825), .ZN(n18821) );
  INV_X1 U11688 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18805) );
  INV_X1 U11689 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18809) );
  INV_X1 U11690 ( .A(n16884), .ZN(n16869) );
  AOI22_X1 U11691 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n15648), .B1(
        n9574), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12876) );
  NOR2_X1 U11692 ( .A1(n16993), .A2(n9734), .ZN(n9731) );
  NOR3_X1 U11693 ( .A1(n16675), .A2(n17038), .A3(n17022), .ZN(n17008) );
  INV_X1 U11694 ( .A(n17138), .ZN(n17103) );
  AND2_X1 U11695 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17167), .ZN(n17164) );
  INV_X1 U11696 ( .A(n17169), .ZN(n17167) );
  INV_X1 U11697 ( .A(n17240), .ZN(n18193) );
  INV_X1 U11698 ( .A(n17184), .ZN(n17191) );
  NOR2_X1 U11699 ( .A1(n9944), .A2(n17726), .ZN(n17599) );
  NAND2_X1 U11700 ( .A1(n17316), .A2(n9797), .ZN(n9796) );
  XNOR2_X1 U11701 ( .A(n10067), .B(n16370), .ZN(n16368) );
  NAND2_X1 U11702 ( .A1(n9805), .A2(n9804), .ZN(n10067) );
  INV_X1 U11703 ( .A(n15797), .ZN(n9804) );
  NOR2_X1 U11704 ( .A1(n18119), .A2(n18608), .ZN(n18048) );
  NAND2_X1 U11705 ( .A1(n18157), .A2(n9586), .ZN(n18107) );
  NAND2_X1 U11706 ( .A1(n11644), .A2(n11643), .ZN(n11674) );
  NAND2_X1 U11707 ( .A1(n11666), .A2(n11642), .ZN(n11644) );
  OAI22_X1 U11708 ( .A1(n10399), .A2(n10543), .B1(n9696), .B2(n12365), .ZN(
        n10528) );
  NAND2_X1 U11709 ( .A1(n10373), .A2(n10374), .ZN(n9903) );
  NOR2_X1 U11710 ( .A1(n17113), .A2(n12812), .ZN(n9788) );
  OAI21_X1 U11711 ( .B1(n11619), .B2(n9954), .A(n11618), .ZN(n9953) );
  INV_X1 U11712 ( .A(n11615), .ZN(n9955) );
  NAND2_X1 U11713 ( .A1(n11503), .A2(n11502), .ZN(n11575) );
  OR2_X1 U11714 ( .A1(n11488), .A2(n11487), .ZN(n11569) );
  NAND2_X1 U11715 ( .A1(n9951), .A2(n14290), .ZN(n9950) );
  AND2_X1 U11716 ( .A1(n13793), .A2(n11336), .ZN(n9951) );
  NAND2_X1 U11717 ( .A1(n11454), .A2(n11346), .ZN(n11443) );
  NAND4_X1 U11718 ( .A1(n19206), .A2(n12592), .A3(n9916), .A4(n10183), .ZN(
        n10211) );
  NAND2_X1 U11719 ( .A1(n10237), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9838) );
  AOI21_X2 U11720 ( .B1(n10868), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n9837), 
        .ZN(n9836) );
  AND2_X1 U11721 ( .A1(n19861), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n9837) );
  OAI21_X1 U11722 ( .B1(n9566), .B2(n10214), .A(n9834), .ZN(n9833) );
  NAND2_X1 U11723 ( .A1(n10509), .A2(n10508), .ZN(n11166) );
  INV_X1 U11724 ( .A(n10244), .ZN(n9917) );
  INV_X1 U11725 ( .A(n10468), .ZN(n11139) );
  NAND2_X1 U11726 ( .A1(n10201), .A2(n9573), .ZN(n10202) );
  NAND2_X1 U11727 ( .A1(n10751), .A2(n9710), .ZN(n10878) );
  NAND2_X1 U11728 ( .A1(n10199), .A2(n10184), .ZN(n9711) );
  OR2_X1 U11729 ( .A1(n10703), .A2(n10702), .ZN(n10704) );
  NAND2_X1 U11730 ( .A1(n12754), .A2(n12753), .ZN(n12733) );
  AOI21_X1 U11731 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18635), .A(
        n12783), .ZN(n12788) );
  NOR2_X1 U11732 ( .A1(n12905), .A2(n12782), .ZN(n12783) );
  AND2_X1 U11733 ( .A1(n9790), .A2(n9787), .ZN(n9786) );
  NOR2_X1 U11734 ( .A1(n9789), .A2(n9788), .ZN(n9787) );
  NAND2_X1 U11735 ( .A1(n17141), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n9790) );
  OAI22_X1 U11736 ( .A1(n17004), .A2(n17035), .B1(n17108), .B2(n17024), .ZN(
        n9789) );
  OR2_X1 U11737 ( .A1(n20122), .A2(n11329), .ZN(n11271) );
  INV_X1 U11738 ( .A(n14401), .ZN(n12040) );
  OR2_X1 U11739 ( .A1(n11855), .A2(n15923), .ZN(n11870) );
  NAND2_X1 U11740 ( .A1(n9661), .A2(n9603), .ZN(n9983) );
  INV_X1 U11741 ( .A(n14082), .ZN(n9984) );
  INV_X1 U11742 ( .A(n13917), .ZN(n11818) );
  AND2_X1 U11743 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n11732), .ZN(
        n11744) );
  NOR2_X1 U11744 ( .A1(n11722), .A2(n13810), .ZN(n11732) );
  NAND2_X1 U11745 ( .A1(n14449), .A2(n14105), .ZN(n9882) );
  OR2_X1 U11746 ( .A1(n11515), .A2(n11514), .ZN(n11609) );
  NAND2_X1 U11747 ( .A1(n14276), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n9870) );
  NAND2_X1 U11748 ( .A1(n13501), .A2(n9872), .ZN(n9871) );
  NAND2_X1 U11749 ( .A1(n14168), .A2(n14838), .ZN(n9873) );
  NAND2_X1 U11750 ( .A1(n13212), .A2(n20102), .ZN(n12217) );
  INV_X1 U11751 ( .A(n11320), .ZN(n13098) );
  AND3_X1 U11752 ( .A1(n11692), .A2(n13216), .A3(n11693), .ZN(n13100) );
  OR2_X1 U11753 ( .A1(n11668), .A2(n11404), .ZN(n11416) );
  OR2_X1 U11754 ( .A1(n11378), .A2(n11377), .ZN(n11380) );
  INV_X1 U11755 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n20888) );
  AND2_X1 U11756 ( .A1(n13213), .A2(n11320), .ZN(n11321) );
  AND3_X1 U11757 ( .A1(n11218), .A2(n11215), .A3(n11214), .ZN(n9714) );
  INV_X1 U11758 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20371) );
  AOI221_X1 U11759 ( .B1(n20763), .B2(n14849), .C1(n13592), .C2(n14849), .A(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n20088) );
  NAND2_X1 U11760 ( .A1(n11522), .A2(n11460), .ZN(n11688) );
  NOR2_X1 U11761 ( .A1(n10883), .A2(n19213), .ZN(n9828) );
  NAND2_X1 U11762 ( .A1(n9901), .A2(n9900), .ZN(n10724) );
  NAND2_X1 U11763 ( .A1(n13035), .A2(n10475), .ZN(n9900) );
  NAND2_X1 U11764 ( .A1(n10701), .A2(n10926), .ZN(n9901) );
  INV_X1 U11765 ( .A(n10655), .ZN(n9907) );
  NOR2_X1 U11766 ( .A1(n9910), .A2(n9909), .ZN(n9908) );
  INV_X1 U11767 ( .A(n10622), .ZN(n9909) );
  NAND2_X1 U11768 ( .A1(n9912), .A2(n9911), .ZN(n9910) );
  NAND2_X1 U11769 ( .A1(n10589), .A2(n10583), .ZN(n10617) );
  AND2_X1 U11770 ( .A1(n10564), .A2(n9650), .ZN(n10585) );
  INV_X1 U11771 ( .A(n15053), .ZN(n10006) );
  INV_X1 U11772 ( .A(n15017), .ZN(n10028) );
  CLKBUF_X1 U11773 ( .A(n10700), .Z(n10880) );
  NOR2_X1 U11774 ( .A1(n9967), .A2(n9965), .ZN(n9964) );
  INV_X1 U11775 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n9965) );
  INV_X1 U11776 ( .A(n10685), .ZN(n9709) );
  AND2_X1 U11777 ( .A1(n14964), .A2(n10039), .ZN(n10038) );
  INV_X1 U11778 ( .A(n13058), .ZN(n10039) );
  OR2_X1 U11779 ( .A1(n14898), .A2(n11175), .ZN(n10686) );
  NAND2_X1 U11780 ( .A1(n9858), .A2(n9860), .ZN(n9852) );
  INV_X1 U11781 ( .A(n15443), .ZN(n9713) );
  INV_X1 U11782 ( .A(n16199), .ZN(n9778) );
  OR2_X1 U11783 ( .A1(n12615), .A2(n9778), .ZN(n9777) );
  OR2_X1 U11784 ( .A1(n9667), .A2(n10002), .ZN(n10001) );
  NOR2_X1 U11785 ( .A1(n13958), .A2(n13957), .ZN(n10036) );
  NOR2_X1 U11786 ( .A1(n12614), .A2(n9780), .ZN(n9779) );
  INV_X1 U11787 ( .A(n15216), .ZN(n9780) );
  NOR2_X1 U11788 ( .A1(n15453), .A2(n10002), .ZN(n13976) );
  NOR2_X1 U11789 ( .A1(n15432), .A2(n10620), .ZN(n9899) );
  INV_X1 U11790 ( .A(n9840), .ZN(n9839) );
  OAI21_X1 U11791 ( .B1(n9654), .B2(n9595), .A(n9842), .ZN(n9840) );
  AND2_X1 U11792 ( .A1(n13655), .A2(n10032), .ZN(n10031) );
  INV_X1 U11793 ( .A(n13684), .ZN(n10032) );
  NOR2_X1 U11794 ( .A1(n13853), .A2(n10013), .ZN(n10012) );
  INV_X1 U11795 ( .A(n15516), .ZN(n10013) );
  NAND2_X1 U11796 ( .A1(n10478), .A2(n18995), .ZN(n10506) );
  OR2_X1 U11797 ( .A1(n10436), .A2(n10435), .ZN(n10935) );
  INV_X1 U11798 ( .A(n13949), .ZN(n9991) );
  AOI22_X1 U11799 ( .A1(n10987), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10315) );
  NOR2_X1 U11800 ( .A1(n10339), .A2(n10338), .ZN(n11141) );
  NAND4_X1 U11801 ( .A1(n10230), .A2(n10229), .A3(n10058), .A4(n10228), .ZN(
        n10257) );
  AND2_X1 U11802 ( .A1(n19213), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12247) );
  INV_X1 U11803 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10074) );
  INV_X1 U11804 ( .A(n10233), .ZN(n13934) );
  NAND2_X1 U11805 ( .A1(n10142), .A2(n10141), .ZN(n10165) );
  NAND2_X1 U11806 ( .A1(n10140), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10141) );
  AND2_X1 U11807 ( .A1(n12246), .A2(n10299), .ZN(n10288) );
  INV_X2 U11808 ( .A(n10165), .ZN(n10889) );
  NAND2_X1 U11809 ( .A1(n10080), .A2(n10079), .ZN(n10081) );
  NAND2_X1 U11810 ( .A1(n10076), .A2(n10075), .ZN(n10082) );
  AND2_X1 U11811 ( .A1(n10713), .A2(n10712), .ZN(n10730) );
  AOI221_X1 U11812 ( .B1(n10697), .B2(n16308), .C1(n10697), .C2(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n10696), .ZN(n10734) );
  NAND2_X1 U11813 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18769), .ZN(
        n12647) );
  INV_X1 U11814 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n20871) );
  INV_X1 U11815 ( .A(n12735), .ZN(n9826) );
  INV_X1 U11816 ( .A(n15716), .ZN(n15705) );
  AND2_X1 U11817 ( .A1(n16496), .A2(n12883), .ZN(n15708) );
  NAND2_X1 U11818 ( .A1(n17486), .A2(n9605), .ZN(n12909) );
  OAI21_X1 U11819 ( .B1(n16402), .B2(n16403), .A(n17734), .ZN(n12756) );
  AOI21_X1 U11820 ( .B1(n12752), .B2(n9819), .A(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n9818) );
  NOR2_X1 U11821 ( .A1(n12881), .A2(n12894), .ZN(n12901) );
  NOR2_X1 U11822 ( .A1(n17408), .A2(n15708), .ZN(n12879) );
  NAND2_X1 U11823 ( .A1(n9794), .A2(n9792), .ZN(n12898) );
  NOR2_X1 U11824 ( .A1(n15723), .A2(n9793), .ZN(n9792) );
  NAND2_X1 U11825 ( .A1(n18175), .A2(n18169), .ZN(n9793) );
  INV_X1 U11826 ( .A(n12892), .ZN(n15711) );
  OAI21_X1 U11827 ( .B1(n12891), .B2(n12890), .A(n12889), .ZN(n12892) );
  AOI211_X1 U11828 ( .C1(n12888), .C2(n18169), .A(n12887), .B(n12902), .ZN(
        n12889) );
  OAI21_X1 U11829 ( .B1(n18193), .B2(n18629), .A(n12882), .ZN(n15710) );
  INV_X1 U11830 ( .A(n18029), .ZN(n18628) );
  NAND2_X1 U11831 ( .A1(n12901), .A2(n18612), .ZN(n14121) );
  AOI211_X1 U11832 ( .C1(n17105), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n12824), .B(n12823), .ZN(n12825) );
  NAND2_X1 U11833 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12804) );
  INV_X1 U11834 ( .A(n12802), .ZN(n12807) );
  OAI211_X1 U11835 ( .C1(n10053), .C2(n18184), .A(n12847), .B(n12846), .ZN(
        n15727) );
  AOI211_X1 U11836 ( .C1(n17131), .C2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n12845), .B(n12844), .ZN(n12846) );
  NAND2_X1 U11837 ( .A1(n18181), .A2(n12901), .ZN(n15706) );
  INV_X1 U11838 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13810) );
  INV_X1 U11839 ( .A(n14168), .ZN(n14277) );
  AND2_X1 U11840 ( .A1(n13364), .A2(n13241), .ZN(n20925) );
  OR2_X1 U11841 ( .A1(n12149), .A2(n12148), .ZN(n12209) );
  AOI21_X1 U11842 ( .B1(n12145), .B2(n12144), .A(n12143), .ZN(n14142) );
  NAND2_X1 U11843 ( .A1(n12124), .A2(n12123), .ZN(n14318) );
  AND2_X1 U11844 ( .A1(n12082), .A2(n12081), .ZN(n14389) );
  AND2_X1 U11845 ( .A1(n14615), .A2(n12142), .ZN(n12056) );
  NOR2_X1 U11846 ( .A1(n12036), .A2(n14622), .ZN(n12037) );
  NOR2_X1 U11847 ( .A1(n11988), .A2(n15983), .ZN(n11989) );
  AND2_X1 U11848 ( .A1(n15980), .A2(n12142), .ZN(n11971) );
  AND2_X1 U11849 ( .A1(n11957), .A2(n11956), .ZN(n14430) );
  OR2_X1 U11850 ( .A1(n11923), .A2(n15880), .ZN(n11954) );
  NAND2_X1 U11851 ( .A1(n11627), .A2(n11626), .ZN(n14627) );
  NAND2_X1 U11852 ( .A1(n11890), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11907) );
  AND2_X1 U11853 ( .A1(n11875), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11890) );
  NOR2_X1 U11854 ( .A1(n13917), .A2(n9983), .ZN(n14048) );
  AND2_X1 U11855 ( .A1(n11811), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11812) );
  NAND2_X1 U11856 ( .A1(n11812), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11855) );
  NOR2_X1 U11857 ( .A1(n11807), .A2(n11806), .ZN(n11811) );
  AND3_X1 U11858 ( .A1(n11781), .A2(n11780), .A3(n11779), .ZN(n13759) );
  NOR2_X1 U11859 ( .A1(n11758), .A2(n11761), .ZN(n11782) );
  INV_X1 U11860 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11761) );
  CLKBUF_X1 U11861 ( .A(n13719), .Z(n13720) );
  OAI211_X1 U11862 ( .C1(n11764), .C2(n11757), .A(n11756), .B(n11755), .ZN(
        n13757) );
  AND2_X1 U11863 ( .A1(n11744), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11754) );
  AOI21_X1 U11864 ( .B1(n11752), .B2(n11887), .A(n11751), .ZN(n13646) );
  INV_X1 U11865 ( .A(n11750), .ZN(n11751) );
  NAND2_X1 U11866 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11722) );
  NOR2_X1 U11867 ( .A1(n11635), .A2(n14556), .ZN(n14545) );
  INV_X1 U11868 ( .A(n11635), .ZN(n11634) );
  NOR2_X1 U11869 ( .A1(n9877), .A2(n9876), .ZN(n14333) );
  NAND2_X1 U11870 ( .A1(n14412), .A2(n14404), .ZN(n14403) );
  NAND2_X1 U11871 ( .A1(n9879), .A2(n9878), .ZN(n14420) );
  INV_X1 U11872 ( .A(n14418), .ZN(n9878) );
  NAND2_X1 U11873 ( .A1(n14627), .A2(n14626), .ZN(n15809) );
  AND2_X1 U11874 ( .A1(n14147), .A2(n14146), .ZN(n14445) );
  NAND2_X1 U11875 ( .A1(n9719), .A2(n14633), .ZN(n14642) );
  NAND2_X1 U11876 ( .A1(n16011), .A2(n9720), .ZN(n9719) );
  INV_X1 U11877 ( .A(n14634), .ZN(n9720) );
  OR2_X1 U11878 ( .A1(n15931), .A2(n14062), .ZN(n14800) );
  INV_X1 U11879 ( .A(n16011), .ZN(n14653) );
  NAND2_X1 U11880 ( .A1(n16012), .A2(n11615), .ZN(n16011) );
  NAND2_X1 U11881 ( .A1(n11613), .A2(n9958), .ZN(n16012) );
  NAND2_X1 U11882 ( .A1(n13925), .A2(n13924), .ZN(n15931) );
  AND2_X1 U11883 ( .A1(n13726), .A2(n13725), .ZN(n13730) );
  NAND2_X1 U11884 ( .A1(n16137), .A2(n16136), .ZN(n16135) );
  AND2_X1 U11885 ( .A1(n13107), .A2(n13089), .ZN(n14692) );
  OAI21_X1 U11886 ( .B1(n20171), .B2(n11678), .A(n11530), .ZN(n13095) );
  NAND2_X1 U11887 ( .A1(n13095), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13097) );
  NOR2_X1 U11888 ( .A1(n20122), .A2(n13385), .ZN(n9725) );
  OR2_X1 U11889 ( .A1(n11668), .A2(n11435), .ZN(n11437) );
  INV_X1 U11890 ( .A(n11334), .ZN(n13072) );
  INV_X1 U11891 ( .A(n13091), .ZN(n14832) );
  AND2_X1 U11892 ( .A1(n13370), .A2(n13369), .ZN(n15765) );
  INV_X1 U11893 ( .A(n20117), .ZN(n20133) );
  INV_X1 U11894 ( .A(n20248), .ZN(n20506) );
  AOI21_X1 U11895 ( .B1(n20536), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20257), 
        .ZN(n20622) );
  NAND2_X1 U11896 ( .A1(n10700), .A2(n10212), .ZN(n12587) );
  CLKBUF_X1 U11897 ( .A(n12416), .Z(n19853) );
  NAND2_X1 U11898 ( .A1(n10670), .A2(n10662), .ZN(n14234) );
  NOR2_X1 U11899 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n10672), .ZN(n10676) );
  NAND2_X1 U11900 ( .A1(n14234), .A2(n10677), .ZN(n10680) );
  NAND2_X1 U11901 ( .A1(n10649), .A2(n9904), .ZN(n10672) );
  NOR2_X1 U11902 ( .A1(n9905), .A2(n10652), .ZN(n9904) );
  NAND2_X1 U11903 ( .A1(n9907), .A2(n9906), .ZN(n9905) );
  NOR2_X1 U11904 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(P2_EBX_REG_24__SCAN_IN), 
        .ZN(n9906) );
  NOR3_X1 U11905 ( .A1(n10654), .A2(n10655), .A3(P2_EBX_REG_24__SCAN_IN), .ZN(
        n10667) );
  NOR2_X1 U11906 ( .A1(n13008), .A2(n15210), .ZN(n13011) );
  NAND2_X1 U11907 ( .A1(n10564), .A2(n9629), .ZN(n10580) );
  NAND2_X1 U11908 ( .A1(n10564), .A2(n9628), .ZN(n10574) );
  NAND2_X1 U11909 ( .A1(n10555), .A2(n10554), .ZN(n10558) );
  NAND2_X1 U11910 ( .A1(n10490), .A2(n10491), .ZN(n10489) );
  NAND2_X1 U11911 ( .A1(n15026), .A2(n14936), .ZN(n15011) );
  OR2_X1 U11912 ( .A1(n12294), .A2(n12293), .ZN(n13994) );
  NAND2_X1 U11913 ( .A1(n10022), .A2(n10021), .ZN(n10020) );
  NAND2_X1 U11914 ( .A1(n14905), .A2(n9672), .ZN(n14873) );
  NAND2_X1 U11915 ( .A1(n14905), .A2(n9671), .ZN(n15050) );
  NAND2_X1 U11916 ( .A1(n14905), .A2(n14214), .ZN(n15052) );
  XNOR2_X1 U11917 ( .A(n12469), .B(n12471), .ZN(n14975) );
  NAND2_X1 U11918 ( .A1(n14975), .A2(n14974), .ZN(n14973) );
  OAI22_X1 U11919 ( .A1(n14988), .A2(n10024), .B1(n9619), .B2(n14980), .ZN(
        n14979) );
  OR2_X1 U11920 ( .A1(n14980), .A2(n14987), .ZN(n10024) );
  OR2_X1 U11921 ( .A1(n14988), .A2(n14987), .ZN(n10025) );
  NAND2_X1 U11922 ( .A1(n14915), .A2(n15335), .ZN(n9994) );
  AND3_X1 U11923 ( .A1(n10999), .A2(n10998), .A3(n10997), .ZN(n15467) );
  AND2_X1 U11924 ( .A1(n19083), .A2(n12605), .ZN(n13255) );
  INV_X1 U11925 ( .A(n10698), .ZN(n13273) );
  INV_X1 U11926 ( .A(n12602), .ZN(n13675) );
  NAND2_X1 U11927 ( .A1(n13049), .A2(n9604), .ZN(n14194) );
  AND2_X1 U11928 ( .A1(n13049), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14195) );
  NOR2_X1 U11929 ( .A1(n13010), .A2(n15190), .ZN(n13012) );
  NOR2_X1 U11930 ( .A1(n15024), .A2(n15023), .ZN(n15026) );
  NOR2_X1 U11931 ( .A1(n13006), .A2(n18917), .ZN(n13009) );
  NAND2_X1 U11932 ( .A1(n13656), .A2(n9627), .ZN(n13753) );
  AND2_X1 U11933 ( .A1(n13003), .A2(n9601), .ZN(n13007) );
  NAND2_X1 U11934 ( .A1(n13003), .A2(n9594), .ZN(n13004) );
  AND2_X1 U11935 ( .A1(n13003), .A2(n9973), .ZN(n13005) );
  NAND2_X1 U11936 ( .A1(n13003), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13002) );
  INV_X1 U11937 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15229) );
  NOR2_X1 U11938 ( .A1(n12998), .A2(n9963), .ZN(n9961) );
  NAND2_X1 U11939 ( .A1(n13543), .A2(n13597), .ZN(n13605) );
  NAND2_X1 U11940 ( .A1(n9643), .A2(n9962), .ZN(n12999) );
  NOR2_X1 U11941 ( .A1(n12998), .A2(n16260), .ZN(n13000) );
  CLKBUF_X2 U11942 ( .A(n10911), .Z(n14248) );
  AND2_X1 U11943 ( .A1(n14905), .A2(n9675), .ZN(n14872) );
  INV_X1 U11944 ( .A(n14874), .ZN(n10004) );
  NOR3_X1 U11945 ( .A1(n10689), .A2(n11175), .A3(n15099), .ZN(n15094) );
  NOR2_X1 U11946 ( .A1(n14880), .A2(n11175), .ZN(n15111) );
  NOR2_X1 U11947 ( .A1(n13057), .A2(n11175), .ZN(n15110) );
  NAND2_X1 U11948 ( .A1(n14965), .A2(n10038), .ZN(n14870) );
  NAND2_X1 U11949 ( .A1(n14965), .A2(n14964), .ZN(n14967) );
  AND2_X1 U11950 ( .A1(n10686), .A2(n15291), .ZN(n15127) );
  AND2_X1 U11951 ( .A1(n10050), .A2(n10049), .ZN(n10048) );
  INV_X1 U11952 ( .A(n14902), .ZN(n10049) );
  CLKBUF_X1 U11953 ( .A(n14209), .Z(n15129) );
  NAND2_X1 U11954 ( .A1(n14922), .A2(n10050), .ZN(n14901) );
  NAND2_X1 U11955 ( .A1(n14922), .A2(n10052), .ZN(n14994) );
  NOR3_X1 U11956 ( .A1(n14932), .A2(n9995), .A3(n9997), .ZN(n15334) );
  AND2_X1 U11957 ( .A1(n10643), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15160) );
  AOI21_X1 U11958 ( .B1(n9929), .B2(n9923), .A(n9927), .ZN(n9922) );
  INV_X1 U11959 ( .A(n15206), .ZN(n9923) );
  INV_X1 U11960 ( .A(n15178), .ZN(n9769) );
  NOR2_X1 U11961 ( .A1(n15453), .A2(n9998), .ZN(n15412) );
  NAND2_X1 U11962 ( .A1(n10000), .A2(n9999), .ZN(n9998) );
  INV_X1 U11963 ( .A(n15411), .ZN(n9999) );
  INV_X1 U11964 ( .A(n10001), .ZN(n10000) );
  NAND2_X1 U11965 ( .A1(n10036), .A2(n10035), .ZN(n15024) );
  INV_X1 U11966 ( .A(n13997), .ZN(n10035) );
  INV_X1 U11967 ( .A(n15400), .ZN(n9892) );
  INV_X1 U11968 ( .A(n10036), .ZN(n13998) );
  OR2_X1 U11969 ( .A1(n16276), .A2(n15350), .ZN(n16261) );
  NAND2_X1 U11970 ( .A1(n12613), .A2(n15216), .ZN(n16202) );
  INV_X1 U11971 ( .A(n13976), .ZN(n15423) );
  NAND2_X1 U11972 ( .A1(n15445), .A2(n15443), .ZN(n9770) );
  NAND2_X1 U11973 ( .A1(n9898), .A2(n9899), .ZN(n16196) );
  NOR2_X1 U11974 ( .A1(n15448), .A2(n15432), .ZN(n15433) );
  NOR2_X1 U11975 ( .A1(n15453), .A2(n15436), .ZN(n15435) );
  NAND2_X1 U11976 ( .A1(n15490), .A2(n9654), .ZN(n9846) );
  AND2_X1 U11977 ( .A1(n13656), .A2(n10031), .ZN(n13707) );
  NAND2_X1 U11978 ( .A1(n13656), .A2(n13655), .ZN(n13683) );
  OR3_X1 U11979 ( .A1(n11176), .A2(n11175), .A3(n11174), .ZN(n11177) );
  XNOR2_X1 U11980 ( .A(n11173), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15500) );
  OR2_X1 U11981 ( .A1(n11176), .A2(n11175), .ZN(n11173) );
  AND2_X1 U11982 ( .A1(n10041), .A2(n10043), .ZN(n10040) );
  NAND2_X1 U11983 ( .A1(n13543), .A2(n10041), .ZN(n13631) );
  NAND2_X1 U11984 ( .A1(n10943), .A2(n10942), .ZN(n15517) );
  NAND2_X1 U11985 ( .A1(n15517), .A2(n15516), .ZN(n15518) );
  NAND2_X1 U11986 ( .A1(n15234), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11165) );
  NAND2_X1 U11987 ( .A1(n15553), .A2(n15549), .ZN(n11163) );
  XNOR2_X1 U11988 ( .A(n10565), .B(n15537), .ZN(n15235) );
  NAND2_X1 U11989 ( .A1(n9831), .A2(n10505), .ZN(n15548) );
  NOR2_X1 U11990 ( .A1(n13281), .A2(n9990), .ZN(n15556) );
  NAND2_X1 U11991 ( .A1(n9992), .A2(n9991), .ZN(n9990) );
  AND2_X1 U11992 ( .A1(n10896), .A2(n16297), .ZN(n13884) );
  NAND2_X1 U11993 ( .A1(n9988), .A2(n10905), .ZN(n13257) );
  NAND2_X1 U11994 ( .A1(n10903), .A2(n10904), .ZN(n9988) );
  INV_X1 U11995 ( .A(n13400), .ZN(n10903) );
  INV_X1 U11996 ( .A(n10183), .ZN(n13229) );
  AOI21_X1 U11997 ( .B1(n15568), .B2(n12629), .A(n12257), .ZN(n13234) );
  NOR2_X1 U11998 ( .A1(n13281), .A2(n10925), .ZN(n13826) );
  CLKBUF_X1 U11999 ( .A(n10316), .Z(n13937) );
  NAND2_X1 U12000 ( .A1(n13324), .A2(n13323), .ZN(n13461) );
  INV_X1 U12001 ( .A(n12266), .ZN(n10015) );
  NAND2_X1 U12002 ( .A1(n19178), .A2(n13911), .ZN(n9829) );
  INV_X1 U12003 ( .A(n10403), .ZN(n19188) );
  INV_X1 U12004 ( .A(n19323), .ZN(n19328) );
  INV_X1 U12005 ( .A(n19383), .ZN(n19319) );
  AND2_X1 U12006 ( .A1(n19235), .A2(n19231), .ZN(n19416) );
  AND2_X1 U12007 ( .A1(n19810), .A2(n19183), .ZN(n19232) );
  INV_X1 U12008 ( .A(n19500), .ZN(n19494) );
  INV_X1 U12009 ( .A(n19353), .ZN(n19352) );
  INV_X1 U12010 ( .A(n19802), .ZN(n19609) );
  NAND2_X1 U12011 ( .A1(n10147), .A2(n10115), .ZN(n10154) );
  NOR2_X1 U12012 ( .A1(n19235), .A2(n19830), .ZN(n19184) );
  CLKBUF_X1 U12013 ( .A(n10469), .Z(n10470) );
  NOR2_X2 U12014 ( .A1(n13674), .A2(n19179), .ZN(n19222) );
  NAND2_X1 U12015 ( .A1(n19805), .A2(n19830), .ZN(n19604) );
  INV_X1 U12016 ( .A(n19221), .ZN(n19217) );
  INV_X1 U12017 ( .A(n19222), .ZN(n19219) );
  INV_X1 U12018 ( .A(n19603), .ZN(n19652) );
  INV_X1 U12019 ( .A(n19656), .ZN(n19421) );
  INV_X1 U12020 ( .A(n10744), .ZN(n16348) );
  OAI22_X1 U12021 ( .A1(n16566), .A2(n9590), .B1(n9590), .B2(n17466), .ZN(
        n16545) );
  INV_X1 U12022 ( .A(n17577), .ZN(n16642) );
  INV_X1 U12023 ( .A(n17602), .ZN(n16665) );
  NAND2_X1 U12024 ( .A1(n17008), .A2(n9732), .ZN(n16963) );
  AND2_X1 U12025 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n9733), .ZN(n9732) );
  NOR2_X1 U12026 ( .A1(n9735), .A2(n9734), .ZN(n9733) );
  INV_X1 U12027 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n9735) );
  CLKBUF_X1 U12028 ( .A(n12670), .Z(n17146) );
  INV_X1 U12029 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16966) );
  NAND2_X1 U12030 ( .A1(n9741), .A2(n18812), .ZN(n15826) );
  OR2_X1 U12031 ( .A1(n15714), .A2(n9742), .ZN(n9741) );
  NOR3_X1 U12032 ( .A1(n14123), .A2(n14124), .A3(n17240), .ZN(n9742) );
  INV_X1 U12033 ( .A(n15827), .ZN(n18629) );
  NOR2_X1 U12034 ( .A1(n12909), .A2(n17823), .ZN(n16381) );
  NOR2_X1 U12035 ( .A1(n17463), .A2(n9752), .ZN(n9751) );
  NAND2_X1 U12036 ( .A1(n17486), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17462) );
  NAND2_X1 U12037 ( .A1(n9592), .A2(n9659), .ZN(n17501) );
  OAI21_X1 U12038 ( .B1(n17823), .B2(n17564), .A(n18313), .ZN(n17617) );
  INV_X1 U12039 ( .A(n9746), .ZN(n17567) );
  NAND2_X1 U12040 ( .A1(n16665), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17577) );
  NOR2_X1 U12041 ( .A1(n12984), .A2(n17618), .ZN(n17614) );
  INV_X1 U12042 ( .A(n18007), .ZN(n17699) );
  NAND2_X1 U12043 ( .A1(n12947), .A2(n17735), .ZN(n17698) );
  NOR2_X1 U12044 ( .A1(n17787), .A2(n17789), .ZN(n16808) );
  NOR2_X1 U12045 ( .A1(n18157), .A2(n18657), .ZN(n9797) );
  AND2_X1 U12046 ( .A1(n12775), .A2(n9945), .ZN(n15797) );
  NOR2_X1 U12047 ( .A1(n9946), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9945) );
  INV_X1 U12048 ( .A(n9947), .ZN(n9946) );
  INV_X1 U12049 ( .A(n17836), .ZN(n17461) );
  INV_X1 U12050 ( .A(n17520), .ZN(n12769) );
  NOR2_X1 U12051 ( .A1(n17632), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17593) );
  INV_X1 U12052 ( .A(n17552), .ZN(n9803) );
  NOR2_X1 U12053 ( .A1(n17733), .A2(n12760), .ZN(n17635) );
  NOR2_X1 U12054 ( .A1(n18007), .A2(n17975), .ZN(n17993) );
  INV_X1 U12055 ( .A(n12899), .ZN(n12970) );
  INV_X1 U12056 ( .A(n9942), .ZN(n17733) );
  NOR2_X1 U12057 ( .A1(n12898), .A2(n12897), .ZN(n12969) );
  AOI21_X1 U12058 ( .B1(n12796), .B2(n12795), .A(n12973), .ZN(n18601) );
  INV_X1 U12059 ( .A(n12896), .ZN(n18610) );
  INV_X1 U12060 ( .A(n18620), .ZN(n18613) );
  NAND2_X1 U12061 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18613), .ZN(
        n18617) );
  NAND3_X1 U12062 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15717) );
  NOR2_X1 U12063 ( .A1(n12816), .A2(n9782), .ZN(n18151) );
  NOR2_X1 U12064 ( .A1(n12856), .A2(n9744), .ZN(n9743) );
  INV_X1 U12065 ( .A(n18508), .ZN(n18312) );
  AOI22_X1 U12066 ( .A1(n18601), .A2(n18597), .B1(n18111), .B2(n18602), .ZN(
        n18606) );
  NAND2_X1 U12067 ( .A1(n13801), .A2(n13799), .ZN(n19901) );
  INV_X1 U12068 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14360) );
  AND2_X1 U12069 ( .A1(n19898), .A2(n13808), .ZN(n19909) );
  NAND2_X1 U12070 ( .A1(n13801), .A2(n13800), .ZN(n19960) );
  AND2_X1 U12071 ( .A1(n19898), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19969) );
  INV_X1 U12072 ( .A(n19923), .ZN(n19977) );
  INV_X1 U12073 ( .A(n19901), .ZN(n19914) );
  CLKBUF_X1 U12074 ( .A(n19923), .Z(n19942) );
  OR2_X1 U12075 ( .A1(n19936), .A2(n13794), .ZN(n19983) );
  INV_X1 U12076 ( .A(n19960), .ZN(n19974) );
  OR2_X1 U12077 ( .A1(n14306), .A2(n14305), .ZN(n14381) );
  INV_X1 U12078 ( .A(n14457), .ZN(n19989) );
  AND2_X1 U12079 ( .A1(n13379), .A2(n13378), .ZN(n19994) );
  NAND2_X1 U12080 ( .A1(n19994), .A2(n13380), .ZN(n14457) );
  INV_X1 U12081 ( .A(n14458), .ZN(n15960) );
  NAND2_X1 U12082 ( .A1(n13393), .A2(n13392), .ZN(n14095) );
  NAND2_X1 U12083 ( .A1(n9726), .A2(n9680), .ZN(n12225) );
  INV_X1 U12084 ( .A(n14095), .ZN(n14542) );
  INV_X1 U12085 ( .A(n15961), .ZN(n14544) );
  NOR2_X1 U12086 ( .A1(n20021), .A2(n20925), .ZN(n20007) );
  CLKBUF_X1 U12087 ( .A(n20007), .Z(n20924) );
  INV_X1 U12088 ( .A(n14417), .ZN(n15973) );
  AOI21_X1 U12089 ( .B1(n14092), .B2(n14091), .A(n14090), .ZN(n16005) );
  INV_X1 U12090 ( .A(n16031), .ZN(n20081) );
  NAND2_X1 U12091 ( .A1(n16139), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n9723) );
  XNOR2_X1 U12092 ( .A(n15995), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16071) );
  NAND2_X1 U12093 ( .A1(n11613), .A2(n11612), .ZN(n14026) );
  NAND2_X1 U12094 ( .A1(n16024), .A2(n11607), .ZN(n13989) );
  NAND2_X1 U12095 ( .A1(n9948), .A2(n11561), .ZN(n13690) );
  NOR2_X1 U12096 ( .A1(n13776), .A2(n16093), .ZN(n20074) );
  INV_X1 U12097 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20536) );
  CLKBUF_X1 U12098 ( .A(n13870), .Z(n20372) );
  CLKBUF_X1 U12099 ( .A(n13571), .Z(n13572) );
  NAND2_X1 U12100 ( .A1(n11554), .A2(n14822), .ZN(n11555) );
  AND2_X1 U12101 ( .A1(n13093), .A2(n13797), .ZN(n14834) );
  INV_X1 U12102 ( .A(n14137), .ZN(n14849) );
  NOR2_X1 U12103 ( .A1(n20841), .A2(n15758), .ZN(n14137) );
  OR2_X1 U12104 ( .A1(n20214), .A2(n20347), .ZN(n20252) );
  OR2_X1 U12105 ( .A1(n20348), .A2(n20424), .ZN(n20370) );
  AND2_X1 U12106 ( .A1(n20564), .A2(n20506), .ZN(n20559) );
  INV_X1 U12107 ( .A(n20441), .ZN(n20629) );
  INV_X1 U12108 ( .A(n20445), .ZN(n20635) );
  INV_X1 U12109 ( .A(n20449), .ZN(n20641) );
  INV_X1 U12110 ( .A(n20453), .ZN(n20647) );
  INV_X1 U12111 ( .A(n20457), .ZN(n20653) );
  INV_X1 U12112 ( .A(n20461), .ZN(n20659) );
  AND2_X1 U12113 ( .A1(n20564), .A2(n20482), .ZN(n20670) );
  INV_X1 U12114 ( .A(n20466), .ZN(n20666) );
  INV_X1 U12115 ( .A(n13364), .ZN(n15758) );
  INV_X2 U12116 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20679) );
  INV_X1 U12117 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20677) );
  NOR2_X1 U12118 ( .A1(n13016), .A2(n14196), .ZN(n14882) );
  NAND2_X1 U12119 ( .A1(n13016), .A2(n15144), .ZN(n9968) );
  NOR2_X1 U12120 ( .A1(n15153), .A2(n14911), .ZN(n9970) );
  NOR2_X1 U12121 ( .A1(n15747), .A2(n13016), .ZN(n13019) );
  NOR2_X1 U12122 ( .A1(n13019), .A2(n15153), .ZN(n13053) );
  INV_X1 U12123 ( .A(n19025), .ZN(n19009) );
  OR2_X1 U12124 ( .A1(n18829), .A2(n13027), .ZN(n18993) );
  INV_X1 U12125 ( .A(n18993), .ZN(n19031) );
  INV_X1 U12126 ( .A(n19720), .ZN(n19002) );
  INV_X1 U12127 ( .A(n19011), .ZN(n19022) );
  OR2_X1 U12128 ( .A1(n11043), .A2(n11042), .ZN(n13751) );
  INV_X1 U12129 ( .A(n15018), .ZN(n15030) );
  AND2_X1 U12130 ( .A1(n13255), .A2(n13674), .ZN(n19052) );
  AND2_X1 U12131 ( .A1(n19083), .A2(n10194), .ZN(n19050) );
  NOR2_X1 U12132 ( .A1(n19100), .A2(n19111), .ZN(n19095) );
  AND2_X1 U12133 ( .A1(n19083), .A2(n12591), .ZN(n19100) );
  INV_X1 U12134 ( .A(n19083), .ZN(n19110) );
  OR2_X1 U12135 ( .A1(n19050), .A2(n13255), .ZN(n19085) );
  AND2_X1 U12136 ( .A1(n13272), .A2(n19854), .ZN(n19144) );
  INV_X1 U12137 ( .A(n19144), .ZN(n19154) );
  INV_X2 U12138 ( .A(n19147), .ZN(n19151) );
  NOR2_X1 U12139 ( .A1(n13121), .A2(n13037), .ZN(n13130) );
  XNOR2_X1 U12140 ( .A(n12992), .B(n12991), .ZN(n14265) );
  NAND2_X1 U12141 ( .A1(n9613), .A2(n9897), .ZN(n9896) );
  INV_X1 U12142 ( .A(n15402), .ZN(n9897) );
  INV_X1 U12143 ( .A(n16269), .ZN(n18912) );
  INV_X1 U12144 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18917) );
  INV_X1 U12145 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16234) );
  INV_X1 U12146 ( .A(n19175), .ZN(n19165) );
  INV_X1 U12147 ( .A(n16259), .ZN(n19166) );
  NAND2_X1 U12148 ( .A1(n9857), .A2(n9864), .ZN(n15142) );
  NAND2_X1 U12149 ( .A1(n15330), .A2(n9866), .ZN(n9857) );
  OAI21_X1 U12150 ( .B1(n15330), .B2(n15328), .A(n15326), .ZN(n15151) );
  NOR2_X1 U12151 ( .A1(n14932), .A2(n14017), .ZN(n14916) );
  INV_X1 U12152 ( .A(n9926), .ZN(n15180) );
  OAI21_X1 U12153 ( .B1(n15197), .B2(n15196), .A(n12617), .ZN(n15189) );
  OAI21_X1 U12154 ( .B1(n15201), .B2(n9893), .A(n9890), .ZN(n15418) );
  NOR2_X1 U12155 ( .A1(n15398), .A2(n16270), .ZN(n9893) );
  AND2_X1 U12156 ( .A1(n15399), .A2(n9891), .ZN(n9890) );
  NAND2_X1 U12157 ( .A1(n9892), .A2(n16267), .ZN(n9891) );
  INV_X1 U12158 ( .A(n9894), .ZN(n15551) );
  NAND2_X1 U12159 ( .A1(n11156), .A2(n11155), .ZN(n15550) );
  NAND2_X1 U12160 ( .A1(n10498), .A2(n13879), .ZN(n13946) );
  NAND2_X1 U12161 ( .A1(n10481), .A2(n11148), .ZN(n9888) );
  INV_X1 U12162 ( .A(n16295), .ZN(n16283) );
  NAND2_X1 U12163 ( .A1(n13237), .A2(n13236), .ZN(n19822) );
  OR2_X1 U12164 ( .A1(n13235), .A2(n13234), .ZN(n13236) );
  INV_X1 U12165 ( .A(n19235), .ZN(n19805) );
  NAND2_X1 U12166 ( .A1(n19023), .A2(n12629), .ZN(n12255) );
  INV_X1 U12167 ( .A(n19822), .ZN(n19183) );
  OAI21_X1 U12168 ( .B1(n13326), .B2(n13325), .A(n13324), .ZN(n19810) );
  AND2_X1 U12169 ( .A1(n13323), .A2(n13322), .ZN(n13326) );
  INV_X1 U12170 ( .A(n16350), .ZN(n15601) );
  CLKBUF_X1 U12171 ( .A(n13168), .Z(n13171) );
  NOR2_X1 U12172 ( .A1(n19237), .A2(n19383), .ZN(n19256) );
  NOR3_X1 U12173 ( .A1(n19292), .A2(P2_STATE2_REG_3__SCAN_IN), .A3(n9697), 
        .ZN(n19293) );
  AND2_X1 U12174 ( .A1(n19388), .A2(n19390), .ZN(n19452) );
  AND2_X1 U12175 ( .A1(n19184), .A2(n19232), .ZN(n19499) );
  INV_X1 U12176 ( .A(n19482), .ZN(n19489) );
  INV_X1 U12177 ( .A(n19704), .ZN(n19545) );
  INV_X1 U12178 ( .A(n19661), .ZN(n19606) );
  INV_X1 U12179 ( .A(n19645), .ZN(n19633) );
  INV_X1 U12180 ( .A(n19693), .ZN(n19634) );
  INV_X1 U12181 ( .A(n19620), .ZN(n19658) );
  INV_X1 U12182 ( .A(n19565), .ZN(n19670) );
  INV_X1 U12183 ( .A(n19709), .ZN(n19677) );
  OAI22_X1 U12184 ( .A1(n14510), .A2(n19219), .B1(n20844), .B2(n19217), .ZN(
        n19684) );
  OAI22_X1 U12185 ( .A1(n14498), .A2(n19219), .B1(n20807), .B2(n19217), .ZN(
        n19696) );
  INV_X1 U12186 ( .A(n19680), .ZN(n19705) );
  OAI22_X1 U12187 ( .A1(n19220), .A2(n19219), .B1(n19218), .B2(n19217), .ZN(
        n19704) );
  AND2_X1 U12188 ( .A1(n16314), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16350) );
  INV_X1 U12189 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n10900) );
  NOR2_X1 U12190 ( .A1(n16558), .A2(n16559), .ZN(n16557) );
  NOR2_X1 U12191 ( .A1(n16566), .A2(n9590), .ZN(n16558) );
  OAI21_X1 U12192 ( .B1(n16590), .B2(n9590), .A(n9602), .ZN(n12985) );
  NOR2_X1 U12193 ( .A1(n16577), .A2(n16578), .ZN(n16576) );
  NOR2_X1 U12194 ( .A1(n16590), .A2(n9590), .ZN(n16577) );
  AND2_X1 U12195 ( .A1(n9750), .A2(n16838), .ZN(n16598) );
  NOR2_X1 U12196 ( .A1(n16620), .A2(n9590), .ZN(n16613) );
  INV_X1 U12197 ( .A(n9750), .ZN(n16612) );
  NOR2_X1 U12198 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16650), .ZN(n16630) );
  NOR2_X1 U12199 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16724), .ZN(n16706) );
  INV_X1 U12200 ( .A(n18660), .ZN(n16824) );
  NAND2_X1 U12201 ( .A1(n12975), .A2(n18652), .ZN(n16830) );
  INV_X1 U12202 ( .A(n16875), .ZN(n16866) );
  NOR2_X2 U12203 ( .A1(n18759), .A2(n16869), .ZN(n16875) );
  INV_X1 U12204 ( .A(n16830), .ZN(n16872) );
  INV_X1 U12205 ( .A(n16833), .ZN(n16881) );
  NAND4_X1 U12206 ( .A1(n18137), .A2(n18821), .A3(n16824), .A4(n12976), .ZN(
        n16884) );
  NOR2_X1 U12207 ( .A1(n16947), .A2(n16920), .ZN(n16928) );
  AND2_X1 U12208 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16946), .ZN(n16941) );
  AND2_X1 U12209 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16962), .ZN(n16946) );
  NOR2_X1 U12210 ( .A1(n16948), .A2(n16947), .ZN(n16962) );
  NAND2_X1 U12211 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16975), .ZN(n16947) );
  NOR2_X1 U12212 ( .A1(n16963), .A2(n17240), .ZN(n16975) );
  NOR2_X1 U12213 ( .A1(n15697), .A2(n14126), .ZN(n17039) );
  OR2_X1 U12214 ( .A1(n9737), .A2(n16725), .ZN(n15697) );
  NAND2_X1 U12215 ( .A1(n17121), .A2(P3_EBX_REG_11__SCAN_IN), .ZN(n17072) );
  AND2_X1 U12216 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17103), .ZN(n17121) );
  NAND2_X1 U12217 ( .A1(n17164), .A2(n9611), .ZN(n17138) );
  NOR2_X1 U12218 ( .A1(n17184), .A2(n17172), .ZN(n17170) );
  NAND2_X1 U12219 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17170), .ZN(n17169) );
  NAND2_X1 U12220 ( .A1(n9740), .A2(n9739), .ZN(n17184) );
  NOR2_X1 U12221 ( .A1(n18157), .A2(n18151), .ZN(n9739) );
  INV_X1 U12222 ( .A(n15826), .ZN(n9740) );
  INV_X1 U12223 ( .A(n17208), .ZN(n17203) );
  NOR2_X1 U12224 ( .A1(n17353), .A2(n17216), .ZN(n17212) );
  INV_X1 U12225 ( .A(n17222), .ZN(n17217) );
  NAND2_X1 U12226 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17217), .ZN(n17216) );
  NOR2_X1 U12227 ( .A1(n17240), .A2(n17235), .ZN(n17231) );
  NOR2_X1 U12228 ( .A1(n17240), .A2(n17275), .ZN(n17269) );
  NAND2_X1 U12229 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17269), .ZN(n17268) );
  INV_X1 U12230 ( .A(n17278), .ZN(n17267) );
  NAND2_X1 U12231 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17279), .ZN(n17275) );
  INV_X1 U12232 ( .A(n17242), .ZN(n17274) );
  NAND2_X1 U12233 ( .A1(n17197), .A2(n10063), .ZN(n17284) );
  NOR2_X1 U12234 ( .A1(n18193), .A2(n17340), .ZN(n17305) );
  INV_X1 U12235 ( .A(n12920), .ZN(n17320) );
  INV_X1 U12236 ( .A(n12919), .ZN(n17327) );
  AOI211_X2 U12237 ( .C1(n17141), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n12710), .B(n12709), .ZN(n17331) );
  AND2_X1 U12238 ( .A1(n12698), .A2(n12697), .ZN(n9940) );
  INV_X1 U12239 ( .A(n12695), .ZN(n12696) );
  INV_X1 U12240 ( .A(n17305), .ZN(n17335) );
  INV_X1 U12241 ( .A(n17341), .ZN(n17339) );
  AOI21_X1 U12242 ( .B1(n17131), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n9939), .ZN(n9938) );
  NOR2_X1 U12243 ( .A1(n12683), .A2(n12682), .ZN(n12684) );
  NOR2_X1 U12244 ( .A1(n9937), .A2(n9936), .ZN(n9935) );
  NAND2_X1 U12245 ( .A1(n9630), .A2(n10056), .ZN(n17826) );
  AND2_X1 U12246 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12742) );
  INV_X1 U12247 ( .A(n17343), .ZN(n17326) );
  NOR2_X1 U12248 ( .A1(n17335), .A2(n18629), .ZN(n17341) );
  NOR2_X1 U12249 ( .A1(n17454), .A2(n18157), .ZN(n17455) );
  INV_X1 U12250 ( .A(n16400), .ZN(n16401) );
  NAND2_X1 U12251 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17824), .ZN(n17666) );
  NAND2_X1 U12252 ( .A1(n16403), .A2(n17820), .ZN(n17737) );
  AOI22_X1 U12253 ( .A1(n17698), .A2(n17816), .B1(n17739), .B2(n17699), .ZN(
        n17726) );
  INV_X1 U12254 ( .A(n9615), .ZN(n17739) );
  NOR2_X1 U12255 ( .A1(n17787), .A2(n17759), .ZN(n9756) );
  NAND2_X1 U12256 ( .A1(n9755), .A2(n9754), .ZN(n17758) );
  INV_X1 U12257 ( .A(n17787), .ZN(n9754) );
  INV_X1 U12258 ( .A(n17827), .ZN(n17786) );
  INV_X1 U12259 ( .A(n18542), .ZN(n18313) );
  NOR2_X1 U12260 ( .A1(n18606), .A2(n9795), .ZN(n17820) );
  INV_X1 U12261 ( .A(n9797), .ZN(n9795) );
  INV_X1 U12262 ( .A(n17816), .ZN(n17832) );
  NAND2_X1 U12263 ( .A1(n12775), .A2(n9947), .ZN(n15741) );
  INV_X2 U12264 ( .A(n18107), .ZN(n18597) );
  AND2_X1 U12265 ( .A1(n12768), .A2(n17525), .ZN(n17521) );
  INV_X1 U12266 ( .A(n17525), .ZN(n17538) );
  NAND2_X1 U12267 ( .A1(n18029), .A2(n18626), .ZN(n18119) );
  AND2_X1 U12268 ( .A1(n9809), .A2(n9810), .ZN(n17605) );
  NAND2_X1 U12269 ( .A1(n12764), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9809) );
  NOR2_X1 U12270 ( .A1(n18116), .A2(n17905), .ZN(n17951) );
  AND2_X1 U12271 ( .A1(n12896), .A2(n9781), .ZN(n18029) );
  NAND2_X1 U12272 ( .A1(n12970), .A2(n18611), .ZN(n9781) );
  CLKBUF_X1 U12273 ( .A(n17732), .Z(n18042) );
  NAND2_X1 U12274 ( .A1(n9814), .A2(n9811), .ZN(n17757) );
  INV_X1 U12275 ( .A(n9813), .ZN(n9811) );
  NAND2_X1 U12276 ( .A1(n9815), .A2(n9625), .ZN(n17771) );
  NOR2_X1 U12277 ( .A1(n17783), .A2(n12752), .ZN(n17772) );
  INV_X1 U12278 ( .A(n18609), .ZN(n18626) );
  NOR3_X1 U12279 ( .A1(n12902), .A2(n15709), .A3(n15731), .ZN(n18111) );
  INV_X1 U12280 ( .A(n18630), .ZN(n18608) );
  NOR2_X1 U12281 ( .A1(n18603), .A2(n18116), .ZN(n18132) );
  INV_X1 U12282 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18640) );
  INV_X1 U12283 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18643) );
  INV_X1 U12284 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18783) );
  AOI21_X1 U12285 ( .B1(n18812), .B2(n18627), .A(n15715), .ZN(n18790) );
  INV_X1 U12286 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18607) );
  INV_X1 U12287 ( .A(n18790), .ZN(n18788) );
  INV_X1 U12288 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18178) );
  INV_X1 U12289 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18244) );
  INV_X1 U12290 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18759) );
  NAND2_X1 U12292 ( .A1(n18682), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18817) );
  AND2_X1 U12293 ( .A1(n12238), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20079)
         );
  AND2_X1 U12295 ( .A1(n13793), .A2(n14290), .ZN(n13158) );
  AOI21_X1 U12296 ( .B1(n14554), .B2(n16031), .A(n14553), .ZN(n14555) );
  OAI21_X1 U12297 ( .B1(n16071), .B2(n16070), .A(n9721), .ZN(P1_U3014) );
  NOR2_X1 U12298 ( .A1(n9724), .A2(n9722), .ZN(n9721) );
  OAI21_X1 U12299 ( .B1(n16069), .B2(n16068), .A(n9723), .ZN(n9722) );
  NOR2_X1 U12300 ( .A1(n16072), .A2(n16073), .ZN(n9724) );
  AOI21_X1 U12301 ( .B1(n14197), .B2(n15087), .A(n19720), .ZN(n14198) );
  AND2_X1 U12302 ( .A1(n12961), .A2(n12960), .ZN(n12962) );
  NAND2_X1 U12303 ( .A1(n15374), .A2(n19167), .ZN(n15176) );
  NAND2_X1 U12304 ( .A1(n10009), .A2(n10007), .ZN(n14260) );
  OR2_X1 U12305 ( .A1(n19045), .A2(n16294), .ZN(n10009) );
  NOR2_X1 U12306 ( .A1(n11137), .A2(n11136), .ZN(n11183) );
  OAI21_X1 U12307 ( .B1(n15273), .B2(n16305), .A(n10046), .ZN(n10045) );
  NAND2_X1 U12308 ( .A1(n17008), .A2(P3_EBX_REG_18__SCAN_IN), .ZN(n16992) );
  NAND2_X1 U12309 ( .A1(n17164), .A2(P3_EBX_REG_7__SCAN_IN), .ZN(n17160) );
  AND3_X1 U12310 ( .A1(n9800), .A2(n9598), .A3(n9799), .ZN(n16369) );
  INV_X1 U12311 ( .A(n16367), .ZN(n9799) );
  OR2_X1 U12312 ( .A1(n16398), .A2(n18772), .ZN(n9919) );
  AOI211_X1 U12313 ( .C1(n16368), .C2(n18033), .A(n16363), .B(n15800), .ZN(
        n15801) );
  AND4_X1 U12314 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A4(n9962), .ZN(n9588) );
  INV_X1 U12315 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16260) );
  NAND2_X1 U12317 ( .A1(n13964), .A2(n9688), .ZN(n13963) );
  AND2_X1 U12318 ( .A1(n9688), .A2(n10028), .ZN(n9591) );
  AND2_X1 U12319 ( .A1(n9746), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9592) );
  AND2_X1 U12320 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9761) );
  AND2_X1 U12321 ( .A1(n14352), .A2(n9980), .ZN(n14415) );
  AND2_X1 U12322 ( .A1(n9973), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9594) );
  NAND2_X1 U12323 ( .A1(n14399), .A2(n9977), .ZN(n14329) );
  OAI211_X1 U12324 ( .C1(n10053), .C2(n18178), .A(n12826), .B(n12825), .ZN(
        n14124) );
  OR2_X1 U12325 ( .A1(n9844), .A2(n15459), .ZN(n9595) );
  AND2_X1 U12326 ( .A1(n12279), .A2(n12280), .ZN(n9596) );
  NAND2_X1 U12327 ( .A1(n12570), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10537) );
  INV_X2 U12328 ( .A(n10537), .ZN(n10423) );
  AND3_X1 U12329 ( .A1(n11216), .A2(n11212), .A3(n11213), .ZN(n9597) );
  OR3_X1 U12330 ( .A1(n17622), .A2(n9798), .A3(n9685), .ZN(n9598) );
  AND2_X1 U12331 ( .A1(n9992), .A2(n9660), .ZN(n9599) );
  AND2_X1 U12332 ( .A1(n9596), .A2(n12281), .ZN(n9600) );
  AND2_X1 U12333 ( .A1(n9594), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9601) );
  INV_X1 U12334 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17789) );
  INV_X1 U12335 ( .A(n10453), .ZN(n10538) );
  OR2_X1 U12336 ( .A1(n9590), .A2(n17504), .ZN(n9602) );
  OR2_X1 U12337 ( .A1(n11817), .A2(n9984), .ZN(n9603) );
  AND2_X1 U12338 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9604) );
  AND2_X1 U12339 ( .A1(n9751), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9605) );
  AND2_X1 U12340 ( .A1(n9964), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9606) );
  AND2_X1 U12341 ( .A1(n16297), .A2(n20859), .ZN(n9607) );
  NAND2_X1 U12342 ( .A1(n17734), .A2(n20916), .ZN(n9608) );
  AND2_X1 U12343 ( .A1(n9604), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9609) );
  AND2_X1 U12344 ( .A1(n11178), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9610) );
  AND2_X1 U12345 ( .A1(n9738), .A2(P3_EBX_REG_9__SCAN_IN), .ZN(n9611) );
  AND2_X1 U12346 ( .A1(n9610), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9612) );
  AND2_X1 U12347 ( .A1(n9899), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9613) );
  OR3_X1 U12348 ( .A1(n14932), .A2(n9995), .A3(n9994), .ZN(n9614) );
  OR2_X1 U12349 ( .A1(n18606), .A2(n9796), .ZN(n9615) );
  INV_X1 U12350 ( .A(n10241), .ZN(n10770) );
  OR2_X1 U12351 ( .A1(n12647), .A2(n16868), .ZN(n9618) );
  INV_X1 U12352 ( .A(n10341), .ZN(n11055) );
  NAND2_X1 U12353 ( .A1(n14995), .A2(n12440), .ZN(n9619) );
  AND2_X1 U12354 ( .A1(n12569), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10987) );
  INV_X1 U12355 ( .A(n12691), .ZN(n12661) );
  NOR2_X2 U12356 ( .A1(n12648), .A2(n12649), .ZN(n12691) );
  XNOR2_X1 U12357 ( .A(n14240), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9620) );
  AND2_X1 U12358 ( .A1(n14352), .A2(n11939), .ZN(n14353) );
  AND2_X1 U12359 ( .A1(n14399), .A2(n12040), .ZN(n14341) );
  OR2_X1 U12360 ( .A1(n9943), .A2(n17952), .ZN(n9621) );
  INV_X1 U12361 ( .A(n14393), .ZN(n9877) );
  OR2_X1 U12362 ( .A1(n12647), .A2(n16867), .ZN(n9622) );
  AND4_X1 U12363 ( .A1(n11270), .A2(n11269), .A3(n11268), .A4(n11267), .ZN(
        n9623) );
  OR2_X1 U12364 ( .A1(n15110), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9624) );
  NOR2_X1 U12365 ( .A1(n12752), .A2(n9819), .ZN(n9625) );
  NOR2_X1 U12366 ( .A1(n13987), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9626) );
  AND2_X1 U12367 ( .A1(n10308), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10453) );
  AND2_X1 U12368 ( .A1(n10031), .A2(n13708), .ZN(n9627) );
  AND2_X1 U12369 ( .A1(n10562), .A2(n10560), .ZN(n9628) );
  AND2_X1 U12370 ( .A1(n9628), .A2(n10793), .ZN(n9629) );
  AND2_X1 U12371 ( .A1(n14399), .A2(n9978), .ZN(n14342) );
  AND4_X1 U12372 ( .A1(n9823), .A2(n12738), .A3(n12739), .A4(n12736), .ZN(
        n9630) );
  AND2_X1 U12373 ( .A1(n15490), .A2(n10573), .ZN(n15469) );
  AND2_X1 U12374 ( .A1(n14352), .A2(n9981), .ZN(n14424) );
  AND4_X1 U12375 ( .A1(n11234), .A2(n11233), .A3(n11232), .A4(n11231), .ZN(
        n9631) );
  NAND2_X1 U12376 ( .A1(n11519), .A2(n11518), .ZN(n11600) );
  OAI211_X1 U12377 ( .C1(n17146), .C2(n20871), .A(n12866), .B(n12865), .ZN(
        n12880) );
  NAND2_X1 U12378 ( .A1(n18151), .A2(n17240), .ZN(n12888) );
  INV_X1 U12379 ( .A(n12888), .ZN(n9794) );
  AND2_X1 U12380 ( .A1(n14922), .A2(n12634), .ZN(n12633) );
  INV_X2 U12381 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10115) );
  OR2_X1 U12382 ( .A1(n14208), .A2(n10693), .ZN(n9632) );
  NOR2_X1 U12383 ( .A1(n9614), .A2(n13040), .ZN(n13039) );
  INV_X1 U12384 ( .A(n19023), .ZN(n10260) );
  AND4_X1 U12385 ( .A1(n12689), .A2(n12688), .A3(n12687), .A4(n12686), .ZN(
        n9633) );
  OR2_X1 U12386 ( .A1(n15965), .A2(n11614), .ZN(n9634) );
  OR3_X1 U12387 ( .A1(n17622), .A2(n9798), .A3(n16360), .ZN(n9635) );
  NOR2_X1 U12388 ( .A1(n12985), .A2(n17491), .ZN(n9636) );
  NOR2_X1 U12389 ( .A1(n16545), .A2(n16546), .ZN(n9637) );
  AND4_X1 U12390 ( .A1(n12610), .A2(n10641), .A3(n12618), .A4(n15205), .ZN(
        n9638) );
  BUF_X1 U12391 ( .A(n10183), .Z(n19213) );
  AND2_X1 U12392 ( .A1(n10090), .A2(n10089), .ZN(n9639) );
  AND2_X1 U12393 ( .A1(n10165), .A2(n10718), .ZN(n9640) );
  AND2_X2 U12394 ( .A1(n10074), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10316) );
  NOR2_X1 U12395 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12401) );
  AND2_X1 U12396 ( .A1(n9632), .A2(n14231), .ZN(n9641) );
  INV_X1 U12397 ( .A(n10371), .ZN(n12389) );
  INV_X1 U12398 ( .A(n12389), .ZN(n12321) );
  AND2_X1 U12399 ( .A1(n11574), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9642) );
  AOI22_X1 U12400 ( .A1(n13410), .A2(n11329), .B1(n11320), .B2(n14276), .ZN(
        n11335) );
  NOR2_X1 U12401 ( .A1(n15448), .A2(n9896), .ZN(n15201) );
  NAND2_X1 U12402 ( .A1(n14872), .A2(n14859), .ZN(n11113) );
  AND2_X1 U12403 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n9643) );
  AND3_X1 U12404 ( .A1(n10283), .A2(n10282), .A3(n10284), .ZN(n9644) );
  NAND2_X1 U12405 ( .A1(n9846), .A2(n10579), .ZN(n15458) );
  OR2_X1 U12406 ( .A1(n11632), .A2(n14736), .ZN(n9645) );
  OAI21_X1 U12407 ( .B1(n14970), .B2(n10020), .A(n10016), .ZN(n12521) );
  AND2_X1 U12408 ( .A1(n14232), .A2(n9849), .ZN(n9646) );
  OR2_X1 U12409 ( .A1(n9565), .A2(n17112), .ZN(n9647) );
  AND2_X1 U12410 ( .A1(n9638), .A2(n10646), .ZN(n9648) );
  INV_X1 U12411 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19819) );
  AND2_X1 U12412 ( .A1(n9627), .A2(n10030), .ZN(n9649) );
  AND2_X1 U12413 ( .A1(n9629), .A2(n13660), .ZN(n9650) );
  NAND2_X1 U12414 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12755), .ZN(
        n9651) );
  AND2_X1 U12415 ( .A1(n9853), .A2(n9852), .ZN(n9652) );
  NAND2_X1 U12416 ( .A1(n19196), .A2(n10900), .ZN(n10975) );
  INV_X2 U12417 ( .A(n10975), .ZN(n10944) );
  NOR2_X1 U12418 ( .A1(n13014), .A2(n15172), .ZN(n12995) );
  AND2_X1 U12419 ( .A1(n12994), .A2(n9964), .ZN(n9653) );
  AND2_X1 U12420 ( .A1(n10573), .A2(n15471), .ZN(n9654) );
  NAND2_X1 U12421 ( .A1(n13462), .A2(n12268), .ZN(n13516) );
  AND2_X1 U12422 ( .A1(n11692), .A2(n11272), .ZN(n13074) );
  AND2_X1 U12423 ( .A1(n10012), .A2(n15480), .ZN(n9655) );
  XNOR2_X1 U12424 ( .A(n10506), .B(n20886), .ZN(n15547) );
  AND2_X1 U12425 ( .A1(n15171), .A2(n15170), .ZN(n9656) );
  INV_X1 U12426 ( .A(n15153), .ZN(n9972) );
  AND2_X1 U12427 ( .A1(n17008), .A2(n9731), .ZN(n9657) );
  OR3_X1 U12428 ( .A1(n14800), .A2(n14079), .A3(n9882), .ZN(n9658) );
  INV_X1 U12429 ( .A(n13661), .ZN(n9874) );
  INV_X1 U12430 ( .A(n14105), .ZN(n9883) );
  AND3_X1 U12431 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n9659) );
  INV_X1 U12432 ( .A(n9582), .ZN(n12592) );
  NAND2_X1 U12433 ( .A1(n13964), .A2(n9591), .ZN(n10029) );
  INV_X1 U12434 ( .A(n15459), .ZN(n9845) );
  OR3_X1 U12435 ( .A1(n10640), .A2(n11175), .A3(n16267), .ZN(n15205) );
  INV_X1 U12436 ( .A(n9879), .ZN(n14427) );
  NOR2_X1 U12437 ( .A1(n14435), .A2(n14428), .ZN(n9879) );
  AND2_X1 U12438 ( .A1(n9991), .A2(n15555), .ZN(n9660) );
  AND2_X1 U12439 ( .A1(n14050), .A2(n14089), .ZN(n9661) );
  OR2_X1 U12440 ( .A1(n11082), .A2(n11081), .ZN(n12281) );
  OR2_X1 U12441 ( .A1(n15453), .A2(n10001), .ZN(n9662) );
  AND2_X1 U12442 ( .A1(n10597), .A2(n15392), .ZN(n15177) );
  INV_X1 U12443 ( .A(n15177), .ZN(n9767) );
  OR2_X1 U12444 ( .A1(n9882), .A2(n14445), .ZN(n9663) );
  OR2_X1 U12445 ( .A1(n9983), .A2(n9982), .ZN(n9664) );
  OR2_X1 U12446 ( .A1(n17528), .A2(n17545), .ZN(n9665) );
  NAND2_X1 U12447 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12998) );
  INV_X1 U12448 ( .A(n12998), .ZN(n9962) );
  AND2_X1 U12449 ( .A1(n12264), .A2(n10015), .ZN(n9666) );
  NAND2_X1 U12450 ( .A1(n17604), .A2(n17734), .ZN(n17525) );
  NAND2_X1 U12451 ( .A1(n13977), .A2(n16262), .ZN(n9667) );
  AND2_X1 U12452 ( .A1(n10025), .A2(n9619), .ZN(n9668) );
  INV_X1 U12453 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11345) );
  INV_X1 U12454 ( .A(n11697), .ZN(n12170) );
  NOR2_X1 U12455 ( .A1(n10925), .A2(n9993), .ZN(n9992) );
  INV_X1 U12456 ( .A(n17888), .ZN(n9944) );
  NAND2_X1 U12457 ( .A1(n13516), .A2(n9596), .ZN(n13837) );
  NAND2_X1 U12458 ( .A1(n16402), .A2(n16403), .ZN(n17734) );
  INV_X1 U12459 ( .A(n17734), .ZN(n17632) );
  NAND2_X1 U12460 ( .A1(n9989), .A2(n9992), .ZN(n13827) );
  NAND2_X1 U12461 ( .A1(n13516), .A2(n12279), .ZN(n13750) );
  NAND2_X1 U12462 ( .A1(n10748), .A2(n9827), .ZN(n11117) );
  AND2_X1 U12463 ( .A1(n17164), .A2(n9738), .ZN(n9669) );
  NAND2_X1 U12464 ( .A1(n14319), .A2(n14182), .ZN(n9670) );
  NOR2_X1 U12465 ( .A1(n13541), .A2(n13542), .ZN(n13543) );
  AND2_X1 U12466 ( .A1(n10006), .A2(n14214), .ZN(n9671) );
  AND2_X1 U12467 ( .A1(n9671), .A2(n10005), .ZN(n9672) );
  NAND2_X1 U12468 ( .A1(n11445), .A2(n11444), .ZN(n20142) );
  OR2_X1 U12469 ( .A1(n9670), .A2(n14391), .ZN(n9673) );
  XOR2_X1 U12470 ( .A(n19007), .B(n13948), .Z(n9674) );
  INV_X1 U12471 ( .A(n13632), .ZN(n10043) );
  INV_X1 U12472 ( .A(n13032), .ZN(n10051) );
  AND2_X1 U12473 ( .A1(n9672), .A2(n10004), .ZN(n9675) );
  AND2_X2 U12474 ( .A1(n13937), .A2(n12401), .ZN(n11071) );
  INV_X1 U12475 ( .A(n9881), .ZN(n13766) );
  NOR2_X1 U12476 ( .A1(n16135), .A2(n13730), .ZN(n9881) );
  INV_X1 U12477 ( .A(n14915), .ZN(n9997) );
  AND2_X1 U12478 ( .A1(n13049), .A2(n9609), .ZN(n9677) );
  AND2_X1 U12479 ( .A1(n10038), .A2(n10037), .ZN(n9678) );
  AND2_X1 U12480 ( .A1(n9609), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9679) );
  INV_X1 U12481 ( .A(n12518), .ZN(n10022) );
  INV_X1 U12482 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n9967) );
  AND3_X1 U12483 ( .A1(n13380), .A2(n11326), .A3(n11695), .ZN(n9680) );
  AND2_X1 U12484 ( .A1(n9612), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9681) );
  NOR2_X1 U12485 ( .A1(n20507), .A2(n20304), .ZN(n9682) );
  NOR2_X1 U12486 ( .A1(n20507), .A2(n20614), .ZN(n9683) );
  AND2_X1 U12487 ( .A1(n9756), .A2(n9755), .ZN(n9684) );
  INV_X1 U12488 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9753) );
  OR3_X1 U12489 ( .A1(n16360), .A2(n16362), .A3(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n9685) );
  NOR2_X1 U12490 ( .A1(n12334), .A2(n12333), .ZN(n9686) );
  AND2_X1 U12491 ( .A1(n14688), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9687) );
  OR2_X1 U12492 ( .A1(n12307), .A2(n12306), .ZN(n9688) );
  INV_X1 U12493 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9752) );
  AND2_X1 U12494 ( .A1(n17486), .A2(n9751), .ZN(n9689) );
  AND2_X1 U12495 ( .A1(n9959), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9690) );
  INV_X1 U12496 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9963) );
  INV_X1 U12497 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9757) );
  INV_X1 U12498 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n9843) );
  INV_X1 U12499 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9966) );
  INV_X1 U12500 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n9734) );
  INV_X1 U12501 ( .A(n17311), .ZN(n17346) );
  AOI22_X2 U12502 ( .A1(DATAI_23_), .A2(n20132), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n20131), .ZN(n20610) );
  AOI22_X2 U12503 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20131), .B1(DATAI_21_), 
        .B2(n20132), .ZN(n20598) );
  AOI22_X2 U12504 ( .A1(DATAI_19_), .A2(n20132), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20131), .ZN(n20590) );
  AOI22_X2 U12505 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19222), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19221), .ZN(n19637) );
  NOR2_X2 U12506 ( .A1(n13675), .A2(n19179), .ZN(n19221) );
  NOR3_X2 U12507 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18502), .A3(
        n18384), .ZN(n18354) );
  NOR3_X4 U12508 ( .A1(n13121), .A2(n19853), .A3(n19865), .ZN(n13199) );
  OR2_X1 U12509 ( .A1(n16310), .A2(n13021), .ZN(n13121) );
  NOR2_X4 U12510 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20771), .ZN(n20731) );
  NOR3_X2 U12511 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20615), .A3(
        n20614), .ZN(n20603) );
  AOI22_X2 U12512 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20131), .B1(DATAI_20_), 
        .B2(n20132), .ZN(n20594) );
  INV_X1 U12513 ( .A(n9698), .ZN(n9691) );
  NAND2_X1 U12514 ( .A1(n9698), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n9692) );
  NAND2_X1 U12515 ( .A1(n19294), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n9693) );
  OAI21_X1 U12516 ( .B1(n10399), .B2(n10272), .A(n9694), .ZN(n10273) );
  NAND2_X1 U12517 ( .A1(n19294), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n9695) );
  INV_X1 U12518 ( .A(n19294), .ZN(n9696) );
  NOR2_X1 U12519 ( .A1(n19294), .A2(n19860), .ZN(n9697) );
  NAND2_X1 U12520 ( .A1(n15547), .A2(n15548), .ZN(n9699) );
  NAND2_X1 U12521 ( .A1(n9699), .A2(n10507), .ZN(n15237) );
  NAND2_X1 U12522 ( .A1(n10556), .A2(n18981), .ZN(n10565) );
  NAND3_X1 U12523 ( .A1(n10480), .A2(n10479), .A3(n10931), .ZN(n11151) );
  NAND2_X2 U12524 ( .A1(n9700), .A2(n10384), .ZN(n10479) );
  NAND3_X1 U12525 ( .A1(n10369), .A2(n10370), .A3(n10368), .ZN(n9701) );
  AND2_X2 U12526 ( .A1(n9702), .A2(n10354), .ZN(n10480) );
  NAND4_X1 U12527 ( .A1(n9703), .A2(n10305), .A3(n10285), .A4(n9644), .ZN(
        n9702) );
  INV_X1 U12528 ( .A(n10304), .ZN(n9703) );
  INV_X1 U12529 ( .A(n9705), .ZN(n9918) );
  NAND2_X1 U12530 ( .A1(n10248), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9704) );
  NAND2_X1 U12531 ( .A1(n9705), .A2(n10244), .ZN(n10245) );
  AND2_X1 U12532 ( .A1(n9850), .A2(n9849), .ZN(n14233) );
  OAI21_X2 U12533 ( .B1(n9708), .B2(n9707), .A(n9706), .ZN(n9850) );
  NAND3_X1 U12534 ( .A1(n10199), .A2(n10184), .A3(n19206), .ZN(n10754) );
  NAND2_X1 U12535 ( .A1(n9711), .A2(n9584), .ZN(n9710) );
  OR2_X2 U12536 ( .A1(n15458), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9772) );
  INV_X2 U12537 ( .A(n11695), .ZN(n11710) );
  NAND2_X2 U12538 ( .A1(n9597), .A2(n9589), .ZN(n11695) );
  AND2_X2 U12539 ( .A1(n11195), .A2(n9715), .ZN(n11251) );
  AND2_X2 U12540 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9715) );
  NOR2_X1 U12541 ( .A1(n9715), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13336) );
  AND2_X1 U12542 ( .A1(n13346), .A2(n9715), .ZN(n11274) );
  NOR2_X1 U12543 ( .A1(n14830), .A2(n9715), .ZN(n14833) );
  AND2_X2 U12544 ( .A1(n11190), .A2(n9715), .ZN(n11419) );
  AND2_X4 U12545 ( .A1(n13345), .A2(n9715), .ZN(n12156) );
  XNOR2_X1 U12546 ( .A(n9715), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14848) );
  MUX2_X1 U12547 ( .A(n13345), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n9715), .Z(n13347) );
  NAND2_X1 U12548 ( .A1(n13773), .A2(n13774), .ZN(n11585) );
  NAND2_X1 U12549 ( .A1(n9718), .A2(n9716), .ZN(n13773) );
  AOI21_X1 U12550 ( .B1(n13689), .B2(n9717), .A(n9642), .ZN(n9716) );
  INV_X1 U12551 ( .A(n11561), .ZN(n9717) );
  NAND3_X1 U12552 ( .A1(n13610), .A2(n13609), .A3(n13689), .ZN(n9718) );
  XNOR2_X1 U12553 ( .A(n11574), .B(n11573), .ZN(n13689) );
  NAND3_X1 U12554 ( .A1(n11340), .A2(n13213), .A3(n13384), .ZN(n9727) );
  INV_X1 U12555 ( .A(n9727), .ZN(n9726) );
  NAND2_X1 U12556 ( .A1(n9727), .A2(n13330), .ZN(n13331) );
  OR2_X2 U12557 ( .A1(n16022), .A2(n16021), .ZN(n16024) );
  INV_X1 U12558 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9730) );
  AND4_X2 U12559 ( .A1(n11184), .A2(n9730), .A3(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A4(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11266) );
  INV_X2 U12560 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18769) );
  INV_X1 U12561 ( .A(n9737), .ZN(n17055) );
  NAND3_X1 U12562 ( .A1(n12855), .A2(n9647), .A3(n9745), .ZN(n9744) );
  AOI21_X1 U12563 ( .B1(n9758), .B2(n10769), .A(n10768), .ZN(n13522) );
  XNOR2_X2 U12564 ( .A(n9758), .B(n10769), .ZN(n10277) );
  NAND2_X1 U12565 ( .A1(n10247), .A2(n10246), .ZN(n9758) );
  NAND3_X1 U12566 ( .A1(n10481), .A2(n11175), .A3(n11148), .ZN(n9920) );
  NAND2_X2 U12567 ( .A1(n10480), .A2(n10479), .ZN(n11148) );
  NAND2_X2 U12568 ( .A1(n9760), .A2(n9759), .ZN(n10481) );
  NOR2_X1 U12569 ( .A1(n9761), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15589) );
  NAND2_X1 U12570 ( .A1(n12401), .A2(n9761), .ZN(n12367) );
  NAND2_X1 U12571 ( .A1(n10091), .A2(n9639), .ZN(n9762) );
  NAND2_X1 U12572 ( .A1(n10086), .A2(n10065), .ZN(n9763) );
  INV_X2 U12573 ( .A(n19206), .ZN(n10883) );
  NAND2_X2 U12574 ( .A1(n9763), .A2(n9762), .ZN(n19206) );
  NAND2_X1 U12575 ( .A1(n10182), .A2(n10883), .ZN(n10749) );
  NAND2_X2 U12576 ( .A1(n13229), .A2(n10469), .ZN(n10182) );
  NAND2_X2 U12577 ( .A1(n9765), .A2(n9764), .ZN(n10469) );
  NAND3_X1 U12578 ( .A1(n12813), .A2(n12814), .A3(n9783), .ZN(n9782) );
  NAND3_X1 U12579 ( .A1(n12815), .A2(n9786), .A3(n9785), .ZN(n9784) );
  NOR2_X1 U12580 ( .A1(n17622), .A2(n16360), .ZN(n17535) );
  INV_X1 U12581 ( .A(n16361), .ZN(n9798) );
  NAND2_X1 U12582 ( .A1(n16368), .A2(n17722), .ZN(n9800) );
  NAND3_X1 U12583 ( .A1(n9802), .A2(n17520), .A3(n9801), .ZN(n17509) );
  AND2_X2 U12584 ( .A1(n9803), .A2(n17525), .ZN(n17595) );
  OR2_X2 U12585 ( .A1(n15742), .A2(n16377), .ZN(n9805) );
  NAND2_X1 U12586 ( .A1(n9942), .A2(n9943), .ZN(n12764) );
  INV_X1 U12587 ( .A(n17773), .ZN(n9819) );
  INV_X1 U12588 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n9820) );
  INV_X2 U12589 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10458) );
  NAND4_X1 U12590 ( .A1(n9828), .A2(n9593), .A3(n10194), .A4(n19852), .ZN(
        n9827) );
  NOR2_X1 U12591 ( .A1(n10286), .A2(n15568), .ZN(n9830) );
  NAND3_X1 U12592 ( .A1(n10498), .A2(n13879), .A3(n9674), .ZN(n9831) );
  NAND4_X1 U12593 ( .A1(n9838), .A2(n9836), .A3(n9835), .A4(n9832), .ZN(n10236) );
  NAND2_X1 U12594 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n9834) );
  NAND2_X1 U12595 ( .A1(n9578), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9835) );
  NAND2_X1 U12596 ( .A1(n9850), .A2(n9646), .ZN(n9848) );
  INV_X1 U12597 ( .A(n9850), .ZN(n15096) );
  INV_X1 U12598 ( .A(n15095), .ZN(n9849) );
  NAND2_X1 U12599 ( .A1(n15330), .A2(n9854), .ZN(n9851) );
  NAND2_X1 U12600 ( .A1(n9851), .A2(n9652), .ZN(n14209) );
  OR2_X2 U12601 ( .A1(n9867), .A2(n9865), .ZN(n9864) );
  NAND3_X1 U12602 ( .A1(n9873), .A2(n9871), .A3(n9870), .ZN(n13499) );
  NOR2_X1 U12603 ( .A1(n14392), .A2(n14391), .ZN(n14393) );
  INV_X1 U12604 ( .A(n14331), .ZN(n9876) );
  NOR2_X2 U12605 ( .A1(n14420), .A2(n14410), .ZN(n14412) );
  INV_X1 U12606 ( .A(n9884), .ZN(n14447) );
  NAND2_X1 U12607 ( .A1(n10264), .A2(n9885), .ZN(n10263) );
  NOR2_X2 U12608 ( .A1(n10259), .A2(n10265), .ZN(n19023) );
  NAND2_X4 U12609 ( .A1(n9886), .A2(n11177), .ZN(n12640) );
  NAND2_X1 U12610 ( .A1(n15501), .A2(n15500), .ZN(n9886) );
  NAND2_X1 U12611 ( .A1(n9888), .A2(n9887), .ZN(n16253) );
  INV_X1 U12612 ( .A(n13887), .ZN(n9887) );
  NAND3_X1 U12613 ( .A1(n15408), .A2(n15409), .A3(n9889), .ZN(P2_U3029) );
  NAND3_X2 U12614 ( .A1(n11156), .A2(n9894), .A3(n11155), .ZN(n15553) );
  NAND2_X1 U12615 ( .A1(n10033), .A2(n15553), .ZN(n9895) );
  OAI211_X2 U12616 ( .C1(n15553), .C2(n11162), .A(n10071), .B(n9895), .ZN(
        n15234) );
  INV_X1 U12617 ( .A(n15448), .ZN(n9898) );
  AND2_X2 U12618 ( .A1(n10564), .A2(n10562), .ZN(n10575) );
  NAND2_X1 U12619 ( .A1(n10649), .A2(n10648), .ZN(n10654) );
  NAND2_X1 U12620 ( .A1(n10623), .A2(n9908), .ZN(n10651) );
  NAND2_X2 U12621 ( .A1(n10623), .A2(n10622), .ZN(n10625) );
  INV_X1 U12622 ( .A(n9914), .ZN(n12749) );
  NOR2_X1 U12623 ( .A1(n17798), .A2(n18093), .ZN(n17797) );
  OR2_X2 U12624 ( .A1(n17804), .A2(n12746), .ZN(n9914) );
  NOR2_X1 U12625 ( .A1(n17806), .A2(n17805), .ZN(n17804) );
  INV_X1 U12626 ( .A(n10183), .ZN(n9915) );
  NAND3_X1 U12627 ( .A1(n16397), .A2(n16396), .A3(n9919), .ZN(P3_U2831) );
  NAND2_X1 U12628 ( .A1(n9920), .A2(n13824), .ZN(n10495) );
  INV_X1 U12629 ( .A(n9921), .ZN(n17755) );
  XNOR2_X2 U12630 ( .A(n12757), .B(n12756), .ZN(n17751) );
  AND2_X2 U12631 ( .A1(n9921), .A2(n9651), .ZN(n12757) );
  OR2_X1 U12632 ( .A1(n15207), .A2(n9925), .ZN(n9924) );
  AND2_X2 U12633 ( .A1(n9924), .A2(n9922), .ZN(n15162) );
  OAI22_X1 U12634 ( .A1(n9565), .A2(n18160), .B1(n12672), .B2(n17113), .ZN(
        n9939) );
  INV_X1 U12635 ( .A(n17732), .ZN(n9941) );
  AND2_X1 U12636 ( .A1(n12775), .A2(n17484), .ZN(n16400) );
  NAND2_X2 U12637 ( .A1(n17492), .A2(n12774), .ZN(n12775) );
  OR2_X2 U12638 ( .A1(n16867), .A2(n12649), .ZN(n17088) );
  INV_X2 U12639 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18777) );
  NAND2_X1 U12640 ( .A1(n13610), .A2(n13609), .ZN(n9948) );
  AND2_X2 U12641 ( .A1(n11202), .A2(n13346), .ZN(n11478) );
  AND2_X2 U12642 ( .A1(n11185), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11202) );
  NAND4_X1 U12643 ( .A1(n9949), .A2(n11335), .A3(n13085), .A4(n11343), .ZN(
        n11391) );
  NAND2_X1 U12644 ( .A1(n14598), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11632) );
  NAND2_X1 U12645 ( .A1(n14627), .A2(n9960), .ZN(n11628) );
  NAND4_X1 U12646 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n9961), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13001) );
  AOI21_X1 U12647 ( .B1(n15747), .B2(n9972), .A(n13016), .ZN(n9971) );
  NAND2_X1 U12648 ( .A1(n9969), .A2(n9968), .ZN(n14910) );
  NAND2_X1 U12649 ( .A1(n15747), .A2(n9970), .ZN(n9969) );
  NAND2_X1 U12650 ( .A1(n13049), .A2(n9679), .ZN(n12992) );
  NAND2_X1 U12651 ( .A1(n12995), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13015) );
  AND3_X2 U12652 ( .A1(n11692), .A2(n11272), .A3(n13242), .ZN(n13212) );
  NAND3_X1 U12653 ( .A1(n11319), .A2(n10073), .A3(n11321), .ZN(n13332) );
  NOR2_X2 U12654 ( .A1(n13917), .A2(n9664), .ZN(n14040) );
  NAND2_X1 U12655 ( .A1(n14141), .A2(n9985), .ZN(n9987) );
  INV_X1 U12656 ( .A(n9987), .ZN(n14300) );
  INV_X1 U12657 ( .A(n13281), .ZN(n9989) );
  NAND2_X1 U12658 ( .A1(n9989), .A2(n9599), .ZN(n15554) );
  NAND2_X1 U12659 ( .A1(n12265), .A2(n12264), .ZN(n10014) );
  NAND2_X1 U12660 ( .A1(n12265), .A2(n9666), .ZN(n12267) );
  NAND2_X1 U12661 ( .A1(n12494), .A2(n10022), .ZN(n10016) );
  NAND2_X1 U12662 ( .A1(n10019), .A2(n10023), .ZN(n10018) );
  OR2_X2 U12663 ( .A1(n14970), .A2(n14969), .ZN(n10023) );
  AND2_X2 U12664 ( .A1(n10018), .A2(n10017), .ZN(n14961) );
  NOR2_X1 U12665 ( .A1(n12494), .A2(n10022), .ZN(n10019) );
  INV_X1 U12666 ( .A(n10023), .ZN(n14968) );
  INV_X1 U12667 ( .A(n10025), .ZN(n14986) );
  AND2_X2 U12668 ( .A1(n13516), .A2(n9600), .ZN(n13995) );
  NOR2_X2 U12669 ( .A1(n13962), .A2(n10026), .ZN(n14019) );
  INV_X1 U12670 ( .A(n10029), .ZN(n14018) );
  AND3_X2 U12672 ( .A1(n10130), .A2(n10129), .A3(n9640), .ZN(n13168) );
  INV_X1 U12673 ( .A(n15549), .ZN(n10034) );
  NAND2_X1 U12674 ( .A1(n13543), .A2(n10040), .ZN(n13642) );
  OAI21_X1 U12675 ( .B1(n15276), .B2(n16274), .A(n10044), .ZN(P2_U3018) );
  OR2_X1 U12676 ( .A1(n15121), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10047) );
  NAND2_X2 U12677 ( .A1(n12640), .A2(n9681), .ZN(n14219) );
  NAND2_X1 U12678 ( .A1(n16395), .A2(n17722), .ZN(n12955) );
  NAND2_X1 U12679 ( .A1(n15091), .A2(n16270), .ZN(n11182) );
  NOR2_X2 U12680 ( .A1(n15967), .A2(n14568), .ZN(n14590) );
  NAND2_X1 U12681 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20536), .ZN(
        n11650) );
  OR2_X1 U12682 ( .A1(n11388), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11389) );
  NOR2_X1 U12683 ( .A1(n13579), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11197) );
  OR2_X1 U12684 ( .A1(n13461), .A2(n13460), .ZN(n13463) );
  NAND2_X1 U12685 ( .A1(n11742), .A2(n11741), .ZN(n13647) );
  INV_X1 U12686 ( .A(n13622), .ZN(n11741) );
  INV_X1 U12687 ( .A(n13525), .ZN(n11742) );
  NAND2_X1 U12688 ( .A1(n12416), .A2(n10200), .ZN(n10201) );
  NAND2_X1 U12689 ( .A1(n12416), .A2(n16322), .ZN(n10700) );
  NAND3_X1 U12690 ( .A1(n10211), .A2(n12416), .A3(n10182), .ZN(n10891) );
  INV_X1 U12691 ( .A(n11151), .ZN(n10509) );
  NAND2_X1 U12692 ( .A1(n14040), .A2(n14098), .ZN(n14099) );
  OR2_X2 U12693 ( .A1(n11327), .A2(n13068), .ZN(n13091) );
  AND3_X1 U12694 ( .A1(n10357), .A2(n10356), .A3(n10355), .ZN(n10370) );
  NOR2_X1 U12695 ( .A1(n13016), .A2(n14887), .ZN(n16161) );
  NAND2_X2 U12696 ( .A1(n13888), .A2(n11147), .ZN(n11152) );
  CLKBUF_X1 U12697 ( .A(n14441), .Z(n14442) );
  NOR2_X1 U12698 ( .A1(n14209), .A2(n10675), .ZN(n15107) );
  OR2_X1 U12699 ( .A1(n10866), .A2(n10865), .ZN(n10867) );
  NAND2_X1 U12700 ( .A1(n14281), .A2(n12227), .ZN(n12245) );
  AND2_X1 U12701 ( .A1(n19196), .A2(n19223), .ZN(n19662) );
  AND2_X1 U12702 ( .A1(n16314), .A2(n19196), .ZN(n13269) );
  NAND3_X1 U12703 ( .A1(n9915), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n19196), 
        .ZN(n12277) );
  NAND2_X1 U12704 ( .A1(n19196), .A2(n19852), .ZN(n10212) );
  NAND2_X1 U12705 ( .A1(n14961), .A2(n14960), .ZN(n14959) );
  OR2_X1 U12706 ( .A1(n12246), .A2(n13911), .ZN(n10279) );
  NAND2_X1 U12707 ( .A1(n10121), .A2(n10115), .ZN(n10128) );
  NAND2_X2 U12708 ( .A1(n10185), .A2(n10754), .ZN(n10877) );
  NAND2_X1 U12709 ( .A1(n11390), .A2(n11389), .ZN(n11393) );
  AOI211_X2 U12710 ( .C1(n16007), .C2(n14578), .A(n14577), .B(n14576), .ZN(
        n14579) );
  BUF_X1 U12711 ( .A(n10237), .Z(n10248) );
  AOI21_X1 U12712 ( .B1(n10308), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n10115), .ZN(n10076) );
  AOI22_X1 U12713 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10123) );
  NAND2_X1 U12714 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10075) );
  OAI21_X1 U12715 ( .B1(n9915), .B2(n10883), .A(n10197), .ZN(n10166) );
  NAND2_X1 U12716 ( .A1(n10883), .A2(n9583), .ZN(n10197) );
  XNOR2_X2 U12717 ( .A(n14241), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14267) );
  NAND2_X1 U12718 ( .A1(n10277), .A2(n12246), .ZN(n10281) );
  OR2_X2 U12719 ( .A1(n10277), .A2(n19023), .ZN(n10286) );
  AND2_X1 U12720 ( .A1(n17240), .A2(n17191), .ZN(n17188) );
  AND3_X1 U12721 ( .A1(n14254), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14253), .ZN(n10054) );
  OR2_X1 U12722 ( .A1(n14458), .A2(n12242), .ZN(n10055) );
  INV_X1 U12723 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11357) );
  NOR2_X1 U12724 ( .A1(n12743), .A2(n12742), .ZN(n10056) );
  INV_X1 U12725 ( .A(n14046), .ZN(n11817) );
  AND2_X1 U12726 ( .A1(n10227), .A2(n10226), .ZN(n10058) );
  AND2_X1 U12727 ( .A1(n15568), .A2(n10260), .ZN(n10059) );
  AND2_X1 U12728 ( .A1(n10184), .A2(n10874), .ZN(n10060) );
  AND2_X1 U12729 ( .A1(n12492), .A2(n12516), .ZN(n10061) );
  AND3_X1 U12730 ( .A1(n12608), .A2(n12607), .A3(n12606), .ZN(n10062) );
  INV_X1 U12731 ( .A(n13836), .ZN(n12280) );
  INV_X1 U12732 ( .A(n18157), .ZN(n18804) );
  INV_X2 U12733 ( .A(n9622), .ZN(n15684) );
  AND3_X1 U12734 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .A3(P3_EAX_REG_14__SCAN_IN), .ZN(n10063) );
  NOR2_X1 U12735 ( .A1(n20507), .A2(n20473), .ZN(n10064) );
  AND2_X1 U12736 ( .A1(n10085), .A2(n10084), .ZN(n10065) );
  OR2_X1 U12737 ( .A1(n12621), .A2(n15177), .ZN(n10066) );
  INV_X1 U12738 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11806) );
  NOR2_X1 U12739 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20481) );
  INV_X1 U12740 ( .A(n20481), .ZN(n20620) );
  OR2_X1 U12741 ( .A1(n9566), .A2(n10240), .ZN(n10068) );
  AND2_X1 U12742 ( .A1(n10242), .A2(n10068), .ZN(n10069) );
  OR2_X1 U12743 ( .A1(n15360), .A2(n16245), .ZN(n10070) );
  OR2_X1 U12744 ( .A1(n15549), .A2(n11167), .ZN(n10071) );
  INV_X1 U12745 ( .A(n11274), .ZN(n13337) );
  AND2_X2 U12746 ( .A1(n11195), .A2(n14830), .ZN(n11420) );
  AND2_X1 U12747 ( .A1(n11318), .A2(n11317), .ZN(n10073) );
  AND2_X1 U12748 ( .A1(n20102), .A2(n20122), .ZN(n11651) );
  INV_X1 U12749 ( .A(n10406), .ZN(n10407) );
  NOR2_X1 U12750 ( .A1(n10405), .A2(n10407), .ZN(n10408) );
  NAND2_X1 U12751 ( .A1(n10414), .A2(n10413), .ZN(n10415) );
  AOI22_X1 U12752 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19323), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10357) );
  NOR3_X1 U12753 ( .A1(n11688), .A2(n13413), .A3(n11659), .ZN(n11669) );
  OR2_X1 U12754 ( .A1(n11668), .A2(n11477), .ZN(n11490) );
  OR2_X1 U12755 ( .A1(n11668), .A2(n11491), .ZN(n11503) );
  INV_X1 U12756 ( .A(n10225), .ZN(n10226) );
  OR2_X1 U12757 ( .A1(n19188), .A2(n13601), .ZN(n10516) );
  NAND2_X1 U12758 ( .A1(n10421), .A2(n10420), .ZN(n10439) );
  INV_X1 U12759 ( .A(n11674), .ZN(n11645) );
  INV_X1 U12760 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11184) );
  AND2_X1 U12761 ( .A1(n11490), .A2(n11489), .ZN(n11562) );
  INV_X1 U12762 ( .A(n12076), .ZN(n12077) );
  OR2_X1 U12763 ( .A1(n11501), .A2(n11500), .ZN(n11589) );
  NAND2_X1 U12764 ( .A1(n11541), .A2(n11452), .ZN(n11554) );
  NAND2_X1 U12765 ( .A1(n9569), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10243) );
  AND4_X1 U12766 ( .A1(n10532), .A2(n10531), .A3(n10530), .A4(n10529), .ZN(
        n10533) );
  INV_X1 U12767 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10083) );
  NAND2_X1 U12768 ( .A1(n12575), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10079) );
  AOI22_X1 U12769 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10119) );
  NOR2_X1 U12770 ( .A1(n12788), .A2(n12787), .ZN(n12784) );
  NOR2_X1 U12771 ( .A1(n11645), .A2(n11673), .ZN(n11646) );
  AND2_X1 U12772 ( .A1(n12077), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12078) );
  INV_X1 U12773 ( .A(n14354), .ZN(n11939) );
  INV_X1 U12774 ( .A(n13722), .ZN(n11767) );
  INV_X1 U12775 ( .A(n11587), .ZN(n11519) );
  OR2_X1 U12776 ( .A1(n11392), .A2(n11387), .ZN(n11442) );
  OR2_X1 U12777 ( .A1(n11403), .A2(n11402), .ZN(n11608) );
  INV_X1 U12778 ( .A(n12470), .ZN(n12471) );
  INV_X1 U12779 ( .A(n15127), .ZN(n10673) );
  AND4_X1 U12780 ( .A1(n10452), .A2(n10451), .A3(n10450), .A4(n10449), .ZN(
        n10455) );
  AOI21_X1 U12781 ( .B1(n17105), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n12737), .ZN(n12738) );
  INV_X1 U12782 ( .A(n17826), .ZN(n12917) );
  AOI21_X1 U12783 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20429), .A(
        n11646), .ZN(n11670) );
  AND4_X1 U12784 ( .A1(n11310), .A2(n11309), .A3(n11308), .A4(n11307), .ZN(
        n11311) );
  NAND2_X1 U12785 ( .A1(n12078), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12119) );
  NOR2_X1 U12786 ( .A1(n20134), .A2(n20679), .ZN(n11713) );
  AND2_X1 U12787 ( .A1(n11617), .A2(n14656), .ZN(n14633) );
  INV_X1 U12788 ( .A(n11380), .ZN(n11545) );
  INV_X1 U12789 ( .A(n11531), .ZN(n13216) );
  OR2_X1 U12790 ( .A1(n11473), .A2(n11472), .ZN(n11565) );
  NAND2_X1 U12791 ( .A1(n10477), .A2(n10476), .ZN(n10483) );
  AND2_X1 U12792 ( .A1(n12493), .A2(n10061), .ZN(n12494) );
  INV_X1 U12793 ( .A(n14264), .ZN(n14256) );
  AND2_X1 U12794 ( .A1(n11086), .A2(n11085), .ZN(n15411) );
  OR2_X1 U12795 ( .A1(n18932), .A2(n11175), .ZN(n10615) );
  NAND2_X1 U12796 ( .A1(n10152), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10153) );
  NOR2_X1 U12797 ( .A1(n20806), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12643) );
  OAI21_X1 U12798 ( .B1(n12885), .B2(n15727), .A(n18163), .ZN(n12881) );
  AND2_X1 U12799 ( .A1(n11683), .A2(n11651), .ZN(n11689) );
  NAND2_X1 U12800 ( .A1(n19898), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13796) );
  INV_X1 U12801 ( .A(n13804), .ZN(n13801) );
  INV_X1 U12802 ( .A(n11743), .ZN(n11752) );
  AND4_X1 U12803 ( .A1(n11290), .A2(n11289), .A3(n11288), .A4(n11287), .ZN(
        n11291) );
  INV_X1 U12804 ( .A(n14834), .ZN(n15760) );
  XNOR2_X1 U12805 ( .A(n12211), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13807) );
  OR2_X1 U12806 ( .A1(n14585), .A2(n12170), .ZN(n12123) );
  NOR2_X1 U12807 ( .A1(n11870), .A2(n14069), .ZN(n11875) );
  AND2_X1 U12808 ( .A1(n20679), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12200) );
  INV_X1 U12809 ( .A(n11651), .ZN(n11678) );
  INV_X2 U12810 ( .A(n10770), .ZN(n10856) );
  AND2_X1 U12811 ( .A1(n12278), .A2(n13518), .ZN(n12279) );
  INV_X1 U12812 ( .A(n14249), .ZN(n14250) );
  NOR2_X1 U12813 ( .A1(n10551), .A2(n10550), .ZN(n10938) );
  INV_X1 U12814 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12991) );
  AOI211_X1 U12815 ( .C1(n14257), .C2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n10054), .B(n14256), .ZN(n14258) );
  XOR2_X1 U12816 ( .A(n10690), .B(n10691), .Z(n14861) );
  OR2_X1 U12817 ( .A1(n10615), .A2(n15432), .ZN(n15443) );
  NAND2_X1 U12818 ( .A1(n10497), .A2(n10496), .ZN(n13879) );
  NAND2_X1 U12819 ( .A1(n12248), .A2(n10900), .ZN(n12263) );
  INV_X1 U12820 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n16335) );
  AOI22_X1 U12821 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n18635), .B2(n18783), .ZN(
        n12905) );
  OAI21_X1 U12822 ( .B1(n10053), .B2(n18160), .A(n12804), .ZN(n12805) );
  NOR2_X1 U12823 ( .A1(n12942), .A2(n18054), .ZN(n12943) );
  NOR2_X1 U12824 ( .A1(n17612), .A2(n17596), .ZN(n17552) );
  NAND2_X1 U12825 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18620) );
  AOI21_X1 U12826 ( .B1(n11688), .B2(n12223), .A(n11687), .ZN(n11691) );
  INV_X1 U12827 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14069) );
  AND2_X1 U12828 ( .A1(n13807), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13792) );
  OR2_X1 U12829 ( .A1(n13796), .A2(n20084), .ZN(n13804) );
  AND2_X1 U12830 ( .A1(n14578), .A2(n12142), .ZN(n12143) );
  OR2_X1 U12831 ( .A1(n13392), .A2(n20079), .ZN(n14458) );
  NOR2_X1 U12832 ( .A1(n13412), .A2(n13411), .ZN(n13414) );
  INV_X1 U12833 ( .A(n12202), .ZN(n12203) );
  OR2_X1 U12834 ( .A1(n11907), .A2(n15891), .ZN(n11923) );
  INV_X1 U12835 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15923) );
  NAND2_X1 U12836 ( .A1(n11782), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11807) );
  NAND2_X1 U12837 ( .A1(n16146), .A2(n20676), .ZN(n12212) );
  INV_X1 U12838 ( .A(n20067), .ZN(n16069) );
  NOR2_X1 U12839 ( .A1(n14805), .A2(n14690), .ZN(n14695) );
  NAND2_X1 U12840 ( .A1(n11446), .A2(n20142), .ZN(n13870) );
  INV_X1 U12841 ( .A(n9587), .ZN(n20082) );
  INV_X1 U12842 ( .A(n20171), .ZN(n20083) );
  INV_X1 U12843 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20615) );
  NAND2_X1 U12844 ( .A1(n10760), .A2(n10717), .ZN(n16314) );
  CLKBUF_X1 U12845 ( .A(n14019), .Z(n15006) );
  AND3_X1 U12846 ( .A1(n10934), .A2(n10933), .A3(n10932), .ZN(n13949) );
  AND2_X1 U12847 ( .A1(n15538), .A2(n11129), .ZN(n15487) );
  AND2_X1 U12848 ( .A1(n11127), .A2(n15559), .ZN(n15538) );
  NAND2_X1 U12849 ( .A1(n19235), .A2(n19830), .ZN(n19383) );
  INV_X1 U12850 ( .A(n19800), .ZN(n19290) );
  OR2_X1 U12851 ( .A1(n19810), .A2(n19822), .ZN(n19353) );
  INV_X1 U12852 ( .A(n19205), .ZN(n19223) );
  NOR2_X1 U12853 ( .A1(n18820), .A2(n14121), .ZN(n18609) );
  NOR2_X1 U12854 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16792), .ZN(n16761) );
  AOI211_X1 U12855 ( .C1(n17131), .C2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n12874), .B(n12873), .ZN(n12875) );
  INV_X1 U12856 ( .A(n17315), .ZN(n17194) );
  INV_X1 U12857 ( .A(n17599), .ZN(n17622) );
  NAND2_X1 U12858 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17633), .ZN(
        n18007) );
  NAND2_X1 U12859 ( .A1(n17664), .A2(n17827), .ZN(n17564) );
  AOI221_X1 U12860 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C1(n15798), .C2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(n12776), .ZN(n12780) );
  NOR2_X1 U12861 ( .A1(n17647), .A2(n17641), .ZN(n17958) );
  NOR2_X1 U12862 ( .A1(n17320), .A2(n12733), .ZN(n16402) );
  NAND2_X1 U12863 ( .A1(n12941), .A2(n17761), .ZN(n17745) );
  NOR2_X1 U12864 ( .A1(n12969), .A2(n12899), .ZN(n18630) );
  AOI21_X1 U12865 ( .B1(n18138), .B2(n18808), .A(n18784), .ZN(n18150) );
  OR2_X1 U12866 ( .A1(n11691), .A2(n11690), .ZN(n13364) );
  AND2_X1 U12867 ( .A1(n19898), .A2(n13792), .ZN(n19936) );
  INV_X1 U12868 ( .A(n19944), .ZN(n19968) );
  INV_X1 U12869 ( .A(n14455), .ZN(n19990) );
  INV_X1 U12870 ( .A(n19994), .ZN(n14438) );
  INV_X1 U12871 ( .A(n15985), .ZN(n15876) );
  OR2_X1 U12872 ( .A1(n15784), .A2(n20676), .ZN(n19873) );
  NAND2_X1 U12873 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n12037), .ZN(
        n12076) );
  NAND2_X1 U12874 ( .A1(n11989), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12036) );
  INV_X1 U12875 ( .A(n14442), .ZN(n14452) );
  INV_X1 U12876 ( .A(n16039), .ZN(n20058) );
  OR2_X1 U12877 ( .A1(n12212), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16041) );
  AND2_X1 U12878 ( .A1(n14700), .A2(n14696), .ZN(n14731) );
  OR2_X1 U12879 ( .A1(n15808), .A2(n14692), .ZN(n14805) );
  INV_X1 U12880 ( .A(n14810), .ZN(n14690) );
  AND2_X1 U12881 ( .A1(n13107), .A2(n14834), .ZN(n15808) );
  INV_X1 U12882 ( .A(n16070), .ZN(n20071) );
  AND2_X1 U12883 ( .A1(n13107), .A2(n13106), .ZN(n20067) );
  INV_X1 U12884 ( .A(n20088), .ZN(n20257) );
  NOR2_X1 U12885 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16146) );
  OR2_X1 U12886 ( .A1(n20172), .A2(n20083), .ZN(n20248) );
  INV_X1 U12887 ( .A(n20217), .ZN(n20245) );
  INV_X1 U12888 ( .A(n20252), .ZN(n20274) );
  INV_X1 U12889 ( .A(n20334), .ZN(n20299) );
  OR2_X1 U12890 ( .A1(n20172), .A2(n20171), .ZN(n20403) );
  NAND2_X1 U12891 ( .A1(n9587), .A2(n14822), .ZN(n20348) );
  INV_X1 U12892 ( .A(n20364), .ZN(n20393) );
  INV_X1 U12893 ( .A(n20472), .ZN(n20427) );
  INV_X1 U12894 ( .A(n20499), .ZN(n20502) );
  AND2_X1 U12895 ( .A1(n20172), .A2(n20083), .ZN(n20482) );
  INV_X1 U12896 ( .A(n20403), .ZN(n20535) );
  INV_X1 U12897 ( .A(n20568), .ZN(n20606) );
  INV_X1 U12898 ( .A(n20425), .ZN(n20618) );
  AND2_X1 U12899 ( .A1(n9587), .A2(n14825), .ZN(n20564) );
  AND2_X1 U12900 ( .A1(n15779), .A2(n15778), .ZN(n15786) );
  INV_X1 U12901 ( .A(n19008), .ZN(n19030) );
  AND2_X1 U12902 ( .A1(n13208), .A2(n13038), .ZN(n19027) );
  INV_X1 U12903 ( .A(n18991), .ZN(n19041) );
  INV_X1 U12904 ( .A(n12281), .ZN(n13956) );
  OR2_X1 U12905 ( .A1(n13653), .A2(n13650), .ZN(n13714) );
  AND2_X1 U12906 ( .A1(n13255), .A2(n13675), .ZN(n19051) );
  AND2_X1 U12907 ( .A1(n19083), .A2(n12592), .ZN(n19111) );
  INV_X1 U12908 ( .A(n13270), .ZN(n13208) );
  AND2_X1 U12909 ( .A1(n13545), .A2(n13544), .ZN(n19001) );
  INV_X1 U12910 ( .A(n16243), .ZN(n19167) );
  AND2_X1 U12911 ( .A1(n13686), .A2(n13685), .ZN(n16219) );
  AND2_X1 U12912 ( .A1(n11181), .A2(n19844), .ZN(n16270) );
  AND2_X1 U12913 ( .A1(n12637), .A2(n18828), .ZN(n19656) );
  INV_X1 U12914 ( .A(n19714), .ZN(n13167) );
  OAI21_X1 U12915 ( .B1(n19193), .B2(n19192), .A(n19191), .ZN(n19226) );
  OR2_X1 U12916 ( .A1(n19267), .A2(n19421), .ZN(n19284) );
  INV_X1 U12917 ( .A(n19318), .ZN(n19308) );
  AND2_X1 U12918 ( .A1(n19416), .A2(n19800), .ZN(n19348) );
  AND2_X1 U12919 ( .A1(n19416), .A2(n19352), .ZN(n19411) );
  NOR2_X1 U12920 ( .A1(n19383), .A2(n19603), .ZN(n19441) );
  AOI21_X1 U12921 ( .B1(n19455), .B2(n19454), .A(n19453), .ZN(n19471) );
  INV_X1 U12922 ( .A(n19232), .ZN(n19237) );
  OAI21_X1 U12923 ( .B1(n19503), .B2(n19518), .A(n19656), .ZN(n19520) );
  NOR2_X2 U12924 ( .A1(n19604), .A2(n19290), .ZN(n19541) );
  AND2_X1 U12925 ( .A1(n19810), .A2(n19822), .ZN(n19800) );
  OR3_X1 U12926 ( .A1(n13699), .A2(n13702), .A3(n13698), .ZN(n19591) );
  OAI21_X1 U12927 ( .B1(n19617), .B2(n19616), .A(n19615), .ZN(n19641) );
  AND2_X1 U12928 ( .A1(n10470), .A2(n19223), .ZN(n19688) );
  OR2_X1 U12929 ( .A1(n19810), .A2(n19183), .ZN(n19603) );
  INV_X1 U12930 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n19712) );
  INV_X1 U12931 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19728) );
  NOR2_X1 U12932 ( .A1(n15705), .A2(n12971), .ZN(n18598) );
  NOR2_X1 U12933 ( .A1(n18735), .A2(n16520), .ZN(n16555) );
  INV_X1 U12934 ( .A(n16880), .ZN(n16849) );
  NOR2_X1 U12935 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16626), .ZN(n16611) );
  NOR2_X1 U12936 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16672), .ZN(n16654) );
  NOR2_X1 U12937 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16695), .ZN(n16676) );
  NOR2_X1 U12938 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16744), .ZN(n16728) );
  NOR2_X1 U12939 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16750), .ZN(n16749) );
  NOR2_X1 U12940 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16814), .ZN(n16795) );
  NOR2_X1 U12941 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16819), .ZN(n16818) );
  AOI211_X1 U12942 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18804), .A(n18652), .B(
        n18823), .ZN(n16863) );
  NAND2_X1 U12943 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17231), .ZN(n17230) );
  NOR2_X1 U12944 ( .A1(n17241), .A2(n17268), .ZN(n17257) );
  NAND2_X1 U12945 ( .A1(n17318), .A2(P3_EAX_REG_8__SCAN_IN), .ZN(n17312) );
  NAND2_X1 U12946 ( .A1(n18812), .A2(n18599), .ZN(n17409) );
  NAND2_X1 U12947 ( .A1(n17888), .A2(n17698), .ZN(n17887) );
  INV_X1 U12948 ( .A(n17737), .ZN(n17722) );
  INV_X1 U12949 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17759) );
  INV_X1 U12950 ( .A(n18051), .ZN(n18033) );
  INV_X1 U12951 ( .A(n18120), .ZN(n18114) );
  NOR2_X1 U12952 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18759), .ZN(
        n18784) );
  NOR2_X1 U12953 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18150), .ZN(n18508) );
  INV_X1 U12954 ( .A(n18495), .ZN(n18498) );
  NOR2_X2 U12955 ( .A1(n18312), .A2(n18505), .ZN(n18542) );
  INV_X1 U12956 ( .A(n18666), .ZN(n18808) );
  NAND2_X1 U12957 ( .A1(n13364), .A2(n13135), .ZN(n13412) );
  INV_X1 U12958 ( .A(n19969), .ZN(n15945) );
  INV_X1 U12959 ( .A(n19936), .ZN(n19946) );
  INV_X1 U12960 ( .A(n19909), .ZN(n19986) );
  INV_X1 U12961 ( .A(n14554), .ZN(n14380) );
  AOI21_X2 U12962 ( .B1(n13368), .B2(n12226), .A(n19873), .ZN(n14540) );
  INV_X1 U12963 ( .A(n20925), .ZN(n20023) );
  INV_X1 U12964 ( .A(n12214), .ZN(n12215) );
  OAI21_X1 U12965 ( .B1(n14090), .B2(n14050), .A(n14049), .ZN(n14663) );
  INV_X1 U12966 ( .A(n16007), .ZN(n16034) );
  NAND2_X1 U12967 ( .A1(n13107), .A2(n13103), .ZN(n16070) );
  INV_X1 U12968 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16150) );
  OR2_X1 U12969 ( .A1(n20214), .A2(n20248), .ZN(n20164) );
  OR2_X1 U12970 ( .A1(n20214), .A2(n20403), .ZN(n20206) );
  OR2_X1 U12971 ( .A1(n20214), .A2(n20424), .ZN(n20242) );
  NAND2_X1 U12972 ( .A1(n20249), .A2(n20506), .ZN(n20303) );
  OR2_X1 U12973 ( .A1(n20348), .A2(n20403), .ZN(n20334) );
  OR2_X1 U12974 ( .A1(n20348), .A2(n20347), .ZN(n20364) );
  NAND2_X1 U12975 ( .A1(n20483), .A2(n20506), .ZN(n20423) );
  NAND2_X1 U12976 ( .A1(n20483), .A2(n20535), .ZN(n20472) );
  NAND2_X1 U12977 ( .A1(n20483), .A2(n20563), .ZN(n20499) );
  NAND2_X1 U12978 ( .A1(n20483), .A2(n20482), .ZN(n20534) );
  NAND2_X1 U12979 ( .A1(n20564), .A2(n20535), .ZN(n20568) );
  NAND2_X1 U12980 ( .A1(n20564), .A2(n20563), .ZN(n20674) );
  AND2_X1 U12981 ( .A1(n20695), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20757) );
  OR2_X1 U12982 ( .A1(n12626), .A2(n12625), .ZN(n18832) );
  INV_X1 U12983 ( .A(n19027), .ZN(n19006) );
  AND2_X2 U12984 ( .A1(n12958), .A2(n13167), .ZN(n15027) );
  NAND2_X1 U12985 ( .A1(n13463), .A2(n13462), .ZN(n19235) );
  AND2_X1 U12986 ( .A1(n12590), .A2(n13167), .ZN(n19083) );
  INV_X1 U12987 ( .A(n19100), .ZN(n19115) );
  NAND2_X1 U12988 ( .A1(n19154), .A2(n19864), .ZN(n19147) );
  INV_X1 U12989 ( .A(n13130), .ZN(n13270) );
  INV_X1 U12990 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16222) );
  INV_X1 U12991 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16251) );
  INV_X1 U12992 ( .A(n16301), .ZN(n16274) );
  INV_X1 U12993 ( .A(n16270), .ZN(n16305) );
  INV_X1 U12994 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16308) );
  INV_X1 U12995 ( .A(n19256), .ZN(n19230) );
  NAND2_X1 U12996 ( .A1(n19232), .A2(n19416), .ZN(n19287) );
  INV_X1 U12997 ( .A(n19348), .ZN(n19326) );
  NAND2_X1 U12998 ( .A1(n19319), .A2(n19800), .ZN(n19318) );
  NAND2_X1 U12999 ( .A1(n19319), .A2(n19352), .ZN(n19372) );
  INV_X1 U13000 ( .A(n19411), .ZN(n19392) );
  INV_X1 U13001 ( .A(n19441), .ZN(n19415) );
  NAND2_X1 U13002 ( .A1(n19652), .A2(n19416), .ZN(n19475) );
  OR2_X1 U13003 ( .A1(n19604), .A2(n19237), .ZN(n19482) );
  INV_X1 U13004 ( .A(n19499), .ZN(n19523) );
  INV_X1 U13005 ( .A(n19696), .ZN(n19538) );
  NAND2_X1 U13006 ( .A1(n19184), .A2(n19800), .ZN(n19579) );
  INV_X1 U13007 ( .A(n19684), .ZN(n19590) );
  INV_X1 U13008 ( .A(n19591), .ZN(n19602) );
  NAND2_X1 U13009 ( .A1(n19184), .A2(n19352), .ZN(n19645) );
  OR2_X1 U13010 ( .A1(n19604), .A2(n19603), .ZN(n19709) );
  INV_X1 U13011 ( .A(n19798), .ZN(n19722) );
  NOR2_X1 U13012 ( .A1(n18598), .A2(n17409), .ZN(n18825) );
  INV_X1 U13013 ( .A(n16863), .ZN(n16833) );
  NOR2_X1 U13014 ( .A1(n17388), .A2(n17304), .ZN(n17309) );
  NAND2_X1 U13015 ( .A1(n17362), .A2(n17406), .ZN(n17357) );
  INV_X1 U13016 ( .A(n17360), .ZN(n17375) );
  OR2_X1 U13017 ( .A1(n17409), .A2(n17348), .ZN(n17406) );
  AOI211_X1 U13018 ( .C1(n18806), .C2(n18804), .A(n17410), .B(n17409), .ZN(
        n17421) );
  INV_X1 U13019 ( .A(n17455), .ZN(n17450) );
  OR3_X1 U13020 ( .A1(n18804), .A2(n17410), .A3(n17409), .ZN(n17457) );
  NAND2_X1 U13021 ( .A1(n16403), .A2(n18132), .ZN(n18051) );
  INV_X1 U13022 ( .A(n18129), .ZN(n18116) );
  INV_X1 U13023 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18635) );
  INV_X1 U13024 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18160) );
  INV_X1 U13025 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18184) );
  INV_X1 U13026 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n20773) );
  INV_X1 U13027 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18228) );
  INV_X1 U13028 ( .A(n18229), .ZN(n18565) );
  INV_X1 U13029 ( .A(n18208), .ZN(n18571) );
  NOR2_X1 U13030 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18666) );
  INV_X1 U13031 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18682) );
  INV_X1 U13032 ( .A(n16456), .ZN(n16461) );
  NAND2_X1 U13033 ( .A1(n12245), .A2(n12244), .ZN(P1_U2873) );
  NAND2_X1 U13034 ( .A1(n12955), .A2(n12954), .ZN(P3_U2799) );
  AND2_X4 U13035 ( .A1(n10739), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10308) );
  AND2_X4 U13036 ( .A1(n10316), .A2(n10458), .ZN(n10310) );
  AND2_X4 U13037 ( .A1(n14004), .A2(n15577), .ZN(n10311) );
  NOR2_X1 U13038 ( .A1(n10082), .A2(n10081), .ZN(n10086) );
  AOI22_X1 U13039 ( .A1(n10306), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10307), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10085) );
  AND2_X4 U13040 ( .A1(n10739), .A2(n15577), .ZN(n12420) );
  AOI22_X1 U13041 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12420), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10084) );
  AOI22_X1 U13042 ( .A1(n10311), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10088) );
  AOI22_X1 U13043 ( .A1(n10306), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10307), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10087) );
  AND3_X1 U13044 ( .A1(n10088), .A2(n10087), .A3(n10115), .ZN(n10091) );
  AOI22_X1 U13045 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12420), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10090) );
  AOI22_X1 U13046 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10089) );
  AOI22_X1 U13047 ( .A1(n10306), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10307), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10094) );
  AOI22_X1 U13048 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10093) );
  AOI22_X1 U13049 ( .A1(n9571), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12420), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10092) );
  NAND3_X1 U13050 ( .A1(n10094), .A2(n10093), .A3(n10092), .ZN(n10097) );
  AOI22_X1 U13051 ( .A1(n10311), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10095) );
  AOI22_X1 U13052 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12420), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10101) );
  AOI22_X1 U13053 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10100) );
  AOI22_X1 U13054 ( .A1(n10306), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10307), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10099) );
  AOI22_X1 U13055 ( .A1(n10311), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10098) );
  NAND4_X1 U13056 ( .A1(n10101), .A2(n10100), .A3(n10099), .A4(n10098), .ZN(
        n10102) );
  AOI22_X1 U13057 ( .A1(n10306), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10307), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10107) );
  AOI22_X1 U13058 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10106) );
  AOI22_X1 U13059 ( .A1(n9571), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12420), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10105) );
  NAND3_X1 U13060 ( .A1(n10107), .A2(n10106), .A3(n10105), .ZN(n10110) );
  AOI22_X1 U13061 ( .A1(n10311), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10108) );
  INV_X1 U13062 ( .A(n10108), .ZN(n10109) );
  AOI22_X1 U13063 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10114) );
  AOI22_X1 U13064 ( .A1(n10311), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10113) );
  AOI22_X1 U13065 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12420), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10112) );
  AOI22_X1 U13066 ( .A1(n10306), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10307), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10111) );
  NAND4_X1 U13067 ( .A1(n10114), .A2(n10113), .A3(n10112), .A4(n10111), .ZN(
        n10116) );
  AOI22_X1 U13068 ( .A1(n10311), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10120) );
  AOI22_X1 U13069 ( .A1(n9571), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12420), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10118) );
  AOI22_X1 U13070 ( .A1(n10306), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10307), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10117) );
  NAND4_X1 U13071 ( .A1(n10120), .A2(n10119), .A3(n10118), .A4(n10117), .ZN(
        n10121) );
  AOI22_X1 U13072 ( .A1(n9571), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12420), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10125) );
  AOI22_X1 U13073 ( .A1(n10306), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10307), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10124) );
  AOI22_X1 U13074 ( .A1(n10311), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10122) );
  NAND4_X1 U13075 ( .A1(n10125), .A2(n10124), .A3(n10123), .A4(n10122), .ZN(
        n10126) );
  NAND2_X1 U13076 ( .A1(n10126), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10127) );
  INV_X1 U13077 ( .A(n10184), .ZN(n10129) );
  AOI22_X1 U13078 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10310), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10135) );
  AOI22_X1 U13079 ( .A1(n10306), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10307), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10134) );
  AOI22_X1 U13080 ( .A1(n10311), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10133) );
  AOI22_X1 U13081 ( .A1(n10308), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12420), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10131) );
  NAND4_X1 U13082 ( .A1(n10135), .A2(n10134), .A3(n10133), .A4(n10132), .ZN(
        n10142) );
  AOI22_X1 U13083 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12420), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10139) );
  AOI22_X1 U13084 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10138) );
  AOI22_X1 U13085 ( .A1(n10306), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10307), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10137) );
  AOI22_X1 U13086 ( .A1(n10311), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10136) );
  AOI22_X1 U13087 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12420), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U13088 ( .A1(n9571), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10145) );
  AOI22_X1 U13089 ( .A1(n10306), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10307), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10144) );
  AOI22_X1 U13090 ( .A1(n10311), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10143) );
  NAND4_X1 U13091 ( .A1(n10146), .A2(n10145), .A3(n10144), .A4(n10143), .ZN(
        n10147) );
  AOI22_X1 U13092 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10151) );
  AOI22_X1 U13093 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12420), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10150) );
  AOI22_X1 U13094 ( .A1(n10306), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10307), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U13095 ( .A1(n10311), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10148) );
  NAND4_X1 U13096 ( .A1(n10151), .A2(n10150), .A3(n10149), .A4(n10148), .ZN(
        n10152) );
  AOI22_X1 U13097 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10158) );
  AOI22_X1 U13098 ( .A1(n9571), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12420), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10157) );
  AOI22_X1 U13099 ( .A1(n10306), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10307), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10156) );
  AOI22_X1 U13100 ( .A1(n10311), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10155) );
  NAND4_X1 U13101 ( .A1(n10158), .A2(n10157), .A3(n10156), .A4(n10155), .ZN(
        n10164) );
  AOI22_X1 U13102 ( .A1(n9571), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10310), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10162) );
  AOI22_X1 U13103 ( .A1(n10311), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10161) );
  AOI22_X1 U13104 ( .A1(n10306), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10307), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10160) );
  AOI22_X1 U13105 ( .A1(n10308), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12420), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10159) );
  NAND4_X1 U13106 ( .A1(n10162), .A2(n10161), .A3(n10160), .A4(n10159), .ZN(
        n10163) );
  MUX2_X2 U13107 ( .A(n10164), .B(n10163), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19852) );
  NOR2_X1 U13108 ( .A1(n13168), .A2(n19852), .ZN(n10168) );
  NAND2_X1 U13109 ( .A1(n10182), .A2(n10889), .ZN(n10203) );
  NAND3_X1 U13110 ( .A1(n10166), .A2(n10203), .A3(n10060), .ZN(n10167) );
  NAND2_X1 U13111 ( .A1(n10168), .A2(n10167), .ZN(n10886) );
  AOI22_X1 U13112 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12420), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U13113 ( .A1(n10306), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10307), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10171) );
  AOI22_X1 U13114 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10170) );
  AOI22_X1 U13115 ( .A1(n10311), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10169) );
  NAND4_X1 U13116 ( .A1(n10172), .A2(n10171), .A3(n10170), .A4(n10169), .ZN(
        n10173) );
  NAND2_X1 U13117 ( .A1(n10173), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10180) );
  AOI22_X1 U13118 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10310), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10177) );
  AOI22_X1 U13119 ( .A1(n10308), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12420), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U13120 ( .A1(n10311), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U13121 ( .A1(n10306), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10307), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10174) );
  NAND4_X1 U13122 ( .A1(n10177), .A2(n10176), .A3(n10175), .A4(n10174), .ZN(
        n10178) );
  NAND2_X4 U13123 ( .A1(n10180), .A2(n10179), .ZN(n19196) );
  NAND2_X1 U13124 ( .A1(n10891), .A2(n16322), .ZN(n10181) );
  NAND2_X1 U13126 ( .A1(n10877), .A2(n10889), .ZN(n10187) );
  NAND2_X1 U13127 ( .A1(n10187), .A2(n10186), .ZN(n10218) );
  NAND2_X1 U13128 ( .A1(n10218), .A2(n10701), .ZN(n10188) );
  NAND2_X1 U13129 ( .A1(n10219), .A2(n10188), .ZN(n10189) );
  NAND2_X1 U13130 ( .A1(n10189), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10193) );
  NAND3_X1 U13131 ( .A1(n16321), .A2(n10874), .A3(n19196), .ZN(n10192) );
  NAND2_X1 U13132 ( .A1(n19852), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10698) );
  NAND2_X2 U13133 ( .A1(n11115), .A2(n13273), .ZN(n10228) );
  NAND2_X1 U13134 ( .A1(n13168), .A2(n16322), .ZN(n10748) );
  INV_X1 U13135 ( .A(n10700), .ZN(n13170) );
  NAND2_X1 U13136 ( .A1(n13170), .A2(n10194), .ZN(n10206) );
  INV_X2 U13137 ( .A(n10879), .ZN(n10892) );
  NAND2_X1 U13138 ( .A1(n10892), .A2(n19213), .ZN(n10195) );
  NOR2_X1 U13139 ( .A1(n10206), .A2(n10195), .ZN(n10196) );
  OR2_X2 U13140 ( .A1(n11117), .A2(n10196), .ZN(n10868) );
  NOR2_X1 U13141 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19861) );
  NOR2_X1 U13142 ( .A1(n19196), .A2(n18828), .ZN(n10205) );
  NAND2_X1 U13143 ( .A1(n11117), .A2(n10205), .ZN(n10209) );
  INV_X1 U13144 ( .A(n10206), .ZN(n10207) );
  NAND3_X1 U13145 ( .A1(n10207), .A2(n10892), .A3(n12247), .ZN(n10208) );
  NOR2_X1 U13146 ( .A1(n12277), .A2(n16322), .ZN(n10210) );
  AND2_X2 U13147 ( .A1(n10744), .A2(n10210), .ZN(n10239) );
  INV_X1 U13148 ( .A(n10211), .ZN(n10881) );
  NOR2_X1 U13149 ( .A1(n10879), .A2(n10212), .ZN(n10213) );
  INV_X1 U13150 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n10214) );
  NAND2_X1 U13151 ( .A1(n10216), .A2(n10215), .ZN(n10217) );
  AND2_X2 U13152 ( .A1(n10236), .A2(n10217), .ZN(n10264) );
  BUF_X1 U13153 ( .A(n10218), .Z(n10890) );
  NAND2_X1 U13154 ( .A1(n10890), .A2(n10891), .ZN(n10220) );
  NAND2_X1 U13155 ( .A1(n10220), .A2(n10219), .ZN(n10221) );
  NAND2_X1 U13156 ( .A1(n10221), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10230) );
  NAND2_X1 U13157 ( .A1(n9569), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10229) );
  INV_X1 U13158 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n10485) );
  AND2_X1 U13159 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10223) );
  NOR2_X1 U13160 ( .A1(n19861), .A2(n10223), .ZN(n10224) );
  NOR2_X1 U13161 ( .A1(n10231), .A2(n13035), .ZN(n10232) );
  OAI22_X1 U13162 ( .A1(n10237), .A2(n10232), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10770), .ZN(n10235) );
  AOI22_X1 U13163 ( .A1(n14003), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19861), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10234) );
  NAND2_X1 U13164 ( .A1(n10235), .A2(n10234), .ZN(n10258) );
  NAND2_X1 U13165 ( .A1(n10263), .A2(n10236), .ZN(n10262) );
  AOI21_X1 U13166 ( .B1(n18828), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10238) );
  AOI22_X1 U13167 ( .A1(n10858), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10242) );
  INV_X1 U13168 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10240) );
  NAND2_X1 U13169 ( .A1(n10243), .A2(n10069), .ZN(n10244) );
  AND2_X2 U13170 ( .A1(n10246), .A2(n10245), .ZN(n10261) );
  NAND2_X1 U13171 ( .A1(n10262), .A2(n10261), .ZN(n10247) );
  NAND2_X1 U13172 ( .A1(n10248), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10250) );
  NAND2_X1 U13173 ( .A1(n19861), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10249) );
  NAND2_X1 U13174 ( .A1(n10250), .A2(n10249), .ZN(n10255) );
  INV_X1 U13175 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10253) );
  NAND2_X1 U13176 ( .A1(n9569), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10252) );
  AOI22_X1 U13177 ( .A1(n10862), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10251) );
  OAI211_X1 U13178 ( .C1(n9580), .C2(n10253), .A(n10252), .B(n10251), .ZN(
        n10254) );
  NAND2_X1 U13179 ( .A1(n10255), .A2(n10254), .ZN(n10256) );
  XNOR2_X2 U13180 ( .A(n10262), .B(n10261), .ZN(n12246) );
  BUF_X1 U13181 ( .A(n10263), .Z(n10267) );
  INV_X1 U13182 ( .A(n10264), .ZN(n10270) );
  NAND2_X1 U13183 ( .A1(n10265), .A2(n10270), .ZN(n10266) );
  NAND2_X1 U13184 ( .A1(n12246), .A2(n15568), .ZN(n10268) );
  NOR2_X2 U13185 ( .A1(n10286), .A2(n10268), .ZN(n19386) );
  INV_X1 U13186 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12299) );
  INV_X1 U13187 ( .A(n10299), .ZN(n10269) );
  BUF_X2 U13188 ( .A(n10277), .Z(n12261) );
  INV_X1 U13189 ( .A(n10290), .ZN(n10271) );
  INV_X1 U13190 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10272) );
  AOI21_X1 U13191 ( .B1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n19386), .A(
        n10273), .ZN(n10285) );
  INV_X1 U13192 ( .A(n12246), .ZN(n19178) );
  INV_X2 U13194 ( .A(n10278), .ZN(n10276) );
  AND2_X2 U13195 ( .A1(n10276), .A2(n10299), .ZN(n10411) );
  INV_X1 U13196 ( .A(n15568), .ZN(n13911) );
  NAND2_X1 U13197 ( .A1(n13911), .A2(n10260), .ZN(n10280) );
  INV_X1 U13198 ( .A(n10280), .ZN(n10275) );
  AND2_X2 U13199 ( .A1(n10276), .A2(n10275), .ZN(n10417) );
  AOI22_X1 U13200 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10411), .B1(
        n10417), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10284) );
  INV_X1 U13201 ( .A(n10281), .ZN(n10300) );
  AOI22_X1 U13202 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10359), .B1(
        n10412), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10283) );
  NOR2_X2 U13203 ( .A1(n10286), .A2(n10279), .ZN(n19262) );
  INV_X1 U13204 ( .A(n19555), .ZN(n19548) );
  AOI22_X1 U13205 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19262), .B1(
        n19548), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10282) );
  INV_X1 U13206 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12429) );
  INV_X1 U13207 ( .A(n12261), .ZN(n10287) );
  NAND2_X2 U13208 ( .A1(n10288), .A2(n10287), .ZN(n10398) );
  INV_X1 U13209 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10289) );
  INV_X1 U13210 ( .A(n12416), .ZN(n13037) );
  OAI21_X1 U13211 ( .B1(n10398), .B2(n10289), .A(n13037), .ZN(n10293) );
  NAND2_X1 U13212 ( .A1(n12246), .A2(n10290), .ZN(n10291) );
  INV_X1 U13213 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10967) );
  NOR2_X1 U13214 ( .A1(n19357), .A2(n10967), .ZN(n10292) );
  NOR2_X1 U13215 ( .A1(n10293), .A2(n10292), .ZN(n10295) );
  NAND2_X1 U13216 ( .A1(n19614), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10294) );
  OAI211_X1 U13217 ( .C1(n19188), .C2(n12429), .A(n10295), .B(n10294), .ZN(
        n10296) );
  INV_X1 U13218 ( .A(n10296), .ZN(n10305) );
  INV_X1 U13219 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10303) );
  NAND2_X1 U13220 ( .A1(n19494), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10302) );
  NAND2_X1 U13221 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10301) );
  OAI211_X1 U13222 ( .C1(n19328), .C2(n10303), .A(n10302), .B(n10301), .ZN(
        n10304) );
  INV_X1 U13223 ( .A(n10308), .ZN(n12399) );
  AND2_X2 U13224 ( .A1(n10308), .A2(n10115), .ZN(n12394) );
  AOI22_X1 U13225 ( .A1(n12383), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12394), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10314) );
  AND2_X2 U13226 ( .A1(n10310), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10422) );
  AOI22_X1 U13227 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10422), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10313) );
  AND2_X1 U13228 ( .A1(n12571), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10371) );
  AOI22_X1 U13229 ( .A1(n12321), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10312) );
  NAND4_X1 U13230 ( .A1(n10315), .A2(n10314), .A3(n10313), .A4(n10312), .ZN(
        n10324) );
  INV_X1 U13231 ( .A(n12401), .ZN(n10317) );
  AOI22_X1 U13232 ( .A1(n11072), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12375), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10322) );
  AOI22_X1 U13233 ( .A1(n11071), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9567), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10321) );
  AOI22_X1 U13234 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10331), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10320) );
  AND2_X1 U13235 ( .A1(n12420), .A2(n10115), .ZN(n10341) );
  AOI22_X1 U13236 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10341), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10319) );
  NAND4_X1 U13237 ( .A1(n10322), .A2(n10321), .A3(n10320), .A4(n10319), .ZN(
        n10323) );
  NAND2_X1 U13238 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10326) );
  NAND2_X1 U13239 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10325) );
  AND2_X1 U13240 ( .A1(n10326), .A2(n10325), .ZN(n10330) );
  AOI22_X1 U13241 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12394), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10329) );
  AOI22_X1 U13242 ( .A1(n10987), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10328) );
  AOI22_X1 U13243 ( .A1(n10371), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10327) );
  NAND4_X1 U13244 ( .A1(n10330), .A2(n10329), .A3(n10328), .A4(n10327), .ZN(
        n10339) );
  AOI22_X1 U13245 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10341), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10337) );
  AOI22_X1 U13246 ( .A1(n11072), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n9567), .ZN(n10333) );
  NAND2_X1 U13247 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10332) );
  AND2_X1 U13248 ( .A1(n10333), .A2(n10332), .ZN(n10336) );
  AOI22_X1 U13249 ( .A1(n11071), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12375), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10335) );
  NAND2_X1 U13250 ( .A1(n10376), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10334) );
  NAND4_X1 U13251 ( .A1(n10337), .A2(n10336), .A3(n10335), .A4(n10334), .ZN(
        n10338) );
  OR2_X1 U13252 ( .A1(n19196), .A2(n11141), .ZN(n10340) );
  OR2_X1 U13253 ( .A1(n13400), .A2(n10340), .ZN(n11138) );
  AOI22_X1 U13254 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n10422), .B1(
        n12393), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10345) );
  AOI22_X1 U13255 ( .A1(n10987), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U13256 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n12383), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10343) );
  AOI22_X1 U13257 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n12394), .B1(
        n10341), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10342) );
  NAND4_X1 U13258 ( .A1(n10345), .A2(n10344), .A3(n10343), .A4(n10342), .ZN(
        n10353) );
  AOI22_X1 U13259 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10351) );
  INV_X1 U13260 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10346) );
  INV_X1 U13261 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10983) );
  OAI22_X1 U13262 ( .A1(n12367), .A2(n10346), .B1(n10983), .B2(n12364), .ZN(
        n10347) );
  AOI21_X1 U13263 ( .B1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B2(n10331), .A(
        n10347), .ZN(n10350) );
  AOI22_X1 U13264 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n11071), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10349) );
  NAND2_X1 U13265 ( .A1(n10376), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10348) );
  NAND4_X1 U13266 ( .A1(n10351), .A2(n10350), .A3(n10349), .A4(n10348), .ZN(
        n10352) );
  NAND2_X1 U13267 ( .A1(n11138), .A2(n11139), .ZN(n10354) );
  AOI22_X1 U13268 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19614), .B1(
        n10412), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10356) );
  AOI22_X1 U13269 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10411), .B1(
        n10417), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10355) );
  INV_X1 U13270 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12476) );
  INV_X1 U13271 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10358) );
  OAI22_X1 U13272 ( .A1(n19500), .A2(n12476), .B1(n10358), .B2(n19555), .ZN(
        n10363) );
  AOI22_X1 U13273 ( .A1(n19262), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n19386), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10361) );
  AOI22_X1 U13274 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n10511), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10360) );
  NAND2_X1 U13275 ( .A1(n10361), .A2(n10360), .ZN(n10362) );
  NOR2_X1 U13276 ( .A1(n10363), .A2(n10362), .ZN(n10369) );
  INV_X1 U13277 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10364) );
  INV_X1 U13278 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11004) );
  OAI22_X1 U13279 ( .A1(n10364), .A2(n10398), .B1(n19357), .B2(n11004), .ZN(
        n10367) );
  INV_X1 U13280 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12326) );
  INV_X1 U13281 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10365) );
  NOR2_X1 U13282 ( .A1(n10367), .A2(n10366), .ZN(n10368) );
  AOI22_X1 U13283 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10341), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10375) );
  AOI22_X1 U13284 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10374) );
  AOI22_X1 U13285 ( .A1(n10987), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12394), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10373) );
  AOI22_X1 U13286 ( .A1(n10371), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10372) );
  AOI22_X1 U13287 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10382) );
  AOI22_X1 U13288 ( .A1(n11072), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9567), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U13289 ( .A1(n11071), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12375), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10378) );
  NAND2_X1 U13290 ( .A1(n10376), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10377) );
  AND2_X1 U13291 ( .A1(n10378), .A2(n10377), .ZN(n10380) );
  NAND2_X1 U13292 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10379) );
  NAND4_X1 U13293 ( .A1(n10382), .A2(n10381), .A3(n10380), .A4(n10379), .ZN(
        n10383) );
  NAND2_X1 U13294 ( .A1(n10472), .A2(n19853), .ZN(n10384) );
  AOI22_X1 U13295 ( .A1(n10987), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10388) );
  AOI22_X1 U13296 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10387) );
  AOI22_X1 U13297 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U13298 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10385) );
  NAND4_X1 U13299 ( .A1(n10388), .A2(n10387), .A3(n10386), .A4(n10385), .ZN(
        n10397) );
  AOI22_X1 U13300 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10341), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10395) );
  INV_X1 U13301 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10390) );
  INV_X1 U13302 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11023) );
  OAI22_X1 U13303 ( .A1(n12367), .A2(n10390), .B1(n12364), .B2(n11023), .ZN(
        n10391) );
  AOI21_X1 U13304 ( .B1(n10376), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n10391), .ZN(n10394) );
  INV_X1 U13305 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n20779) );
  AOI22_X1 U13306 ( .A1(n11071), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10393) );
  NAND2_X1 U13307 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10392) );
  NAND4_X1 U13308 ( .A1(n10395), .A2(n10394), .A3(n10393), .A4(n10392), .ZN(
        n10396) );
  INV_X1 U13309 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10400) );
  INV_X1 U13310 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10428) );
  OAI22_X1 U13311 ( .A1(n10400), .A2(n10398), .B1(n10399), .B2(n10428), .ZN(
        n10402) );
  INV_X1 U13312 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11036) );
  INV_X1 U13313 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12351) );
  NOR2_X1 U13314 ( .A1(n10402), .A2(n10401), .ZN(n10410) );
  AOI22_X1 U13315 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19323), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10409) );
  INV_X1 U13316 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10404) );
  INV_X1 U13317 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12524) );
  OAI22_X1 U13318 ( .A1(n10404), .A2(n19555), .B1(n19500), .B2(n12524), .ZN(
        n10405) );
  AOI22_X1 U13319 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19386), .B1(
        n19262), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10406) );
  NAND3_X1 U13320 ( .A1(n10410), .A2(n10409), .A3(n10408), .ZN(n10416) );
  AOI22_X1 U13321 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19614), .B1(
        n10411), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10414) );
  AOI22_X1 U13322 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n10511), .B1(
        n13740), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10413) );
  INV_X1 U13323 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10418) );
  INV_X1 U13324 ( .A(n10359), .ZN(n10513) );
  INV_X1 U13325 ( .A(n10417), .ZN(n10520) );
  INV_X1 U13326 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12522) );
  OAI22_X1 U13327 ( .A1(n10418), .A2(n10513), .B1(n10520), .B2(n12522), .ZN(
        n10419) );
  INV_X1 U13328 ( .A(n10419), .ZN(n10420) );
  AOI22_X1 U13329 ( .A1(n10987), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10427) );
  AOI22_X1 U13330 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10426) );
  AOI22_X1 U13331 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10425) );
  AOI22_X1 U13332 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10424) );
  NAND4_X1 U13333 ( .A1(n10427), .A2(n10426), .A3(n10425), .A4(n10424), .ZN(
        n10436) );
  AOI22_X1 U13334 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10341), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10434) );
  INV_X1 U13335 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10429) );
  OAI22_X1 U13336 ( .A1(n12367), .A2(n10429), .B1(n12364), .B2(n10428), .ZN(
        n10430) );
  AOI21_X1 U13337 ( .B1(n10376), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n10430), .ZN(n10433) );
  AOI22_X1 U13338 ( .A1(n11071), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10432) );
  NAND2_X1 U13339 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10431) );
  NAND4_X1 U13340 ( .A1(n10434), .A2(n10433), .A3(n10432), .A4(n10431), .ZN(
        n10435) );
  INV_X1 U13341 ( .A(n10935), .ZN(n10437) );
  NAND2_X1 U13342 ( .A1(n19853), .A2(n10437), .ZN(n10438) );
  XNOR2_X1 U13343 ( .A(n11151), .B(n10508), .ZN(n11157) );
  NAND2_X1 U13344 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10443) );
  NAND2_X1 U13345 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10442) );
  NAND2_X1 U13346 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10441) );
  NAND2_X1 U13347 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10440) );
  INV_X1 U13348 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10444) );
  INV_X1 U13349 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12384) );
  OAI22_X1 U13350 ( .A1(n12367), .A2(n10444), .B1(n12384), .B2(n12364), .ZN(
        n10445) );
  AOI21_X1 U13351 ( .B1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n10331), .A(
        n10445), .ZN(n10448) );
  AOI22_X1 U13352 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n11071), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10447) );
  NAND2_X1 U13353 ( .A1(n10376), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10446) );
  NAND2_X1 U13354 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10452) );
  NAND2_X1 U13355 ( .A1(n12321), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10451) );
  NAND2_X1 U13356 ( .A1(n10423), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10450) );
  NAND2_X1 U13357 ( .A1(n12383), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10449) );
  AOI22_X1 U13358 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10341), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10454) );
  NAND4_X1 U13359 ( .A1(n10457), .A2(n10456), .A3(n10455), .A4(n10454), .ZN(
        n10559) );
  NAND2_X1 U13360 ( .A1(n11157), .A2(n11175), .ZN(n10478) );
  MUX2_X1 U13361 ( .A(n19819), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        n10458), .Z(n10466) );
  INV_X1 U13362 ( .A(n10466), .ZN(n10461) );
  NAND2_X1 U13363 ( .A1(n19828), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10460) );
  NAND2_X1 U13364 ( .A1(n10077), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10459) );
  NAND2_X1 U13365 ( .A1(n10460), .A2(n10459), .ZN(n10703) );
  NAND2_X1 U13366 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19837), .ZN(
        n10702) );
  NAND2_X1 U13367 ( .A1(n10704), .A2(n10460), .ZN(n10467) );
  NAND2_X1 U13368 ( .A1(n10461), .A2(n10467), .ZN(n10463) );
  NAND2_X1 U13369 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19819), .ZN(
        n10462) );
  INV_X1 U13370 ( .A(n10474), .ZN(n10464) );
  MUX2_X1 U13371 ( .A(n16335), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        n10115), .Z(n10473) );
  NAND3_X1 U13372 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10697), .A3(
        n16308), .ZN(n10713) );
  MUX2_X1 U13373 ( .A(n10713), .B(n10931), .S(n10701), .Z(n10725) );
  INV_X1 U13374 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n10774) );
  MUX2_X1 U13375 ( .A(n10725), .B(n10774), .S(n14236), .Z(n10499) );
  XNOR2_X1 U13376 ( .A(n10467), .B(n10466), .ZN(n10731) );
  MUX2_X1 U13377 ( .A(n10468), .B(n10731), .S(n13035), .Z(n10720) );
  MUX2_X1 U13378 ( .A(n10720), .B(n10240), .S(n14236), .Z(n10490) );
  OR2_X1 U13379 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(
        n10471) );
  MUX2_X1 U13380 ( .A(n10471), .B(n11141), .S(n10470), .Z(n10487) );
  XNOR2_X1 U13381 ( .A(n10474), .B(n10473), .ZN(n10712) );
  INV_X1 U13382 ( .A(n10712), .ZN(n10475) );
  AND2_X2 U13383 ( .A1(n10499), .A2(n10482), .ZN(n10555) );
  INV_X1 U13384 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n18994) );
  MUX2_X1 U13385 ( .A(n10935), .B(n18994), .S(n14236), .Z(n10554) );
  XNOR2_X1 U13386 ( .A(n10555), .B(n10554), .ZN(n18995) );
  INV_X1 U13387 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n20886) );
  INV_X1 U13388 ( .A(n10482), .ZN(n10501) );
  NAND2_X1 U13389 ( .A1(n10489), .A2(n10483), .ZN(n10484) );
  NAND2_X1 U13390 ( .A1(n10501), .A2(n10484), .ZN(n13824) );
  NAND2_X1 U13391 ( .A1(n10495), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13878) );
  OAI21_X1 U13392 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19837), .A(
        n10702), .ZN(n10737) );
  MUX2_X1 U13393 ( .A(n10737), .B(n13400), .S(n10701), .Z(n10723) );
  MUX2_X1 U13394 ( .A(n10723), .B(n10485), .S(n14236), .Z(n19028) );
  INV_X1 U13395 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13404) );
  NOR2_X1 U13396 ( .A1(n19028), .A2(n13404), .ZN(n13403) );
  INV_X1 U13397 ( .A(n13403), .ZN(n15243) );
  NAND3_X1 U13398 ( .A1(n14236), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n10486) );
  NAND2_X1 U13399 ( .A1(n10487), .A2(n10486), .ZN(n15244) );
  NOR2_X1 U13400 ( .A1(n15243), .A2(n15244), .ZN(n10488) );
  NAND2_X1 U13401 ( .A1(n15243), .A2(n15244), .ZN(n15242) );
  OAI21_X1 U13402 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10488), .A(
        n15242), .ZN(n13289) );
  OAI21_X1 U13403 ( .B1(n10491), .B2(n10490), .A(n10489), .ZN(n13865) );
  INV_X1 U13404 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13297) );
  XNOR2_X1 U13405 ( .A(n13865), .B(n13297), .ZN(n13288) );
  OR2_X1 U13406 ( .A1(n13289), .A2(n13288), .ZN(n13286) );
  INV_X1 U13407 ( .A(n13865), .ZN(n10492) );
  NAND2_X1 U13408 ( .A1(n10492), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10493) );
  NAND2_X1 U13409 ( .A1(n13286), .A2(n10493), .ZN(n13880) );
  INV_X1 U13410 ( .A(n13880), .ZN(n10494) );
  NAND2_X1 U13411 ( .A1(n13878), .A2(n10494), .ZN(n10498) );
  INV_X1 U13412 ( .A(n10495), .ZN(n10497) );
  INV_X1 U13413 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10496) );
  INV_X1 U13414 ( .A(n10555), .ZN(n10503) );
  INV_X1 U13415 ( .A(n10499), .ZN(n10500) );
  NAND2_X1 U13416 ( .A1(n10501), .A2(n10500), .ZN(n10502) );
  NAND2_X1 U13417 ( .A1(n10503), .A2(n10502), .ZN(n19007) );
  INV_X1 U13418 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13948) );
  INV_X1 U13419 ( .A(n19007), .ZN(n10504) );
  NAND2_X1 U13420 ( .A1(n10504), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10505) );
  NAND2_X1 U13421 ( .A1(n10506), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10507) );
  INV_X1 U13422 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10510) );
  INV_X1 U13423 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12541) );
  OAI22_X1 U13424 ( .A1(n10510), .A2(n19555), .B1(n19500), .B2(n12541), .ZN(
        n10515) );
  INV_X1 U13425 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11056) );
  INV_X1 U13426 ( .A(n10511), .ZN(n19647) );
  INV_X1 U13427 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10512) );
  OAI22_X1 U13428 ( .A1(n11056), .A2(n19647), .B1(n10513), .B2(n10512), .ZN(
        n10514) );
  NOR2_X1 U13429 ( .A1(n10515), .A2(n10514), .ZN(n10536) );
  INV_X1 U13430 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10544) );
  INV_X1 U13431 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13601) );
  INV_X1 U13432 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10519) );
  INV_X1 U13433 ( .A(n19614), .ZN(n19611) );
  INV_X1 U13434 ( .A(n13740), .ZN(n13733) );
  INV_X1 U13435 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10518) );
  OAI22_X1 U13436 ( .A1(n10519), .A2(n19611), .B1(n13733), .B2(n10518), .ZN(
        n10524) );
  INV_X1 U13437 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10522) );
  INV_X1 U13438 ( .A(n10411), .ZN(n10521) );
  INV_X1 U13439 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12539) );
  OAI22_X1 U13440 ( .A1(n10522), .A2(n10521), .B1(n10520), .B2(n12539), .ZN(
        n10523) );
  NOR2_X1 U13441 ( .A1(n10524), .A2(n10523), .ZN(n10534) );
  INV_X1 U13442 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10526) );
  INV_X1 U13443 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10525) );
  OAI22_X1 U13444 ( .A1(n10526), .A2(n10398), .B1(n19357), .B2(n10525), .ZN(
        n10527) );
  INV_X1 U13445 ( .A(n10527), .ZN(n10532) );
  INV_X1 U13446 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10543) );
  INV_X1 U13447 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12365) );
  INV_X1 U13448 ( .A(n10528), .ZN(n10531) );
  NAND2_X1 U13449 ( .A1(n19386), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10530) );
  NAND2_X1 U13450 ( .A1(n19262), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10529) );
  NAND4_X1 U13451 ( .A1(n10536), .A2(n10535), .A3(n10534), .A4(n10533), .ZN(
        n10553) );
  AOI22_X1 U13452 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n10422), .B1(
        n10987), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10542) );
  AOI22_X1 U13453 ( .A1(n12321), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U13454 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10341), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10540) );
  AOI22_X1 U13455 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12394), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10539) );
  NAND4_X1 U13456 ( .A1(n10542), .A2(n10541), .A3(n10540), .A4(n10539), .ZN(
        n10551) );
  AOI22_X1 U13457 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10549) );
  OAI22_X1 U13458 ( .A1(n12367), .A2(n10544), .B1(n10543), .B2(n12364), .ZN(
        n10545) );
  AOI21_X1 U13459 ( .B1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B2(n10376), .A(
        n10545), .ZN(n10548) );
  AOI22_X1 U13460 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n11071), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10547) );
  NAND2_X1 U13461 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10546) );
  NAND4_X1 U13462 ( .A1(n10549), .A2(n10548), .A3(n10547), .A4(n10546), .ZN(
        n10550) );
  NAND2_X1 U13463 ( .A1(n10938), .A2(n12416), .ZN(n10552) );
  NAND2_X1 U13464 ( .A1(n11160), .A2(n11175), .ZN(n10556) );
  MUX2_X1 U13465 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n10938), .S(n10470), .Z(
        n10557) );
  XNOR2_X1 U13466 ( .A(n10558), .B(n10557), .ZN(n18981) );
  INV_X1 U13467 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15537) );
  NOR2_X2 U13468 ( .A1(n10558), .A2(n10557), .ZN(n10564) );
  INV_X1 U13469 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10786) );
  MUX2_X1 U13470 ( .A(n10786), .B(n10559), .S(n10470), .Z(n10562) );
  NAND2_X1 U13471 ( .A1(n14236), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10560) );
  OR2_X1 U13472 ( .A1(n10575), .A2(n10560), .ZN(n10561) );
  NAND2_X1 U13473 ( .A1(n10574), .A2(n10561), .ZN(n13860) );
  NOR2_X1 U13474 ( .A1(n13860), .A2(n11175), .ZN(n10569) );
  NAND2_X1 U13475 ( .A1(n10569), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15507) );
  INV_X1 U13476 ( .A(n10562), .ZN(n10563) );
  XNOR2_X1 U13477 ( .A(n10564), .B(n10563), .ZN(n18974) );
  NAND2_X1 U13478 ( .A1(n18974), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15508) );
  AND2_X1 U13479 ( .A1(n15507), .A2(n15508), .ZN(n10566) );
  NAND2_X1 U13480 ( .A1(n10565), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15226) );
  AND2_X1 U13481 ( .A1(n10566), .A2(n15226), .ZN(n10567) );
  NAND2_X1 U13482 ( .A1(n14236), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10568) );
  XNOR2_X1 U13483 ( .A(n10574), .B(n10568), .ZN(n18964) );
  NAND2_X1 U13484 ( .A1(n18964), .A2(n14239), .ZN(n10578) );
  INV_X1 U13485 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15486) );
  AND2_X1 U13486 ( .A1(n10578), .A2(n15486), .ZN(n15493) );
  INV_X1 U13487 ( .A(n15493), .ZN(n10572) );
  INV_X1 U13488 ( .A(n10569), .ZN(n10570) );
  INV_X1 U13489 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11174) );
  NAND2_X1 U13490 ( .A1(n10570), .A2(n11174), .ZN(n15506) );
  INV_X1 U13491 ( .A(n18974), .ZN(n10571) );
  INV_X1 U13492 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15520) );
  NAND2_X1 U13493 ( .A1(n10571), .A2(n15520), .ZN(n15510) );
  AND2_X1 U13494 ( .A1(n15506), .A2(n15510), .ZN(n15489) );
  AND2_X1 U13495 ( .A1(n10572), .A2(n15489), .ZN(n10573) );
  NAND2_X2 U13496 ( .A1(n10575), .A2(n10470), .ZN(n10670) );
  NAND3_X1 U13497 ( .A1(n10580), .A2(n14236), .A3(P2_EBX_REG_10__SCAN_IN), 
        .ZN(n10576) );
  OAI211_X1 U13498 ( .C1(n10580), .C2(P2_EBX_REG_10__SCAN_IN), .A(n10670), .B(
        n10576), .ZN(n18950) );
  INV_X1 U13499 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n20795) );
  OAI21_X1 U13500 ( .B1(n18950), .B2(n11175), .A(n20795), .ZN(n15471) );
  NAND2_X1 U13501 ( .A1(n14239), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10577) );
  OR2_X1 U13502 ( .A1(n18950), .A2(n10577), .ZN(n15470) );
  OR2_X1 U13503 ( .A1(n10578), .A2(n15486), .ZN(n15488) );
  AND2_X1 U13504 ( .A1(n15470), .A2(n15488), .ZN(n10579) );
  INV_X1 U13505 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n18944) );
  NAND2_X1 U13506 ( .A1(n14236), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10583) );
  INV_X1 U13507 ( .A(n10581), .ZN(n10582) );
  OR2_X1 U13508 ( .A1(n10583), .A2(n10582), .ZN(n10584) );
  NAND2_X1 U13509 ( .A1(n10617), .A2(n10584), .ZN(n18932) );
  INV_X1 U13510 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15432) );
  INV_X1 U13511 ( .A(n10585), .ZN(n10586) );
  NAND2_X1 U13512 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n10586), .ZN(n10587) );
  NOR2_X1 U13513 ( .A1(n10470), .A2(n10587), .ZN(n10588) );
  OR2_X1 U13514 ( .A1(n10589), .A2(n10588), .ZN(n18941) );
  NOR2_X1 U13515 ( .A1(n18941), .A2(n11175), .ZN(n15459) );
  INV_X1 U13516 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10805) );
  NOR2_X1 U13517 ( .A1(n10470), .A2(n10805), .ZN(n10616) );
  OR2_X2 U13518 ( .A1(n10617), .A2(n10616), .ZN(n10619) );
  INV_X1 U13519 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n13979) );
  NOR2_X1 U13520 ( .A1(n10470), .A2(n13979), .ZN(n10612) );
  NOR2_X2 U13521 ( .A1(n10619), .A2(n10612), .ZN(n10610) );
  NAND2_X1 U13522 ( .A1(n14236), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10608) );
  NAND2_X1 U13523 ( .A1(n10610), .A2(n10608), .ZN(n10604) );
  OR2_X2 U13524 ( .A1(n10604), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10605) );
  NAND2_X2 U13525 ( .A1(n10605), .A2(n10670), .ZN(n10623) );
  NAND2_X1 U13526 ( .A1(n14236), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10622) );
  NOR2_X1 U13527 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(P2_EBX_REG_18__SCAN_IN), 
        .ZN(n10590) );
  NOR2_X1 U13528 ( .A1(n10470), .A2(n10590), .ZN(n10591) );
  INV_X1 U13529 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n18859) );
  NAND2_X1 U13530 ( .A1(n14236), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10592) );
  NOR2_X1 U13531 ( .A1(n10629), .A2(n10592), .ZN(n10593) );
  OR2_X1 U13532 ( .A1(n18860), .A2(n11175), .ZN(n10594) );
  INV_X1 U13533 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15352) );
  NAND2_X1 U13534 ( .A1(n10594), .A2(n15352), .ZN(n12611) );
  NAND2_X1 U13535 ( .A1(n14236), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10595) );
  MUX2_X1 U13536 ( .A(n14236), .B(n10595), .S(n10625), .Z(n10596) );
  OR2_X1 U13537 ( .A1(n10625), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10599) );
  NAND2_X1 U13538 ( .A1(n10596), .A2(n10599), .ZN(n14935) );
  OR2_X1 U13539 ( .A1(n14935), .A2(n11175), .ZN(n10597) );
  INV_X1 U13540 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15392) );
  INV_X1 U13541 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n10827) );
  NOR2_X1 U13542 ( .A1(n10470), .A2(n10827), .ZN(n10598) );
  NAND2_X1 U13543 ( .A1(n10599), .A2(n10598), .ZN(n10600) );
  NAND2_X1 U13544 ( .A1(n10600), .A2(n10630), .ZN(n18872) );
  OR2_X1 U13545 ( .A1(n18872), .A2(n11175), .ZN(n10601) );
  INV_X1 U13546 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n20881) );
  NAND2_X1 U13547 ( .A1(n10601), .A2(n20881), .ZN(n15171) );
  INV_X1 U13548 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n18899) );
  NOR2_X1 U13549 ( .A1(n10470), .A2(n18899), .ZN(n10603) );
  INV_X1 U13550 ( .A(n10670), .ZN(n10602) );
  AOI21_X1 U13551 ( .B1(n10604), .B2(n10603), .A(n10602), .ZN(n10606) );
  NAND2_X1 U13552 ( .A1(n10606), .A2(n10605), .ZN(n18896) );
  OR2_X1 U13553 ( .A1(n18896), .A2(n11175), .ZN(n10607) );
  XNOR2_X1 U13554 ( .A(n10607), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12616) );
  INV_X1 U13555 ( .A(n10608), .ZN(n10609) );
  XNOR2_X1 U13556 ( .A(n10610), .B(n10609), .ZN(n18910) );
  NAND2_X1 U13557 ( .A1(n18910), .A2(n14239), .ZN(n10611) );
  INV_X1 U13558 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16267) );
  NAND2_X1 U13559 ( .A1(n10611), .A2(n16267), .ZN(n15206) );
  INV_X1 U13560 ( .A(n10612), .ZN(n10613) );
  XNOR2_X1 U13561 ( .A(n10619), .B(n10613), .ZN(n13981) );
  NAND2_X1 U13562 ( .A1(n13981), .A2(n14239), .ZN(n10614) );
  INV_X1 U13563 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16278) );
  NAND2_X1 U13564 ( .A1(n10614), .A2(n16278), .ZN(n16200) );
  NAND2_X1 U13565 ( .A1(n10615), .A2(n15432), .ZN(n15442) );
  NAND2_X1 U13566 ( .A1(n10617), .A2(n10616), .ZN(n10618) );
  NAND2_X1 U13567 ( .A1(n10619), .A2(n10618), .ZN(n18918) );
  OR2_X1 U13568 ( .A1(n18918), .A2(n11175), .ZN(n10621) );
  INV_X1 U13569 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10620) );
  NAND2_X1 U13570 ( .A1(n10621), .A2(n10620), .ZN(n15216) );
  AND4_X1 U13571 ( .A1(n15206), .A2(n16200), .A3(n15442), .A4(n15216), .ZN(
        n10627) );
  OR2_X1 U13572 ( .A1(n10623), .A2(n10622), .ZN(n10624) );
  AND2_X1 U13573 ( .A1(n10625), .A2(n10624), .ZN(n18880) );
  NAND2_X1 U13574 ( .A1(n18880), .A2(n14239), .ZN(n10626) );
  INV_X1 U13575 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15410) );
  NAND2_X1 U13576 ( .A1(n10626), .A2(n15410), .ZN(n12619) );
  NAND4_X1 U13577 ( .A1(n15171), .A2(n12616), .A3(n10627), .A4(n12619), .ZN(
        n10628) );
  NOR2_X1 U13578 ( .A1(n15177), .A2(n10628), .ZN(n10634) );
  INV_X1 U13579 ( .A(n10629), .ZN(n10633) );
  NAND2_X1 U13580 ( .A1(n14236), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10631) );
  MUX2_X1 U13581 ( .A(n14236), .B(n10631), .S(n10630), .Z(n10632) );
  NAND2_X1 U13582 ( .A1(n14927), .A2(n14239), .ZN(n10642) );
  INV_X1 U13583 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15364) );
  NAND2_X1 U13584 ( .A1(n10642), .A2(n15364), .ZN(n15158) );
  NAND3_X1 U13585 ( .A1(n12611), .A2(n10634), .A3(n15158), .ZN(n10635) );
  NAND2_X1 U13586 ( .A1(n14239), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10636) );
  OR2_X1 U13587 ( .A1(n18860), .A2(n10636), .ZN(n12610) );
  INV_X1 U13588 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n20859) );
  OR3_X1 U13589 ( .A1(n18896), .A2(n11175), .A3(n20859), .ZN(n12617) );
  AND2_X1 U13590 ( .A1(n14239), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10637) );
  NAND2_X1 U13591 ( .A1(n13981), .A2(n10637), .ZN(n16199) );
  NAND2_X1 U13592 ( .A1(n14239), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10638) );
  OR2_X1 U13593 ( .A1(n18918), .A2(n10638), .ZN(n15215) );
  AND3_X1 U13594 ( .A1(n12617), .A2(n16199), .A3(n15215), .ZN(n10641) );
  AND2_X1 U13595 ( .A1(n14239), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10639) );
  NAND2_X1 U13596 ( .A1(n18880), .A2(n10639), .ZN(n12618) );
  INV_X1 U13597 ( .A(n18910), .ZN(n10640) );
  INV_X1 U13598 ( .A(n10642), .ZN(n10643) );
  NAND2_X1 U13599 ( .A1(n14239), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10644) );
  NAND2_X1 U13600 ( .A1(n14239), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10645) );
  OR2_X1 U13601 ( .A1(n18872), .A2(n10645), .ZN(n15170) );
  NAND2_X1 U13602 ( .A1(n15178), .A2(n15170), .ZN(n12620) );
  NAND2_X1 U13603 ( .A1(n14236), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10648) );
  INV_X1 U13604 ( .A(n10648), .ZN(n10652) );
  INV_X1 U13605 ( .A(n10654), .ZN(n10650) );
  AOI21_X1 U13606 ( .B1(n10652), .B2(n10651), .A(n10650), .ZN(n15750) );
  AOI21_X1 U13607 ( .B1(n15750), .B2(n14239), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15328) );
  NAND3_X1 U13608 ( .A1(n15750), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n14239), .ZN(n15326) );
  INV_X1 U13609 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10839) );
  NOR2_X1 U13610 ( .A1(n10470), .A2(n10839), .ZN(n10655) );
  INV_X1 U13611 ( .A(n10661), .ZN(n10653) );
  AOI21_X1 U13612 ( .B1(n10655), .B2(n10654), .A(n10653), .ZN(n13028) );
  NAND2_X1 U13613 ( .A1(n13028), .A2(n14239), .ZN(n10656) );
  XNOR2_X1 U13614 ( .A(n10656), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15150) );
  INV_X1 U13615 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15315) );
  NOR2_X1 U13616 ( .A1(n11175), .A2(n15315), .ZN(n10657) );
  INV_X1 U13617 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10658) );
  NAND2_X1 U13618 ( .A1(n14236), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10659) );
  MUX2_X1 U13619 ( .A(P2_EBX_REG_24__SCAN_IN), .B(n10659), .S(n10661), .Z(
        n10660) );
  NAND2_X1 U13620 ( .A1(n10660), .A2(n10670), .ZN(n14906) );
  NOR2_X1 U13621 ( .A1(n14906), .A2(n11175), .ZN(n15140) );
  INV_X1 U13622 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14976) );
  INV_X1 U13623 ( .A(n10676), .ZN(n10662) );
  NAND2_X1 U13624 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n10672), .ZN(n10663) );
  NOR2_X1 U13625 ( .A1(n10470), .A2(n10663), .ZN(n10664) );
  NOR2_X1 U13626 ( .A1(n14234), .A2(n10664), .ZN(n16165) );
  INV_X1 U13627 ( .A(n16165), .ZN(n10665) );
  NOR2_X1 U13628 ( .A1(n10665), .A2(n11175), .ZN(n10666) );
  NAND3_X1 U13629 ( .A1(n16165), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14239), .ZN(n10688) );
  OAI21_X1 U13630 ( .B1(n10666), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n10688), .ZN(n15131) );
  NOR2_X1 U13631 ( .A1(n10667), .A2(n14976), .ZN(n10668) );
  NAND2_X1 U13632 ( .A1(n14236), .A2(n10668), .ZN(n10669) );
  AND2_X1 U13633 ( .A1(n10670), .A2(n10669), .ZN(n10671) );
  NAND2_X1 U13634 ( .A1(n10672), .A2(n10671), .ZN(n14898) );
  INV_X1 U13635 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15291) );
  NAND2_X1 U13636 ( .A1(n14236), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10677) );
  OR2_X1 U13637 ( .A1(n10677), .A2(n10676), .ZN(n10678) );
  NAND2_X1 U13638 ( .A1(n10680), .A2(n10678), .ZN(n13057) );
  INV_X1 U13639 ( .A(n10680), .ZN(n10682) );
  INV_X1 U13640 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n14877) );
  NOR2_X1 U13641 ( .A1(n10470), .A2(n14877), .ZN(n10679) );
  INV_X1 U13642 ( .A(n10679), .ZN(n10681) );
  OAI21_X1 U13643 ( .B1(n10682), .B2(n10681), .A(n10691), .ZN(n14880) );
  OAI21_X1 U13644 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n15111), .ZN(n10685) );
  INV_X1 U13645 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10684) );
  INV_X1 U13646 ( .A(n15111), .ZN(n10683) );
  INV_X1 U13647 ( .A(n10686), .ZN(n10687) );
  NAND2_X1 U13648 ( .A1(n10687), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15128) );
  NAND2_X1 U13649 ( .A1(n15128), .A2(n10688), .ZN(n15106) );
  INV_X1 U13650 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n10861) );
  NOR2_X1 U13651 ( .A1(n10470), .A2(n10861), .ZN(n10690) );
  AOI21_X1 U13652 ( .B1(n14861), .B2(n14239), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15095) );
  INV_X1 U13653 ( .A(n14861), .ZN(n10689) );
  INV_X1 U13654 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15099) );
  NOR2_X1 U13655 ( .A1(n14233), .A2(n15094), .ZN(n10695) );
  INV_X1 U13656 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n14201) );
  NOR2_X1 U13657 ( .A1(n10470), .A2(n14201), .ZN(n10692) );
  XNOR2_X1 U13658 ( .A(n14235), .B(n10692), .ZN(n14208) );
  NAND2_X1 U13659 ( .A1(n14239), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10693) );
  INV_X1 U13660 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11180) );
  OAI21_X1 U13661 ( .B1(n14208), .B2(n11175), .A(n11180), .ZN(n14232) );
  NAND2_X1 U13662 ( .A1(n9632), .A2(n14232), .ZN(n10694) );
  XNOR2_X1 U13663 ( .A(n10695), .B(n10694), .ZN(n15093) );
  INV_X1 U13664 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15824) );
  NOR2_X1 U13665 ( .A1(n15824), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10696) );
  INV_X1 U13666 ( .A(n10734), .ZN(n10728) );
  NAND2_X1 U13667 ( .A1(n10698), .A2(n13037), .ZN(n10699) );
  MUX2_X1 U13668 ( .A(n10699), .B(n13035), .S(n10731), .Z(n10711) );
  INV_X1 U13669 ( .A(n10731), .ZN(n10709) );
  OAI21_X1 U13670 ( .B1(n10737), .B2(n10703), .A(n10701), .ZN(n10708) );
  INV_X1 U13671 ( .A(n10737), .ZN(n10706) );
  NAND2_X1 U13672 ( .A1(n10703), .A2(n10702), .ZN(n10719) );
  NAND2_X1 U13673 ( .A1(n10704), .A2(n10719), .ZN(n10732) );
  INV_X1 U13674 ( .A(n10732), .ZN(n10705) );
  OAI211_X1 U13675 ( .C1(n19196), .C2(n10706), .A(n16322), .B(n10705), .ZN(
        n10707) );
  OAI211_X1 U13676 ( .C1(n10880), .C2(n10709), .A(n10708), .B(n10707), .ZN(
        n10710) );
  NAND2_X1 U13677 ( .A1(n10711), .A2(n10710), .ZN(n10714) );
  MUX2_X1 U13678 ( .A(n13035), .B(n10714), .S(n10730), .Z(n10715) );
  NAND2_X1 U13679 ( .A1(n10728), .A2(n10715), .ZN(n10716) );
  MUX2_X1 U13680 ( .A(n10716), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18828), .Z(n10760) );
  NAND2_X1 U13681 ( .A1(n10734), .A2(n13273), .ZN(n10717) );
  NAND2_X1 U13682 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19711) );
  INV_X1 U13683 ( .A(n19711), .ZN(n19865) );
  NAND2_X1 U13684 ( .A1(n19728), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19869) );
  INV_X2 U13685 ( .A(n19869), .ZN(n19868) );
  NAND2_X2 U13686 ( .A1(n19868), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19790) );
  NOR2_X1 U13687 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19723) );
  INV_X1 U13688 ( .A(n19723), .ZN(n19733) );
  NAND3_X1 U13689 ( .A1(n19728), .A2(n19790), .A3(n19733), .ZN(n19727) );
  NOR2_X1 U13690 ( .A1(n19865), .A2(n19727), .ZN(n16316) );
  NAND3_X1 U13691 ( .A1(n13269), .A2(n16316), .A3(n10718), .ZN(n10765) );
  INV_X1 U13692 ( .A(n10719), .ZN(n10722) );
  INV_X1 U13693 ( .A(n10720), .ZN(n10721) );
  OAI21_X1 U13694 ( .B1(n10723), .B2(n10722), .A(n10721), .ZN(n10727) );
  INV_X1 U13695 ( .A(n10724), .ZN(n10726) );
  NAND3_X1 U13696 ( .A1(n10727), .A2(n10726), .A3(n10725), .ZN(n10729) );
  AND2_X1 U13697 ( .A1(n10729), .A2(n10728), .ZN(n19841) );
  NAND2_X1 U13698 ( .A1(n19853), .A2(n19852), .ZN(n19851) );
  NOR2_X1 U13699 ( .A1(n16321), .A2(n19851), .ZN(n19844) );
  NAND2_X1 U13700 ( .A1(n10731), .A2(n10730), .ZN(n10736) );
  NOR2_X1 U13701 ( .A1(n10732), .A2(n10736), .ZN(n10733) );
  OR2_X1 U13702 ( .A1(n10734), .A2(n10733), .ZN(n16310) );
  INV_X1 U13703 ( .A(n16310), .ZN(n10735) );
  OAI21_X1 U13704 ( .B1(n10737), .B2(n10736), .A(n10735), .ZN(n10738) );
  INV_X1 U13705 ( .A(n10738), .ZN(n10741) );
  NAND2_X1 U13706 ( .A1(n10739), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10740) );
  NAND2_X1 U13707 ( .A1(n10740), .A2(n16308), .ZN(n13169) );
  INV_X1 U13708 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n18833) );
  OAI21_X1 U13709 ( .B1(n10389), .B2(n13169), .A(n18833), .ZN(n19833) );
  MUX2_X1 U13710 ( .A(n10741), .B(n19833), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n16346) );
  NAND2_X1 U13711 ( .A1(n16346), .A2(n13037), .ZN(n10742) );
  NOR2_X1 U13712 ( .A1(n16321), .A2(n10742), .ZN(n10743) );
  AOI21_X1 U13713 ( .B1(n19841), .B2(n19844), .A(n10743), .ZN(n12626) );
  NAND2_X1 U13714 ( .A1(n10744), .A2(n16316), .ZN(n10745) );
  OR2_X1 U13715 ( .A1(n16310), .A2(n10745), .ZN(n10756) );
  OAI21_X1 U13716 ( .B1(n19206), .B2(n13037), .A(n16322), .ZN(n10746) );
  AOI21_X1 U13717 ( .B1(n10746), .B2(n9583), .A(n10718), .ZN(n10747) );
  NOR2_X1 U13718 ( .A1(n10747), .A2(n10892), .ZN(n10753) );
  NAND2_X1 U13719 ( .A1(n10749), .A2(n10874), .ZN(n10750) );
  NAND2_X1 U13720 ( .A1(n10748), .A2(n10750), .ZN(n10752) );
  INV_X1 U13721 ( .A(n19851), .ZN(n10751) );
  AND4_X1 U13722 ( .A1(n10754), .A2(n10753), .A3(n10752), .A4(n10878), .ZN(
        n10755) );
  NAND2_X1 U13723 ( .A1(n10756), .A2(n10755), .ZN(n13161) );
  MUX2_X1 U13724 ( .A(n10744), .B(n10718), .S(n19853), .Z(n10757) );
  NAND2_X1 U13725 ( .A1(n10757), .A2(n19711), .ZN(n10758) );
  NOR2_X1 U13726 ( .A1(n16310), .A2(n10758), .ZN(n10759) );
  NOR2_X1 U13727 ( .A1(n13161), .A2(n10759), .ZN(n10764) );
  INV_X1 U13728 ( .A(n13269), .ZN(n10762) );
  AOI21_X1 U13729 ( .B1(n10760), .B2(n16322), .A(n19206), .ZN(n10761) );
  NAND2_X1 U13730 ( .A1(n10762), .A2(n10761), .ZN(n10763) );
  NAND4_X1 U13731 ( .A1(n10765), .A2(n12626), .A3(n10764), .A4(n10763), .ZN(
        n10766) );
  NAND3_X1 U13732 ( .A1(n19712), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n19714) );
  NOR2_X1 U13733 ( .A1(n16321), .A2(n13035), .ZN(n19842) );
  INV_X1 U13734 ( .A(n10767), .ZN(n10768) );
  NAND2_X1 U13735 ( .A1(n10771), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10773) );
  AOI22_X1 U13736 ( .A1(n14242), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10772) );
  OAI211_X1 U13737 ( .C1(n10774), .C2(n10856), .A(n10773), .B(n10772), .ZN(
        n13521) );
  NAND2_X1 U13738 ( .A1(n13522), .A2(n13521), .ZN(n13541) );
  NAND2_X1 U13739 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10776) );
  NAND2_X1 U13740 ( .A1(n10858), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n10775) );
  OAI211_X1 U13741 ( .C1(n10856), .C2(n18994), .A(n10776), .B(n10775), .ZN(
        n10777) );
  AOI21_X1 U13742 ( .B1(n10771), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n10777), .ZN(n13542) );
  NAND2_X1 U13743 ( .A1(n10771), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10783) );
  INV_X1 U13744 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n10780) );
  NAND2_X1 U13745 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10779) );
  NAND2_X1 U13746 ( .A1(n10862), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n10778) );
  OAI211_X1 U13747 ( .C1(n10856), .C2(n10780), .A(n10779), .B(n10778), .ZN(
        n10781) );
  INV_X1 U13748 ( .A(n10781), .ZN(n10782) );
  NAND2_X1 U13749 ( .A1(n10783), .A2(n10782), .ZN(n13597) );
  NAND2_X1 U13750 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10785) );
  NAND2_X1 U13751 ( .A1(n14242), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n10784) );
  OAI211_X1 U13752 ( .C1(n10856), .C2(n10786), .A(n10785), .B(n10784), .ZN(
        n10787) );
  AOI21_X1 U13753 ( .B1(n10771), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n10787), .ZN(n13604) );
  INV_X1 U13754 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n13855) );
  NAND2_X1 U13755 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10789) );
  NAND2_X1 U13756 ( .A1(n10858), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10788) );
  OAI211_X1 U13757 ( .C1(n10856), .C2(n13855), .A(n10789), .B(n10788), .ZN(
        n10790) );
  AOI21_X1 U13758 ( .B1(n10771), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n10790), .ZN(n13632) );
  INV_X1 U13759 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10793) );
  NAND2_X1 U13760 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10792) );
  NAND2_X1 U13761 ( .A1(n10862), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10791) );
  OAI211_X1 U13762 ( .C1(n10856), .C2(n10793), .A(n10792), .B(n10791), .ZN(
        n10794) );
  AOI21_X1 U13763 ( .B1(n10771), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n10794), .ZN(n13641) );
  INV_X1 U13764 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13660) );
  NAND2_X1 U13765 ( .A1(n10771), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10796) );
  AOI22_X1 U13766 ( .A1(n14242), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10795) );
  OAI211_X1 U13767 ( .C1(n13660), .C2(n10856), .A(n10796), .B(n10795), .ZN(
        n13655) );
  NAND2_X1 U13768 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10798) );
  NAND2_X1 U13769 ( .A1(n10858), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n10797) );
  OAI211_X1 U13770 ( .C1(n10856), .C2(n18944), .A(n10798), .B(n10797), .ZN(
        n10799) );
  AOI21_X1 U13771 ( .B1(n10771), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n10799), .ZN(n13684) );
  INV_X1 U13772 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n10802) );
  NAND2_X1 U13773 ( .A1(n10771), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10801) );
  AOI22_X1 U13774 ( .A1(n10862), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n10800) );
  OAI211_X1 U13775 ( .C1(n10802), .C2(n10856), .A(n10801), .B(n10800), .ZN(
        n13708) );
  NAND2_X1 U13776 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10804) );
  NAND2_X1 U13777 ( .A1(n14242), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n10803) );
  OAI211_X1 U13778 ( .C1(n10856), .C2(n10805), .A(n10804), .B(n10803), .ZN(
        n10806) );
  AOI21_X1 U13779 ( .B1(n10771), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n10806), .ZN(n13754) );
  NAND2_X1 U13780 ( .A1(n10771), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10811) );
  NAND2_X1 U13781 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10808) );
  NAND2_X1 U13782 ( .A1(n10858), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n10807) );
  OAI211_X1 U13783 ( .C1(n10856), .C2(n13979), .A(n10808), .B(n10807), .ZN(
        n10809) );
  INV_X1 U13784 ( .A(n10809), .ZN(n10810) );
  NAND2_X1 U13785 ( .A1(n10811), .A2(n10810), .ZN(n13834) );
  NAND2_X1 U13786 ( .A1(n13833), .A2(n13834), .ZN(n13958) );
  INV_X1 U13787 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10814) );
  NAND2_X1 U13788 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10813) );
  NAND2_X1 U13789 ( .A1(n10862), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n10812) );
  OAI211_X1 U13790 ( .C1(n10856), .C2(n10814), .A(n10813), .B(n10812), .ZN(
        n10815) );
  AOI21_X1 U13791 ( .B1(n10771), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n10815), .ZN(n13957) );
  NAND2_X1 U13792 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10817) );
  NAND2_X1 U13793 ( .A1(n14242), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10816) );
  OAI211_X1 U13794 ( .C1(n10856), .C2(n18899), .A(n10817), .B(n10816), .ZN(
        n10818) );
  AOI21_X1 U13795 ( .B1(n10771), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10818), .ZN(n13997) );
  INV_X1 U13796 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10821) );
  NAND2_X1 U13797 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10820) );
  NAND2_X1 U13798 ( .A1(n10858), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n10819) );
  OAI211_X1 U13799 ( .C1(n10856), .C2(n10821), .A(n10820), .B(n10819), .ZN(
        n10822) );
  AOI21_X1 U13800 ( .B1(n10771), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10822), .ZN(n15023) );
  INV_X1 U13801 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n14941) );
  NAND2_X1 U13802 ( .A1(n10771), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10824) );
  AOI22_X1 U13803 ( .A1(n10862), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n10823) );
  OAI211_X1 U13804 ( .C1(n10856), .C2(n14941), .A(n10824), .B(n10823), .ZN(
        n14936) );
  NAND2_X1 U13805 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10826) );
  NAND2_X1 U13806 ( .A1(n14242), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n10825) );
  OAI211_X1 U13807 ( .C1(n10856), .C2(n10827), .A(n10826), .B(n10825), .ZN(
        n10828) );
  AOI21_X1 U13808 ( .B1(n10771), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n10828), .ZN(n15010) );
  INV_X1 U13809 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10831) );
  NAND2_X1 U13810 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10830) );
  NAND2_X1 U13811 ( .A1(n10858), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n10829) );
  OAI211_X1 U13812 ( .C1(n10856), .C2(n10831), .A(n10830), .B(n10829), .ZN(
        n10832) );
  AOI21_X1 U13813 ( .B1(n10771), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n10832), .ZN(n14921) );
  NAND2_X1 U13814 ( .A1(n10771), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10834) );
  AOI22_X1 U13815 ( .A1(n10862), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n10833) );
  OAI211_X1 U13816 ( .C1(n10856), .C2(n18859), .A(n10834), .B(n10833), .ZN(
        n12634) );
  INV_X1 U13817 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15752) );
  NAND2_X1 U13818 ( .A1(n10771), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10836) );
  AOI22_X1 U13819 ( .A1(n14242), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n10835) );
  OAI211_X1 U13820 ( .C1(n10856), .C2(n15752), .A(n10836), .B(n10835), .ZN(
        n14992) );
  NAND2_X1 U13821 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10838) );
  NAND2_X1 U13822 ( .A1(n10858), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n10837) );
  OAI211_X1 U13823 ( .C1(n10856), .C2(n10839), .A(n10838), .B(n10837), .ZN(
        n10840) );
  AOI21_X1 U13824 ( .B1(n10771), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n10840), .ZN(n13032) );
  INV_X1 U13825 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n14983) );
  NAND2_X1 U13826 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10842) );
  NAND2_X1 U13827 ( .A1(n10862), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n10841) );
  OAI211_X1 U13828 ( .C1(n10856), .C2(n14983), .A(n10842), .B(n10841), .ZN(
        n10843) );
  AOI21_X1 U13829 ( .B1(n10771), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n10843), .ZN(n14902) );
  NAND2_X1 U13830 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10845) );
  NAND2_X1 U13831 ( .A1(n14242), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n10844) );
  OAI211_X1 U13832 ( .C1(n10856), .C2(n14976), .A(n10845), .B(n10844), .ZN(
        n10846) );
  AOI21_X1 U13833 ( .B1(n10771), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n10846), .ZN(n14212) );
  INV_X1 U13834 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n10849) );
  NAND2_X1 U13835 ( .A1(n10771), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10848) );
  AOI22_X1 U13836 ( .A1(n10858), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n10847) );
  OAI211_X1 U13837 ( .C1(n10856), .C2(n10849), .A(n10848), .B(n10847), .ZN(
        n14964) );
  INV_X1 U13838 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n10852) );
  NAND2_X1 U13839 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10851) );
  NAND2_X1 U13840 ( .A1(n10862), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n10850) );
  OAI211_X1 U13841 ( .C1(n10856), .C2(n10852), .A(n10851), .B(n10850), .ZN(
        n10853) );
  AOI21_X1 U13842 ( .B1(n10771), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10853), .ZN(n13058) );
  NAND2_X1 U13843 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10855) );
  NAND2_X1 U13844 ( .A1(n14242), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n10854) );
  OAI211_X1 U13845 ( .C1(n10856), .C2(n14877), .A(n10855), .B(n10854), .ZN(
        n10857) );
  AOI21_X1 U13846 ( .B1(n10771), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n10857), .ZN(n14871) );
  NAND2_X1 U13847 ( .A1(n10771), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10860) );
  AOI22_X1 U13848 ( .A1(n10858), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10859) );
  OAI211_X1 U13849 ( .C1(n10856), .C2(n10861), .A(n10860), .B(n10859), .ZN(
        n14858) );
  NAND2_X1 U13850 ( .A1(n10771), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10864) );
  AOI22_X1 U13851 ( .A1(n10862), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n10863) );
  OAI211_X1 U13852 ( .C1(n10856), .C2(n14201), .A(n10864), .B(n10863), .ZN(
        n10865) );
  INV_X1 U13853 ( .A(n14003), .ZN(n10870) );
  NAND2_X1 U13854 ( .A1(n10868), .A2(n12416), .ZN(n10869) );
  NAND2_X1 U13855 ( .A1(n10870), .A2(n10869), .ZN(n10871) );
  NAND2_X1 U13856 ( .A1(n11181), .A2(n10871), .ZN(n16295) );
  NAND2_X1 U13857 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15449) );
  NAND2_X1 U13858 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16277) );
  INV_X1 U13859 ( .A(n16277), .ZN(n15349) );
  NAND3_X1 U13860 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n15349), .ZN(n10872) );
  NOR2_X1 U13861 ( .A1(n15449), .A2(n10872), .ZN(n15385) );
  NAND3_X1 U13862 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15386) );
  NOR2_X1 U13863 ( .A1(n15392), .A2(n15386), .ZN(n15351) );
  AND2_X1 U13864 ( .A1(n15385), .A2(n15351), .ZN(n15366) );
  AND3_X1 U13865 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10873) );
  AND2_X1 U13866 ( .A1(n15366), .A2(n10873), .ZN(n11178) );
  INV_X1 U13867 ( .A(n11178), .ZN(n11130) );
  NAND2_X1 U13868 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15531) );
  INV_X1 U13869 ( .A(n15531), .ZN(n15558) );
  NAND2_X1 U13870 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15558), .ZN(
        n11122) );
  AND3_X1 U13871 ( .A1(n12416), .A2(n10874), .A3(n10470), .ZN(n10875) );
  AND2_X1 U13872 ( .A1(n13934), .A2(n10875), .ZN(n16309) );
  NAND2_X1 U13873 ( .A1(n11181), .A2(n16309), .ZN(n13277) );
  NAND2_X1 U13874 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15571) );
  INV_X1 U13875 ( .A(n15571), .ZN(n13293) );
  NAND2_X1 U13876 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13293), .ZN(
        n10876) );
  NOR2_X1 U13877 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13293), .ZN(
        n11123) );
  AOI21_X1 U13878 ( .B1(n13277), .B2(n10876), .A(n11123), .ZN(n10896) );
  NAND2_X1 U13879 ( .A1(n10877), .A2(n13037), .ZN(n13933) );
  NAND2_X1 U13880 ( .A1(n13933), .A2(n10878), .ZN(n10888) );
  NOR2_X1 U13881 ( .A1(n10880), .A2(n10879), .ZN(n10882) );
  NAND2_X1 U13882 ( .A1(n10882), .A2(n10881), .ZN(n12589) );
  INV_X1 U13883 ( .A(n12587), .ZN(n13118) );
  OAI21_X1 U13884 ( .B1(n10892), .B2(n10883), .A(n13118), .ZN(n10885) );
  NAND2_X1 U13885 ( .A1(n19852), .A2(n10718), .ZN(n10884) );
  NAND4_X1 U13886 ( .A1(n10886), .A2(n12589), .A3(n10885), .A4(n10884), .ZN(
        n10887) );
  AOI21_X1 U13887 ( .B1(n10889), .B2(n10888), .A(n10887), .ZN(n10894) );
  NAND3_X1 U13888 ( .A1(n10890), .A2(n10892), .A3(n10891), .ZN(n10893) );
  AND2_X1 U13889 ( .A1(n10894), .A2(n10893), .ZN(n13932) );
  INV_X1 U13890 ( .A(n14002), .ZN(n12957) );
  NAND2_X1 U13891 ( .A1(n13932), .A2(n12957), .ZN(n10895) );
  NAND2_X1 U13892 ( .A1(n11181), .A2(n10895), .ZN(n15400) );
  NAND2_X1 U13893 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13884), .ZN(
        n15557) );
  NOR2_X1 U13894 ( .A1(n11122), .A2(n15557), .ZN(n15521) );
  NAND3_X1 U13895 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n15521), .ZN(n15482) );
  NOR2_X1 U13896 ( .A1(n11130), .A2(n15482), .ZN(n15337) );
  INV_X1 U13897 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15342) );
  NOR2_X1 U13898 ( .A1(n15315), .A2(n15342), .ZN(n15314) );
  AND2_X1 U13899 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15314), .ZN(
        n10897) );
  AND2_X1 U13900 ( .A1(n15337), .A2(n10897), .ZN(n15288) );
  NAND2_X1 U13901 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11179) );
  INV_X1 U13902 ( .A(n11179), .ZN(n15290) );
  NAND2_X1 U13903 ( .A1(n15288), .A2(n15290), .ZN(n15252) );
  INV_X1 U13904 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15253) );
  OR2_X1 U13905 ( .A1(n15252), .A2(n15253), .ZN(n15268) );
  NAND2_X1 U13906 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10898) );
  NOR2_X1 U13907 ( .A1(n15268), .A2(n10898), .ZN(n14254) );
  NOR2_X2 U13908 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19802) );
  NAND2_X1 U13909 ( .A1(n19802), .A2(n19712), .ZN(n18827) );
  INV_X1 U13910 ( .A(n18827), .ZN(n13116) );
  NAND2_X1 U13911 ( .A1(n13116), .A2(n18828), .ZN(n18992) );
  INV_X2 U13912 ( .A(n18992), .ZN(n19155) );
  INV_X1 U13913 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n10899) );
  NOR2_X1 U13914 ( .A1(n16264), .A2(n10899), .ZN(n15086) );
  AOI21_X1 U13915 ( .B1(n14254), .B2(n11180), .A(n15086), .ZN(n11121) );
  AND2_X2 U13916 ( .A1(n10194), .A2(n10902), .ZN(n10910) );
  NOR2_X1 U13917 ( .A1(n9583), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10911) );
  AOI222_X1 U13918 ( .A1(n10910), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n14248), 
        .B2(P2_EAX_REG_30__SCAN_IN), .C1(n10944), .C2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11114) );
  MUX2_X1 U13919 ( .A(n9583), .B(n19837), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10901) );
  INV_X1 U13920 ( .A(n10182), .ZN(n12591) );
  NAND2_X1 U13921 ( .A1(n12591), .A2(n10944), .ZN(n10919) );
  AND2_X1 U13922 ( .A1(n10901), .A2(n10919), .ZN(n10905) );
  INV_X1 U13923 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18848) );
  NAND2_X1 U13924 ( .A1(n10910), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10909) );
  INV_X1 U13925 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13263) );
  NAND2_X1 U13926 ( .A1(n19196), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10906) );
  OAI211_X1 U13927 ( .C1(n9584), .C2(n13263), .A(n10906), .B(n10900), .ZN(
        n10907) );
  INV_X1 U13928 ( .A(n10907), .ZN(n10908) );
  NAND2_X1 U13929 ( .A1(n10909), .A2(n10908), .ZN(n13258) );
  INV_X1 U13930 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19740) );
  NAND2_X1 U13931 ( .A1(n10910), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10913) );
  AOI22_X1 U13932 ( .A1(n10911), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n10944), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10912) );
  NAND2_X1 U13933 ( .A1(n10913), .A2(n10912), .ZN(n10916) );
  XNOR2_X1 U13934 ( .A(n13256), .B(n10916), .ZN(n13550) );
  NAND2_X1 U13935 ( .A1(n10182), .A2(n9584), .ZN(n10914) );
  MUX2_X1 U13936 ( .A(n10914), .B(n19828), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10915) );
  OAI21_X1 U13937 ( .B1(n11141), .B2(n11063), .A(n10915), .ZN(n13549) );
  NOR2_X1 U13938 ( .A1(n13550), .A2(n13549), .ZN(n10918) );
  NOR2_X1 U13939 ( .A1(n13256), .A2(n10916), .ZN(n10917) );
  NAND2_X1 U13940 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10920) );
  OAI211_X1 U13941 ( .C1(n11063), .C2(n11139), .A(n10920), .B(n10919), .ZN(
        n10923) );
  XNOR2_X1 U13942 ( .A(n10924), .B(n10923), .ZN(n13280) );
  NAND2_X1 U13943 ( .A1(n10910), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U13944 ( .A1(n14248), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n10944), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10921) );
  NAND2_X1 U13945 ( .A1(n10922), .A2(n10921), .ZN(n13279) );
  NOR2_X1 U13946 ( .A1(n13280), .A2(n13279), .ZN(n13281) );
  NOR2_X1 U13947 ( .A1(n10924), .A2(n10923), .ZN(n10925) );
  NAND2_X1 U13948 ( .A1(n10910), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10930) );
  AOI22_X1 U13949 ( .A1(n10944), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n10929) );
  OR2_X1 U13950 ( .A1(n11063), .A2(n10926), .ZN(n10928) );
  NAND2_X1 U13951 ( .A1(n14248), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10927) );
  NAND4_X1 U13952 ( .A1(n10930), .A2(n10929), .A3(n10928), .A4(n10927), .ZN(
        n13825) );
  NAND2_X1 U13953 ( .A1(n10910), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U13954 ( .A1(n14248), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n10944), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10933) );
  INV_X1 U13955 ( .A(n10931), .ZN(n11149) );
  OR2_X1 U13956 ( .A1(n11063), .A2(n11149), .ZN(n10932) );
  AOI22_X1 U13957 ( .A1(n10904), .A2(n10935), .B1(n10910), .B2(
        P2_REIP_REG_5__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U13958 ( .A1(n14248), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n10944), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10936) );
  NAND2_X1 U13959 ( .A1(n10937), .A2(n10936), .ZN(n15555) );
  OR2_X1 U13960 ( .A1(n11063), .A2(n10938), .ZN(n10939) );
  NAND2_X1 U13961 ( .A1(n10910), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U13962 ( .A1(n14248), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n10944), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10940) );
  NAND2_X1 U13963 ( .A1(n10941), .A2(n10940), .ZN(n15532) );
  NAND2_X1 U13964 ( .A1(n15533), .A2(n15532), .ZN(n10943) );
  OR2_X1 U13965 ( .A1(n11063), .A2(n11175), .ZN(n10942) );
  NAND2_X1 U13966 ( .A1(n10910), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n10946) );
  AOI22_X1 U13967 ( .A1(n14248), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n10944), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10945) );
  NAND2_X1 U13968 ( .A1(n10946), .A2(n10945), .ZN(n15516) );
  INV_X1 U13969 ( .A(n12387), .ZN(n10962) );
  AOI22_X1 U13970 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10950) );
  AOI22_X1 U13971 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10949) );
  AOI22_X1 U13972 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10948) );
  AOI22_X1 U13973 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12394), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10947) );
  NAND4_X1 U13974 ( .A1(n10950), .A2(n10949), .A3(n10948), .A4(n10947), .ZN(
        n10959) );
  AOI22_X1 U13975 ( .A1(n10341), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10957) );
  INV_X1 U13976 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10952) );
  INV_X1 U13977 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10951) );
  OAI22_X1 U13978 ( .A1(n12367), .A2(n10952), .B1(n12364), .B2(n10951), .ZN(
        n10953) );
  AOI21_X1 U13979 ( .B1(n10376), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A(
        n10953), .ZN(n10956) );
  AOI22_X1 U13980 ( .A1(n11071), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10955) );
  NAND2_X1 U13981 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10954) );
  NAND4_X1 U13982 ( .A1(n10957), .A2(n10956), .A3(n10955), .A4(n10954), .ZN(
        n10958) );
  NOR2_X1 U13983 ( .A1(n10959), .A2(n10958), .ZN(n13636) );
  AOI22_X1 U13984 ( .A1(n14248), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n10944), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10960) );
  OAI21_X1 U13985 ( .B1(n13636), .B2(n11063), .A(n10960), .ZN(n10961) );
  AOI21_X1 U13986 ( .B1(n10910), .B2(P2_REIP_REG_8__SCAN_IN), .A(n10961), .ZN(
        n13853) );
  AOI22_X1 U13987 ( .A1(n10910), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n14248), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n10978) );
  AOI22_X1 U13988 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10966) );
  AOI22_X1 U13989 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10965) );
  AOI22_X1 U13990 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10964) );
  AOI22_X1 U13991 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12394), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10963) );
  NAND4_X1 U13992 ( .A1(n10966), .A2(n10965), .A3(n10964), .A4(n10963), .ZN(
        n10974) );
  AOI22_X1 U13993 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10341), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10972) );
  INV_X1 U13994 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12431) );
  OAI22_X1 U13995 ( .A1(n12367), .A2(n10967), .B1(n12431), .B2(n12364), .ZN(
        n10968) );
  AOI21_X1 U13996 ( .B1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n10376), .A(
        n10968), .ZN(n10971) );
  AOI22_X1 U13997 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11071), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10970) );
  NAND2_X1 U13998 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10969) );
  NAND4_X1 U13999 ( .A1(n10972), .A2(n10971), .A3(n10970), .A4(n10969), .ZN(
        n10973) );
  OR2_X1 U14000 ( .A1(n10974), .A2(n10973), .ZN(n12270) );
  INV_X1 U14001 ( .A(n12270), .ZN(n13652) );
  OAI22_X1 U14002 ( .A1(n11063), .A2(n13652), .B1(n10975), .B2(n15486), .ZN(
        n10976) );
  INV_X1 U14003 ( .A(n10976), .ZN(n10977) );
  NAND2_X1 U14004 ( .A1(n10978), .A2(n10977), .ZN(n15480) );
  NAND2_X1 U14005 ( .A1(n10910), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n10999) );
  AOI22_X1 U14006 ( .A1(n14248), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U14007 ( .A1(n11071), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__2__SCAN_IN), .B2(n12375), .ZN(n10982) );
  AOI22_X1 U14008 ( .A1(n11072), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n9567), .ZN(n10981) );
  NAND2_X1 U14009 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10980) );
  NAND2_X1 U14010 ( .A1(n10376), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10979) );
  NAND4_X1 U14011 ( .A1(n10982), .A2(n10981), .A3(n10980), .A4(n10979), .ZN(
        n10986) );
  INV_X1 U14012 ( .A(n10389), .ZN(n11057) );
  INV_X1 U14013 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10984) );
  OAI22_X1 U14014 ( .A1(n11057), .A2(n10984), .B1(n10538), .B2(n10983), .ZN(
        n10985) );
  NOR2_X1 U14015 ( .A1(n10986), .A2(n10985), .ZN(n10996) );
  INV_X1 U14016 ( .A(n10987), .ZN(n12387) );
  INV_X1 U14017 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10988) );
  INV_X1 U14018 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12450) );
  OAI22_X1 U14019 ( .A1(n12387), .A2(n10988), .B1(n12389), .B2(n12450), .ZN(
        n10992) );
  INV_X1 U14020 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10990) );
  INV_X1 U14021 ( .A(n12394), .ZN(n15595) );
  INV_X1 U14022 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10989) );
  OAI22_X1 U14023 ( .A1(n10990), .A2(n15595), .B1(n10537), .B2(n10989), .ZN(
        n10991) );
  NOR2_X1 U14024 ( .A1(n10992), .A2(n10991), .ZN(n10995) );
  AOI22_X1 U14025 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10341), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U14026 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10993) );
  NAND4_X1 U14027 ( .A1(n10996), .A2(n10995), .A3(n10994), .A4(n10993), .ZN(
        n12271) );
  INV_X1 U14028 ( .A(n12271), .ZN(n13651) );
  OR2_X1 U14029 ( .A1(n11063), .A2(n13651), .ZN(n10997) );
  AOI22_X1 U14030 ( .A1(n10910), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n14248), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n11013) );
  AOI22_X1 U14031 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11003) );
  AOI22_X1 U14032 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11002) );
  AOI22_X1 U14033 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11001) );
  AOI22_X1 U14034 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11000) );
  NAND4_X1 U14035 ( .A1(n11003), .A2(n11002), .A3(n11001), .A4(n11000), .ZN(
        n11011) );
  AOI22_X1 U14036 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10341), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11009) );
  INV_X1 U14037 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12484) );
  OAI22_X1 U14038 ( .A1(n12367), .A2(n11004), .B1(n12364), .B2(n12484), .ZN(
        n11005) );
  AOI21_X1 U14039 ( .B1(n10376), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n11005), .ZN(n11008) );
  AOI22_X1 U14040 ( .A1(n11071), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11007) );
  NAND2_X1 U14041 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11006) );
  NAND4_X1 U14042 ( .A1(n11009), .A2(n11008), .A3(n11007), .A4(n11006), .ZN(
        n11010) );
  OR2_X1 U14043 ( .A1(n11011), .A2(n11010), .ZN(n13682) );
  AOI22_X1 U14044 ( .A1(n10904), .A2(n13682), .B1(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n10944), .ZN(n11012) );
  NAND2_X1 U14045 ( .A1(n11013), .A2(n11012), .ZN(n15454) );
  NAND2_X1 U14046 ( .A1(n15455), .A2(n15454), .ZN(n15453) );
  INV_X1 U14047 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11015) );
  INV_X1 U14048 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11014) );
  OAI22_X1 U14049 ( .A1(n11057), .A2(n11015), .B1(n10537), .B2(n11014), .ZN(
        n11018) );
  INV_X1 U14050 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11016) );
  INV_X1 U14051 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12500) );
  OAI22_X1 U14052 ( .A1(n12387), .A2(n11016), .B1(n12389), .B2(n12500), .ZN(
        n11017) );
  NOR2_X1 U14053 ( .A1(n11018), .A2(n11017), .ZN(n11029) );
  AOI22_X1 U14054 ( .A1(n11071), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12375), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U14055 ( .A1(n11072), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9567), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11021) );
  NAND2_X1 U14056 ( .A1(n10376), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11020) );
  NAND2_X1 U14057 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11019) );
  NAND4_X1 U14058 ( .A1(n11022), .A2(n11021), .A3(n11020), .A4(n11019), .ZN(
        n11025) );
  INV_X1 U14059 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12498) );
  OAI22_X1 U14060 ( .A1(n11055), .A2(n12498), .B1(n10538), .B2(n11023), .ZN(
        n11024) );
  NOR2_X1 U14061 ( .A1(n11025), .A2(n11024), .ZN(n11028) );
  AOI22_X1 U14062 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10422), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U14063 ( .A1(n12383), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12394), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11026) );
  NAND4_X1 U14064 ( .A1(n11029), .A2(n11028), .A3(n11027), .A4(n11026), .ZN(
        n12269) );
  INV_X1 U14065 ( .A(n12269), .ZN(n13712) );
  AOI22_X1 U14066 ( .A1(n14248), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11030) );
  OAI21_X1 U14067 ( .B1(n13712), .B2(n11063), .A(n11030), .ZN(n11031) );
  AOI21_X1 U14068 ( .B1(n10910), .B2(P2_REIP_REG_12__SCAN_IN), .A(n11031), 
        .ZN(n15436) );
  AOI22_X1 U14069 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11035) );
  AOI22_X1 U14070 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11034) );
  AOI22_X1 U14071 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11033) );
  AOI22_X1 U14072 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11032) );
  NAND4_X1 U14073 ( .A1(n11035), .A2(n11034), .A3(n11033), .A4(n11032), .ZN(
        n11043) );
  AOI22_X1 U14074 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10341), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11041) );
  INV_X1 U14075 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12531) );
  OAI22_X1 U14076 ( .A1(n12367), .A2(n11036), .B1(n12364), .B2(n12531), .ZN(
        n11037) );
  AOI21_X1 U14077 ( .B1(n10376), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n11037), .ZN(n11040) );
  AOI22_X1 U14078 ( .A1(n11071), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11039) );
  NAND2_X1 U14079 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11038) );
  NAND4_X1 U14080 ( .A1(n11041), .A2(n11040), .A3(n11039), .A4(n11038), .ZN(
        n11042) );
  INV_X1 U14081 ( .A(n13751), .ZN(n11046) );
  NAND2_X1 U14082 ( .A1(n10910), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11045) );
  AOI22_X1 U14083 ( .A1(n14248), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11044) );
  OAI211_X1 U14084 ( .C1(n11063), .C2(n11046), .A(n11045), .B(n11044), .ZN(
        n15422) );
  AOI22_X1 U14085 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11050) );
  AOI22_X1 U14086 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__6__SCAN_IN), .B2(n10423), .ZN(n11049) );
  AOI22_X1 U14087 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11048) );
  AOI22_X1 U14088 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12394), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11047) );
  NAND4_X1 U14089 ( .A1(n11050), .A2(n11049), .A3(n11048), .A4(n11047), .ZN(
        n11061) );
  AOI22_X1 U14090 ( .A1(n11071), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__6__SCAN_IN), .B2(n12375), .ZN(n11054) );
  AOI22_X1 U14091 ( .A1(n11072), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n9567), .ZN(n11053) );
  NAND2_X1 U14092 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11052) );
  NAND2_X1 U14093 ( .A1(n10376), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11051) );
  NAND4_X1 U14094 ( .A1(n11054), .A2(n11053), .A3(n11052), .A4(n11051), .ZN(
        n11059) );
  OAI22_X1 U14095 ( .A1(n11057), .A2(n11056), .B1(n11055), .B2(n12539), .ZN(
        n11058) );
  OR2_X1 U14096 ( .A1(n11059), .A2(n11058), .ZN(n11060) );
  NOR2_X1 U14097 ( .A1(n11061), .A2(n11060), .ZN(n13836) );
  AOI22_X1 U14098 ( .A1(n14248), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11062) );
  OAI21_X1 U14099 ( .B1(n13836), .B2(n11063), .A(n11062), .ZN(n11064) );
  AOI21_X1 U14100 ( .B1(P2_REIP_REG_14__SCAN_IN), .B2(n10910), .A(n11064), 
        .ZN(n13978) );
  INV_X1 U14101 ( .A(n13978), .ZN(n13977) );
  AOI22_X1 U14102 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11068) );
  AOI22_X1 U14103 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11067) );
  AOI22_X1 U14104 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U14105 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n12394), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11065) );
  NAND4_X1 U14106 ( .A1(n11068), .A2(n11067), .A3(n11066), .A4(n11065), .ZN(
        n11082) );
  AOI22_X1 U14107 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10341), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11080) );
  INV_X1 U14108 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11069) );
  INV_X1 U14109 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12568) );
  OAI22_X1 U14110 ( .A1(n12367), .A2(n11069), .B1(n12568), .B2(n12364), .ZN(
        n11070) );
  AOI21_X1 U14111 ( .B1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n10376), .A(
        n11070), .ZN(n11079) );
  INV_X1 U14112 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11075) );
  INV_X1 U14113 ( .A(n11071), .ZN(n11074) );
  INV_X1 U14114 ( .A(n11072), .ZN(n11073) );
  OAI22_X1 U14115 ( .A1(n11075), .A2(n11074), .B1(n11073), .B2(n10444), .ZN(
        n11076) );
  INV_X1 U14116 ( .A(n11076), .ZN(n11078) );
  NAND2_X1 U14117 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11077) );
  NAND4_X1 U14118 ( .A1(n11080), .A2(n11079), .A3(n11078), .A4(n11077), .ZN(
        n11081) );
  AOI22_X1 U14119 ( .A1(n10904), .A2(n12281), .B1(n10910), .B2(
        P2_REIP_REG_15__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U14120 ( .A1(n14248), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11083) );
  NAND2_X1 U14121 ( .A1(n11084), .A2(n11083), .ZN(n16262) );
  NAND2_X1 U14122 ( .A1(n10910), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11086) );
  AOI22_X1 U14123 ( .A1(n14248), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11085) );
  NAND2_X1 U14124 ( .A1(n10910), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11088) );
  AOI22_X1 U14125 ( .A1(n14248), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11087) );
  NAND2_X1 U14126 ( .A1(n11088), .A2(n11087), .ZN(n13966) );
  NAND2_X1 U14127 ( .A1(n15412), .A2(n13966), .ZN(n13965) );
  NAND2_X1 U14128 ( .A1(n10910), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11090) );
  AOI22_X1 U14129 ( .A1(n14248), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11089) );
  AND2_X1 U14130 ( .A1(n11090), .A2(n11089), .ZN(n14934) );
  NAND2_X1 U14131 ( .A1(n10910), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11092) );
  AOI22_X1 U14132 ( .A1(n14248), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11091) );
  NAND2_X1 U14133 ( .A1(n10910), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11094) );
  AOI22_X1 U14134 ( .A1(n14248), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11093) );
  NAND2_X1 U14135 ( .A1(n11094), .A2(n11093), .ZN(n14915) );
  NAND2_X1 U14136 ( .A1(n10910), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11096) );
  AOI22_X1 U14137 ( .A1(n14248), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11095) );
  NAND2_X1 U14138 ( .A1(n11096), .A2(n11095), .ZN(n15078) );
  NAND2_X1 U14139 ( .A1(n10910), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U14140 ( .A1(n14248), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11097) );
  NAND2_X1 U14141 ( .A1(n11098), .A2(n11097), .ZN(n15335) );
  NAND2_X1 U14142 ( .A1(n10910), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11100) );
  AOI22_X1 U14143 ( .A1(n14248), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11099) );
  AND2_X1 U14144 ( .A1(n11100), .A2(n11099), .ZN(n13040) );
  NAND2_X1 U14145 ( .A1(n10910), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11102) );
  AOI22_X1 U14146 ( .A1(n14248), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11101) );
  NAND2_X1 U14147 ( .A1(n11102), .A2(n11101), .ZN(n14903) );
  NAND2_X1 U14148 ( .A1(n10910), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11104) );
  AOI22_X1 U14149 ( .A1(n14248), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11103) );
  NAND2_X1 U14150 ( .A1(n11104), .A2(n11103), .ZN(n14214) );
  NAND2_X1 U14151 ( .A1(n10910), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11106) );
  AOI22_X1 U14152 ( .A1(n14248), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11105) );
  AND2_X1 U14153 ( .A1(n11106), .A2(n11105), .ZN(n15053) );
  NAND2_X1 U14154 ( .A1(n10910), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11108) );
  AOI22_X1 U14155 ( .A1(n14248), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11107) );
  AND2_X1 U14156 ( .A1(n11108), .A2(n11107), .ZN(n13060) );
  NAND2_X1 U14157 ( .A1(n10910), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11110) );
  AOI22_X1 U14158 ( .A1(n14248), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11109) );
  AND2_X1 U14159 ( .A1(n11110), .A2(n11109), .ZN(n14874) );
  NAND2_X1 U14160 ( .A1(n10910), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11112) );
  AOI22_X1 U14161 ( .A1(n14248), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n10944), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11111) );
  NAND2_X1 U14162 ( .A1(n11112), .A2(n11111), .ZN(n14859) );
  AOI21_X1 U14163 ( .B1(n11114), .B2(n11113), .A(n14251), .ZN(n14205) );
  INV_X1 U14164 ( .A(n11115), .ZN(n11116) );
  AND2_X1 U14165 ( .A1(n11116), .A2(n13934), .ZN(n16311) );
  INV_X1 U14166 ( .A(n11117), .ZN(n12586) );
  NOR2_X1 U14167 ( .A1(n12586), .A2(n12416), .ZN(n11118) );
  OR2_X1 U14168 ( .A1(n16311), .A2(n11118), .ZN(n11119) );
  NAND2_X1 U14169 ( .A1(n11181), .A2(n11119), .ZN(n16294) );
  NAND2_X1 U14170 ( .A1(n14205), .A2(n16280), .ZN(n11120) );
  OAI211_X1 U14171 ( .C1(n14202), .C2(n16295), .A(n11121), .B(n11120), .ZN(
        n11137) );
  NAND3_X1 U14172 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11135) );
  INV_X1 U14173 ( .A(n16297), .ZN(n15384) );
  NAND2_X1 U14174 ( .A1(n16297), .A2(n11122), .ZN(n11127) );
  INV_X1 U14175 ( .A(n11123), .ZN(n11124) );
  NOR2_X1 U14176 ( .A1(n13277), .A2(n11124), .ZN(n13292) );
  AND2_X1 U14177 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13293), .ZN(
        n11125) );
  NOR2_X1 U14178 ( .A1(n15400), .A2(n11125), .ZN(n13294) );
  NOR2_X1 U14179 ( .A1(n11181), .A2(n19155), .ZN(n16296) );
  NOR3_X1 U14180 ( .A1(n13292), .A2(n13294), .A3(n16296), .ZN(n13882) );
  OAI21_X1 U14181 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15384), .A(
        n13882), .ZN(n11126) );
  INV_X1 U14182 ( .A(n11126), .ZN(n15559) );
  NOR2_X1 U14183 ( .A1(n11174), .A2(n15520), .ZN(n15503) );
  INV_X1 U14184 ( .A(n15503), .ZN(n11128) );
  NAND2_X1 U14185 ( .A1(n16297), .A2(n11128), .ZN(n11129) );
  NAND2_X1 U14186 ( .A1(n16297), .A2(n11130), .ZN(n11131) );
  NAND2_X1 U14187 ( .A1(n15487), .A2(n11131), .ZN(n15357) );
  INV_X1 U14188 ( .A(n15314), .ZN(n11133) );
  AND2_X1 U14189 ( .A1(n16297), .A2(n11133), .ZN(n11132) );
  OR2_X1 U14190 ( .A1(n15357), .A2(n11132), .ZN(n15310) );
  NOR2_X1 U14191 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n11133), .ZN(
        n11134) );
  AND2_X1 U14192 ( .A1(n15337), .A2(n11134), .ZN(n15303) );
  NOR2_X1 U14193 ( .A1(n15310), .A2(n15303), .ZN(n14211) );
  OAI21_X1 U14194 ( .B1(n15290), .B2(n15384), .A(n14211), .ZN(n15277) );
  AOI21_X1 U14195 ( .B1(n11135), .B2(n16297), .A(n15277), .ZN(n14252) );
  NOR2_X1 U14196 ( .A1(n14252), .A2(n11180), .ZN(n11136) );
  XOR2_X1 U14197 ( .A(n11139), .B(n11138), .Z(n13285) );
  OR2_X1 U14198 ( .A1(n13400), .A2(n19196), .ZN(n11140) );
  NAND2_X1 U14199 ( .A1(n11140), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13402) );
  XNOR2_X1 U14200 ( .A(n13400), .B(n11141), .ZN(n11142) );
  NOR2_X1 U14201 ( .A1(n13402), .A2(n11142), .ZN(n11143) );
  INV_X1 U14202 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15248) );
  XNOR2_X1 U14203 ( .A(n13402), .B(n11142), .ZN(n15247) );
  NOR2_X1 U14204 ( .A1(n15248), .A2(n15247), .ZN(n15246) );
  NOR2_X1 U14205 ( .A1(n11143), .A2(n15246), .ZN(n11144) );
  XOR2_X1 U14206 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11144), .Z(
        n13284) );
  NOR2_X1 U14207 ( .A1(n13285), .A2(n13284), .ZN(n13283) );
  NOR2_X1 U14208 ( .A1(n11144), .A2(n13297), .ZN(n11145) );
  OR2_X1 U14209 ( .A1(n13283), .A2(n11145), .ZN(n11146) );
  XNOR2_X1 U14210 ( .A(n11146), .B(n10496), .ZN(n13887) );
  NAND2_X1 U14211 ( .A1(n11146), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11147) );
  NAND2_X1 U14212 ( .A1(n11148), .A2(n11149), .ZN(n11150) );
  XNOR2_X2 U14213 ( .A(n11152), .B(n11153), .ZN(n13945) );
  NAND2_X1 U14214 ( .A1(n13945), .A2(n13948), .ZN(n11156) );
  INV_X1 U14215 ( .A(n11152), .ZN(n11154) );
  NAND2_X1 U14216 ( .A1(n11154), .A2(n11153), .ZN(n11155) );
  INV_X1 U14217 ( .A(n11159), .ZN(n11158) );
  NAND2_X1 U14218 ( .A1(n11159), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15549) );
  INV_X1 U14219 ( .A(n11162), .ZN(n11161) );
  NAND2_X1 U14220 ( .A1(n11163), .A2(n11162), .ZN(n11164) );
  INV_X1 U14221 ( .A(n11166), .ZN(n11168) );
  XNOR2_X1 U14222 ( .A(n11176), .B(n11175), .ZN(n11169) );
  XNOR2_X1 U14223 ( .A(n11169), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15224) );
  NAND2_X1 U14224 ( .A1(n15225), .A2(n15224), .ZN(n11172) );
  INV_X1 U14225 ( .A(n11169), .ZN(n11170) );
  NAND2_X1 U14226 ( .A1(n11170), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11171) );
  NOR2_X4 U14227 ( .A1(n15134), .A2(n15253), .ZN(n15121) );
  NAND2_X2 U14228 ( .A1(n15121), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15116) );
  XNOR2_X1 U14229 ( .A(n15098), .B(n11180), .ZN(n15091) );
  OAI211_X1 U14230 ( .C1(n15093), .C2(n16274), .A(n11183), .B(n11182), .ZN(
        P2_U3016) );
  AND2_X2 U14231 ( .A1(n11202), .A2(n11195), .ZN(n11819) );
  NAND2_X1 U14232 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11189) );
  NOR2_X2 U14233 ( .A1(n11184), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11190) );
  AND2_X2 U14234 ( .A1(n11190), .A2(n14830), .ZN(n11422) );
  NAND2_X1 U14235 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11188) );
  NAND2_X1 U14236 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11187) );
  INV_X1 U14237 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11185) );
  AND2_X2 U14238 ( .A1(n11190), .A2(n11196), .ZN(n11461) );
  NAND2_X1 U14239 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11186) );
  NAND2_X1 U14240 ( .A1(n11419), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11194) );
  NOR2_X4 U14241 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13345) );
  AND2_X2 U14242 ( .A1(n11202), .A2(n13345), .ZN(n11273) );
  NAND2_X1 U14243 ( .A1(n11273), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11193) );
  NAND2_X1 U14244 ( .A1(n11251), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11192) );
  NAND2_X1 U14245 ( .A1(n11274), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11191) );
  NAND2_X1 U14246 ( .A1(n11420), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11201) );
  NAND2_X1 U14247 ( .A1(n11467), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11200) );
  INV_X2 U14248 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13579) );
  NAND2_X1 U14249 ( .A1(n11421), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11199) );
  NAND2_X1 U14250 ( .A1(n12014), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11198) );
  NAND2_X1 U14252 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11206) );
  AND2_X2 U14253 ( .A1(n14830), .A2(n13345), .ZN(n11372) );
  NAND2_X1 U14254 ( .A1(n11372), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11205) );
  NAND2_X1 U14255 ( .A1(n12156), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11204) );
  NAND2_X1 U14256 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11203) );
  NAND4_X4 U14257 ( .A1(n11210), .A2(n11209), .A3(n11208), .A4(n11207), .ZN(
        n20122) );
  AOI22_X1 U14258 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11214) );
  AOI22_X1 U14259 ( .A1(n11273), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11251), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11213) );
  AOI22_X1 U14260 ( .A1(n11420), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12156), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14261 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11274), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11211) );
  AOI22_X1 U14262 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11461), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11218) );
  AOI22_X1 U14263 ( .A1(n11467), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11217) );
  AOI22_X1 U14264 ( .A1(n11419), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11372), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11216) );
  AOI22_X1 U14265 ( .A1(n11421), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11266), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11215) );
  NAND2_X1 U14266 ( .A1(n11323), .A2(n11695), .ZN(n11229) );
  AOI22_X1 U14267 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11251), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11222) );
  AOI22_X1 U14268 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11467), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11221) );
  BUF_X4 U14269 ( .A(n11266), .Z(n12174) );
  AOI22_X1 U14270 ( .A1(n11421), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11220) );
  AOI22_X1 U14271 ( .A1(n12184), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12156), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11219) );
  NAND4_X1 U14272 ( .A1(n11222), .A2(n11221), .A3(n11220), .A4(n11219), .ZN(
        n11228) );
  AOI22_X1 U14273 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11419), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11226) );
  AOI22_X1 U14274 ( .A1(n11273), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11420), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11225) );
  AOI22_X1 U14275 ( .A1(n11372), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11224) );
  AOI22_X1 U14276 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11274), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11223) );
  NAND4_X1 U14277 ( .A1(n11226), .A2(n11225), .A3(n11224), .A4(n11223), .ZN(
        n11227) );
  OR2_X2 U14278 ( .A1(n11228), .A2(n11227), .ZN(n20134) );
  AND2_X2 U14279 ( .A1(n11229), .A2(n20134), .ZN(n11337) );
  NAND2_X1 U14280 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11234) );
  NAND2_X1 U14281 ( .A1(n11467), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11233) );
  NAND2_X1 U14282 ( .A1(n11372), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11232) );
  NAND2_X1 U14283 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11231) );
  NAND2_X1 U14284 ( .A1(n11419), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11238) );
  NAND2_X1 U14285 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11237) );
  NAND2_X1 U14286 ( .A1(n11251), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11236) );
  NAND2_X1 U14287 ( .A1(n12156), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11235) );
  NAND2_X1 U14288 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11242) );
  NAND2_X1 U14289 ( .A1(n11420), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11241) );
  NAND2_X1 U14290 ( .A1(n12014), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11240) );
  NAND2_X1 U14291 ( .A1(n11421), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11239) );
  NAND2_X1 U14292 ( .A1(n11273), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11246) );
  NAND2_X1 U14293 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11245) );
  NAND2_X1 U14294 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11244) );
  NAND2_X1 U14295 ( .A1(n11274), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11243) );
  AND4_X4 U14296 ( .A1(n9631), .A2(n11249), .A3(n11248), .A4(n11247), .ZN(
        n11326) );
  NAND2_X1 U14297 ( .A1(n11710), .A2(n11320), .ZN(n11250) );
  AND2_X2 U14298 ( .A1(n11337), .A2(n11250), .ZN(n11692) );
  AOI22_X1 U14299 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11251), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11255) );
  AOI22_X1 U14300 ( .A1(n12184), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11467), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14301 ( .A1(n11421), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11253) );
  AOI22_X1 U14302 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12156), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11252) );
  NAND4_X1 U14303 ( .A1(n11255), .A2(n11254), .A3(n11253), .A4(n11252), .ZN(
        n11261) );
  AOI22_X1 U14304 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11461), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11259) );
  AOI22_X1 U14305 ( .A1(n11420), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11372), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11258) );
  AOI22_X1 U14306 ( .A1(n11419), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11257) );
  AOI22_X1 U14307 ( .A1(n11273), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11274), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11256) );
  NAND4_X1 U14308 ( .A1(n11259), .A2(n11258), .A3(n11257), .A4(n11256), .ZN(
        n11260) );
  AOI22_X1 U14309 ( .A1(n11273), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11461), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11265) );
  AOI22_X1 U14310 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11251), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11264) );
  AOI22_X1 U14311 ( .A1(n11419), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12156), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11263) );
  AOI22_X1 U14312 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11274), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11262) );
  AOI22_X1 U14313 ( .A1(n12184), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11420), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11270) );
  AOI22_X1 U14314 ( .A1(n11467), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11372), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11269) );
  AOI22_X1 U14315 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11268) );
  AOI22_X1 U14316 ( .A1(n11421), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11266), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11267) );
  NAND2_X2 U14317 ( .A1(n10072), .A2(n9623), .ZN(n20112) );
  INV_X1 U14318 ( .A(n11326), .ZN(n11329) );
  NOR2_X2 U14319 ( .A1(n11531), .A2(n11271), .ZN(n11272) );
  NAND2_X1 U14320 ( .A1(n11273), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11278) );
  NAND2_X1 U14321 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11277) );
  NAND2_X1 U14322 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11276) );
  NAND2_X1 U14323 ( .A1(n11274), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11275) );
  NAND2_X1 U14324 ( .A1(n11419), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11282) );
  NAND2_X1 U14325 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11281) );
  NAND2_X1 U14326 ( .A1(n11251), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11280) );
  NAND2_X1 U14327 ( .A1(n12156), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11279) );
  BUF_X4 U14328 ( .A(n11478), .Z(n12101) );
  NAND2_X1 U14329 ( .A1(n12101), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11286) );
  NAND2_X1 U14330 ( .A1(n11420), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11285) );
  NAND2_X1 U14331 ( .A1(n12014), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11284) );
  NAND2_X1 U14332 ( .A1(n11421), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11283) );
  NAND2_X1 U14333 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11290) );
  NAND2_X1 U14334 ( .A1(n11467), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11289) );
  NAND2_X1 U14335 ( .A1(n11372), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11288) );
  NAND2_X1 U14336 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11287) );
  AND4_X4 U14337 ( .A1(n11294), .A2(n11293), .A3(n11292), .A4(n11291), .ZN(
        n20084) );
  NAND2_X1 U14338 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11298) );
  NAND2_X1 U14339 ( .A1(n12101), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11297) );
  NAND2_X1 U14340 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11296) );
  NAND2_X1 U14341 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11295) );
  AND4_X2 U14342 ( .A1(n11298), .A2(n11297), .A3(n11296), .A4(n11295), .ZN(
        n11314) );
  NAND2_X1 U14343 ( .A1(n11419), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11302) );
  NAND2_X1 U14344 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11301) );
  NAND2_X1 U14345 ( .A1(n11251), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11300) );
  NAND2_X1 U14346 ( .A1(n11274), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11299) );
  NAND2_X1 U14347 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11306) );
  NAND2_X1 U14348 ( .A1(n11273), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11305) );
  NAND2_X1 U14349 ( .A1(n11467), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11304) );
  NAND2_X1 U14350 ( .A1(n12156), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11303) );
  NAND2_X1 U14351 ( .A1(n11420), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11310) );
  NAND2_X1 U14352 ( .A1(n11372), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11309) );
  NAND2_X1 U14353 ( .A1(n11421), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11308) );
  NAND2_X1 U14354 ( .A1(n12014), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11307) );
  NAND2_X1 U14355 ( .A1(n11329), .A2(n20134), .ZN(n11327) );
  NAND2_X1 U14356 ( .A1(n11327), .A2(n13385), .ZN(n11315) );
  NAND2_X1 U14357 ( .A1(n13068), .A2(n20112), .ZN(n11336) );
  NAND2_X1 U14358 ( .A1(n13098), .A2(n20107), .ZN(n11318) );
  AND2_X1 U14359 ( .A1(n20122), .A2(n11695), .ZN(n11316) );
  INV_X1 U14360 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n11322) );
  XNOR2_X1 U14361 ( .A(n11322), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n13075) );
  NOR2_X2 U14362 ( .A1(n20112), .A2(n20107), .ZN(n11340) );
  NAND2_X2 U14363 ( .A1(n11348), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11386) );
  NAND2_X1 U14364 ( .A1(n11692), .A2(n11326), .ZN(n13071) );
  NAND2_X1 U14365 ( .A1(n13071), .A2(n13091), .ZN(n11331) );
  AND2_X4 U14366 ( .A1(n20112), .A2(n11328), .ZN(n14276) );
  NAND2_X1 U14367 ( .A1(n13242), .A2(n20107), .ZN(n13330) );
  INV_X1 U14368 ( .A(n11340), .ZN(n13335) );
  AND2_X1 U14369 ( .A1(n13330), .A2(n13335), .ZN(n11330) );
  NAND2_X1 U14370 ( .A1(n20084), .A2(n20102), .ZN(n13358) );
  NAND4_X1 U14371 ( .A1(n11331), .A2(n11335), .A3(n11330), .A4(n13358), .ZN(
        n11332) );
  INV_X1 U14372 ( .A(n11460), .ZN(n11381) );
  AOI22_X2 U14373 ( .A1(n11332), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11381), 
        .B2(n11334), .ZN(n11384) );
  NAND2_X1 U14374 ( .A1(n11334), .A2(n20084), .ZN(n13085) );
  NAND3_X1 U14375 ( .A1(n13071), .A2(n20102), .A3(n13091), .ZN(n11344) );
  INV_X1 U14376 ( .A(n13213), .ZN(n13793) );
  INV_X1 U14377 ( .A(n11337), .ZN(n11338) );
  NAND2_X1 U14378 ( .A1(n13410), .A2(n11338), .ZN(n11339) );
  NAND4_X1 U14379 ( .A1(n11339), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n16146), 
        .A4(n13358), .ZN(n11342) );
  NAND2_X1 U14380 ( .A1(n11340), .A2(n11710), .ZN(n11341) );
  NAND2_X1 U14381 ( .A1(n11341), .A2(n13330), .ZN(n13088) );
  NOR2_X1 U14382 ( .A1(n11342), .A2(n13088), .ZN(n11343) );
  NOR2_X1 U14383 ( .A1(n11392), .A2(n11345), .ZN(n11346) );
  NAND2_X1 U14384 ( .A1(n20677), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15784) );
  INV_X1 U14385 ( .A(n15784), .ZN(n15791) );
  MUX2_X1 U14386 ( .A(n12212), .B(n15791), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11387) );
  NAND2_X1 U14387 ( .A1(n11443), .A2(n11442), .ZN(n11356) );
  NAND2_X1 U14388 ( .A1(n20615), .A2(n20536), .ZN(n20507) );
  NAND2_X1 U14389 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20611) );
  NAND2_X1 U14390 ( .A1(n20507), .A2(n20611), .ZN(n20430) );
  NAND2_X1 U14391 ( .A1(n15784), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11358) );
  OAI21_X1 U14392 ( .B1(n12212), .B2(n20430), .A(n11358), .ZN(n11349) );
  OR2_X1 U14393 ( .A1(n11349), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11351) );
  AND2_X1 U14394 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n11351), .ZN(n11347) );
  NAND2_X1 U14395 ( .A1(n11348), .A2(n11347), .ZN(n11354) );
  INV_X1 U14396 ( .A(n11349), .ZN(n11350) );
  NAND2_X1 U14397 ( .A1(n11384), .A2(n11350), .ZN(n11352) );
  NAND2_X1 U14398 ( .A1(n11352), .A2(n11351), .ZN(n11353) );
  NAND2_X1 U14399 ( .A1(n11354), .A2(n11353), .ZN(n11355) );
  XNOR2_X2 U14400 ( .A(n11355), .B(n11386), .ZN(n20210) );
  INV_X1 U14401 ( .A(n11386), .ZN(n11360) );
  NAND2_X1 U14402 ( .A1(n11358), .A2(n11357), .ZN(n11359) );
  NAND2_X1 U14403 ( .A1(n11360), .A2(n11359), .ZN(n11365) );
  NAND2_X1 U14404 ( .A1(n11446), .A2(n11365), .ZN(n11363) );
  XNOR2_X1 U14405 ( .A(n20611), .B(n20371), .ZN(n20095) );
  NOR2_X1 U14406 ( .A1(n20095), .A2(n12212), .ZN(n11361) );
  NAND2_X1 U14407 ( .A1(n15784), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11364) );
  NAND2_X1 U14408 ( .A1(n11366), .A2(n11364), .ZN(n11362) );
  NAND4_X1 U14409 ( .A1(n11446), .A2(n11366), .A3(n11365), .A4(n11364), .ZN(
        n11367) );
  NAND2_X1 U14410 ( .A1(n11453), .A2(n11367), .ZN(n13571) );
  INV_X1 U14411 ( .A(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n20870) );
  AOI22_X1 U14412 ( .A1(n12183), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11371) );
  AOI22_X1 U14413 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11370) );
  AOI22_X1 U14414 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12156), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11369) );
  INV_X2 U14415 ( .A(n13337), .ZN(n12177) );
  AOI22_X1 U14416 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11368) );
  NAND4_X1 U14417 ( .A1(n11371), .A2(n11370), .A3(n11369), .A4(n11368), .ZN(
        n11378) );
  AOI22_X1 U14418 ( .A1(n12101), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11376) );
  AOI22_X1 U14419 ( .A1(n9576), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14420 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11374) );
  AOI22_X1 U14421 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11373) );
  NAND4_X1 U14422 ( .A1(n11376), .A2(n11375), .A3(n11374), .A4(n11373), .ZN(
        n11377) );
  AOI22_X1 U14423 ( .A1(n11683), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11381), .B2(n11380), .ZN(n11382) );
  AND2_X1 U14424 ( .A1(n11384), .A2(n11387), .ZN(n11385) );
  NAND2_X1 U14425 ( .A1(n11386), .A2(n11385), .ZN(n11390) );
  INV_X1 U14426 ( .A(n11387), .ZN(n11388) );
  INV_X1 U14427 ( .A(n11391), .ZN(n11392) );
  XNOR2_X2 U14428 ( .A(n11393), .B(n11391), .ZN(n11712) );
  NAND2_X1 U14429 ( .A1(n11712), .A2(n20676), .ZN(n11526) );
  AOI22_X1 U14430 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14431 ( .A1(n12184), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U14432 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12156), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14433 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11394) );
  NAND4_X1 U14434 ( .A1(n11397), .A2(n11396), .A3(n11395), .A4(n11394), .ZN(
        n11403) );
  AOI22_X1 U14435 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12183), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14436 ( .A1(n9576), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U14437 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11399) );
  BUF_X1 U14438 ( .A(n11421), .Z(n12175) );
  AOI22_X1 U14439 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11398) );
  NAND4_X1 U14440 ( .A1(n11401), .A2(n11400), .A3(n11399), .A4(n11398), .ZN(
        n11402) );
  INV_X1 U14441 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11404) );
  AOI22_X1 U14442 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11408) );
  AOI22_X1 U14443 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9576), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11407) );
  AOI22_X1 U14444 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11406) );
  AOI22_X1 U14445 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11405) );
  NAND4_X1 U14446 ( .A1(n11408), .A2(n11407), .A3(n11406), .A4(n11405), .ZN(
        n11414) );
  AOI22_X1 U14447 ( .A1(n12184), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11412) );
  AOI22_X1 U14448 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11411) );
  AOI22_X1 U14449 ( .A1(n12183), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12156), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14451 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11409) );
  NAND4_X1 U14452 ( .A1(n11412), .A2(n11411), .A3(n11410), .A4(n11409), .ZN(
        n11413) );
  OR2_X1 U14453 ( .A1(n11448), .A2(n11460), .ZN(n11415) );
  OAI211_X1 U14454 ( .C1(n11522), .C2(n11608), .A(n11416), .B(n11415), .ZN(
        n11438) );
  INV_X1 U14455 ( .A(n11438), .ZN(n11417) );
  AOI22_X1 U14456 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12013), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14457 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9576), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11426) );
  AOI22_X1 U14458 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U14459 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12156), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11424) );
  NAND4_X1 U14460 ( .A1(n11427), .A2(n11426), .A3(n11425), .A4(n11424), .ZN(
        n11434) );
  AOI22_X1 U14461 ( .A1(n12182), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11432) );
  AOI22_X1 U14462 ( .A1(n12184), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U14463 ( .A1(n12183), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11430) );
  AOI22_X1 U14464 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11429) );
  NAND4_X1 U14465 ( .A1(n11432), .A2(n11431), .A3(n11430), .A4(n11429), .ZN(
        n11433) );
  INV_X1 U14466 ( .A(n11542), .ZN(n11523) );
  INV_X1 U14467 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11435) );
  AOI21_X1 U14468 ( .B1(n11326), .B2(n11608), .A(n20676), .ZN(n11436) );
  AND2_X1 U14469 ( .A1(n11438), .A2(n11527), .ZN(n11440) );
  INV_X1 U14470 ( .A(n11522), .ZN(n11439) );
  NAND2_X1 U14471 ( .A1(n11440), .A2(n11439), .ZN(n11441) );
  INV_X1 U14472 ( .A(n20210), .ZN(n11445) );
  AND2_X1 U14473 ( .A1(n11443), .A2(n11442), .ZN(n11444) );
  OR2_X1 U14474 ( .A1(n11448), .A2(n11522), .ZN(n11449) );
  NAND2_X2 U14475 ( .A1(n11450), .A2(n11449), .ZN(n11705) );
  OAI21_X2 U14476 ( .B1(n11704), .B2(n11705), .A(n11451), .ZN(n11540) );
  INV_X1 U14477 ( .A(n11540), .ZN(n11452) );
  INV_X1 U14478 ( .A(n11554), .ZN(n11476) );
  NAND2_X1 U14479 ( .A1(n11454), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11459) );
  OAI21_X1 U14480 ( .B1(n20611), .B2(n20371), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11456) );
  INV_X1 U14481 ( .A(n20611), .ZN(n20207) );
  INV_X1 U14482 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20429) );
  NAND2_X1 U14483 ( .A1(n20429), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20304) );
  INV_X1 U14484 ( .A(n20304), .ZN(n11455) );
  NAND2_X1 U14485 ( .A1(n20207), .A2(n11455), .ZN(n20340) );
  NAND2_X1 U14486 ( .A1(n11456), .A2(n20340), .ZN(n20373) );
  INV_X1 U14487 ( .A(n12212), .ZN(n11457) );
  AOI22_X1 U14488 ( .A1(n20373), .A2(n11457), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15784), .ZN(n11458) );
  AOI22_X1 U14489 ( .A1(n12183), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11466) );
  AOI22_X1 U14490 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11465) );
  AOI22_X1 U14491 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12156), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U14492 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11463) );
  NAND4_X1 U14493 ( .A1(n11466), .A2(n11465), .A3(n11464), .A4(n11463), .ZN(
        n11473) );
  AOI22_X1 U14494 ( .A1(n12101), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U14495 ( .A1(n9576), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11470) );
  AOI22_X1 U14496 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11469) );
  AOI22_X1 U14497 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11468) );
  NAND4_X1 U14498 ( .A1(n11471), .A2(n11470), .A3(n11469), .A4(n11468), .ZN(
        n11472) );
  AOI22_X1 U14499 ( .A1(n11683), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11688), .B2(n11565), .ZN(n11474) );
  INV_X1 U14500 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11477) );
  AOI22_X1 U14501 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12059), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U14502 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9576), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U14503 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14504 ( .A1(n12183), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11479) );
  NAND4_X1 U14505 ( .A1(n11482), .A2(n11481), .A3(n11480), .A4(n11479), .ZN(
        n11488) );
  AOI22_X1 U14506 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20932), .B1(
        n11835), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11486) );
  AOI22_X1 U14507 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14508 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12013), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11484) );
  AOI22_X1 U14509 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12155), .B1(
        n12156), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11483) );
  NAND4_X1 U14510 ( .A1(n11486), .A2(n11485), .A3(n11484), .A4(n11483), .ZN(
        n11487) );
  NAND2_X1 U14511 ( .A1(n11688), .A2(n11569), .ZN(n11489) );
  INV_X1 U14512 ( .A(n11577), .ZN(n11504) );
  INV_X1 U14513 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U14514 ( .A1(n12183), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11495) );
  AOI22_X1 U14515 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11494) );
  AOI22_X1 U14516 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12156), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11493) );
  AOI22_X1 U14517 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11492) );
  NAND4_X1 U14518 ( .A1(n11495), .A2(n11494), .A3(n11493), .A4(n11492), .ZN(
        n11501) );
  AOI22_X1 U14519 ( .A1(n12101), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11499) );
  AOI22_X1 U14520 ( .A1(n9576), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11498) );
  INV_X1 U14521 ( .A(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n20905) );
  AOI22_X1 U14522 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11497) );
  AOI22_X1 U14523 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11496) );
  NAND4_X1 U14524 ( .A1(n11499), .A2(n11498), .A3(n11497), .A4(n11496), .ZN(
        n11500) );
  NAND2_X1 U14525 ( .A1(n11688), .A2(n11589), .ZN(n11502) );
  NAND2_X1 U14526 ( .A1(n11504), .A2(n11575), .ZN(n11587) );
  INV_X1 U14527 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U14528 ( .A1(n12101), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12183), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11509) );
  AOI22_X1 U14529 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12013), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U14530 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9576), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U14531 ( .A1(n12182), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11506) );
  NAND4_X1 U14532 ( .A1(n11509), .A2(n11508), .A3(n11507), .A4(n11506), .ZN(
        n11515) );
  AOI22_X1 U14533 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U14534 ( .A1(n12155), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14535 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U14536 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11510) );
  NAND4_X1 U14537 ( .A1(n11513), .A2(n11512), .A3(n11511), .A4(n11510), .ZN(
        n11514) );
  NAND2_X1 U14538 ( .A1(n11688), .A2(n11609), .ZN(n11516) );
  NAND2_X1 U14539 ( .A1(n11651), .A2(n11608), .ZN(n11520) );
  NOR2_X1 U14540 ( .A1(n11520), .A2(n11522), .ZN(n11521) );
  NAND2_X4 U14541 ( .A1(n11600), .A2(n11521), .ZN(n15965) );
  XNOR2_X1 U14542 ( .A(n11523), .B(n11608), .ZN(n11524) );
  NAND2_X1 U14543 ( .A1(n11439), .A2(n11524), .ZN(n11525) );
  NAND2_X1 U14544 ( .A1(n11526), .A2(n11525), .ZN(n11528) );
  INV_X1 U14545 ( .A(n13410), .ZN(n20765) );
  NAND2_X1 U14546 ( .A1(n20084), .A2(n20112), .ZN(n11546) );
  OAI21_X1 U14547 ( .B1(n20765), .B2(n11542), .A(n11546), .ZN(n11529) );
  INV_X1 U14548 ( .A(n11529), .ZN(n11530) );
  OR2_X1 U14549 ( .A1(n11705), .A2(n13413), .ZN(n11535) );
  XNOR2_X1 U14550 ( .A(n11543), .B(n11542), .ZN(n11532) );
  OAI211_X1 U14551 ( .C1(n11532), .C2(n20765), .A(n13216), .B(n20122), .ZN(
        n11533) );
  INV_X1 U14552 ( .A(n11533), .ZN(n11534) );
  NAND2_X1 U14553 ( .A1(n11535), .A2(n11534), .ZN(n11536) );
  XNOR2_X1 U14554 ( .A(n13097), .B(n11536), .ZN(n13455) );
  NAND2_X1 U14555 ( .A1(n13455), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11539) );
  INV_X1 U14556 ( .A(n11536), .ZN(n11537) );
  OR2_X1 U14557 ( .A1(n13097), .A2(n11537), .ZN(n11538) );
  NAND2_X1 U14558 ( .A1(n11539), .A2(n11538), .ZN(n11551) );
  INV_X1 U14559 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13498) );
  XNOR2_X1 U14560 ( .A(n11551), .B(n13498), .ZN(n13492) );
  NAND2_X1 U14561 ( .A1(n9587), .A2(n11651), .ZN(n11550) );
  NAND2_X1 U14562 ( .A1(n11543), .A2(n11542), .ZN(n11544) );
  NAND2_X1 U14563 ( .A1(n11544), .A2(n11545), .ZN(n11566) );
  OAI21_X1 U14564 ( .B1(n11545), .B2(n11544), .A(n11566), .ZN(n11548) );
  INV_X1 U14565 ( .A(n11546), .ZN(n11547) );
  AOI21_X1 U14566 ( .B1(n11548), .B2(n13410), .A(n11547), .ZN(n11549) );
  NAND2_X1 U14567 ( .A1(n11550), .A2(n11549), .ZN(n13491) );
  NAND2_X1 U14568 ( .A1(n13492), .A2(n13491), .ZN(n11553) );
  NAND2_X1 U14569 ( .A1(n11551), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11552) );
  INV_X1 U14570 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13775) );
  INV_X1 U14571 ( .A(n14825), .ZN(n14822) );
  OR2_X1 U14572 ( .A1(n11720), .A2(n11678), .ZN(n11559) );
  INV_X1 U14573 ( .A(n11565), .ZN(n11556) );
  XNOR2_X1 U14574 ( .A(n11566), .B(n11556), .ZN(n11557) );
  NAND2_X1 U14575 ( .A1(n11557), .A2(n13410), .ZN(n11558) );
  NAND2_X1 U14576 ( .A1(n11559), .A2(n11558), .ZN(n13609) );
  NAND2_X1 U14577 ( .A1(n11560), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11561) );
  NAND2_X1 U14578 ( .A1(n11563), .A2(n11562), .ZN(n11564) );
  AND2_X1 U14579 ( .A1(n11577), .A2(n11564), .ZN(n11740) );
  NAND2_X1 U14580 ( .A1(n11740), .A2(n11651), .ZN(n11572) );
  NAND2_X1 U14581 ( .A1(n11566), .A2(n11565), .ZN(n11568) );
  INV_X1 U14582 ( .A(n11568), .ZN(n11570) );
  INV_X1 U14583 ( .A(n11569), .ZN(n11567) );
  OR2_X1 U14584 ( .A1(n11568), .A2(n11567), .ZN(n11588) );
  OAI211_X1 U14585 ( .C1(n11570), .C2(n11569), .A(n13410), .B(n11588), .ZN(
        n11571) );
  NAND2_X1 U14586 ( .A1(n11572), .A2(n11571), .ZN(n11574) );
  INV_X1 U14587 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11573) );
  INV_X1 U14588 ( .A(n11575), .ZN(n11576) );
  NAND2_X1 U14589 ( .A1(n11577), .A2(n11576), .ZN(n11578) );
  NAND2_X1 U14590 ( .A1(n11587), .A2(n11578), .ZN(n11743) );
  OR2_X1 U14591 ( .A1(n11743), .A2(n11678), .ZN(n11581) );
  XNOR2_X1 U14592 ( .A(n11588), .B(n11589), .ZN(n11579) );
  NAND2_X1 U14593 ( .A1(n11579), .A2(n13410), .ZN(n11580) );
  NAND2_X1 U14594 ( .A1(n11581), .A2(n11580), .ZN(n11583) );
  INV_X1 U14595 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11582) );
  XNOR2_X1 U14596 ( .A(n11583), .B(n11582), .ZN(n13774) );
  NAND2_X1 U14597 ( .A1(n11583), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11584) );
  NAND2_X1 U14598 ( .A1(n11585), .A2(n11584), .ZN(n16030) );
  NAND2_X1 U14599 ( .A1(n11587), .A2(n11586), .ZN(n11753) );
  NAND3_X1 U14600 ( .A1(n11600), .A2(n11753), .A3(n11651), .ZN(n11593) );
  INV_X1 U14601 ( .A(n11588), .ZN(n11590) );
  NAND2_X1 U14602 ( .A1(n11590), .A2(n11589), .ZN(n11601) );
  XNOR2_X1 U14603 ( .A(n11601), .B(n11609), .ZN(n11591) );
  NAND2_X1 U14604 ( .A1(n11591), .A2(n13410), .ZN(n11592) );
  AND2_X1 U14605 ( .A1(n11593), .A2(n11592), .ZN(n11594) );
  INV_X1 U14606 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16129) );
  NAND2_X1 U14607 ( .A1(n11594), .A2(n16129), .ZN(n16028) );
  NAND2_X1 U14608 ( .A1(n16030), .A2(n16028), .ZN(n11596) );
  INV_X1 U14609 ( .A(n11594), .ZN(n11595) );
  NAND2_X1 U14610 ( .A1(n11595), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16027) );
  NAND2_X1 U14611 ( .A1(n11596), .A2(n16027), .ZN(n16022) );
  INV_X1 U14612 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11598) );
  NAND2_X1 U14613 ( .A1(n11688), .A2(n11608), .ZN(n11597) );
  OAI21_X1 U14614 ( .B1(n11668), .B2(n11598), .A(n11597), .ZN(n11599) );
  NAND2_X1 U14615 ( .A1(n11766), .A2(n11651), .ZN(n11605) );
  INV_X1 U14616 ( .A(n11601), .ZN(n11610) );
  NAND2_X1 U14617 ( .A1(n11610), .A2(n11609), .ZN(n11602) );
  XNOR2_X1 U14618 ( .A(n11602), .B(n11608), .ZN(n11603) );
  NAND2_X1 U14619 ( .A1(n11603), .A2(n13410), .ZN(n11604) );
  NAND2_X1 U14620 ( .A1(n11605), .A2(n11604), .ZN(n11606) );
  XNOR2_X1 U14621 ( .A(n11606), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16021) );
  OR2_X1 U14622 ( .A1(n11606), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11607) );
  NAND4_X1 U14623 ( .A1(n11610), .A2(n13410), .A3(n11609), .A4(n11608), .ZN(
        n11611) );
  NAND2_X1 U14624 ( .A1(n15965), .A2(n11611), .ZN(n13987) );
  NAND2_X1 U14625 ( .A1(n13987), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11612) );
  INV_X1 U14626 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11614) );
  NAND2_X1 U14627 ( .A1(n15965), .A2(n11614), .ZN(n11615) );
  INV_X1 U14628 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11624) );
  NAND2_X1 U14629 ( .A1(n15965), .A2(n11624), .ZN(n14655) );
  NAND2_X1 U14630 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11616) );
  NAND2_X1 U14631 ( .A1(n15965), .A2(n11616), .ZN(n14652) );
  AND2_X1 U14632 ( .A1(n14655), .A2(n14652), .ZN(n11617) );
  XNOR2_X1 U14633 ( .A(n15965), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14656) );
  XNOR2_X1 U14634 ( .A(n15965), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15990) );
  INV_X1 U14635 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16077) );
  NAND2_X1 U14636 ( .A1(n15965), .A2(n16077), .ZN(n14782) );
  INV_X1 U14637 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16085) );
  NAND2_X1 U14638 ( .A1(n15965), .A2(n16085), .ZN(n14635) );
  NAND4_X1 U14639 ( .A1(n14633), .A2(n15990), .A3(n14782), .A4(n14635), .ZN(
        n11619) );
  OAI21_X1 U14640 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(n16013), .ZN(n11618) );
  INV_X1 U14641 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11620) );
  NAND2_X1 U14642 ( .A1(n15965), .A2(n11620), .ZN(n11621) );
  NAND2_X1 U14643 ( .A1(n11622), .A2(n11621), .ZN(n11627) );
  INV_X1 U14644 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14643) );
  NAND2_X1 U14645 ( .A1(n14643), .A2(n16085), .ZN(n11623) );
  NAND2_X1 U14646 ( .A1(n16013), .A2(n11623), .ZN(n14779) );
  NAND2_X1 U14647 ( .A1(n16013), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14783) );
  NAND2_X1 U14648 ( .A1(n14779), .A2(n14783), .ZN(n14637) );
  NOR2_X1 U14649 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14650) );
  AND2_X1 U14650 ( .A1(n14650), .A2(n11624), .ZN(n11625) );
  NOR2_X1 U14651 ( .A1(n15965), .A2(n11625), .ZN(n14634) );
  NOR2_X1 U14652 ( .A1(n14637), .A2(n14634), .ZN(n11626) );
  XNOR2_X1 U14653 ( .A(n15965), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14626) );
  NAND2_X1 U14654 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14767) );
  INV_X1 U14655 ( .A(n14767), .ZN(n14688) );
  NAND2_X1 U14656 ( .A1(n11628), .A2(n15965), .ZN(n14617) );
  NAND2_X1 U14657 ( .A1(n14617), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11631) );
  INV_X1 U14658 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16067) );
  INV_X1 U14659 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15806) );
  NAND2_X1 U14660 ( .A1(n16067), .A2(n15806), .ZN(n11629) );
  OR2_X2 U14661 ( .A1(n14627), .A2(n11629), .ZN(n15812) );
  INV_X1 U14662 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14772) );
  INV_X1 U14663 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15822) );
  NAND2_X1 U14664 ( .A1(n14772), .A2(n15822), .ZN(n11630) );
  OAI21_X1 U14665 ( .B1(n15812), .B2(n11630), .A(n16013), .ZN(n14618) );
  NAND2_X1 U14666 ( .A1(n11631), .A2(n14618), .ZN(n15967) );
  INV_X1 U14667 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16047) );
  INV_X1 U14668 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14609) );
  INV_X1 U14669 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14741) );
  NAND3_X1 U14670 ( .A1(n16047), .A2(n14609), .A3(n14741), .ZN(n14568) );
  NOR2_X1 U14671 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14720) );
  NAND2_X1 U14672 ( .A1(n11631), .A2(n15965), .ZN(n14598) );
  NAND3_X1 U14673 ( .A1(n14590), .A2(n14720), .A3(n11632), .ZN(n14547) );
  AND2_X1 U14674 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14742) );
  NAND2_X1 U14675 ( .A1(n14742), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14736) );
  NAND2_X1 U14676 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14698) );
  INV_X1 U14677 ( .A(n14698), .ZN(n11633) );
  AOI21_X1 U14678 ( .B1(n16013), .B2(n14547), .A(n11634), .ZN(n14558) );
  INV_X1 U14679 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14697) );
  NAND2_X1 U14680 ( .A1(n16013), .A2(n14697), .ZN(n14557) );
  NOR2_X1 U14681 ( .A1(n14557), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11636) );
  NAND2_X1 U14682 ( .A1(n15965), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14556) );
  AOI22_X1 U14683 ( .A1(n14558), .A2(n11636), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14545), .ZN(n11637) );
  NAND2_X1 U14684 ( .A1(n20615), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11639) );
  NAND2_X1 U14685 ( .A1(n11357), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11638) );
  NAND2_X1 U14686 ( .A1(n11639), .A2(n11638), .ZN(n11648) );
  NAND2_X1 U14687 ( .A1(n20888), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11641) );
  NAND2_X1 U14688 ( .A1(n11643), .A2(n11641), .ZN(n11665) );
  INV_X1 U14689 ( .A(n11665), .ZN(n11642) );
  XNOR2_X1 U14690 ( .A(n13579), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11673) );
  AOI222_X1 U14691 ( .A1(n11670), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .B1(n11670), .B2(n16150), .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .C2(n16150), .ZN(n12223) );
  INV_X1 U14692 ( .A(n11650), .ZN(n11647) );
  XNOR2_X1 U14693 ( .A(n11648), .B(n11647), .ZN(n12221) );
  NAND2_X1 U14694 ( .A1(n13384), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11658) );
  NAND2_X1 U14695 ( .A1(n11688), .A2(n20102), .ZN(n11649) );
  OAI211_X1 U14696 ( .C1(n11668), .C2(n12221), .A(n11658), .B(n11649), .ZN(
        n11660) );
  INV_X1 U14697 ( .A(n11660), .ZN(n11664) );
  OAI21_X1 U14698 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20536), .A(
        n11650), .ZN(n11655) );
  INV_X1 U14699 ( .A(n11655), .ZN(n11652) );
  AOI21_X1 U14700 ( .B1(n11652), .B2(n11688), .A(n11689), .ZN(n11657) );
  OR2_X1 U14701 ( .A1(n20084), .A2(n20122), .ZN(n11653) );
  NAND2_X1 U14702 ( .A1(n11653), .A2(n13413), .ZN(n11675) );
  OAI21_X1 U14703 ( .B1(n13098), .B2(n20084), .A(n11675), .ZN(n11654) );
  NOR2_X1 U14704 ( .A1(n11655), .A2(n11654), .ZN(n11656) );
  NOR2_X1 U14705 ( .A1(n11657), .A2(n11656), .ZN(n11661) );
  INV_X1 U14706 ( .A(n11661), .ZN(n11663) );
  INV_X1 U14707 ( .A(n11658), .ZN(n11659) );
  OAI22_X1 U14708 ( .A1(n11661), .A2(n11660), .B1(n11669), .B2(n12221), .ZN(
        n11662) );
  OAI21_X1 U14709 ( .B1(n11664), .B2(n11663), .A(n11662), .ZN(n11682) );
  XNOR2_X1 U14710 ( .A(n11666), .B(n11665), .ZN(n12220) );
  NAND2_X1 U14711 ( .A1(n11688), .A2(n12220), .ZN(n11667) );
  OAI211_X1 U14712 ( .C1(n11668), .C2(n12220), .A(n11675), .B(n11667), .ZN(
        n11681) );
  INV_X1 U14713 ( .A(n11669), .ZN(n11672) );
  AND2_X1 U14714 ( .A1(n16150), .A2(n11670), .ZN(n11671) );
  NAND2_X1 U14715 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n11671), .ZN(
        n12222) );
  NOR2_X1 U14716 ( .A1(n11672), .A2(n12222), .ZN(n11680) );
  XNOR2_X1 U14717 ( .A(n11674), .B(n11673), .ZN(n12219) );
  INV_X1 U14718 ( .A(n11675), .ZN(n11676) );
  NAND3_X1 U14719 ( .A1(n11676), .A2(n11688), .A3(n12220), .ZN(n11677) );
  OAI21_X1 U14720 ( .B1(n12219), .B2(n11678), .A(n11677), .ZN(n11679) );
  AOI211_X1 U14721 ( .C1(n11682), .C2(n11681), .A(n11680), .B(n11679), .ZN(
        n11685) );
  AOI21_X1 U14722 ( .B1(n12222), .B2(n12219), .A(n11683), .ZN(n11684) );
  OR2_X1 U14723 ( .A1(n11685), .A2(n11684), .ZN(n11686) );
  AND2_X1 U14724 ( .A1(n12223), .A2(n11689), .ZN(n11690) );
  NAND2_X1 U14725 ( .A1(n13091), .A2(n20084), .ZN(n11693) );
  NAND2_X1 U14726 ( .A1(n13100), .A2(n11320), .ZN(n15776) );
  NOR2_X1 U14727 ( .A1(n15776), .A2(n19873), .ZN(n11694) );
  NOR2_X2 U14728 ( .A1(n11695), .A2(n20679), .ZN(n11887) );
  NAND2_X1 U14729 ( .A1(n11696), .A2(n11887), .ZN(n11702) );
  INV_X1 U14730 ( .A(n13385), .ZN(n12241) );
  NAND2_X1 U14731 ( .A1(n12241), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11726) );
  NOR2_X1 U14732 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11697) );
  XNOR2_X1 U14733 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14365) );
  AOI21_X1 U14734 ( .B1(n11697), .B2(n14365), .A(n12200), .ZN(n11699) );
  NAND2_X1 U14735 ( .A1(n12201), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11698) );
  OAI211_X1 U14736 ( .C1(n11726), .C2(n20888), .A(n11699), .B(n11698), .ZN(
        n11700) );
  INV_X1 U14737 ( .A(n11700), .ZN(n11701) );
  NAND2_X1 U14738 ( .A1(n11702), .A2(n11701), .ZN(n11703) );
  NAND2_X1 U14739 ( .A1(n12200), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11719) );
  XNOR2_X2 U14740 ( .A(n11705), .B(n11704), .ZN(n20172) );
  NAND2_X1 U14741 ( .A1(n20172), .A2(n11887), .ZN(n11709) );
  AOI22_X1 U14742 ( .A1(n12201), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20679), .ZN(n11707) );
  INV_X1 U14743 ( .A(n11726), .ZN(n11730) );
  NAND2_X1 U14744 ( .A1(n11730), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11706) );
  AND2_X1 U14745 ( .A1(n11707), .A2(n11706), .ZN(n11708) );
  NAND2_X1 U14746 ( .A1(n11709), .A2(n11708), .ZN(n13374) );
  NAND2_X1 U14747 ( .A1(n20171), .A2(n11710), .ZN(n11711) );
  NAND2_X1 U14748 ( .A1(n11711), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13395) );
  NAND2_X1 U14749 ( .A1(n11713), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11715) );
  NAND2_X1 U14750 ( .A1(n20679), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11714) );
  OAI211_X1 U14751 ( .C1(n11726), .C2(n11345), .A(n11715), .B(n11714), .ZN(
        n11716) );
  AOI21_X1 U14752 ( .B1(n11712), .B2(n11887), .A(n11716), .ZN(n13394) );
  OR2_X1 U14753 ( .A1(n13395), .A2(n13394), .ZN(n13397) );
  INV_X1 U14754 ( .A(n13394), .ZN(n11717) );
  OR2_X1 U14755 ( .A1(n11717), .A2(n12170), .ZN(n11718) );
  NAND2_X1 U14756 ( .A1(n13397), .A2(n11718), .ZN(n13373) );
  NAND2_X1 U14757 ( .A1(n13374), .A2(n13373), .ZN(n13511) );
  NAND2_X1 U14758 ( .A1(n9676), .A2(n13513), .ZN(n13512) );
  INV_X1 U14759 ( .A(n11720), .ZN(n11721) );
  NAND2_X1 U14760 ( .A1(n11721), .A2(n11887), .ZN(n11729) );
  INV_X1 U14761 ( .A(n11722), .ZN(n11723) );
  INV_X1 U14762 ( .A(n11732), .ZN(n11733) );
  OAI21_X1 U14763 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11723), .A(
        n11733), .ZN(n13806) );
  AOI22_X1 U14764 ( .A1(n12142), .A2(n13806), .B1(n12200), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11725) );
  NAND2_X1 U14765 ( .A1(n12201), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11724) );
  OAI211_X1 U14766 ( .C1(n11726), .C2(n13579), .A(n11725), .B(n11724), .ZN(
        n11727) );
  INV_X1 U14767 ( .A(n11727), .ZN(n11728) );
  NAND2_X1 U14768 ( .A1(n11730), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11738) );
  INV_X1 U14769 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11734) );
  AOI21_X1 U14770 ( .B1(n11734), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11731) );
  AOI21_X1 U14771 ( .B1(n12201), .B2(P1_EAX_REG_4__SCAN_IN), .A(n11731), .ZN(
        n11737) );
  INV_X1 U14772 ( .A(n11744), .ZN(n11745) );
  NAND2_X1 U14773 ( .A1(n11734), .A2(n11733), .ZN(n11735) );
  NAND2_X1 U14774 ( .A1(n11745), .A2(n11735), .ZN(n19987) );
  NOR2_X1 U14775 ( .A1(n19987), .A2(n12170), .ZN(n11736) );
  AOI21_X1 U14776 ( .B1(n11738), .B2(n11737), .A(n11736), .ZN(n11739) );
  AOI21_X1 U14777 ( .B1(n11740), .B2(n11887), .A(n11739), .ZN(n13622) );
  INV_X1 U14778 ( .A(n11887), .ZN(n11873) );
  INV_X1 U14779 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16040) );
  INV_X1 U14780 ( .A(n12200), .ZN(n11815) );
  INV_X1 U14781 ( .A(n11754), .ZN(n11747) );
  NAND2_X1 U14782 ( .A1(n11745), .A2(n16040), .ZN(n11746) );
  NAND2_X1 U14783 ( .A1(n11747), .A2(n11746), .ZN(n19957) );
  NAND2_X1 U14784 ( .A1(n19957), .A2(n11697), .ZN(n11748) );
  OAI21_X1 U14785 ( .B1(n16040), .B2(n11815), .A(n11748), .ZN(n11749) );
  AOI21_X1 U14786 ( .B1(n12201), .B2(P1_EAX_REG_5__SCAN_IN), .A(n11749), .ZN(
        n11750) );
  INV_X1 U14787 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11757) );
  NAND2_X1 U14788 ( .A1(n11753), .A2(n11887), .ZN(n11756) );
  OAI21_X1 U14789 ( .B1(n11754), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n11758), .ZN(n19945) );
  INV_X1 U14790 ( .A(n12170), .ZN(n12142) );
  AOI22_X1 U14791 ( .A1(n19945), .A2(n12142), .B1(n12200), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11755) );
  NAND2_X1 U14792 ( .A1(n13648), .A2(n13757), .ZN(n13721) );
  INV_X1 U14793 ( .A(n13721), .ZN(n11768) );
  INV_X1 U14794 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13748) );
  NAND2_X1 U14795 ( .A1(n11758), .A2(n11761), .ZN(n11760) );
  INV_X1 U14796 ( .A(n11782), .ZN(n11759) );
  NAND2_X1 U14797 ( .A1(n11760), .A2(n11759), .ZN(n19934) );
  NOR2_X1 U14798 ( .A1(n11815), .A2(n11761), .ZN(n11762) );
  AOI21_X1 U14799 ( .B1(n19934), .B2(n12142), .A(n11762), .ZN(n11763) );
  OAI21_X1 U14800 ( .B1(n11764), .B2(n13748), .A(n11763), .ZN(n11765) );
  AOI21_X1 U14801 ( .B1(n11766), .B2(n11887), .A(n11765), .ZN(n13722) );
  NAND2_X1 U14802 ( .A1(n11768), .A2(n11767), .ZN(n13719) );
  AOI22_X1 U14803 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11772) );
  AOI22_X1 U14804 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11771) );
  AOI22_X1 U14805 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11770) );
  AOI22_X1 U14806 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11769) );
  NAND4_X1 U14807 ( .A1(n11772), .A2(n11771), .A3(n11770), .A4(n11769), .ZN(
        n11778) );
  AOI22_X1 U14808 ( .A1(n12101), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U14809 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U14810 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9576), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U14811 ( .A1(n12183), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11773) );
  NAND4_X1 U14812 ( .A1(n11776), .A2(n11775), .A3(n11774), .A4(n11773), .ZN(
        n11777) );
  OAI21_X1 U14813 ( .B1(n11778), .B2(n11777), .A(n11887), .ZN(n11781) );
  NAND2_X1 U14814 ( .A1(n12201), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11780) );
  XNOR2_X1 U14815 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11782), .ZN(
        n19917) );
  AOI22_X1 U14816 ( .A1(n12142), .A2(n19917), .B1(n12200), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11779) );
  XOR2_X1 U14817 ( .A(n11806), .B(n11807), .Z(n19908) );
  AOI22_X1 U14818 ( .A1(n12101), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U14819 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11785) );
  AOI22_X1 U14820 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11784) );
  AOI22_X1 U14821 ( .A1(n12183), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11783) );
  NAND4_X1 U14822 ( .A1(n11786), .A2(n11785), .A3(n11784), .A4(n11783), .ZN(
        n11792) );
  AOI22_X1 U14823 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9576), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11790) );
  AOI22_X1 U14824 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11789) );
  AOI22_X1 U14825 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U14826 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11787) );
  NAND4_X1 U14827 ( .A1(n11790), .A2(n11789), .A3(n11788), .A4(n11787), .ZN(
        n11791) );
  OR2_X1 U14828 ( .A1(n11792), .A2(n11791), .ZN(n11793) );
  AOI22_X1 U14829 ( .A1(n11887), .A2(n11793), .B1(n12200), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11795) );
  NAND2_X1 U14830 ( .A1(n12201), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11794) );
  OAI211_X1 U14831 ( .C1(n19908), .C2(n12170), .A(n11795), .B(n11794), .ZN(
        n13893) );
  AOI22_X1 U14832 ( .A1(n12183), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U14833 ( .A1(n12101), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9576), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U14834 ( .A1(n11421), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U14835 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11796) );
  NAND4_X1 U14836 ( .A1(n11799), .A2(n11798), .A3(n11797), .A4(n11796), .ZN(
        n11805) );
  AOI22_X1 U14837 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11803) );
  AOI22_X1 U14838 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U14839 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U14840 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11800) );
  NAND4_X1 U14841 ( .A1(n11803), .A2(n11802), .A3(n11801), .A4(n11800), .ZN(
        n11804) );
  NOR2_X1 U14842 ( .A1(n11805), .A2(n11804), .ZN(n11810) );
  XNOR2_X1 U14843 ( .A(n11811), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15941) );
  NAND2_X1 U14844 ( .A1(n15941), .A2(n11697), .ZN(n11809) );
  AOI22_X1 U14845 ( .A1(n12201), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12200), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11808) );
  OAI211_X1 U14846 ( .C1(n11810), .C2(n11873), .A(n11809), .B(n11808), .ZN(
        n13918) );
  INV_X1 U14847 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11814) );
  OAI21_X1 U14848 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11812), .A(
        n11855), .ZN(n16020) );
  NAND2_X1 U14849 ( .A1(n16020), .A2(n12142), .ZN(n11813) );
  OAI21_X1 U14850 ( .B1(n11815), .B2(n11814), .A(n11813), .ZN(n11816) );
  AOI21_X1 U14851 ( .B1(n12201), .B2(P1_EAX_REG_11__SCAN_IN), .A(n11816), .ZN(
        n14046) );
  AOI22_X1 U14852 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11823) );
  AOI22_X1 U14853 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12013), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11822) );
  AOI22_X1 U14854 ( .A1(n12182), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11821) );
  AOI22_X1 U14855 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11820) );
  NAND4_X1 U14856 ( .A1(n11823), .A2(n11822), .A3(n11821), .A4(n11820), .ZN(
        n11829) );
  AOI22_X1 U14857 ( .A1(n12101), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9576), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U14858 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U14859 ( .A1(n12183), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U14860 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11824) );
  NAND4_X1 U14861 ( .A1(n11827), .A2(n11826), .A3(n11825), .A4(n11824), .ZN(
        n11828) );
  OR2_X1 U14862 ( .A1(n11829), .A2(n11828), .ZN(n11830) );
  NAND2_X1 U14863 ( .A1(n11887), .A2(n11830), .ZN(n14082) );
  XOR2_X1 U14864 ( .A(n14069), .B(n11870), .Z(n14658) );
  AOI22_X1 U14865 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12183), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11834) );
  AOI22_X1 U14866 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U14867 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11832) );
  AOI22_X1 U14868 ( .A1(n12101), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11831) );
  NAND4_X1 U14869 ( .A1(n11834), .A2(n11833), .A3(n11832), .A4(n11831), .ZN(
        n11841) );
  AOI22_X1 U14870 ( .A1(n12182), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U14871 ( .A1(n9576), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U14872 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U14873 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11836) );
  NAND4_X1 U14874 ( .A1(n11839), .A2(n11838), .A3(n11837), .A4(n11836), .ZN(
        n11840) );
  OR2_X1 U14875 ( .A1(n11841), .A2(n11840), .ZN(n11842) );
  AOI22_X1 U14876 ( .A1(n11887), .A2(n11842), .B1(n12200), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11844) );
  NAND2_X1 U14877 ( .A1(n12201), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11843) );
  OAI211_X1 U14878 ( .C1(n14658), .C2(n12170), .A(n11844), .B(n11843), .ZN(
        n14050) );
  AOI22_X1 U14879 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U14880 ( .A1(n12059), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9576), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U14881 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U14882 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11845) );
  NAND4_X1 U14883 ( .A1(n11848), .A2(n11847), .A3(n11846), .A4(n11845), .ZN(
        n11854) );
  AOI22_X1 U14884 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12182), .B1(
        n12183), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11852) );
  AOI22_X1 U14885 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12013), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11851) );
  AOI22_X1 U14886 ( .A1(n12155), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U14887 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11849) );
  NAND4_X1 U14888 ( .A1(n11852), .A2(n11851), .A3(n11850), .A4(n11849), .ZN(
        n11853) );
  NOR2_X1 U14889 ( .A1(n11854), .A2(n11853), .ZN(n11859) );
  XOR2_X1 U14890 ( .A(n15923), .B(n11855), .Z(n16006) );
  INV_X1 U14891 ( .A(n16006), .ZN(n11856) );
  AOI22_X1 U14892 ( .A1(n12200), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n11697), .B2(n11856), .ZN(n11858) );
  NAND2_X1 U14893 ( .A1(n12201), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11857) );
  OAI211_X1 U14894 ( .C1(n11873), .C2(n11859), .A(n11858), .B(n11857), .ZN(
        n14089) );
  AOI22_X1 U14895 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11863) );
  AOI22_X1 U14896 ( .A1(n12059), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11862) );
  AOI22_X1 U14897 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U14898 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11860) );
  NAND4_X1 U14899 ( .A1(n11863), .A2(n11862), .A3(n11861), .A4(n11860), .ZN(
        n11869) );
  AOI22_X1 U14900 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12183), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U14901 ( .A1(n9576), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11866) );
  AOI22_X1 U14902 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U14903 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11864) );
  NAND4_X1 U14904 ( .A1(n11867), .A2(n11866), .A3(n11865), .A4(n11864), .ZN(
        n11868) );
  NOR2_X1 U14905 ( .A1(n11869), .A2(n11868), .ZN(n11874) );
  XNOR2_X1 U14906 ( .A(n11875), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15916) );
  NAND2_X1 U14907 ( .A1(n15916), .A2(n12142), .ZN(n11872) );
  AOI22_X1 U14908 ( .A1(n12201), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n12200), 
        .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11871) );
  OAI211_X1 U14909 ( .C1(n11874), .C2(n11873), .A(n11872), .B(n11871), .ZN(
        n14041) );
  XOR2_X1 U14910 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n11890), .Z(
        n16000) );
  AOI22_X1 U14911 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12183), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U14912 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U14913 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U14914 ( .A1(n12059), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11876) );
  NAND4_X1 U14915 ( .A1(n11879), .A2(n11878), .A3(n11877), .A4(n11876), .ZN(
        n11885) );
  AOI22_X1 U14916 ( .A1(n12182), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9576), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11883) );
  AOI22_X1 U14917 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U14918 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11881) );
  AOI22_X1 U14919 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11880) );
  NAND4_X1 U14920 ( .A1(n11883), .A2(n11882), .A3(n11881), .A4(n11880), .ZN(
        n11884) );
  OR2_X1 U14921 ( .A1(n11885), .A2(n11884), .ZN(n11886) );
  AOI22_X1 U14922 ( .A1(n11887), .A2(n11886), .B1(n12200), .B2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11889) );
  NAND2_X1 U14923 ( .A1(n12201), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11888) );
  OAI211_X1 U14924 ( .C1(n16000), .C2(n12170), .A(n11889), .B(n11888), .ZN(
        n14098) );
  XNOR2_X1 U14925 ( .A(n11907), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15897) );
  NAND2_X1 U14926 ( .A1(n15897), .A2(n12142), .ZN(n11906) );
  AOI22_X1 U14927 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U14928 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9576), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U14929 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12014), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U14930 ( .A1(n12059), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11891) );
  NAND4_X1 U14931 ( .A1(n11894), .A2(n11893), .A3(n11892), .A4(n11891), .ZN(
        n11902) );
  AOI22_X1 U14932 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12013), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11900) );
  AOI22_X1 U14933 ( .A1(n12155), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U14934 ( .A1(n12183), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11898) );
  NAND2_X1 U14935 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11896) );
  NAND2_X1 U14936 ( .A1(n12177), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11895) );
  AND3_X1 U14937 ( .A1(n11896), .A2(n12170), .A3(n11895), .ZN(n11897) );
  NAND4_X1 U14938 ( .A1(n11900), .A2(n11899), .A3(n11898), .A4(n11897), .ZN(
        n11901) );
  NAND2_X1 U14939 ( .A1(n12167), .A2(n12170), .ZN(n12002) );
  OAI21_X1 U14940 ( .B1(n11902), .B2(n11901), .A(n12002), .ZN(n11904) );
  AOI22_X1 U14941 ( .A1(n12201), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20679), .ZN(n11903) );
  NAND2_X1 U14942 ( .A1(n11904), .A2(n11903), .ZN(n11905) );
  NAND2_X1 U14943 ( .A1(n11906), .A2(n11905), .ZN(n14451) );
  NOR2_X2 U14944 ( .A1(n14099), .A2(n14451), .ZN(n14441) );
  INV_X1 U14945 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15880) );
  INV_X1 U14946 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15891) );
  XOR2_X1 U14947 ( .A(n15880), .B(n11923), .Z(n15996) );
  INV_X1 U14948 ( .A(n15996), .ZN(n11921) );
  AOI22_X1 U14949 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12013), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U14950 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U14951 ( .A1(n11421), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12014), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U14952 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11908) );
  NAND4_X1 U14953 ( .A1(n11911), .A2(n11910), .A3(n11909), .A4(n11908), .ZN(
        n11917) );
  AOI22_X1 U14954 ( .A1(n12059), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U14955 ( .A1(n9576), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U14956 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U14957 ( .A1(n12183), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11912) );
  NAND4_X1 U14958 ( .A1(n11915), .A2(n11914), .A3(n11913), .A4(n11912), .ZN(
        n11916) );
  NOR2_X1 U14959 ( .A1(n11917), .A2(n11916), .ZN(n11919) );
  AOI22_X1 U14960 ( .A1(n12201), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n12200), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11918) );
  OAI21_X1 U14961 ( .B1(n12167), .B2(n11919), .A(n11918), .ZN(n11920) );
  AOI21_X1 U14962 ( .B1(n11921), .B2(n12142), .A(n11920), .ZN(n14444) );
  INV_X1 U14963 ( .A(n14444), .ZN(n11922) );
  XNOR2_X1 U14964 ( .A(n11954), .B(n14360), .ZN(n14629) );
  AOI22_X1 U14965 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12013), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11927) );
  AOI22_X1 U14966 ( .A1(n12182), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U14967 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12014), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U14968 ( .A1(n12155), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11924) );
  NAND4_X1 U14969 ( .A1(n11927), .A2(n11926), .A3(n11925), .A4(n11924), .ZN(
        n11935) );
  AOI22_X1 U14970 ( .A1(n12059), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11423), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U14971 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9576), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11932) );
  AOI22_X1 U14972 ( .A1(n12183), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11931) );
  NAND2_X1 U14973 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11929) );
  NAND2_X1 U14974 ( .A1(n12177), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11928) );
  AND3_X1 U14975 ( .A1(n11929), .A2(n12170), .A3(n11928), .ZN(n11930) );
  NAND4_X1 U14976 ( .A1(n11933), .A2(n11932), .A3(n11931), .A4(n11930), .ZN(
        n11934) );
  OAI21_X1 U14977 ( .B1(n11935), .B2(n11934), .A(n12002), .ZN(n11937) );
  AOI22_X1 U14978 ( .A1(n12201), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20679), .ZN(n11936) );
  NAND2_X1 U14979 ( .A1(n11937), .A2(n11936), .ZN(n11938) );
  OAI21_X1 U14980 ( .B1(n14629), .B2(n12170), .A(n11938), .ZN(n14354) );
  AOI22_X1 U14981 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12183), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U14982 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11942) );
  AOI22_X1 U14983 ( .A1(n12059), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9576), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11941) );
  AOI22_X1 U14984 ( .A1(n12182), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11940) );
  NAND4_X1 U14985 ( .A1(n11943), .A2(n11942), .A3(n11941), .A4(n11940), .ZN(
        n11949) );
  AOI22_X1 U14986 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11947) );
  AOI22_X1 U14987 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11946) );
  AOI22_X1 U14988 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12156), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U14989 ( .A1(n11421), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12014), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11944) );
  NAND4_X1 U14990 ( .A1(n11947), .A2(n11946), .A3(n11945), .A4(n11944), .ZN(
        n11948) );
  NOR2_X1 U14991 ( .A1(n11949), .A2(n11948), .ZN(n11953) );
  INV_X1 U14992 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20777) );
  OAI21_X1 U14993 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20777), .A(
        n20679), .ZN(n11950) );
  INV_X1 U14994 ( .A(n11950), .ZN(n11951) );
  AOI21_X1 U14995 ( .B1(n12201), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11951), .ZN(
        n11952) );
  OAI21_X1 U14996 ( .B1(n12167), .B2(n11953), .A(n11952), .ZN(n11957) );
  OAI21_X1 U14997 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n11955), .A(
        n11988), .ZN(n15989) );
  OR2_X1 U14998 ( .A1(n12170), .A2(n15989), .ZN(n11956) );
  AOI22_X1 U14999 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12182), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U15000 ( .A1(n12059), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U15001 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12156), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11961) );
  NAND2_X1 U15002 ( .A1(n12177), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11959) );
  NAND2_X1 U15003 ( .A1(n12014), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11958) );
  AND3_X1 U15004 ( .A1(n11959), .A2(n11958), .A3(n12170), .ZN(n11960) );
  NAND4_X1 U15005 ( .A1(n11963), .A2(n11962), .A3(n11961), .A4(n11960), .ZN(
        n11969) );
  AOI22_X1 U15006 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11835), .B1(
        n12013), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U15007 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12183), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U15008 ( .A1(n9576), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12175), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11965) );
  AOI22_X1 U15009 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11964) );
  NAND4_X1 U15010 ( .A1(n11967), .A2(n11966), .A3(n11965), .A4(n11964), .ZN(
        n11968) );
  OR2_X1 U15011 ( .A1(n11969), .A2(n11968), .ZN(n11970) );
  NAND2_X1 U15012 ( .A1(n12002), .A2(n11970), .ZN(n11973) );
  AOI22_X1 U15013 ( .A1(n12201), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20679), .ZN(n11972) );
  XNOR2_X1 U15014 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n11988), .ZN(
        n15980) );
  AOI21_X1 U15015 ( .B1(n11973), .B2(n11972), .A(n11971), .ZN(n14426) );
  AOI22_X1 U15016 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12013), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U15017 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U15018 ( .A1(n11421), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12014), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U15019 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12156), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11974) );
  NAND4_X1 U15020 ( .A1(n11977), .A2(n11976), .A3(n11975), .A4(n11974), .ZN(
        n11983) );
  AOI22_X1 U15021 ( .A1(n12059), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11981) );
  AOI22_X1 U15022 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9576), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11980) );
  AOI22_X1 U15023 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11979) );
  AOI22_X1 U15024 ( .A1(n12183), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11978) );
  NAND4_X1 U15025 ( .A1(n11981), .A2(n11980), .A3(n11979), .A4(n11978), .ZN(
        n11982) );
  NOR2_X1 U15026 ( .A1(n11983), .A2(n11982), .ZN(n11987) );
  NAND2_X1 U15027 ( .A1(n20679), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11984) );
  NAND2_X1 U15028 ( .A1(n12170), .A2(n11984), .ZN(n11985) );
  AOI21_X1 U15029 ( .B1(n11713), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11985), .ZN(
        n11986) );
  OAI21_X1 U15030 ( .B1(n12167), .B2(n11987), .A(n11986), .ZN(n11991) );
  INV_X1 U15031 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15983) );
  OAI21_X1 U15032 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n11989), .A(
        n12036), .ZN(n15976) );
  OR2_X1 U15033 ( .A1(n12170), .A2(n15976), .ZN(n11990) );
  AOI22_X1 U15034 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11835), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11995) );
  AOI22_X1 U15035 ( .A1(n12101), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12175), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11994) );
  AOI22_X1 U15036 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U15037 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12156), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11992) );
  NAND4_X1 U15038 ( .A1(n11995), .A2(n11994), .A3(n11993), .A4(n11992), .ZN(
        n12004) );
  AOI22_X1 U15039 ( .A1(n12183), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U15040 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9576), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U15041 ( .A1(n12182), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11999) );
  NAND2_X1 U15042 ( .A1(n12177), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11997) );
  NAND2_X1 U15043 ( .A1(n12014), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11996) );
  AND3_X1 U15044 ( .A1(n11997), .A2(n11996), .A3(n12170), .ZN(n11998) );
  NAND4_X1 U15045 ( .A1(n12001), .A2(n12000), .A3(n11999), .A4(n11998), .ZN(
        n12003) );
  OAI21_X1 U15046 ( .B1(n12004), .B2(n12003), .A(n12002), .ZN(n12006) );
  AOI22_X1 U15047 ( .A1(n12201), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20679), .ZN(n12005) );
  NAND2_X1 U15048 ( .A1(n12006), .A2(n12005), .ZN(n12008) );
  XNOR2_X1 U15049 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B(n12036), .ZN(
        n15847) );
  NAND2_X1 U15050 ( .A1(n15847), .A2(n12142), .ZN(n12007) );
  NAND2_X1 U15051 ( .A1(n12008), .A2(n12007), .ZN(n14408) );
  AOI22_X1 U15052 ( .A1(n12059), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U15053 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12011) );
  AOI22_X1 U15054 ( .A1(n12182), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U15055 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12009) );
  NAND4_X1 U15056 ( .A1(n12012), .A2(n12011), .A3(n12010), .A4(n12009), .ZN(
        n12021) );
  AOI22_X1 U15057 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12013), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U15058 ( .A1(n11273), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U15059 ( .A1(n11421), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12014), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U15060 ( .A1(n9576), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12016) );
  NAND4_X1 U15061 ( .A1(n12019), .A2(n12018), .A3(n12017), .A4(n12016), .ZN(
        n12020) );
  NOR2_X1 U15062 ( .A1(n12021), .A2(n12020), .ZN(n12042) );
  AOI22_X1 U15063 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12183), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12025) );
  AOI22_X1 U15064 ( .A1(n12101), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11421), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12024) );
  AOI22_X1 U15065 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12023) );
  AOI22_X1 U15066 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12022) );
  NAND4_X1 U15067 ( .A1(n12025), .A2(n12024), .A3(n12023), .A4(n12022), .ZN(
        n12031) );
  AOI22_X1 U15068 ( .A1(n12182), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U15069 ( .A1(n9576), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U15070 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U15071 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12026) );
  NAND4_X1 U15072 ( .A1(n12029), .A2(n12028), .A3(n12027), .A4(n12026), .ZN(
        n12030) );
  NOR2_X1 U15073 ( .A1(n12031), .A2(n12030), .ZN(n12041) );
  XNOR2_X1 U15074 ( .A(n12042), .B(n12041), .ZN(n12035) );
  INV_X1 U15075 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12032) );
  AOI21_X1 U15076 ( .B1(n12032), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12033) );
  AOI21_X1 U15077 ( .B1(n11713), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12033), .ZN(
        n12034) );
  OAI21_X1 U15078 ( .B1(n12167), .B2(n12035), .A(n12034), .ZN(n12039) );
  INV_X1 U15079 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14622) );
  OAI21_X1 U15080 ( .B1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n12037), .A(
        n12076), .ZN(n15971) );
  OR2_X1 U15081 ( .A1(n15971), .A2(n12170), .ZN(n12038) );
  NAND2_X1 U15082 ( .A1(n12039), .A2(n12038), .ZN(n14401) );
  NOR2_X1 U15083 ( .A1(n12042), .A2(n12041), .ZN(n12071) );
  AOI22_X1 U15084 ( .A1(n11273), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U15085 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U15086 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12044) );
  AOI22_X1 U15087 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12043) );
  NAND4_X1 U15088 ( .A1(n12046), .A2(n12045), .A3(n12044), .A4(n12043), .ZN(
        n12052) );
  AOI22_X1 U15089 ( .A1(n12101), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15090 ( .A1(n9576), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12049) );
  AOI22_X1 U15091 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12048) );
  AOI22_X1 U15092 ( .A1(n11421), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12047) );
  NAND4_X1 U15093 ( .A1(n12050), .A2(n12049), .A3(n12048), .A4(n12047), .ZN(
        n12051) );
  OR2_X1 U15094 ( .A1(n12052), .A2(n12051), .ZN(n12070) );
  INV_X1 U15095 ( .A(n12070), .ZN(n12053) );
  XNOR2_X1 U15096 ( .A(n12071), .B(n12053), .ZN(n12054) );
  INV_X1 U15097 ( .A(n12167), .ZN(n12193) );
  NAND2_X1 U15098 ( .A1(n12054), .A2(n12193), .ZN(n12058) );
  INV_X1 U15099 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14611) );
  OAI21_X1 U15100 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14611), .A(n12170), 
        .ZN(n12055) );
  AOI21_X1 U15101 ( .B1(n11713), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12055), .ZN(
        n12057) );
  XNOR2_X1 U15102 ( .A(n12076), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14615) );
  AOI21_X1 U15103 ( .B1(n12058), .B2(n12057), .A(n12056), .ZN(n14344) );
  AOI22_X1 U15104 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12063) );
  AOI22_X1 U15105 ( .A1(n12059), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12175), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15106 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12061) );
  AOI22_X1 U15107 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12060) );
  NAND4_X1 U15108 ( .A1(n12063), .A2(n12062), .A3(n12061), .A4(n12060), .ZN(
        n12069) );
  AOI22_X1 U15109 ( .A1(n11273), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U15110 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U15111 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12156), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U15112 ( .A1(n9576), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12064) );
  NAND4_X1 U15113 ( .A1(n12067), .A2(n12066), .A3(n12065), .A4(n12064), .ZN(
        n12068) );
  NOR2_X1 U15114 ( .A1(n12069), .A2(n12068), .ZN(n12084) );
  NAND2_X1 U15115 ( .A1(n12071), .A2(n12070), .ZN(n12083) );
  XNOR2_X1 U15116 ( .A(n12084), .B(n12083), .ZN(n12075) );
  NAND2_X1 U15117 ( .A1(n20679), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12072) );
  NAND2_X1 U15118 ( .A1(n12170), .A2(n12072), .ZN(n12073) );
  AOI21_X1 U15119 ( .B1(n11713), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12073), .ZN(
        n12074) );
  OAI21_X1 U15120 ( .B1(n12075), .B2(n12167), .A(n12074), .ZN(n12082) );
  INV_X1 U15121 ( .A(n12078), .ZN(n12079) );
  INV_X1 U15122 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14603) );
  NAND2_X1 U15123 ( .A1(n12079), .A2(n14603), .ZN(n12080) );
  AND2_X1 U15124 ( .A1(n12119), .A2(n12080), .ZN(n15830) );
  NAND2_X1 U15125 ( .A1(n15830), .A2(n12142), .ZN(n12081) );
  NOR2_X1 U15126 ( .A1(n12084), .A2(n12083), .ZN(n12114) );
  AOI22_X1 U15127 ( .A1(n11273), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12088) );
  AOI22_X1 U15128 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12087) );
  AOI22_X1 U15129 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U15130 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12085) );
  NAND4_X1 U15131 ( .A1(n12088), .A2(n12087), .A3(n12086), .A4(n12085), .ZN(
        n12094) );
  AOI22_X1 U15132 ( .A1(n12184), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U15133 ( .A1(n9576), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U15134 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12090) );
  AOI22_X1 U15135 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12089) );
  NAND4_X1 U15136 ( .A1(n12092), .A2(n12091), .A3(n12090), .A4(n12089), .ZN(
        n12093) );
  OR2_X1 U15137 ( .A1(n12094), .A2(n12093), .ZN(n12113) );
  XNOR2_X1 U15138 ( .A(n12114), .B(n12113), .ZN(n12098) );
  NAND2_X1 U15139 ( .A1(n20679), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12095) );
  NAND2_X1 U15140 ( .A1(n12170), .A2(n12095), .ZN(n12096) );
  AOI21_X1 U15141 ( .B1(n11713), .B2(P1_EAX_REG_26__SCAN_IN), .A(n12096), .ZN(
        n12097) );
  OAI21_X1 U15142 ( .B1(n12098), .B2(n12167), .A(n12097), .ZN(n12100) );
  XNOR2_X1 U15143 ( .A(n12119), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14592) );
  NAND2_X1 U15144 ( .A1(n14592), .A2(n12142), .ZN(n12099) );
  NAND2_X1 U15145 ( .A1(n12100), .A2(n12099), .ZN(n14330) );
  AOI22_X1 U15146 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12182), .B1(
        n12183), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U15147 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9576), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U15148 ( .A1(n12101), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12103) );
  AOI22_X1 U15149 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12102) );
  NAND4_X1 U15150 ( .A1(n12105), .A2(n12104), .A3(n12103), .A4(n12102), .ZN(
        n12112) );
  AOI22_X1 U15151 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12110) );
  AOI22_X1 U15152 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U15153 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12156), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15154 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12015), .B1(
        n11421), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12107) );
  NAND4_X1 U15155 ( .A1(n12110), .A2(n12109), .A3(n12108), .A4(n12107), .ZN(
        n12111) );
  NOR2_X1 U15156 ( .A1(n12112), .A2(n12111), .ZN(n12127) );
  NAND2_X1 U15157 ( .A1(n12114), .A2(n12113), .ZN(n12126) );
  XNOR2_X1 U15158 ( .A(n12127), .B(n12126), .ZN(n12118) );
  NAND2_X1 U15159 ( .A1(n20679), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12115) );
  NAND2_X1 U15160 ( .A1(n12170), .A2(n12115), .ZN(n12116) );
  AOI21_X1 U15161 ( .B1(n11713), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12116), .ZN(
        n12117) );
  OAI21_X1 U15162 ( .B1(n12118), .B2(n12167), .A(n12117), .ZN(n12124) );
  INV_X1 U15163 ( .A(n12119), .ZN(n12120) );
  NAND2_X1 U15164 ( .A1(n12120), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12121) );
  INV_X1 U15165 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14322) );
  NAND2_X1 U15166 ( .A1(n12121), .A2(n14322), .ZN(n12122) );
  NAND2_X1 U15167 ( .A1(n12146), .A2(n12122), .ZN(n14585) );
  INV_X1 U15168 ( .A(n14318), .ZN(n12125) );
  NOR2_X1 U15169 ( .A1(n12127), .A2(n12126), .ZN(n12164) );
  AOI22_X1 U15170 ( .A1(n11273), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U15171 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12130) );
  AOI22_X1 U15172 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U15173 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12128) );
  NAND4_X1 U15174 ( .A1(n12131), .A2(n12130), .A3(n12129), .A4(n12128), .ZN(
        n12137) );
  AOI22_X1 U15175 ( .A1(n12184), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U15176 ( .A1(n9576), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U15177 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15178 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12132) );
  NAND4_X1 U15179 ( .A1(n12135), .A2(n12134), .A3(n12133), .A4(n12132), .ZN(
        n12136) );
  OR2_X1 U15180 ( .A1(n12137), .A2(n12136), .ZN(n12163) );
  INV_X1 U15181 ( .A(n12163), .ZN(n12138) );
  XNOR2_X1 U15182 ( .A(n12164), .B(n12138), .ZN(n12139) );
  NAND2_X1 U15183 ( .A1(n12139), .A2(n12193), .ZN(n12145) );
  NAND2_X1 U15184 ( .A1(n20679), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12140) );
  NAND2_X1 U15185 ( .A1(n12170), .A2(n12140), .ZN(n12141) );
  AOI21_X1 U15186 ( .B1(n11713), .B2(P1_EAX_REG_28__SCAN_IN), .A(n12141), .ZN(
        n12144) );
  XNOR2_X1 U15187 ( .A(n12146), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14578) );
  INV_X1 U15188 ( .A(n12146), .ZN(n12147) );
  NAND2_X1 U15189 ( .A1(n12147), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12149) );
  INV_X1 U15190 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12148) );
  NAND2_X1 U15191 ( .A1(n12149), .A2(n12148), .ZN(n12150) );
  NAND2_X1 U15192 ( .A1(n12209), .A2(n12150), .ZN(n14561) );
  AOI22_X1 U15193 ( .A1(n12184), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U15194 ( .A1(n11419), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12153) );
  AOI22_X1 U15195 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9576), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U15196 ( .A1(n11273), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12151) );
  NAND4_X1 U15197 ( .A1(n12154), .A2(n12153), .A3(n12152), .A4(n12151), .ZN(
        n12162) );
  AOI22_X1 U15198 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12160) );
  AOI22_X1 U15199 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15200 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12156), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15201 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12157) );
  NAND4_X1 U15202 ( .A1(n12160), .A2(n12159), .A3(n12158), .A4(n12157), .ZN(
        n12161) );
  NOR2_X1 U15203 ( .A1(n12162), .A2(n12161), .ZN(n12172) );
  NAND2_X1 U15204 ( .A1(n12164), .A2(n12163), .ZN(n12171) );
  XNOR2_X1 U15205 ( .A(n12172), .B(n12171), .ZN(n12168) );
  AOI21_X1 U15206 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20679), .A(
        n11697), .ZN(n12166) );
  NAND2_X1 U15207 ( .A1(n12201), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12165) );
  OAI211_X1 U15208 ( .C1(n12168), .C2(n12167), .A(n12166), .B(n12165), .ZN(
        n12169) );
  OAI21_X1 U15209 ( .B1(n12170), .B2(n14561), .A(n12169), .ZN(n14302) );
  NOR2_X1 U15210 ( .A1(n12172), .A2(n12171), .ZN(n12192) );
  AOI22_X1 U15211 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15212 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15213 ( .A1(n12013), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15214 ( .A1(n12155), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12177), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12178) );
  NAND4_X1 U15215 ( .A1(n12181), .A2(n12180), .A3(n12179), .A4(n12178), .ZN(
        n12190) );
  AOI22_X1 U15216 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12182), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U15217 ( .A1(n20932), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12183), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12187) );
  AOI22_X1 U15218 ( .A1(n12184), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9576), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U15219 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12185) );
  NAND4_X1 U15220 ( .A1(n12188), .A2(n12187), .A3(n12186), .A4(n12185), .ZN(
        n12189) );
  NOR2_X1 U15221 ( .A1(n12190), .A2(n12189), .ZN(n12191) );
  XNOR2_X1 U15222 ( .A(n12192), .B(n12191), .ZN(n12194) );
  NAND2_X1 U15223 ( .A1(n12194), .A2(n12193), .ZN(n12199) );
  INV_X1 U15224 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12195) );
  AOI21_X1 U15225 ( .B1(n12195), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12196) );
  AOI21_X1 U15226 ( .B1(n11713), .B2(P1_EAX_REG_30__SCAN_IN), .A(n12196), .ZN(
        n12198) );
  XNOR2_X1 U15227 ( .A(n12209), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14549) );
  AOI21_X1 U15228 ( .B1(n12199), .B2(n12198), .A(n12197), .ZN(n14287) );
  NAND2_X1 U15229 ( .A1(n14300), .A2(n14287), .ZN(n12204) );
  AOI22_X1 U15230 ( .A1(n12201), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12200), .ZN(n12202) );
  AND2_X1 U15231 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12206) );
  NOR2_X1 U15232 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20620), .ZN(n12205) );
  NAND2_X1 U15233 ( .A1(n14281), .A2(n16031), .ZN(n12216) );
  INV_X1 U15234 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n20885) );
  NAND2_X1 U15235 ( .A1(n12212), .A2(n20620), .ZN(n20758) );
  NAND2_X1 U15236 ( .A1(n20758), .A2(n20676), .ZN(n12207) );
  NAND2_X1 U15237 ( .A1(n20676), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15785) );
  NAND2_X1 U15238 ( .A1(n20777), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12208) );
  NAND2_X1 U15239 ( .A1(n15785), .A2(n12208), .ZN(n20057) );
  INV_X1 U15240 ( .A(n12209), .ZN(n12210) );
  NAND2_X1 U15241 ( .A1(n12210), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12211) );
  NAND2_X1 U15242 ( .A1(n16007), .A2(n13807), .ZN(n12213) );
  INV_X2 U15243 ( .A(n16041), .ZN(n16139) );
  NAND2_X1 U15244 ( .A1(n16139), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14670) );
  OAI211_X1 U15245 ( .C1(n20885), .C2(n16039), .A(n12213), .B(n14670), .ZN(
        n12214) );
  OAI211_X1 U15246 ( .C1(n9563), .C2(n19879), .A(n12216), .B(n12215), .ZN(
        P1_U2968) );
  NAND2_X1 U15247 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20691) );
  INV_X1 U15248 ( .A(n20691), .ZN(n20762) );
  NAND2_X1 U15249 ( .A1(n13100), .A2(n13213), .ZN(n13344) );
  OAI21_X1 U15250 ( .B1(n12217), .B2(n20762), .A(n13344), .ZN(n12218) );
  NAND2_X1 U15251 ( .A1(n13364), .A2(n12218), .ZN(n13368) );
  INV_X1 U15252 ( .A(n13332), .ZN(n13588) );
  AND3_X1 U15253 ( .A1(n12221), .A2(n12220), .A3(n12219), .ZN(n12224) );
  OAI21_X1 U15254 ( .B1(n12224), .B2(n12223), .A(n12222), .ZN(n13219) );
  NAND3_X1 U15255 ( .A1(n13588), .A2(n13219), .A3(n20691), .ZN(n13365) );
  INV_X1 U15256 ( .A(n20134), .ZN(n13380) );
  AND2_X1 U15257 ( .A1(n13365), .A2(n12225), .ZN(n12226) );
  AND2_X1 U15258 ( .A1(n14540), .A2(n13380), .ZN(n12227) );
  NOR4_X1 U15259 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n12231) );
  NOR4_X1 U15260 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n12230) );
  NOR4_X1 U15261 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n12229) );
  NOR4_X1 U15262 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n12228) );
  AND4_X1 U15263 ( .A1(n12231), .A2(n12230), .A3(n12229), .A4(n12228), .ZN(
        n12237) );
  NOR4_X1 U15264 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12235) );
  NOR4_X1 U15265 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n12234) );
  NOR4_X1 U15266 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n12233) );
  INV_X1 U15267 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n12232) );
  AND4_X1 U15268 ( .A1(n12235), .A2(n12234), .A3(n12233), .A4(n12232), .ZN(
        n12236) );
  NAND2_X1 U15269 ( .A1(n12237), .A2(n12236), .ZN(n12238) );
  INV_X2 U15270 ( .A(n20079), .ZN(n20080) );
  NOR2_X1 U15271 ( .A1(n13385), .A2(n20080), .ZN(n12239) );
  NAND2_X1 U15272 ( .A1(n14540), .A2(n12239), .ZN(n15964) );
  INV_X1 U15273 ( .A(n15964), .ZN(n12240) );
  AOI22_X1 U15274 ( .A1(n12240), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n15957), .ZN(n12243) );
  NAND2_X1 U15275 ( .A1(n14540), .A2(n12241), .ZN(n13392) );
  INV_X1 U15276 ( .A(DATAI_31_), .ZN(n12242) );
  AND2_X1 U15277 ( .A1(n12243), .A2(n10055), .ZN(n12244) );
  NAND2_X1 U15278 ( .A1(n12246), .A2(n12629), .ZN(n12251) );
  INV_X1 U15279 ( .A(n12247), .ZN(n12248) );
  AND2_X1 U15280 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19388) );
  NOR2_X1 U15281 ( .A1(n19819), .A2(n19828), .ZN(n19605) );
  NAND2_X1 U15282 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19605), .ZN(
        n19186) );
  OAI21_X1 U15283 ( .B1(n19388), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n19186), .ZN(n19321) );
  NOR2_X1 U15284 ( .A1(n19321), .A2(n19609), .ZN(n12249) );
  AOI21_X1 U15285 ( .B1(n12263), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12249), .ZN(n12250) );
  NAND2_X1 U15286 ( .A1(n12251), .A2(n12250), .ZN(n12253) );
  INV_X1 U15287 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12456) );
  NOR2_X1 U15288 ( .A1(n12277), .A2(n12456), .ZN(n12252) );
  NAND2_X1 U15289 ( .A1(n12253), .A2(n12252), .ZN(n13323) );
  AOI22_X1 U15290 ( .A1(n12263), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19802), .B2(n19837), .ZN(n12254) );
  INV_X1 U15291 ( .A(n12277), .ZN(n12516) );
  NAND2_X1 U15292 ( .A1(n12516), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12258) );
  XNOR2_X1 U15293 ( .A(n15584), .B(n12258), .ZN(n13235) );
  NAND2_X1 U15294 ( .A1(n12263), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12256) );
  NAND2_X1 U15295 ( .A1(n19828), .A2(n19837), .ZN(n19445) );
  INV_X1 U15296 ( .A(n19445), .ZN(n19322) );
  NOR2_X1 U15297 ( .A1(n19388), .A2(n19322), .ZN(n19320) );
  NAND2_X1 U15298 ( .A1(n19320), .A2(n19802), .ZN(n19496) );
  NAND2_X1 U15299 ( .A1(n12256), .A2(n19496), .ZN(n12257) );
  NAND2_X1 U15300 ( .A1(n13235), .A2(n13234), .ZN(n13237) );
  INV_X1 U15301 ( .A(n15584), .ZN(n12259) );
  NAND2_X1 U15302 ( .A1(n12259), .A2(n12258), .ZN(n12260) );
  NAND3_X1 U15303 ( .A1(n13322), .A2(n13323), .A3(n13325), .ZN(n13324) );
  NOR2_X1 U15304 ( .A1(n19819), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19390) );
  INV_X1 U15305 ( .A(n19452), .ZN(n19449) );
  NAND2_X1 U15306 ( .A1(n19186), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12262) );
  AOI21_X1 U15307 ( .B1(n19449), .B2(n12262), .A(n19609), .ZN(n19546) );
  AOI21_X1 U15308 ( .B1(n12263), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19546), .ZN(n12264) );
  INV_X1 U15309 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12482) );
  NOR2_X1 U15310 ( .A1(n12277), .A2(n12482), .ZN(n12266) );
  AND2_X2 U15311 ( .A1(n12267), .A2(n12268), .ZN(n13460) );
  NAND2_X1 U15312 ( .A1(n13461), .A2(n13460), .ZN(n13462) );
  INV_X1 U15313 ( .A(n13636), .ZN(n13638) );
  NAND2_X1 U15314 ( .A1(n12269), .A2(n13682), .ZN(n12272) );
  NAND2_X1 U15315 ( .A1(n12271), .A2(n12270), .ZN(n13650) );
  NOR2_X1 U15316 ( .A1(n12272), .A2(n13650), .ZN(n12273) );
  AND2_X1 U15317 ( .A1(n13638), .A2(n12273), .ZN(n13710) );
  AND2_X1 U15318 ( .A1(n13751), .A2(n13710), .ZN(n12276) );
  INV_X1 U15319 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12274) );
  OR2_X1 U15320 ( .A1(n12274), .A2(n13601), .ZN(n12275) );
  INV_X1 U15321 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13539) );
  NOR2_X1 U15322 ( .A1(n12275), .A2(n13539), .ZN(n13634) );
  AND2_X1 U15323 ( .A1(n12276), .A2(n13634), .ZN(n12278) );
  INV_X1 U15324 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12506) );
  NOR2_X1 U15325 ( .A1(n12277), .A2(n12506), .ZN(n13518) );
  AOI22_X1 U15326 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12285) );
  AOI22_X1 U15327 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12284) );
  AOI22_X1 U15328 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12283) );
  AOI22_X1 U15329 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12282) );
  NAND4_X1 U15330 ( .A1(n12285), .A2(n12284), .A3(n12283), .A4(n12282), .ZN(
        n12294) );
  AOI22_X1 U15331 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10341), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12292) );
  INV_X1 U15332 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12287) );
  INV_X1 U15333 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12286) );
  OAI22_X1 U15334 ( .A1(n12367), .A2(n12287), .B1(n12364), .B2(n12286), .ZN(
        n12288) );
  AOI21_X1 U15335 ( .B1(n10376), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n12288), .ZN(n12291) );
  AOI22_X1 U15336 ( .A1(n11071), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12290) );
  NAND2_X1 U15337 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12289) );
  NAND4_X1 U15338 ( .A1(n12292), .A2(n12291), .A3(n12290), .A4(n12289), .ZN(
        n12293) );
  NAND2_X1 U15339 ( .A1(n13995), .A2(n13994), .ZN(n13962) );
  AOI22_X1 U15340 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15341 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U15342 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12296) );
  AOI22_X1 U15343 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n12394), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12295) );
  NAND4_X1 U15344 ( .A1(n12298), .A2(n12297), .A3(n12296), .A4(n12295), .ZN(
        n12307) );
  AOI22_X1 U15345 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10341), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12305) );
  INV_X1 U15346 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12300) );
  OAI22_X1 U15347 ( .A1(n12367), .A2(n12300), .B1(n12299), .B2(n12364), .ZN(
        n12301) );
  AOI21_X1 U15348 ( .B1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n10376), .A(
        n12301), .ZN(n12304) );
  AOI22_X1 U15349 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11071), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12303) );
  NAND2_X1 U15350 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12302) );
  NAND4_X1 U15351 ( .A1(n12305), .A2(n12304), .A3(n12303), .A4(n12302), .ZN(
        n12306) );
  AOI22_X1 U15352 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U15353 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12310) );
  AOI22_X1 U15354 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U15355 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n12394), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12308) );
  NAND4_X1 U15356 ( .A1(n12311), .A2(n12310), .A3(n12309), .A4(n12308), .ZN(
        n12320) );
  AOI22_X1 U15357 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10341), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12318) );
  INV_X1 U15358 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12313) );
  INV_X1 U15359 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12312) );
  OAI22_X1 U15360 ( .A1(n12367), .A2(n12313), .B1(n12312), .B2(n12364), .ZN(
        n12314) );
  AOI21_X1 U15361 ( .B1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B2(n10376), .A(
        n12314), .ZN(n12317) );
  AOI22_X1 U15362 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11071), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12316) );
  NAND2_X1 U15363 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12315) );
  NAND4_X1 U15364 ( .A1(n12318), .A2(n12317), .A3(n12316), .A4(n12315), .ZN(
        n12319) );
  NOR2_X1 U15365 ( .A1(n12320), .A2(n12319), .ZN(n15017) );
  AOI22_X1 U15366 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12325) );
  AOI22_X1 U15367 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12324) );
  AOI22_X1 U15368 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12323) );
  AOI22_X1 U15369 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12322) );
  NAND4_X1 U15370 ( .A1(n12325), .A2(n12324), .A3(n12323), .A4(n12322), .ZN(
        n12334) );
  AOI22_X1 U15371 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10341), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12332) );
  INV_X1 U15372 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12327) );
  OAI22_X1 U15373 ( .A1(n12367), .A2(n12327), .B1(n12364), .B2(n12326), .ZN(
        n12328) );
  AOI21_X1 U15374 ( .B1(n10376), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n12328), .ZN(n12331) );
  AOI22_X1 U15375 ( .A1(n11071), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12330) );
  NAND2_X1 U15376 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12329) );
  NAND4_X1 U15377 ( .A1(n12332), .A2(n12331), .A3(n12330), .A4(n12329), .ZN(
        n12333) );
  AOI22_X1 U15378 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U15379 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U15380 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U15381 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12335) );
  NAND4_X1 U15382 ( .A1(n12338), .A2(n12337), .A3(n12336), .A4(n12335), .ZN(
        n12346) );
  AOI22_X1 U15383 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10341), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12344) );
  INV_X1 U15384 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12339) );
  OAI22_X1 U15385 ( .A1(n12367), .A2(n12339), .B1(n12364), .B2(n20779), .ZN(
        n12340) );
  AOI21_X1 U15386 ( .B1(n10376), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n12340), .ZN(n12343) );
  AOI22_X1 U15387 ( .A1(n11071), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12342) );
  NAND2_X1 U15388 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12341) );
  NAND4_X1 U15389 ( .A1(n12344), .A2(n12343), .A3(n12342), .A4(n12341), .ZN(
        n12345) );
  OR2_X1 U15390 ( .A1(n12346), .A2(n12345), .ZN(n15005) );
  NAND2_X1 U15391 ( .A1(n14019), .A2(n15005), .ZN(n15000) );
  AOI22_X1 U15392 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12350) );
  AOI22_X1 U15393 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12349) );
  AOI22_X1 U15394 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12348) );
  AOI22_X1 U15395 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12347) );
  NAND4_X1 U15396 ( .A1(n12350), .A2(n12349), .A3(n12348), .A4(n12347), .ZN(
        n12359) );
  AOI22_X1 U15397 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10341), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12357) );
  INV_X1 U15398 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12352) );
  OAI22_X1 U15399 ( .A1(n12367), .A2(n12352), .B1(n12364), .B2(n12351), .ZN(
        n12353) );
  AOI21_X1 U15400 ( .B1(n10376), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n12353), .ZN(n12356) );
  AOI22_X1 U15401 ( .A1(n11071), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12355) );
  NAND2_X1 U15402 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12354) );
  NAND4_X1 U15403 ( .A1(n12357), .A2(n12356), .A3(n12355), .A4(n12354), .ZN(
        n12358) );
  NOR2_X1 U15404 ( .A1(n12359), .A2(n12358), .ZN(n15001) );
  OR2_X2 U15405 ( .A1(n15000), .A2(n15001), .ZN(n15003) );
  AOI22_X1 U15406 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12363) );
  AOI22_X1 U15407 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U15408 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U15409 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12394), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12360) );
  NAND4_X1 U15410 ( .A1(n12363), .A2(n12362), .A3(n12361), .A4(n12360), .ZN(
        n12374) );
  AOI22_X1 U15411 ( .A1(n10389), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10341), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12372) );
  INV_X1 U15412 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12366) );
  OAI22_X1 U15413 ( .A1(n12367), .A2(n12366), .B1(n12365), .B2(n12364), .ZN(
        n12368) );
  AOI21_X1 U15414 ( .B1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B2(n10376), .A(
        n12368), .ZN(n12371) );
  AOI22_X1 U15415 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11071), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12370) );
  NAND2_X1 U15416 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12369) );
  NAND4_X1 U15417 ( .A1(n12372), .A2(n12371), .A3(n12370), .A4(n12369), .ZN(
        n12373) );
  NOR2_X1 U15418 ( .A1(n12374), .A2(n12373), .ZN(n14996) );
  NOR2_X4 U15419 ( .A1(n15003), .A2(n14996), .ZN(n14995) );
  AOI22_X1 U15420 ( .A1(n11071), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n12375), .ZN(n12379) );
  AOI22_X1 U15421 ( .A1(n11072), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n9567), .ZN(n12378) );
  NAND2_X1 U15422 ( .A1(n10376), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12377) );
  NAND2_X1 U15423 ( .A1(n10331), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12376) );
  NAND4_X1 U15424 ( .A1(n12379), .A2(n12378), .A3(n12377), .A4(n12376), .ZN(
        n12382) );
  INV_X1 U15425 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12380) );
  OAI22_X1 U15426 ( .A1(n12380), .A2(n11055), .B1(n10538), .B2(n12568), .ZN(
        n12381) );
  NOR2_X1 U15427 ( .A1(n12382), .A2(n12381), .ZN(n12398) );
  INV_X1 U15428 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12386) );
  INV_X1 U15429 ( .A(n12383), .ZN(n12385) );
  OAI22_X1 U15430 ( .A1(n12387), .A2(n12386), .B1(n12385), .B2(n12384), .ZN(
        n12392) );
  INV_X1 U15431 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12390) );
  INV_X1 U15432 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12388) );
  OAI22_X1 U15433 ( .A1(n12390), .A2(n12389), .B1(n10537), .B2(n12388), .ZN(
        n12391) );
  NOR2_X1 U15434 ( .A1(n12392), .A2(n12391), .ZN(n12397) );
  AOI22_X1 U15435 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n12393), .B1(
        n10389), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12396) );
  AOI22_X1 U15436 ( .A1(n10422), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12394), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12395) );
  NAND4_X1 U15437 ( .A1(n12398), .A2(n12397), .A3(n12396), .A4(n12395), .ZN(
        n12419) );
  AOI22_X1 U15438 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12569), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12407) );
  AOI22_X1 U15439 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12406) );
  AOI22_X1 U15440 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12420), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12405) );
  INV_X1 U15441 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n19526) );
  INV_X1 U15442 ( .A(n12575), .ZN(n12547) );
  INV_X1 U15443 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12400) );
  OR2_X1 U15444 ( .A1(n12547), .A2(n12400), .ZN(n12402) );
  AOI21_X1 U15445 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n12401), .ZN(n12565) );
  OAI211_X1 U15446 ( .C1(n12399), .C2(n19526), .A(n12402), .B(n12565), .ZN(
        n12403) );
  INV_X1 U15447 ( .A(n12403), .ZN(n12404) );
  NAND4_X1 U15448 ( .A1(n12407), .A2(n12406), .A3(n12405), .A4(n12404), .ZN(
        n12415) );
  AOI22_X1 U15449 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12569), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12413) );
  AOI22_X1 U15450 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12412) );
  AOI22_X1 U15451 ( .A1(n10308), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12420), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12411) );
  NAND2_X1 U15452 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12409) );
  AOI21_X1 U15453 ( .B1(n12575), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        n12565), .ZN(n12408) );
  AND2_X1 U15454 ( .A1(n12409), .A2(n12408), .ZN(n12410) );
  NAND4_X1 U15455 ( .A1(n12413), .A2(n12412), .A3(n12411), .A4(n12410), .ZN(
        n12414) );
  NAND2_X1 U15456 ( .A1(n12415), .A2(n12414), .ZN(n12442) );
  NOR2_X1 U15457 ( .A1(n12416), .A2(n12442), .ZN(n12417) );
  XOR2_X1 U15458 ( .A(n12419), .B(n12417), .Z(n12440) );
  INV_X1 U15459 ( .A(n12442), .ZN(n12418) );
  NAND2_X1 U15460 ( .A1(n19853), .A2(n12418), .ZN(n14987) );
  NAND2_X1 U15461 ( .A1(n12419), .A2(n12418), .ZN(n12445) );
  AOI22_X1 U15462 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12569), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12428) );
  AOI22_X1 U15463 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12427) );
  AOI22_X1 U15464 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12426) );
  INV_X1 U15465 ( .A(n12420), .ZN(n12578) );
  INV_X1 U15466 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12423) );
  INV_X1 U15467 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12421) );
  OR2_X1 U15468 ( .A1(n12547), .A2(n12421), .ZN(n12422) );
  OAI211_X1 U15469 ( .C1(n12578), .C2(n12423), .A(n12422), .B(n12565), .ZN(
        n12424) );
  INV_X1 U15470 ( .A(n12424), .ZN(n12425) );
  NAND4_X1 U15471 ( .A1(n12428), .A2(n12427), .A3(n12426), .A4(n12425), .ZN(
        n12438) );
  AOI22_X1 U15472 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12569), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U15473 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12435) );
  AOI22_X1 U15474 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12434) );
  OR2_X1 U15475 ( .A1(n12547), .A2(n12429), .ZN(n12430) );
  INV_X1 U15476 ( .A(n12565), .ZN(n12574) );
  OAI211_X1 U15477 ( .C1(n12578), .C2(n12431), .A(n12430), .B(n12574), .ZN(
        n12432) );
  INV_X1 U15478 ( .A(n12432), .ZN(n12433) );
  NAND4_X1 U15479 ( .A1(n12436), .A2(n12435), .A3(n12434), .A4(n12433), .ZN(
        n12437) );
  NAND2_X1 U15480 ( .A1(n12438), .A2(n12437), .ZN(n12441) );
  XOR2_X1 U15481 ( .A(n12445), .B(n12441), .Z(n12439) );
  NAND2_X1 U15482 ( .A1(n12439), .A2(n12516), .ZN(n14980) );
  INV_X1 U15483 ( .A(n12440), .ZN(n12443) );
  INV_X1 U15484 ( .A(n12441), .ZN(n12446) );
  NAND2_X1 U15485 ( .A1(n19853), .A2(n12446), .ZN(n14982) );
  NOR3_X1 U15486 ( .A1(n12443), .A2(n12442), .A3(n14982), .ZN(n12444) );
  INV_X1 U15487 ( .A(n12445), .ZN(n12447) );
  AND2_X1 U15488 ( .A1(n12447), .A2(n12446), .ZN(n12466) );
  AOI22_X1 U15489 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12569), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U15490 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U15491 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12453) );
  INV_X1 U15492 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12448) );
  OR2_X1 U15493 ( .A1(n12547), .A2(n12448), .ZN(n12449) );
  OAI211_X1 U15494 ( .C1(n12578), .C2(n12450), .A(n12449), .B(n12565), .ZN(
        n12451) );
  INV_X1 U15495 ( .A(n12451), .ZN(n12452) );
  NAND4_X1 U15496 ( .A1(n12455), .A2(n12454), .A3(n12453), .A4(n12452), .ZN(
        n12465) );
  AOI22_X1 U15497 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12569), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12463) );
  AOI22_X1 U15498 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12462) );
  AOI22_X1 U15499 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12461) );
  INV_X1 U15500 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12458) );
  OR2_X1 U15501 ( .A1(n12547), .A2(n12456), .ZN(n12457) );
  OAI211_X1 U15502 ( .C1(n12578), .C2(n12458), .A(n12457), .B(n12574), .ZN(
        n12459) );
  INV_X1 U15503 ( .A(n12459), .ZN(n12460) );
  NAND4_X1 U15504 ( .A1(n12463), .A2(n12462), .A3(n12461), .A4(n12460), .ZN(
        n12464) );
  AND2_X1 U15505 ( .A1(n12465), .A2(n12464), .ZN(n12467) );
  NAND2_X1 U15506 ( .A1(n12466), .A2(n12467), .ZN(n12495) );
  OAI211_X1 U15507 ( .C1(n12466), .C2(n12467), .A(n12516), .B(n12495), .ZN(
        n12470) );
  INV_X1 U15508 ( .A(n12467), .ZN(n12468) );
  NOR2_X1 U15509 ( .A1(n13037), .A2(n12468), .ZN(n14974) );
  INV_X1 U15510 ( .A(n12469), .ZN(n12472) );
  AOI22_X1 U15511 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12569), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12481) );
  AOI22_X1 U15512 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12480) );
  AOI22_X1 U15513 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12479) );
  INV_X1 U15514 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12474) );
  OR2_X1 U15515 ( .A1(n12547), .A2(n12474), .ZN(n12475) );
  OAI211_X1 U15516 ( .C1(n12578), .C2(n12476), .A(n12475), .B(n12565), .ZN(
        n12477) );
  INV_X1 U15517 ( .A(n12477), .ZN(n12478) );
  NAND4_X1 U15518 ( .A1(n12481), .A2(n12480), .A3(n12479), .A4(n12478), .ZN(
        n12491) );
  AOI22_X1 U15519 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12569), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12489) );
  AOI22_X1 U15520 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12488) );
  AOI22_X1 U15521 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12487) );
  OR2_X1 U15522 ( .A1(n12547), .A2(n12482), .ZN(n12483) );
  OAI211_X1 U15523 ( .C1(n12578), .C2(n12484), .A(n12483), .B(n12574), .ZN(
        n12485) );
  INV_X1 U15524 ( .A(n12485), .ZN(n12486) );
  NAND4_X1 U15525 ( .A1(n12489), .A2(n12488), .A3(n12487), .A4(n12486), .ZN(
        n12490) );
  AND2_X1 U15526 ( .A1(n12491), .A2(n12490), .ZN(n12496) );
  XNOR2_X1 U15527 ( .A(n12495), .B(n12496), .ZN(n12492) );
  XNOR2_X2 U15528 ( .A(n12493), .B(n10061), .ZN(n14970) );
  NAND2_X1 U15529 ( .A1(n19853), .A2(n12496), .ZN(n14969) );
  INV_X1 U15530 ( .A(n12495), .ZN(n12497) );
  AND2_X1 U15531 ( .A1(n12497), .A2(n12496), .ZN(n12517) );
  AOI22_X1 U15532 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12569), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12505) );
  AOI22_X1 U15533 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12504) );
  AOI22_X1 U15534 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12503) );
  OR2_X1 U15535 ( .A1(n12547), .A2(n12498), .ZN(n12499) );
  OAI211_X1 U15536 ( .C1(n12578), .C2(n12500), .A(n12499), .B(n12565), .ZN(
        n12501) );
  INV_X1 U15537 ( .A(n12501), .ZN(n12502) );
  NAND4_X1 U15538 ( .A1(n12505), .A2(n12504), .A3(n12503), .A4(n12502), .ZN(
        n12515) );
  AOI22_X1 U15539 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12569), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12513) );
  AOI22_X1 U15540 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12512) );
  AOI22_X1 U15541 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12511) );
  INV_X1 U15542 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12508) );
  OR2_X1 U15543 ( .A1(n12547), .A2(n12506), .ZN(n12507) );
  OAI211_X1 U15544 ( .C1(n12578), .C2(n12508), .A(n12507), .B(n12574), .ZN(
        n12509) );
  INV_X1 U15545 ( .A(n12509), .ZN(n12510) );
  NAND4_X1 U15546 ( .A1(n12513), .A2(n12512), .A3(n12511), .A4(n12510), .ZN(
        n12514) );
  AND2_X1 U15547 ( .A1(n12515), .A2(n12514), .ZN(n12519) );
  NAND2_X1 U15548 ( .A1(n12517), .A2(n12519), .ZN(n14954) );
  OAI211_X1 U15549 ( .C1(n12517), .C2(n12519), .A(n14954), .B(n12516), .ZN(
        n12518) );
  INV_X1 U15550 ( .A(n12519), .ZN(n12520) );
  NOR2_X1 U15551 ( .A1(n13037), .A2(n12520), .ZN(n14960) );
  AOI22_X1 U15552 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12569), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12529) );
  AOI22_X1 U15553 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12528) );
  AOI22_X1 U15554 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12527) );
  OR2_X1 U15555 ( .A1(n12547), .A2(n12522), .ZN(n12523) );
  OAI211_X1 U15556 ( .C1(n12578), .C2(n12524), .A(n12523), .B(n12565), .ZN(
        n12525) );
  INV_X1 U15557 ( .A(n12525), .ZN(n12526) );
  NAND4_X1 U15558 ( .A1(n12529), .A2(n12528), .A3(n12527), .A4(n12526), .ZN(
        n12538) );
  AOI22_X1 U15559 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12569), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12536) );
  AOI22_X1 U15560 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12535) );
  AOI22_X1 U15561 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12534) );
  OR2_X1 U15562 ( .A1(n12547), .A2(n13539), .ZN(n12530) );
  OAI211_X1 U15563 ( .C1(n12578), .C2(n12531), .A(n12530), .B(n12574), .ZN(
        n12532) );
  INV_X1 U15564 ( .A(n12532), .ZN(n12533) );
  NAND4_X1 U15565 ( .A1(n12536), .A2(n12535), .A3(n12534), .A4(n12533), .ZN(
        n12537) );
  NAND2_X1 U15566 ( .A1(n12538), .A2(n12537), .ZN(n12557) );
  AOI21_X2 U15567 ( .B1(n14959), .B2(n10017), .A(n12557), .ZN(n14950) );
  AOI22_X1 U15568 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12569), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12546) );
  AOI22_X1 U15569 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12545) );
  AOI22_X1 U15570 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12544) );
  OR2_X1 U15571 ( .A1(n12547), .A2(n12539), .ZN(n12540) );
  OAI211_X1 U15572 ( .C1(n12578), .C2(n12541), .A(n12540), .B(n12565), .ZN(
        n12542) );
  INV_X1 U15573 ( .A(n12542), .ZN(n12543) );
  NAND4_X1 U15574 ( .A1(n12546), .A2(n12545), .A3(n12544), .A4(n12543), .ZN(
        n12556) );
  AOI22_X1 U15575 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12571), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12554) );
  AOI22_X1 U15576 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12553) );
  AOI22_X1 U15577 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12552) );
  INV_X1 U15578 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12549) );
  OR2_X1 U15579 ( .A1(n12547), .A2(n13601), .ZN(n12548) );
  OAI211_X1 U15580 ( .C1(n12578), .C2(n12549), .A(n12548), .B(n12574), .ZN(
        n12550) );
  INV_X1 U15581 ( .A(n12550), .ZN(n12551) );
  NAND4_X1 U15582 ( .A1(n12554), .A2(n12553), .A3(n12552), .A4(n12551), .ZN(
        n12555) );
  NAND2_X1 U15583 ( .A1(n12556), .A2(n12555), .ZN(n12560) );
  INV_X1 U15584 ( .A(n12557), .ZN(n14955) );
  NAND2_X1 U15585 ( .A1(n19196), .A2(n14955), .ZN(n12558) );
  OR2_X1 U15586 ( .A1(n14954), .A2(n12558), .ZN(n12559) );
  NOR2_X1 U15587 ( .A1(n12559), .A2(n12560), .ZN(n12561) );
  AOI21_X1 U15588 ( .B1(n12560), .B2(n12559), .A(n12561), .ZN(n14949) );
  NAND2_X1 U15589 ( .A1(n14950), .A2(n14949), .ZN(n14951) );
  INV_X1 U15590 ( .A(n12561), .ZN(n12562) );
  NAND2_X1 U15591 ( .A1(n14951), .A2(n12562), .ZN(n12585) );
  AOI22_X1 U15592 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12571), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U15593 ( .A1(n10308), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12563) );
  NAND2_X1 U15594 ( .A1(n12564), .A2(n12563), .ZN(n12583) );
  AOI22_X1 U15595 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10310), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12567) );
  AOI21_X1 U15596 ( .B1(n12575), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n12565), .ZN(n12566) );
  OAI211_X1 U15597 ( .C1(n12578), .C2(n12568), .A(n12567), .B(n12566), .ZN(
        n12582) );
  AOI22_X1 U15598 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12569), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12573) );
  AOI22_X1 U15599 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12572) );
  NAND2_X1 U15600 ( .A1(n12573), .A2(n12572), .ZN(n12581) );
  INV_X1 U15601 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12579) );
  AOI22_X1 U15602 ( .A1(n10310), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10308), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12577) );
  AOI21_X1 U15603 ( .B1(n12575), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n12574), .ZN(n12576) );
  OAI211_X1 U15604 ( .C1(n12579), .C2(n12578), .A(n12577), .B(n12576), .ZN(
        n12580) );
  OAI22_X1 U15605 ( .A1(n12583), .A2(n12582), .B1(n12581), .B2(n12580), .ZN(
        n12584) );
  XNOR2_X1 U15606 ( .A(n12585), .B(n12584), .ZN(n12959) );
  OR2_X1 U15607 ( .A1(n16310), .A2(n12586), .ZN(n16318) );
  NAND2_X1 U15608 ( .A1(n12587), .A2(n19711), .ZN(n16315) );
  NOR2_X1 U15609 ( .A1(n16318), .A2(n16315), .ZN(n12588) );
  AOI21_X1 U15610 ( .B1(n16314), .B2(n16309), .A(n12588), .ZN(n13164) );
  NAND2_X1 U15611 ( .A1(n13164), .A2(n12589), .ZN(n12590) );
  NAND2_X1 U15612 ( .A1(n12959), .A2(n19100), .ZN(n12609) );
  AOI22_X1 U15613 ( .A1(n14205), .A2(n19111), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n19110), .ZN(n12608) );
  NOR4_X1 U15614 ( .A1(P2_ADDRESS_REG_16__SCAN_IN), .A2(
        P2_ADDRESS_REG_15__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n12596) );
  NOR4_X1 U15615 ( .A1(P2_ADDRESS_REG_21__SCAN_IN), .A2(
        P2_ADDRESS_REG_20__SCAN_IN), .A3(P2_ADDRESS_REG_19__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n12595) );
  NOR4_X1 U15616 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_6__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12594) );
  NOR4_X1 U15617 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n12593) );
  NAND4_X1 U15618 ( .A1(n12596), .A2(n12595), .A3(n12594), .A4(n12593), .ZN(
        n12601) );
  NOR4_X1 U15619 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n12599) );
  NOR4_X1 U15620 ( .A1(P2_ADDRESS_REG_25__SCAN_IN), .A2(
        P2_ADDRESS_REG_24__SCAN_IN), .A3(P2_ADDRESS_REG_23__SCAN_IN), .A4(
        P2_ADDRESS_REG_22__SCAN_IN), .ZN(n12598) );
  NOR4_X1 U15621 ( .A1(P2_ADDRESS_REG_4__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_27__SCAN_IN), .A4(
        P2_ADDRESS_REG_26__SCAN_IN), .ZN(n12597) );
  INV_X1 U15622 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19745) );
  NAND4_X1 U15623 ( .A1(n12599), .A2(n12598), .A3(n12597), .A4(n19745), .ZN(
        n12600) );
  OAI21_X1 U15624 ( .B1(n12601), .B2(n12600), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12602) );
  NAND2_X1 U15625 ( .A1(n13674), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12604) );
  INV_X1 U15626 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14042) );
  OR2_X1 U15627 ( .A1(n13674), .A2(n14042), .ZN(n12603) );
  NAND2_X1 U15628 ( .A1(n12604), .A2(n12603), .ZN(n19063) );
  NAND2_X1 U15629 ( .A1(n19050), .A2(n19063), .ZN(n12607) );
  AND2_X1 U15630 ( .A1(n19213), .A2(n9583), .ZN(n12605) );
  AOI22_X1 U15631 ( .A1(n19052), .A2(BUF2_REG_30__SCAN_IN), .B1(n19051), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n12606) );
  NAND2_X1 U15632 ( .A1(n12609), .A2(n10062), .ZN(P2_U2889) );
  NAND2_X1 U15633 ( .A1(n12611), .A2(n12610), .ZN(n12624) );
  NAND2_X1 U15634 ( .A1(n15217), .A2(n15215), .ZN(n12613) );
  INV_X1 U15635 ( .A(n16200), .ZN(n12614) );
  INV_X1 U15636 ( .A(n15205), .ZN(n12615) );
  INV_X1 U15637 ( .A(n12616), .ZN(n15196) );
  NAND2_X1 U15638 ( .A1(n12619), .A2(n12618), .ZN(n15188) );
  INV_X1 U15639 ( .A(n12620), .ZN(n12622) );
  INV_X1 U15640 ( .A(n15171), .ZN(n12621) );
  XOR2_X1 U15641 ( .A(n12624), .B(n12623), .Z(n15347) );
  AND2_X1 U15642 ( .A1(n19852), .A2(n13167), .ZN(n13020) );
  INV_X1 U15643 ( .A(n13020), .ZN(n12625) );
  INV_X1 U15644 ( .A(n18832), .ZN(n12627) );
  NAND2_X1 U15645 ( .A1(n12627), .A2(n13037), .ZN(n16243) );
  NAND2_X1 U15646 ( .A1(n15347), .A2(n19167), .ZN(n12642) );
  NAND2_X1 U15647 ( .A1(n19712), .A2(n10900), .ZN(n15600) );
  INV_X1 U15648 ( .A(n15600), .ZN(n19801) );
  OR2_X1 U15649 ( .A1(n19802), .A2(n19801), .ZN(n19820) );
  NAND2_X1 U15650 ( .A1(n19820), .A2(n18828), .ZN(n12628) );
  INV_X1 U15651 ( .A(n12629), .ZN(n12631) );
  INV_X1 U15652 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19446) );
  NAND2_X1 U15653 ( .A1(n19446), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12630) );
  NAND2_X1 U15654 ( .A1(n12631), .A2(n12630), .ZN(n13407) );
  INV_X1 U15655 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12632) );
  NOR2_X2 U15656 ( .A1(n13001), .A2(n15229), .ZN(n13003) );
  NAND2_X1 U15657 ( .A1(n13009), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13008) );
  INV_X1 U15658 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15210) );
  NAND2_X1 U15659 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n13011), .ZN(
        n13010) );
  INV_X1 U15660 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15190) );
  INV_X1 U15661 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15172) );
  NOR2_X2 U15662 ( .A1(n13015), .A2(n12632), .ZN(n12994) );
  AOI21_X1 U15663 ( .B1(n12632), .B2(n13015), .A(n12994), .ZN(n18856) );
  NAND2_X1 U15664 ( .A1(n19155), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15354) );
  OAI21_X1 U15665 ( .B1(n16259), .B2(n12632), .A(n15354), .ZN(n12639) );
  NOR2_X1 U15666 ( .A1(n14922), .A2(n12634), .ZN(n12635) );
  OR2_X1 U15667 ( .A1(n12633), .A2(n12635), .ZN(n18862) );
  NOR2_X1 U15668 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19857) );
  INV_X1 U15669 ( .A(n19857), .ZN(n13025) );
  NAND2_X1 U15670 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n13274) );
  NAND2_X1 U15671 ( .A1(n13025), .A2(n13274), .ZN(n12636) );
  NOR2_X1 U15672 ( .A1(n18862), .A2(n19179), .ZN(n12638) );
  AOI211_X1 U15673 ( .C1(n19175), .C2(n18856), .A(n12639), .B(n12638), .ZN(
        n12641) );
  AND2_X1 U15674 ( .A1(n12640), .A2(n15366), .ZN(n15181) );
  NAND2_X1 U15675 ( .A1(n15181), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15169) );
  NOR2_X1 U15676 ( .A1(n15169), .A2(n15364), .ZN(n15163) );
  OAI21_X1 U15677 ( .B1(n15163), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15333), .ZN(n15360) );
  NOR2_X2 U15678 ( .A1(n18832), .A2(n13037), .ZN(n19169) );
  NAND3_X1 U15679 ( .A1(n12642), .A2(n12641), .A3(n10070), .ZN(P2_U2993) );
  INV_X1 U15680 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16377) );
  INV_X1 U15681 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17067) );
  AOI22_X1 U15682 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12658) );
  INV_X1 U15683 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18190) );
  AOI22_X1 U15684 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17056), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12646) );
  AOI22_X1 U15685 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12645) );
  OAI211_X1 U15686 ( .C1(n9565), .C2(n18190), .A(n12646), .B(n12645), .ZN(
        n12656) );
  AOI22_X1 U15687 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12654) );
  INV_X2 U15688 ( .A(n9616), .ZN(n17122) );
  AOI22_X1 U15689 ( .A1(n17122), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12653) );
  INV_X2 U15690 ( .A(n9564), .ZN(n17044) );
  AOI22_X1 U15691 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12652) );
  NAND2_X1 U15692 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12651) );
  NAND4_X1 U15693 ( .A1(n12654), .A2(n12653), .A3(n12652), .A4(n12651), .ZN(
        n12655) );
  AOI211_X1 U15694 ( .C1(n17105), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n12656), .B(n12655), .ZN(n12657) );
  OAI211_X1 U15695 ( .C1(n17108), .C2(n17067), .A(n12658), .B(n12657), .ZN(
        n12920) );
  INV_X1 U15696 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n20874) );
  AOI22_X1 U15697 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12669) );
  AOI22_X1 U15698 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12660) );
  AOI22_X1 U15699 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12659) );
  OAI211_X1 U15700 ( .C1(n9565), .C2(n18178), .A(n12660), .B(n12659), .ZN(
        n12667) );
  AOI22_X1 U15701 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17056), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12665) );
  AOI22_X1 U15702 ( .A1(n17122), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12691), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12664) );
  AOI22_X1 U15703 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17131), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12663) );
  NAND2_X1 U15704 ( .A1(n12701), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12662) );
  NAND4_X1 U15705 ( .A1(n12665), .A2(n12664), .A3(n12663), .A4(n12662), .ZN(
        n12666) );
  AOI211_X1 U15706 ( .C1(n17105), .C2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n12667), .B(n12666), .ZN(n12668) );
  OAI211_X1 U15707 ( .C1(n16980), .C2(n20874), .A(n12669), .B(n12668), .ZN(
        n12919) );
  INV_X1 U15708 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12672) );
  INV_X2 U15709 ( .A(n12670), .ZN(n17105) );
  AOI22_X1 U15710 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12671) );
  AOI22_X1 U15711 ( .A1(n17122), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12674) );
  AOI22_X1 U15712 ( .A1(n9579), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12691), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12673) );
  AOI22_X1 U15713 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12676) );
  INV_X1 U15714 ( .A(n12676), .ZN(n12683) );
  INV_X1 U15715 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15608) );
  AOI22_X1 U15716 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12677) );
  OAI21_X1 U15717 ( .B1(n9622), .B2(n15608), .A(n12677), .ZN(n12678) );
  INV_X1 U15718 ( .A(n12678), .ZN(n12681) );
  INV_X1 U15719 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17128) );
  INV_X2 U15720 ( .A(n9616), .ZN(n17147) );
  AOI22_X1 U15721 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12689) );
  AOI22_X1 U15722 ( .A1(n9579), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17056), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12688) );
  AOI22_X1 U15723 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12687) );
  NAND2_X1 U15724 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12686) );
  AOI22_X1 U15725 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9574), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12698) );
  AOI22_X1 U15726 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12694) );
  AOI22_X1 U15727 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12693) );
  OAI211_X1 U15728 ( .C1(n17090), .C2(n18228), .A(n12694), .B(n12693), .ZN(
        n12695) );
  NAND2_X1 U15729 ( .A1(n12932), .A2(n12918), .ZN(n12747) );
  AOI22_X1 U15730 ( .A1(n9579), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17056), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12699) );
  OAI21_X1 U15731 ( .B1(n17088), .B2(n20809), .A(n12699), .ZN(n12710) );
  INV_X1 U15732 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17089) );
  AOI22_X1 U15733 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9574), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12708) );
  AOI22_X1 U15734 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12702) );
  OAI21_X1 U15735 ( .B1(n17113), .B2(n20871), .A(n12702), .ZN(n12706) );
  INV_X1 U15736 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18172) );
  AOI22_X1 U15737 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12691), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12704) );
  AOI22_X1 U15738 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12703) );
  OAI211_X1 U15739 ( .C1(n9565), .C2(n18172), .A(n12704), .B(n12703), .ZN(
        n12705) );
  AOI211_X1 U15740 ( .C1(n12701), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n12706), .B(n12705), .ZN(n12707) );
  OAI211_X1 U15741 ( .C1(n12700), .C2(n17089), .A(n12708), .B(n12707), .ZN(
        n12709) );
  AOI22_X1 U15742 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12711) );
  OAI21_X1 U15743 ( .B1(n10053), .B2(n16966), .A(n12711), .ZN(n12720) );
  INV_X1 U15744 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15671) );
  AOI22_X1 U15745 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12718) );
  AOI22_X1 U15746 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12712) );
  OAI21_X1 U15747 ( .B1(n9565), .B2(n18184), .A(n12712), .ZN(n12716) );
  INV_X1 U15748 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15686) );
  AOI22_X1 U15749 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15684), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12714) );
  AOI22_X1 U15750 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12713) );
  OAI211_X1 U15751 ( .C1(n17108), .C2(n15686), .A(n12714), .B(n12713), .ZN(
        n12715) );
  AOI211_X1 U15752 ( .C1(n12701), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n12716), .B(n12715), .ZN(n12717) );
  OAI211_X1 U15753 ( .C1(n17113), .C2(n15671), .A(n12718), .B(n12717), .ZN(
        n12719) );
  INV_X1 U15754 ( .A(n17323), .ZN(n12753) );
  INV_X1 U15755 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17041) );
  INV_X1 U15756 ( .A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15636) );
  OAI22_X1 U15757 ( .A1(n12721), .A2(n17041), .B1(n16980), .B2(n15636), .ZN(
        n12732) );
  AOI22_X1 U15758 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12730) );
  INV_X2 U15759 ( .A(n9618), .ZN(n17032) );
  AOI22_X1 U15760 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17032), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U15761 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12722) );
  INV_X1 U15762 ( .A(n12722), .ZN(n12727) );
  AOI22_X1 U15763 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15684), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12725) );
  AOI22_X1 U15764 ( .A1(n9568), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12724) );
  AOI22_X1 U15765 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12723) );
  NAND3_X1 U15766 ( .A1(n12725), .A2(n12724), .A3(n12723), .ZN(n12726) );
  AOI211_X1 U15767 ( .C1(n17131), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n12727), .B(n12726), .ZN(n12728) );
  NAND3_X1 U15768 ( .A1(n12730), .A2(n12729), .A3(n12728), .ZN(n12731) );
  INV_X1 U15769 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18054) );
  XOR2_X1 U15770 ( .A(n12733), .B(n17320), .Z(n12755) );
  XOR2_X1 U15771 ( .A(n12734), .B(n17327), .Z(n12751) );
  INV_X1 U15772 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17024) );
  AOI22_X1 U15773 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12740) );
  AOI22_X1 U15774 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12736) );
  AOI22_X1 U15775 ( .A1(n9579), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12691), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12735) );
  AOI22_X1 U15776 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12739) );
  INV_X1 U15777 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18154) );
  INV_X1 U15778 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15615) );
  AOI22_X1 U15779 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17056), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12741) );
  OAI21_X1 U15780 ( .B1(n10053), .B2(n15615), .A(n12741), .ZN(n12743) );
  NAND2_X1 U15781 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17826), .ZN(
        n17825) );
  INV_X1 U15782 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18771) );
  NOR2_X1 U15783 ( .A1(n17825), .A2(n17818), .ZN(n17817) );
  NOR2_X1 U15784 ( .A1(n12932), .A2(n18771), .ZN(n12744) );
  XOR2_X1 U15785 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12745), .Z(
        n17805) );
  INV_X1 U15786 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18103) );
  NOR2_X1 U15787 ( .A1(n18103), .A2(n12745), .ZN(n12746) );
  XNOR2_X1 U15788 ( .A(n12747), .B(n17331), .ZN(n12748) );
  NOR2_X1 U15789 ( .A1(n12749), .A2(n12748), .ZN(n12750) );
  INV_X1 U15790 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18093) );
  INV_X1 U15791 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18081) );
  XOR2_X1 U15792 ( .A(n18081), .B(n12751), .Z(n17784) );
  XNOR2_X1 U15793 ( .A(n12754), .B(n12753), .ZN(n17773) );
  INV_X1 U15794 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18055) );
  XOR2_X1 U15795 ( .A(n18055), .B(n12755), .Z(n17756) );
  NOR2_X2 U15796 ( .A1(n18054), .A2(n17751), .ZN(n17750) );
  NOR2_X1 U15797 ( .A1(n12757), .A2(n12756), .ZN(n12758) );
  NOR2_X2 U15798 ( .A1(n17750), .A2(n12758), .ZN(n12915) );
  INV_X1 U15799 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12759) );
  INV_X1 U15800 ( .A(n12762), .ZN(n12760) );
  NAND2_X1 U15801 ( .A1(n17611), .A2(n12762), .ZN(n17732) );
  INV_X1 U15802 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17641) );
  NAND2_X1 U15803 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18014) );
  INV_X1 U15804 ( .A(n18014), .ZN(n17697) );
  NAND2_X1 U15805 ( .A1(n17697), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17989) );
  INV_X1 U15806 ( .A(n17989), .ZN(n18006) );
  NAND2_X1 U15807 ( .A1(n18006), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17975) );
  INV_X1 U15808 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17654) );
  NOR2_X1 U15809 ( .A1(n17975), .A2(n17654), .ZN(n17977) );
  NAND2_X1 U15810 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17977), .ZN(
        n17960) );
  NOR2_X1 U15811 ( .A1(n17641), .A2(n17960), .ZN(n17888) );
  NOR3_X1 U15812 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17634) );
  NOR2_X1 U15813 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17639) );
  NAND4_X1 U15814 ( .A1(n17634), .A2(n17639), .A3(n17654), .A4(n17641), .ZN(
        n12761) );
  INV_X1 U15815 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17952) );
  INV_X1 U15816 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17943) );
  NAND2_X1 U15817 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17596) );
  NAND2_X1 U15818 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17559) );
  INV_X1 U15819 ( .A(n17559), .ZN(n17894) );
  NAND3_X1 U15820 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n17894), .ZN(n17897) );
  INV_X1 U15821 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17896) );
  NOR2_X1 U15822 ( .A1(n17897), .A2(n17896), .ZN(n15736) );
  NAND2_X1 U15823 ( .A1(n15736), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17851) );
  NOR2_X1 U15824 ( .A1(n17596), .A2(n17851), .ZN(n17497) );
  INV_X1 U15825 ( .A(n17497), .ZN(n17506) );
  INV_X1 U15826 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17922) );
  NAND2_X1 U15827 ( .A1(n17593), .A2(n17922), .ZN(n12766) );
  INV_X1 U15828 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17906) );
  INV_X1 U15829 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17878) );
  INV_X1 U15830 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17855) );
  NOR2_X1 U15831 ( .A1(n17632), .A2(n12769), .ZN(n17508) );
  INV_X1 U15832 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17843) );
  INV_X1 U15833 ( .A(n17509), .ZN(n12772) );
  INV_X1 U15834 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17484) );
  INV_X1 U15835 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n20916) );
  NOR2_X1 U15836 ( .A1(n17632), .A2(n15797), .ZN(n12776) );
  INV_X1 U15837 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18772) );
  AOI22_X1 U15838 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17734), .B1(
        n17632), .B2(n18772), .ZN(n12779) );
  NOR2_X1 U15839 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18772), .ZN(
        n16387) );
  AOI211_X1 U15840 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n18772), .A(
        n15798), .B(n12776), .ZN(n12777) );
  OAI21_X1 U15841 ( .B1(n16387), .B2(n12777), .A(n12779), .ZN(n12778) );
  OAI21_X1 U15842 ( .B1(n12780), .B2(n12779), .A(n12778), .ZN(n16395) );
  AOI21_X1 U15843 ( .B1(n20806), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n12906), .ZN(n12907) );
  INV_X1 U15844 ( .A(n12907), .ZN(n12781) );
  NOR2_X1 U15845 ( .A1(n12781), .A2(n12905), .ZN(n12796) );
  INV_X1 U15846 ( .A(n12906), .ZN(n12782) );
  OAI22_X1 U15847 ( .A1(n18777), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18640), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12787) );
  AOI22_X1 U15848 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18607), .B1(
        n12785), .B2(n18769), .ZN(n12789) );
  NOR2_X1 U15849 ( .A1(n12785), .A2(n18769), .ZN(n12790) );
  NAND2_X1 U15850 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18607), .ZN(
        n12786) );
  OAI22_X1 U15851 ( .A1(n12789), .A2(n18643), .B1(n12790), .B2(n12786), .ZN(
        n12793) );
  INV_X1 U15852 ( .A(n12793), .ZN(n12795) );
  XNOR2_X1 U15853 ( .A(n12788), .B(n12787), .ZN(n12794) );
  OAI21_X1 U15854 ( .B1(n18643), .B2(n12790), .A(n12789), .ZN(n12791) );
  OAI21_X1 U15855 ( .B1(n18607), .B2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n12791), .ZN(n12792) );
  INV_X1 U15856 ( .A(n12792), .ZN(n12904) );
  INV_X1 U15857 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14111) );
  AOI22_X1 U15858 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12797) );
  OAI21_X1 U15859 ( .B1(n9565), .B2(n14111), .A(n12797), .ZN(n12801) );
  INV_X1 U15860 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17124) );
  AOI22_X1 U15861 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n15684), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12799) );
  AOI22_X1 U15862 ( .A1(n9579), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12798) );
  OAI211_X1 U15863 ( .C1(n17108), .C2(n17124), .A(n12799), .B(n12798), .ZN(
        n12800) );
  AOI211_X1 U15864 ( .C1(n12701), .C2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n12801), .B(n12800), .ZN(n12809) );
  AOI22_X1 U15865 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12691), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12802) );
  INV_X1 U15866 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17134) );
  AOI22_X1 U15867 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12803) );
  OAI21_X1 U15868 ( .B1(n17088), .B2(n17134), .A(n12803), .ZN(n12806) );
  AOI22_X1 U15869 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12691), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12810) );
  OAI21_X1 U15870 ( .B1(n12700), .B2(n20773), .A(n12810), .ZN(n12816) );
  INV_X1 U15871 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17035) );
  INV_X2 U15872 ( .A(n17088), .ZN(n15648) );
  AOI22_X1 U15873 ( .A1(n17122), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15648), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12815) );
  INV_X1 U15874 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12812) );
  AOI22_X1 U15875 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12811) );
  AOI22_X1 U15876 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15684), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12814) );
  AOI22_X1 U15877 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12813) );
  INV_X1 U15878 ( .A(n12883), .ZN(n12900) );
  NAND2_X1 U15879 ( .A1(n18157), .A2(n16820), .ZN(n15707) );
  NAND2_X1 U15880 ( .A1(n12900), .A2(n15707), .ZN(n18820) );
  AOI22_X1 U15881 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9574), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12826) );
  INV_X1 U15882 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17083) );
  AOI22_X1 U15883 ( .A1(n17122), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17056), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12818) );
  AOI22_X1 U15884 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12817) );
  OAI211_X1 U15885 ( .C1(n17090), .C2(n17083), .A(n12818), .B(n12817), .ZN(
        n12824) );
  AOI22_X1 U15886 ( .A1(n9568), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15648), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12822) );
  AOI22_X1 U15887 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12821) );
  AOI22_X1 U15888 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12820) );
  NAND2_X1 U15889 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12819) );
  NAND4_X1 U15890 ( .A1(n12822), .A2(n12821), .A3(n12820), .A4(n12819), .ZN(
        n12823) );
  INV_X1 U15891 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16951) );
  AOI22_X1 U15892 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12837) );
  INV_X1 U15893 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17060) );
  AOI22_X1 U15894 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12691), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12828) );
  AOI22_X1 U15895 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12827) );
  OAI211_X1 U15896 ( .C1(n9565), .C2(n17060), .A(n12828), .B(n12827), .ZN(
        n12835) );
  AOI22_X1 U15897 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U15898 ( .A1(n9579), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12832) );
  AOI22_X1 U15899 ( .A1(n15684), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15648), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12831) );
  NAND2_X1 U15900 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12830) );
  NAND4_X1 U15901 ( .A1(n12833), .A2(n12832), .A3(n12831), .A4(n12830), .ZN(
        n12834) );
  AOI211_X2 U15902 ( .C1(n17105), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n12835), .B(n12834), .ZN(n12836) );
  OAI211_X2 U15903 ( .C1(n17108), .C2(n16951), .A(n12837), .B(n12836), .ZN(
        n17199) );
  NOR2_X1 U15904 ( .A1(n14124), .A2(n17199), .ZN(n12885) );
  AOI22_X1 U15905 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15684), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12847) );
  AOI22_X1 U15906 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12839) );
  AOI22_X1 U15907 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12838) );
  OAI211_X1 U15908 ( .C1(n17090), .C2(n16966), .A(n12839), .B(n12838), .ZN(
        n12845) );
  AOI22_X1 U15909 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12843) );
  AOI22_X1 U15910 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15648), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12842) );
  AOI22_X1 U15911 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12841) );
  NAND2_X1 U15912 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12840) );
  NAND4_X1 U15913 ( .A1(n12843), .A2(n12842), .A3(n12841), .A4(n12840), .ZN(
        n12844) );
  AOI22_X1 U15914 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9579), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12848) );
  OAI21_X1 U15915 ( .B1(n9616), .B2(n20864), .A(n12848), .ZN(n12856) );
  INV_X1 U15916 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17112) );
  AOI22_X1 U15917 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12855) );
  INV_X1 U15918 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15643) );
  INV_X1 U15919 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17118) );
  OAI22_X1 U15920 ( .A1(n17113), .A2(n15643), .B1(n9622), .B2(n17118), .ZN(
        n12853) );
  AOI22_X1 U15921 ( .A1(n9568), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15648), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12851) );
  AOI22_X1 U15922 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12850) );
  AOI22_X1 U15923 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12849) );
  NAND3_X1 U15924 ( .A1(n12851), .A2(n12850), .A3(n12849), .ZN(n12852) );
  AOI211_X1 U15925 ( .C1(n17100), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n12853), .B(n12852), .ZN(n12854) );
  AOI22_X1 U15926 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12866) );
  AOI22_X1 U15927 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12858) );
  AOI22_X1 U15928 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15684), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12857) );
  OAI211_X1 U15929 ( .C1(n17108), .C2(n20809), .A(n12858), .B(n12857), .ZN(
        n12864) );
  AOI22_X1 U15930 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17032), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12862) );
  AOI22_X1 U15931 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12861) );
  AOI22_X1 U15932 ( .A1(n17122), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15648), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12860) );
  NAND2_X1 U15933 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12859) );
  NAND4_X1 U15934 ( .A1(n12862), .A2(n12861), .A3(n12860), .A4(n12859), .ZN(
        n12863) );
  INV_X1 U15935 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U15936 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12868) );
  AOI22_X1 U15937 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12867) );
  OAI211_X1 U15938 ( .C1(n9565), .C2(n17043), .A(n12868), .B(n12867), .ZN(
        n12874) );
  AOI22_X1 U15939 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n15684), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n9568), .ZN(n12872) );
  AOI22_X1 U15940 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17143), .B1(
        n17032), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12871) );
  AOI22_X1 U15941 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n12701), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n17105), .ZN(n12870) );
  NAND2_X1 U15942 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17149), .ZN(
        n12869) );
  NAND4_X1 U15943 ( .A1(n12872), .A2(n12871), .A3(n12870), .A4(n12869), .ZN(
        n12873) );
  NAND2_X1 U15944 ( .A1(n12880), .A2(n17240), .ZN(n12894) );
  INV_X1 U15945 ( .A(n14124), .ZN(n18175) );
  NOR2_X1 U15946 ( .A1(n18175), .A2(n17199), .ZN(n18612) );
  INV_X2 U15947 ( .A(n12890), .ZN(n15723) );
  NAND3_X1 U15948 ( .A1(n18181), .A2(n18611), .A3(n17199), .ZN(n14123) );
  INV_X1 U15949 ( .A(n14123), .ZN(n12877) );
  NAND3_X1 U15950 ( .A1(n9794), .A2(n18157), .A3(n12877), .ZN(n12878) );
  NAND2_X1 U15951 ( .A1(n12879), .A2(n12878), .ZN(n12899) );
  INV_X1 U15952 ( .A(n12879), .ZN(n12971) );
  NOR2_X1 U15953 ( .A1(n18157), .A2(n12971), .ZN(n12895) );
  INV_X1 U15954 ( .A(n12880), .ZN(n18169) );
  INV_X1 U15955 ( .A(n12881), .ZN(n12893) );
  NAND2_X1 U15956 ( .A1(n15727), .A2(n18187), .ZN(n15827) );
  INV_X1 U15957 ( .A(n15707), .ZN(n12882) );
  NOR2_X1 U15958 ( .A1(n12883), .A2(n15724), .ZN(n12891) );
  OAI21_X1 U15959 ( .B1(n15724), .B2(n16820), .A(n15827), .ZN(n12884) );
  OAI21_X1 U15960 ( .B1(n12890), .B2(n12885), .A(n12884), .ZN(n12886) );
  INV_X1 U15961 ( .A(n12886), .ZN(n12887) );
  AOI21_X1 U15962 ( .B1(n17240), .B2(n15723), .A(n18175), .ZN(n12902) );
  OAI211_X1 U15963 ( .C1(n18169), .C2(n12893), .A(n15710), .B(n15711), .ZN(
        n12897) );
  AOI21_X1 U15964 ( .B1(n12895), .B2(n12894), .A(n12897), .ZN(n12896) );
  NAND2_X1 U15965 ( .A1(n12901), .A2(n12900), .ZN(n15709) );
  NOR2_X1 U15966 ( .A1(n18157), .A2(n15724), .ZN(n15726) );
  NAND2_X1 U15967 ( .A1(n15726), .A2(n17199), .ZN(n15731) );
  NAND2_X1 U15968 ( .A1(n12906), .A2(n12905), .ZN(n12903) );
  OAI211_X1 U15969 ( .C1(n12906), .C2(n12905), .A(n12904), .B(n12903), .ZN(
        n12972) );
  OAI21_X1 U15970 ( .B1(n12907), .B2(n12972), .A(n12973), .ZN(n18602) );
  NOR3_X1 U15971 ( .A1(n18809), .A2(n18805), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n18812) );
  INV_X1 U15972 ( .A(n18812), .ZN(n18657) );
  NAND2_X1 U15973 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18138) );
  NAND2_X1 U15974 ( .A1(n18759), .A2(n18138), .ZN(n18811) );
  INV_X1 U15975 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18770) );
  INV_X1 U15976 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16500) );
  NOR2_X1 U15977 ( .A1(n18770), .A2(n16500), .ZN(n17788) );
  NOR2_X2 U15978 ( .A1(n17786), .A2(n17788), .ZN(n17824) );
  INV_X1 U15979 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16534) );
  INV_X1 U15980 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17823) );
  NAND2_X1 U15981 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17787) );
  INV_X1 U15982 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16748) );
  NAND4_X1 U15983 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16738) );
  NOR2_X1 U15984 ( .A1(n16748), .A2(n16738), .ZN(n17648) );
  NAND2_X1 U15985 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16701) );
  INV_X1 U15986 ( .A(n16701), .ZN(n17660) );
  NAND2_X1 U15987 ( .A1(n17660), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17618) );
  NAND3_X1 U15988 ( .A1(n17614), .A2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17602) );
  INV_X1 U15989 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17566) );
  NAND2_X1 U15990 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17502) );
  NAND2_X1 U15991 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17463) );
  NAND2_X1 U15992 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16381), .ZN(
        n12908) );
  XOR2_X2 U15993 ( .A(n16534), .B(n12908), .Z(n16838) );
  NOR2_X1 U15994 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18786) );
  NAND2_X1 U15995 ( .A1(n18805), .A2(n18786), .ZN(n18818) );
  OR2_X2 U15996 ( .A1(n18818), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18137) );
  NAND2_X1 U15997 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n9577), .ZN(n16396) );
  INV_X1 U15998 ( .A(n16396), .ZN(n12914) );
  INV_X1 U15999 ( .A(n12909), .ZN(n12910) );
  NAND2_X1 U16000 ( .A1(n18809), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17828) );
  INV_X1 U16001 ( .A(n17828), .ZN(n17664) );
  NAND3_X1 U16002 ( .A1(n18805), .A2(n18759), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18505) );
  NAND2_X1 U16003 ( .A1(n12910), .A2(n17617), .ZN(n16366) );
  XNOR2_X1 U16004 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12912) );
  NOR2_X1 U16005 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17564), .ZN(
        n16382) );
  NOR2_X1 U16006 ( .A1(n17823), .A2(n17462), .ZN(n12978) );
  INV_X1 U16007 ( .A(n12978), .ZN(n16524) );
  OR2_X1 U16008 ( .A1(n16524), .A2(n17463), .ZN(n16522) );
  NOR2_X1 U16009 ( .A1(n18313), .A2(n12910), .ZN(n16371) );
  AOI211_X1 U16010 ( .C1(n16522), .C2(n17664), .A(n17786), .B(n16371), .ZN(
        n12911) );
  INV_X1 U16011 ( .A(n12911), .ZN(n16372) );
  NOR2_X1 U16012 ( .A1(n16382), .A2(n16372), .ZN(n16365) );
  OAI22_X1 U16013 ( .A1(n16366), .A2(n12912), .B1(n16365), .B2(n16534), .ZN(
        n12913) );
  AOI211_X1 U16014 ( .C1(n17682), .C2(n16838), .A(n12914), .B(n12913), .ZN(
        n12953) );
  NAND2_X1 U16015 ( .A1(n12915), .A2(n17734), .ZN(n17633) );
  NAND3_X1 U16016 ( .A1(n17993), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17647) );
  INV_X1 U16017 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17870) );
  NOR4_X1 U16018 ( .A1(n17870), .A2(n17878), .A3(n17855), .A4(n17843), .ZN(
        n16361) );
  NAND2_X1 U16019 ( .A1(n15736), .A2(n16361), .ZN(n16410) );
  NOR2_X1 U16020 ( .A1(n17596), .A2(n16410), .ZN(n12949) );
  NAND2_X1 U16021 ( .A1(n17958), .A2(n12949), .ZN(n16374) );
  NOR2_X1 U16022 ( .A1(n20916), .A2(n17484), .ZN(n16375) );
  NAND2_X1 U16023 ( .A1(n16375), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16362) );
  NAND2_X1 U16024 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16359), .ZN(
        n12916) );
  XOR2_X1 U16025 ( .A(n18772), .B(n12916), .Z(n16388) );
  NOR2_X1 U16026 ( .A1(n17347), .A2(n12917), .ZN(n12928) );
  NOR2_X1 U16027 ( .A1(n12928), .A2(n12918), .ZN(n12926) );
  NOR2_X1 U16028 ( .A1(n17331), .A2(n12926), .ZN(n12925) );
  NAND2_X1 U16029 ( .A1(n12925), .A2(n12919), .ZN(n12923) );
  NOR2_X1 U16030 ( .A1(n17323), .A2(n12923), .ZN(n12922) );
  NAND2_X1 U16031 ( .A1(n12922), .A2(n12920), .ZN(n12921) );
  NOR2_X1 U16032 ( .A1(n17316), .A2(n12921), .ZN(n12946) );
  XOR2_X1 U16033 ( .A(n17316), .B(n12921), .Z(n17744) );
  XNOR2_X1 U16034 ( .A(n17320), .B(n12922), .ZN(n12939) );
  XOR2_X1 U16035 ( .A(n17323), .B(n12923), .Z(n12924) );
  NAND2_X1 U16036 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12924), .ZN(
        n12938) );
  XOR2_X1 U16037 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n12924), .Z(
        n17769) );
  XNOR2_X1 U16038 ( .A(n17327), .B(n12925), .ZN(n12936) );
  XOR2_X1 U16039 ( .A(n12926), .B(n17331), .Z(n12927) );
  NAND2_X1 U16040 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12927), .ZN(
        n12934) );
  XOR2_X1 U16041 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n12927), .Z(
        n17796) );
  XNOR2_X1 U16042 ( .A(n17336), .B(n12928), .ZN(n12929) );
  OR2_X1 U16043 ( .A1(n18103), .A2(n12929), .ZN(n12933) );
  XOR2_X1 U16044 ( .A(n18103), .B(n12929), .Z(n17809) );
  AOI21_X1 U16045 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12932), .A(
        n17826), .ZN(n12931) );
  INV_X1 U16046 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18787) );
  NOR2_X1 U16047 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12932), .ZN(
        n12930) );
  AOI221_X1 U16048 ( .B1(n17826), .B2(n12932), .C1(n12931), .C2(n18787), .A(
        n12930), .ZN(n17808) );
  NAND2_X1 U16049 ( .A1(n17809), .A2(n17808), .ZN(n17807) );
  NAND2_X1 U16050 ( .A1(n12933), .A2(n17807), .ZN(n17795) );
  NAND2_X1 U16051 ( .A1(n17796), .A2(n17795), .ZN(n17794) );
  NAND2_X1 U16052 ( .A1(n12934), .A2(n17794), .ZN(n12935) );
  NAND2_X1 U16053 ( .A1(n12936), .A2(n12935), .ZN(n12937) );
  XOR2_X1 U16054 ( .A(n12936), .B(n12935), .Z(n17781) );
  NAND2_X1 U16055 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17781), .ZN(
        n17780) );
  NAND2_X1 U16056 ( .A1(n12937), .A2(n17780), .ZN(n17768) );
  NAND2_X1 U16057 ( .A1(n17769), .A2(n17768), .ZN(n17767) );
  NAND2_X1 U16058 ( .A1(n12938), .A2(n17767), .ZN(n12940) );
  NAND2_X1 U16059 ( .A1(n12939), .A2(n12940), .ZN(n12941) );
  XOR2_X1 U16060 ( .A(n12940), .B(n12939), .Z(n17762) );
  NAND2_X1 U16061 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17762), .ZN(
        n17761) );
  NAND2_X1 U16062 ( .A1(n12946), .A2(n12943), .ZN(n12947) );
  INV_X1 U16063 ( .A(n12943), .ZN(n12945) );
  NAND2_X1 U16064 ( .A1(n17744), .A2(n17745), .ZN(n17743) );
  NAND2_X1 U16065 ( .A1(n12946), .A2(n12945), .ZN(n12944) );
  OAI211_X1 U16066 ( .C1(n12946), .C2(n12945), .A(n17743), .B(n12944), .ZN(
        n17736) );
  NAND2_X1 U16067 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17736), .ZN(
        n17735) );
  INV_X1 U16068 ( .A(n17887), .ZN(n12948) );
  NAND2_X1 U16069 ( .A1(n12949), .A2(n12948), .ZN(n17836) );
  INV_X1 U16070 ( .A(n16362), .ZN(n16390) );
  NAND3_X1 U16071 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17461), .A3(
        n16390), .ZN(n12950) );
  XNOR2_X1 U16072 ( .A(n18772), .B(n12950), .ZN(n16393) );
  NOR2_X1 U16073 ( .A1(n16393), .A2(n17832), .ZN(n12951) );
  AOI21_X1 U16074 ( .B1(n16388), .B2(n17739), .A(n12951), .ZN(n12952) );
  AND2_X1 U16075 ( .A1(n12953), .A2(n12952), .ZN(n12954) );
  INV_X1 U16076 ( .A(n16314), .ZN(n12956) );
  NAND2_X1 U16077 ( .A1(n12956), .A2(n16311), .ZN(n13162) );
  NAND2_X1 U16078 ( .A1(n13162), .A2(n12957), .ZN(n12958) );
  NAND2_X1 U16079 ( .A1(n12959), .A2(n15018), .ZN(n12963) );
  NAND2_X1 U16080 ( .A1(n15022), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12960) );
  NAND2_X1 U16081 ( .A1(n12963), .A2(n12962), .ZN(P2_U2857) );
  NOR2_X1 U16082 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12965) );
  NOR4_X1 U16083 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12964) );
  NAND4_X1 U16084 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12965), .A4(n12964), .ZN(n12968) );
  NOR2_X1 U16085 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12968), .ZN(n16488)
         );
  INV_X1 U16086 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20792) );
  NOR3_X1 U16087 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20792), .ZN(n12967) );
  NOR4_X1 U16088 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12966) );
  NAND4_X1 U16089 ( .A1(n20079), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12967), .A4(
        n12966), .ZN(U214) );
  NOR2_X1 U16090 ( .A1(n13674), .A2(n12968), .ZN(n16420) );
  NAND2_X1 U16091 ( .A1(n16420), .A2(U214), .ZN(U212) );
  NOR3_X1 U16092 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16850) );
  INV_X1 U16093 ( .A(n16850), .ZN(n16836) );
  NOR2_X1 U16094 ( .A1(n16836), .A2(P3_EBX_REG_3__SCAN_IN), .ZN(n16835) );
  INV_X1 U16095 ( .A(n16835), .ZN(n16819) );
  INV_X1 U16096 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16815) );
  NAND2_X1 U16097 ( .A1(n16818), .A2(n16815), .ZN(n16814) );
  INV_X1 U16098 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17163) );
  NAND2_X1 U16099 ( .A1(n16795), .A2(n17163), .ZN(n16792) );
  INV_X1 U16100 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16762) );
  NAND2_X1 U16101 ( .A1(n16761), .A2(n16762), .ZN(n16750) );
  INV_X1 U16102 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16745) );
  NAND2_X1 U16103 ( .A1(n16749), .A2(n16745), .ZN(n16744) );
  INV_X1 U16104 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16725) );
  NAND2_X1 U16105 ( .A1(n16728), .A2(n16725), .ZN(n16724) );
  INV_X1 U16106 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16696) );
  NAND2_X1 U16107 ( .A1(n16706), .A2(n16696), .ZN(n16695) );
  INV_X1 U16108 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16675) );
  NAND2_X1 U16109 ( .A1(n16676), .A2(n16675), .ZN(n16672) );
  INV_X1 U16110 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16993) );
  NAND2_X1 U16111 ( .A1(n16654), .A2(n16993), .ZN(n16650) );
  INV_X1 U16112 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16977) );
  NAND2_X1 U16113 ( .A1(n16630), .A2(n16977), .ZN(n16626) );
  INV_X1 U16114 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16605) );
  NAND2_X1 U16115 ( .A1(n16611), .A2(n16605), .ZN(n16604) );
  NOR2_X1 U16116 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16604), .ZN(n16589) );
  INV_X1 U16117 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16584) );
  NAND2_X1 U16118 ( .A1(n16589), .A2(n16584), .ZN(n16583) );
  NOR2_X1 U16119 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16583), .ZN(n16572) );
  NAND2_X1 U16120 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18814) );
  NAND2_X1 U16121 ( .A1(n12970), .A2(n12969), .ZN(n15716) );
  NAND2_X1 U16122 ( .A1(n12973), .A2(n12972), .ZN(n18599) );
  NAND2_X1 U16123 ( .A1(n18825), .A2(n16820), .ZN(n18823) );
  NAND2_X1 U16124 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18804), .ZN(n12974) );
  AOI211_X4 U16125 ( .C1(n16500), .C2(n18814), .A(n18823), .B(n12974), .ZN(
        n16880) );
  AOI211_X1 U16126 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16583), .A(n16572), .B(
        n16849), .ZN(n12990) );
  INV_X1 U16127 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18735) );
  INV_X1 U16128 ( .A(n18823), .ZN(n12975) );
  NAND2_X1 U16129 ( .A1(n18800), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18747) );
  OAI211_X1 U16130 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18682), .B(n18739), .ZN(n18675) );
  INV_X1 U16131 ( .A(n18814), .ZN(n18806) );
  AOI211_X1 U16132 ( .C1(n18675), .C2(n18157), .A(n18806), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18652) );
  INV_X1 U16133 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18733) );
  INV_X1 U16134 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18730) );
  INV_X1 U16135 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18726) );
  INV_X1 U16136 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18707) );
  INV_X1 U16137 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18700) );
  INV_X1 U16138 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18691) );
  NAND3_X1 U16139 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16840) );
  NOR2_X1 U16140 ( .A1(n18691), .A2(n16840), .ZN(n16807) );
  NAND2_X1 U16141 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16807), .ZN(n16787) );
  NAND2_X1 U16142 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n16788) );
  NOR3_X1 U16143 ( .A1(n18700), .A2(n16787), .A3(n16788), .ZN(n16755) );
  NAND4_X1 U16144 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16755), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n16732) );
  NOR2_X1 U16145 ( .A1(n18707), .A2(n16732), .ZN(n16708) );
  NAND3_X1 U16146 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n16708), .ZN(n16677) );
  INV_X1 U16147 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18718) );
  NAND2_X1 U16148 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16679) );
  NOR2_X1 U16149 ( .A1(n18718), .A2(n16679), .ZN(n16641) );
  NAND3_X1 U16150 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16641), .A3(
        P3_REIP_REG_18__SCAN_IN), .ZN(n16637) );
  NOR2_X1 U16151 ( .A1(n16677), .A2(n16637), .ZN(n16636) );
  NAND2_X1 U16152 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16636), .ZN(n16619) );
  NOR2_X1 U16153 ( .A1(n18726), .A2(n16619), .ZN(n16610) );
  NAND2_X1 U16154 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16610), .ZN(n16601) );
  NOR2_X1 U16155 ( .A1(n18730), .A2(n16601), .ZN(n16599) );
  NAND2_X1 U16156 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16599), .ZN(n16580) );
  NOR2_X1 U16157 ( .A1(n18733), .A2(n16580), .ZN(n12977) );
  NAND2_X1 U16158 ( .A1(n16872), .A2(n12977), .ZN(n16520) );
  NOR3_X1 U16159 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n18665) );
  NAND2_X1 U16160 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18665), .ZN(n16843) );
  INV_X1 U16161 ( .A(n16843), .ZN(n18660) );
  NAND3_X1 U16162 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .A3(n18666), .ZN(n12976) );
  OAI221_X1 U16163 ( .B1(n16830), .B2(P3_REIP_REG_26__SCAN_IN), .C1(n16830), 
        .C2(n12977), .A(n16884), .ZN(n16525) );
  INV_X1 U16164 ( .A(n16525), .ZN(n16575) );
  AOI21_X1 U16165 ( .B1(n18735), .B2(n16520), .A(n16575), .ZN(n12989) );
  INV_X1 U16166 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16618) );
  NAND3_X1 U16167 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9592), .A3(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12982) );
  NOR2_X1 U16168 ( .A1(n16618), .A2(n12982), .ZN(n17499) );
  NAND2_X1 U16169 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17499), .ZN(
        n12980) );
  OR2_X1 U16170 ( .A1(n17502), .A2(n12980), .ZN(n17459) );
  AOI21_X1 U16171 ( .B1(n9752), .B2(n17459), .A(n12978), .ZN(n17491) );
  INV_X1 U16172 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17517) );
  NOR2_X1 U16173 ( .A1(n17517), .A2(n12980), .ZN(n12979) );
  OAI21_X1 U16174 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n12979), .A(
        n17459), .ZN(n17504) );
  INV_X1 U16175 ( .A(n17504), .ZN(n16578) );
  AOI21_X1 U16176 ( .B1(n17517), .B2(n12980), .A(n12979), .ZN(n17513) );
  OAI21_X1 U16177 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17499), .A(
        n12980), .ZN(n12981) );
  INV_X1 U16178 ( .A(n12981), .ZN(n17528) );
  AOI21_X1 U16179 ( .B1(n16618), .B2(n12982), .A(n17499), .ZN(n17545) );
  AND2_X1 U16180 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9592), .ZN(
        n12983) );
  OAI21_X1 U16181 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n12983), .A(
        n12982), .ZN(n17555) );
  INV_X1 U16182 ( .A(n17555), .ZN(n16622) );
  NOR2_X1 U16183 ( .A1(n17823), .A2(n17567), .ZN(n17543) );
  INV_X1 U16184 ( .A(n17543), .ZN(n16644) );
  AOI21_X1 U16185 ( .B1(n17566), .B2(n16644), .A(n12983), .ZN(n17570) );
  INV_X1 U16186 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17630) );
  INV_X1 U16187 ( .A(n12984), .ZN(n17661) );
  NAND2_X1 U16188 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17661), .ZN(
        n17663) );
  NOR2_X1 U16189 ( .A1(n17618), .A2(n17663), .ZN(n17616) );
  INV_X1 U16190 ( .A(n17616), .ZN(n16703) );
  NOR2_X1 U16191 ( .A1(n17630), .A2(n16703), .ZN(n16681) );
  INV_X1 U16192 ( .A(n16681), .ZN(n16688) );
  NOR2_X1 U16193 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16688), .ZN(
        n16643) );
  AOI21_X1 U16194 ( .B1(n17543), .B2(n16643), .A(n9590), .ZN(n16632) );
  NOR2_X1 U16195 ( .A1(n17570), .A2(n16632), .ZN(n16631) );
  NOR2_X1 U16196 ( .A1(n16631), .A2(n9590), .ZN(n16621) );
  NOR2_X1 U16197 ( .A1(n16622), .A2(n16621), .ZN(n16620) );
  NOR2_X1 U16198 ( .A1(n16597), .A2(n9590), .ZN(n16591) );
  NOR2_X1 U16199 ( .A1(n17513), .A2(n16591), .ZN(n16590) );
  AOI211_X1 U16200 ( .C1(n17491), .C2(n12985), .A(n9636), .B(n16824), .ZN(
        n12988) );
  AOI22_X1 U16201 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16875), .B1(
        n16881), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n12986) );
  INV_X1 U16202 ( .A(n12986), .ZN(n12987) );
  OR4_X1 U16203 ( .A1(n12990), .A2(n12989), .A3(n12988), .A4(n12987), .ZN(
        P3_U2645) );
  AOI21_X1 U16204 ( .B1(n12993), .B2(n9967), .A(n9653), .ZN(n15153) );
  INV_X1 U16205 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14893) );
  INV_X1 U16206 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15100) );
  INV_X1 U16207 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14253) );
  OAI22_X2 U16208 ( .A1(n14265), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n18828), 
        .B2(n14253), .ZN(n13017) );
  OAI21_X1 U16209 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12994), .A(
        n12993), .ZN(n16195) );
  INV_X1 U16210 ( .A(n16195), .ZN(n15749) );
  AOI21_X1 U16211 ( .B1(n15172), .B2(n13014), .A(n12995), .ZN(n18870) );
  INV_X1 U16212 ( .A(n13010), .ZN(n12997) );
  INV_X1 U16213 ( .A(n13012), .ZN(n12996) );
  OAI21_X1 U16214 ( .B1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n12997), .A(
        n12996), .ZN(n18887) );
  AOI21_X1 U16215 ( .B1(n15210), .B2(n13008), .A(n13011), .ZN(n15209) );
  AOI21_X1 U16216 ( .B1(n18917), .B2(n13006), .A(n13009), .ZN(n18923) );
  AOI21_X1 U16217 ( .B1(n16222), .B2(n13004), .A(n13007), .ZN(n18939) );
  AOI21_X1 U16218 ( .B1(n16234), .B2(n13002), .A(n13005), .ZN(n18962) );
  AOI21_X1 U16219 ( .B1(n15229), .B2(n13001), .A(n13003), .ZN(n18972) );
  AOI21_X1 U16220 ( .B1(n16251), .B2(n12999), .A(n9588), .ZN(n19000) );
  AOI21_X1 U16221 ( .B1(n16260), .B2(n12998), .A(n13000), .ZN(n16252) );
  OAI22_X1 U16222 ( .A1(n18828), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n13931) );
  INV_X1 U16223 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15241) );
  OAI22_X1 U16224 ( .A1(n18828), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n15241), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13913) );
  AND2_X1 U16225 ( .A1(n13931), .A2(n13913), .ZN(n13861) );
  OAI21_X1 U16226 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12998), .ZN(n19171) );
  NAND2_X1 U16227 ( .A1(n13861), .A2(n19171), .ZN(n13819) );
  NOR2_X1 U16228 ( .A1(n16252), .A2(n13819), .ZN(n19014) );
  OAI21_X1 U16229 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13000), .A(
        n12999), .ZN(n19164) );
  NAND2_X1 U16230 ( .A1(n19014), .A2(n19164), .ZN(n18998) );
  NOR2_X1 U16231 ( .A1(n19000), .A2(n18998), .ZN(n18983) );
  OAI21_X1 U16232 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9588), .A(
        n13001), .ZN(n18985) );
  NAND2_X1 U16233 ( .A1(n18983), .A2(n18985), .ZN(n18971) );
  NOR2_X1 U16234 ( .A1(n18972), .A2(n18971), .ZN(n13850) );
  OAI21_X1 U16235 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13003), .A(
        n13002), .ZN(n16242) );
  NAND2_X1 U16236 ( .A1(n13850), .A2(n16242), .ZN(n18961) );
  NOR2_X1 U16237 ( .A1(n18962), .A2(n18961), .ZN(n18952) );
  OAI21_X1 U16238 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13005), .A(
        n13004), .ZN(n18954) );
  NAND2_X1 U16239 ( .A1(n18952), .A2(n18954), .ZN(n18938) );
  NOR2_X1 U16240 ( .A1(n18939), .A2(n18938), .ZN(n18928) );
  OAI21_X1 U16241 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n13007), .A(
        n13006), .ZN(n18929) );
  NAND2_X1 U16242 ( .A1(n18928), .A2(n18929), .ZN(n18921) );
  NOR2_X1 U16243 ( .A1(n18923), .A2(n18921), .ZN(n13973) );
  OAI21_X1 U16244 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n13009), .A(
        n13008), .ZN(n16208) );
  NAND2_X1 U16245 ( .A1(n13973), .A2(n16208), .ZN(n18907) );
  NOR2_X1 U16246 ( .A1(n15209), .A2(n18907), .ZN(n18893) );
  OAI21_X1 U16247 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n13011), .A(
        n13010), .ZN(n18894) );
  AND2_X1 U16248 ( .A1(n18893), .A2(n18894), .ZN(n18888) );
  AND2_X1 U16249 ( .A1(n18887), .A2(n18888), .ZN(n14939) );
  OR2_X1 U16250 ( .A1(n13012), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13013) );
  NAND2_X1 U16251 ( .A1(n13014), .A2(n13013), .ZN(n15185) );
  NAND2_X1 U16252 ( .A1(n14939), .A2(n15185), .ZN(n18868) );
  NOR2_X1 U16253 ( .A1(n18870), .A2(n18868), .ZN(n14920) );
  OAI21_X1 U16254 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12995), .A(
        n13015), .ZN(n15164) );
  AND2_X1 U16255 ( .A1(n14920), .A2(n15164), .ZN(n18858) );
  INV_X1 U16256 ( .A(n18855), .ZN(n13018) );
  NAND2_X1 U16257 ( .A1(n18856), .A2(n13017), .ZN(n18857) );
  NAND2_X1 U16258 ( .A1(n13018), .A2(n18857), .ZN(n15748) );
  NOR2_X1 U16259 ( .A1(n15749), .A2(n15748), .ZN(n15747) );
  INV_X1 U16260 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19860) );
  NAND4_X1 U16261 ( .A1(n18828), .A2(n19860), .A3(n19446), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19720) );
  AOI211_X1 U16262 ( .C1(n15153), .C2(n13019), .A(n13053), .B(n19720), .ZN(
        n13046) );
  NAND2_X1 U16263 ( .A1(n10744), .A2(n13020), .ZN(n13021) );
  NAND2_X1 U16264 ( .A1(n19446), .A2(n19711), .ZN(n13034) );
  INV_X1 U16265 ( .A(n13034), .ZN(n13022) );
  OAI21_X1 U16266 ( .B1(P2_EBX_REG_31__SCAN_IN), .B2(n13022), .A(n13037), .ZN(
        n13023) );
  NAND2_X1 U16267 ( .A1(n19446), .A2(n16316), .ZN(n16347) );
  NAND2_X1 U16268 ( .A1(n13023), .A2(n16347), .ZN(n13024) );
  NOR2_X2 U16269 ( .A1(n13121), .A2(n13024), .ZN(n19025) );
  INV_X1 U16270 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19777) );
  NOR3_X1 U16271 ( .A1(n18828), .A2(n10900), .A3(n13025), .ZN(n16343) );
  NOR2_X1 U16272 ( .A1(n16343), .A2(n19002), .ZN(n13026) );
  NAND2_X1 U16273 ( .A1(n16264), .A2(n13026), .ZN(n13027) );
  OAI22_X1 U16274 ( .A1(n10839), .A2(n19009), .B1(n19777), .B2(n18993), .ZN(
        n13045) );
  INV_X1 U16275 ( .A(n13028), .ZN(n13031) );
  NAND2_X1 U16276 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13034), .ZN(n13029) );
  NOR2_X1 U16277 ( .A1(n13035), .A2(n13029), .ZN(n13030) );
  NAND2_X1 U16278 ( .A1(n18829), .A2(n13030), .ZN(n19008) );
  NAND2_X1 U16279 ( .A1(n18993), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18991) );
  OAI22_X1 U16280 ( .A1(n13031), .A2(n19008), .B1(n18991), .B2(n9967), .ZN(
        n13044) );
  INV_X1 U16281 ( .A(n14994), .ZN(n13033) );
  OAI21_X1 U16282 ( .B1(n13033), .B2(n10051), .A(n14901), .ZN(n15321) );
  NOR2_X1 U16283 ( .A1(n13035), .A2(n13034), .ZN(n13036) );
  NAND2_X1 U16284 ( .A1(n18829), .A2(n13036), .ZN(n19011) );
  INV_X1 U16285 ( .A(n16347), .ZN(n13038) );
  AND2_X1 U16286 ( .A1(n9614), .A2(n13040), .ZN(n13041) );
  NOR2_X1 U16287 ( .A1(n13039), .A2(n13041), .ZN(n15318) );
  INV_X1 U16288 ( .A(n15318), .ZN(n13042) );
  OAI22_X1 U16289 ( .A1(n15321), .A2(n19011), .B1(n19006), .B2(n13042), .ZN(
        n13043) );
  OR4_X1 U16290 ( .A1(n13046), .A2(n13045), .A3(n13044), .A4(n13043), .ZN(
        P2_U2832) );
  INV_X1 U16291 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13056) );
  INV_X1 U16292 ( .A(n13049), .ZN(n13047) );
  AOI21_X1 U16293 ( .B1(n13056), .B2(n13047), .A(n14195), .ZN(n15122) );
  NOR2_X1 U16294 ( .A1(n13051), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13048) );
  OR2_X1 U16295 ( .A1(n13049), .A2(n13048), .ZN(n15133) );
  INV_X1 U16296 ( .A(n15133), .ZN(n16162) );
  AND2_X1 U16297 ( .A1(n13052), .A2(n14893), .ZN(n13050) );
  NOR2_X1 U16298 ( .A1(n13051), .A2(n13050), .ZN(n14888) );
  OAI21_X1 U16299 ( .B1(n9653), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n13052), .ZN(n15144) );
  INV_X1 U16300 ( .A(n15144), .ZN(n14911) );
  NOR2_X1 U16301 ( .A1(n13016), .A2(n14910), .ZN(n14889) );
  NOR2_X1 U16302 ( .A1(n14888), .A2(n14889), .ZN(n14887) );
  NOR2_X1 U16303 ( .A1(n16162), .A2(n16161), .ZN(n16160) );
  NOR2_X1 U16304 ( .A1(n13016), .A2(n16160), .ZN(n13054) );
  NOR2_X1 U16305 ( .A1(n15122), .A2(n13054), .ZN(n14196) );
  AOI211_X1 U16306 ( .C1(n15122), .C2(n13054), .A(n14196), .B(n19720), .ZN(
        n13066) );
  AOI22_X1 U16307 ( .A1(P2_EBX_REG_27__SCAN_IN), .A2(n19025), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19031), .ZN(n13055) );
  INV_X1 U16308 ( .A(n13055), .ZN(n13065) );
  OAI22_X1 U16309 ( .A1(n13057), .A2(n19008), .B1(n18991), .B2(n13056), .ZN(
        n13064) );
  NAND2_X1 U16310 ( .A1(n14967), .A2(n13058), .ZN(n13059) );
  NAND2_X1 U16311 ( .A1(n14870), .A2(n13059), .ZN(n15283) );
  NAND2_X1 U16312 ( .A1(n15050), .A2(n13060), .ZN(n13061) );
  AND2_X1 U16313 ( .A1(n14873), .A2(n13061), .ZN(n15280) );
  INV_X1 U16314 ( .A(n15280), .ZN(n13062) );
  OAI22_X1 U16315 ( .A1(n15283), .A2(n19011), .B1(n13062), .B2(n19006), .ZN(
        n13063) );
  OR4_X1 U16316 ( .A1(n13066), .A2(n13065), .A3(n13064), .A4(n13063), .ZN(
        P2_U2828) );
  NAND2_X1 U16317 ( .A1(n14832), .A2(n20102), .ZN(n13067) );
  OAI21_X1 U16318 ( .B1(n13068), .B2(n13413), .A(n13242), .ZN(n13069) );
  INV_X1 U16319 ( .A(n13069), .ZN(n13070) );
  NAND2_X1 U16320 ( .A1(n13071), .A2(n13070), .ZN(n13087) );
  AND2_X1 U16321 ( .A1(n13087), .A2(n13100), .ZN(n13073) );
  AND2_X1 U16322 ( .A1(n13072), .A2(n11320), .ZN(n13093) );
  AND2_X1 U16323 ( .A1(n13093), .A2(n20084), .ZN(n13220) );
  NOR2_X1 U16324 ( .A1(n13073), .A2(n13220), .ZN(n13361) );
  NOR2_X1 U16325 ( .A1(n13357), .A2(n13361), .ZN(n13082) );
  INV_X1 U16326 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20695) );
  AND2_X1 U16327 ( .A1(n13075), .A2(n20695), .ZN(n15804) );
  OAI21_X1 U16328 ( .B1(n20102), .B2(n15804), .A(n20691), .ZN(n13795) );
  INV_X1 U16329 ( .A(n13795), .ZN(n13076) );
  NAND2_X1 U16330 ( .A1(n13074), .A2(n13076), .ZN(n13077) );
  NAND3_X1 U16331 ( .A1(n13077), .A2(n13242), .A3(n13385), .ZN(n13078) );
  NAND2_X1 U16332 ( .A1(n13364), .A2(n13078), .ZN(n13080) );
  OAI211_X1 U16333 ( .C1(n13413), .C2(n15804), .A(n13219), .B(n20691), .ZN(
        n13079) );
  MUX2_X1 U16334 ( .A(n13080), .B(n13079), .S(n20107), .Z(n13081) );
  NOR2_X1 U16335 ( .A1(n11692), .A2(n14290), .ZN(n13084) );
  OAI22_X1 U16336 ( .A1(n14168), .A2(n13216), .B1(n11320), .B2(n13358), .ZN(
        n13083) );
  NOR2_X1 U16337 ( .A1(n13084), .A2(n13083), .ZN(n13086) );
  NAND3_X1 U16338 ( .A1(n13087), .A2(n13086), .A3(n13085), .ZN(n13329) );
  OR2_X1 U16339 ( .A1(n13329), .A2(n13088), .ZN(n13089) );
  INV_X1 U16340 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14837) );
  AND2_X1 U16341 ( .A1(n14692), .A2(n14837), .ZN(n13493) );
  NAND3_X1 U16342 ( .A1(n13242), .A2(n14276), .A3(n13359), .ZN(n13090) );
  NOR2_X1 U16343 ( .A1(n13091), .A2(n13090), .ZN(n13342) );
  NAND2_X1 U16344 ( .A1(n13107), .A2(n13342), .ZN(n14810) );
  NOR2_X1 U16345 ( .A1(n14810), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13092) );
  OR2_X1 U16346 ( .A1(n13493), .A2(n13092), .ZN(n13457) );
  INV_X1 U16347 ( .A(n13358), .ZN(n13797) );
  INV_X1 U16348 ( .A(n15808), .ZN(n13497) );
  NOR2_X1 U16349 ( .A1(n16139), .A2(n13107), .ZN(n13494) );
  INV_X1 U16350 ( .A(n13494), .ZN(n13094) );
  AOI21_X1 U16351 ( .B1(n13497), .B2(n13094), .A(n14837), .ZN(n13114) );
  OR2_X1 U16352 ( .A1(n13095), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13096) );
  NAND2_X1 U16353 ( .A1(n13097), .A2(n13096), .ZN(n20056) );
  INV_X1 U16354 ( .A(n13104), .ZN(n13102) );
  NAND2_X1 U16355 ( .A1(n13793), .A2(n13098), .ZN(n13099) );
  NAND2_X1 U16356 ( .A1(n13100), .A2(n13099), .ZN(n13218) );
  OAI211_X1 U16357 ( .C1(n11326), .C2(n13102), .A(n13101), .B(n13218), .ZN(
        n13103) );
  NAND2_X1 U16358 ( .A1(n13074), .A2(n13410), .ZN(n15782) );
  NAND2_X1 U16359 ( .A1(n13104), .A2(n11326), .ZN(n13105) );
  NAND2_X1 U16360 ( .A1(n15782), .A2(n13105), .ZN(n13106) );
  INV_X1 U16361 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13109) );
  NAND2_X1 U16362 ( .A1(n14276), .A2(n13109), .ZN(n13108) );
  OAI21_X1 U16363 ( .B1(n9581), .B2(n13109), .A(n13108), .ZN(n13382) );
  INV_X1 U16364 ( .A(n13382), .ZN(n13111) );
  NAND2_X1 U16365 ( .A1(n14168), .A2(n14837), .ZN(n13110) );
  AND2_X1 U16366 ( .A1(n13111), .A2(n13110), .ZN(n13841) );
  NAND2_X1 U16367 ( .A1(n20067), .A2(n13841), .ZN(n13112) );
  INV_X1 U16368 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13848) );
  OR2_X1 U16369 ( .A1(n16041), .A2(n13848), .ZN(n20062) );
  OAI211_X1 U16370 ( .C1(n20056), .C2(n16070), .A(n13112), .B(n20062), .ZN(
        n13113) );
  OR3_X1 U16371 ( .A1(n13457), .A2(n13114), .A3(n13113), .ZN(P1_U3031) );
  OR2_X1 U16372 ( .A1(n10748), .A2(n19714), .ZN(n13267) );
  NOR2_X1 U16373 ( .A1(n16310), .A2(n13267), .ZN(n19039) );
  INV_X1 U16374 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13115) );
  OAI211_X1 U16375 ( .C1(n19039), .C2(n13115), .A(n13121), .B(n18827), .ZN(
        P2_U2814) );
  INV_X1 U16376 ( .A(n18829), .ZN(n19862) );
  OAI21_X1 U16377 ( .B1(P2_READREQUEST_REG_SCAN_IN), .B2(n13116), .A(n19862), 
        .ZN(n13117) );
  OAI21_X1 U16378 ( .B1(n13118), .B2(n19862), .A(n13117), .ZN(P2_U3612) );
  INV_X1 U16379 ( .A(n13121), .ZN(n13120) );
  NAND2_X1 U16380 ( .A1(n19196), .A2(n19865), .ZN(n13119) );
  NAND2_X2 U16381 ( .A1(n13120), .A2(n13119), .ZN(n13207) );
  AOI22_X1 U16382 ( .A1(P2_EAX_REG_29__SCAN_IN), .A2(n13130), .B1(n13207), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13125) );
  INV_X1 U16383 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14051) );
  OR2_X1 U16384 ( .A1(n13674), .A2(n14051), .ZN(n13123) );
  NAND2_X1 U16385 ( .A1(n13674), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13122) );
  AND2_X1 U16386 ( .A1(n13123), .A2(n13122), .ZN(n19066) );
  INV_X1 U16387 ( .A(n19066), .ZN(n13124) );
  NAND2_X1 U16388 ( .A1(n13199), .A2(n13124), .ZN(n13195) );
  NAND2_X1 U16389 ( .A1(n13125), .A2(n13195), .ZN(P2_U2965) );
  AOI22_X1 U16390 ( .A1(P2_EAX_REG_25__SCAN_IN), .A2(n13130), .B1(n13207), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13129) );
  INV_X1 U16391 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13895) );
  OR2_X1 U16392 ( .A1(n13674), .A2(n13895), .ZN(n13127) );
  NAND2_X1 U16393 ( .A1(n13674), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13126) );
  AND2_X1 U16394 ( .A1(n13127), .A2(n13126), .ZN(n19077) );
  INV_X1 U16395 ( .A(n19077), .ZN(n13128) );
  NAND2_X1 U16396 ( .A1(n13199), .A2(n13128), .ZN(n13192) );
  NAND2_X1 U16397 ( .A1(n13129), .A2(n13192), .ZN(P2_U2961) );
  AOI22_X1 U16398 ( .A1(P2_EAX_REG_27__SCAN_IN), .A2(n13130), .B1(n13207), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13134) );
  INV_X1 U16399 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n14083) );
  OR2_X1 U16400 ( .A1(n13674), .A2(n14083), .ZN(n13132) );
  NAND2_X1 U16401 ( .A1(n13674), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13131) );
  AND2_X1 U16402 ( .A1(n13132), .A2(n13131), .ZN(n19072) );
  INV_X1 U16403 ( .A(n19072), .ZN(n13133) );
  NAND2_X1 U16404 ( .A1(n13199), .A2(n13133), .ZN(n13197) );
  NAND2_X1 U16405 ( .A1(n13134), .A2(n13197), .ZN(P2_U2963) );
  INV_X1 U16406 ( .A(n19873), .ZN(n13239) );
  AND2_X1 U16407 ( .A1(n13212), .A2(n13239), .ZN(n13135) );
  AND2_X1 U16408 ( .A1(n13220), .A2(n13219), .ZN(n13211) );
  NAND2_X1 U16409 ( .A1(n13211), .A2(n13239), .ZN(n13156) );
  NAND2_X1 U16410 ( .A1(n20677), .A2(n20481), .ZN(n19876) );
  INV_X1 U16411 ( .A(n19876), .ZN(n14067) );
  AOI21_X1 U16412 ( .B1(n13156), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n14067), 
        .ZN(n13136) );
  NAND2_X1 U16413 ( .A1(n13412), .A2(n13136), .ZN(P1_U2801) );
  INV_X1 U16414 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n20883) );
  NAND2_X1 U16415 ( .A1(n13674), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13138) );
  INV_X1 U16416 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16442) );
  OR2_X1 U16417 ( .A1(n13674), .A2(n16442), .ZN(n13137) );
  NAND2_X1 U16418 ( .A1(n13138), .A2(n13137), .ZN(n19069) );
  NAND2_X1 U16419 ( .A1(n13199), .A2(n19069), .ZN(n13149) );
  NAND2_X1 U16420 ( .A1(n13207), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13139) );
  OAI211_X1 U16421 ( .C1(n20883), .C2(n13270), .A(n13149), .B(n13139), .ZN(
        P2_U2964) );
  INV_X1 U16422 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19123) );
  NAND2_X1 U16423 ( .A1(n13199), .A2(n19063), .ZN(n13142) );
  NAND2_X1 U16424 ( .A1(n13207), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13140) );
  OAI211_X1 U16425 ( .C1(n19123), .C2(n13270), .A(n13142), .B(n13140), .ZN(
        P2_U2981) );
  INV_X1 U16426 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13321) );
  NAND2_X1 U16427 ( .A1(n13207), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13141) );
  OAI211_X1 U16428 ( .C1(n13321), .C2(n13270), .A(n13142), .B(n13141), .ZN(
        P2_U2966) );
  INV_X1 U16429 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13314) );
  NAND2_X1 U16430 ( .A1(n13674), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13144) );
  INV_X1 U16431 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16445) );
  OR2_X1 U16432 ( .A1(n13674), .A2(n16445), .ZN(n13143) );
  NAND2_X1 U16433 ( .A1(n13144), .A2(n13143), .ZN(n19074) );
  NAND2_X1 U16434 ( .A1(n13199), .A2(n19074), .ZN(n13147) );
  NAND2_X1 U16435 ( .A1(n13207), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13145) );
  OAI211_X1 U16436 ( .C1(n13314), .C2(n13270), .A(n13147), .B(n13145), .ZN(
        P2_U2962) );
  INV_X1 U16437 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19131) );
  NAND2_X1 U16438 ( .A1(n13207), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13146) );
  OAI211_X1 U16439 ( .C1(n19131), .C2(n13270), .A(n13147), .B(n13146), .ZN(
        P2_U2977) );
  INV_X1 U16440 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19127) );
  NAND2_X1 U16441 ( .A1(n13207), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13148) );
  OAI211_X1 U16442 ( .C1(n19127), .C2(n13270), .A(n13149), .B(n13148), .ZN(
        P2_U2979) );
  INV_X1 U16443 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13151) );
  INV_X1 U16444 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13150) );
  INV_X1 U16445 ( .A(n13207), .ZN(n13153) );
  INV_X1 U16446 ( .A(n13199), .ZN(n13155) );
  AOI22_X1 U16447 ( .A1(n13675), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13674), .ZN(n19060) );
  OAI222_X1 U16448 ( .A1(n13151), .A2(n13270), .B1(n13150), .B2(n13153), .C1(
        n13155), .C2(n19060), .ZN(P2_U2982) );
  INV_X1 U16449 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n13152) );
  OAI22_X1 U16450 ( .A1(n13674), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13675), .ZN(n13703) );
  OAI222_X1 U16451 ( .A1(n13263), .A2(n13270), .B1(n13152), .B2(n13153), .C1(
        n13155), .C2(n13703), .ZN(P2_U2967) );
  INV_X1 U16452 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13311) );
  INV_X1 U16453 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13154) );
  OAI222_X1 U16454 ( .A1(n13155), .A2(n13703), .B1(n13270), .B2(n13311), .C1(
        n13154), .C2(n13153), .ZN(P2_U2952) );
  OAI21_X1 U16455 ( .B1(n14067), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n20760), 
        .ZN(n13157) );
  OAI21_X1 U16456 ( .B1(n13158), .B2(n20760), .A(n13157), .ZN(P1_U3487) );
  INV_X1 U16457 ( .A(n16316), .ZN(n13159) );
  NOR2_X1 U16458 ( .A1(n10748), .A2(n13159), .ZN(n13160) );
  NAND2_X1 U16459 ( .A1(n13269), .A2(n13160), .ZN(n13165) );
  INV_X1 U16460 ( .A(n13161), .ZN(n13163) );
  NAND4_X1 U16461 ( .A1(n13165), .A2(n13164), .A3(n13163), .A4(n13162), .ZN(
        n16306) );
  NOR2_X1 U16462 ( .A1(n18828), .A2(n13274), .ZN(n16345) );
  AOI21_X1 U16463 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n18828), .A(n16345), 
        .ZN(n16357) );
  AOI21_X1 U16464 ( .B1(n18833), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16357), 
        .ZN(n13166) );
  AOI21_X1 U16465 ( .B1(n16306), .B2(n13167), .A(n13166), .ZN(n15602) );
  INV_X1 U16466 ( .A(n15602), .ZN(n13173) );
  NAND3_X1 U16467 ( .A1(n13171), .A2(n13170), .A3(n13169), .ZN(n16319) );
  OR3_X1 U16468 ( .A1(n15602), .A2(n15600), .A3(n16319), .ZN(n13172) );
  OAI21_X1 U16469 ( .B1(n13173), .B2(n16308), .A(n13172), .ZN(P2_U3595) );
  AOI22_X1 U16470 ( .A1(n13208), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13207), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13174) );
  AOI22_X1 U16471 ( .A1(n13675), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13674), .ZN(n19210) );
  INV_X1 U16472 ( .A(n19210), .ZN(n19086) );
  NAND2_X1 U16473 ( .A1(n13199), .A2(n19086), .ZN(n13181) );
  NAND2_X1 U16474 ( .A1(n13174), .A2(n13181), .ZN(P2_U2957) );
  AOI22_X1 U16475 ( .A1(n13208), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13207), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13175) );
  AOI22_X1 U16476 ( .A1(n13675), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13674), .ZN(n19197) );
  INV_X1 U16477 ( .A(n19197), .ZN(n13967) );
  NAND2_X1 U16478 ( .A1(n13199), .A2(n13967), .ZN(n13183) );
  NAND2_X1 U16479 ( .A1(n13175), .A2(n13183), .ZN(P2_U2953) );
  AOI22_X1 U16480 ( .A1(n13208), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13207), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13177) );
  AOI22_X1 U16481 ( .A1(n13675), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13674), .ZN(n19202) );
  INV_X1 U16482 ( .A(n19202), .ZN(n13176) );
  NAND2_X1 U16483 ( .A1(n13199), .A2(n13176), .ZN(n13179) );
  NAND2_X1 U16484 ( .A1(n13177), .A2(n13179), .ZN(P2_U2955) );
  AOI22_X1 U16485 ( .A1(n13208), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n13207), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n13178) );
  AOI22_X1 U16486 ( .A1(n13675), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13674), .ZN(n19225) );
  INV_X1 U16487 ( .A(n19225), .ZN(n15071) );
  NAND2_X1 U16488 ( .A1(n13199), .A2(n15071), .ZN(n13186) );
  NAND2_X1 U16489 ( .A1(n13178), .A2(n13186), .ZN(P2_U2974) );
  AOI22_X1 U16490 ( .A1(n13208), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n13207), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13180) );
  NAND2_X1 U16491 ( .A1(n13180), .A2(n13179), .ZN(P2_U2970) );
  AOI22_X1 U16492 ( .A1(n13208), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13207), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n13182) );
  NAND2_X1 U16493 ( .A1(n13182), .A2(n13181), .ZN(P2_U2972) );
  AOI22_X1 U16494 ( .A1(n13208), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n13207), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13184) );
  NAND2_X1 U16495 ( .A1(n13184), .A2(n13183), .ZN(P2_U2968) );
  AOI22_X1 U16496 ( .A1(n13208), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13207), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13185) );
  OAI22_X1 U16497 ( .A1(n13674), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13675), .ZN(n13678) );
  INV_X1 U16498 ( .A(n13678), .ZN(n16184) );
  NAND2_X1 U16499 ( .A1(n13199), .A2(n16184), .ZN(n13209) );
  NAND2_X1 U16500 ( .A1(n13185), .A2(n13209), .ZN(P2_U2969) );
  AOI22_X1 U16501 ( .A1(n13208), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13207), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13187) );
  NAND2_X1 U16502 ( .A1(n13187), .A2(n13186), .ZN(P2_U2959) );
  AOI22_X1 U16503 ( .A1(n13208), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n13207), .B2(
        P2_LWORD_REG_8__SCAN_IN), .ZN(n13191) );
  INV_X1 U16504 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n13769) );
  OR2_X1 U16505 ( .A1(n13674), .A2(n13769), .ZN(n13189) );
  NAND2_X1 U16506 ( .A1(n13674), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13188) );
  AND2_X1 U16507 ( .A1(n13189), .A2(n13188), .ZN(n19080) );
  INV_X1 U16508 ( .A(n19080), .ZN(n13190) );
  NAND2_X1 U16509 ( .A1(n13199), .A2(n13190), .ZN(n13205) );
  NAND2_X1 U16510 ( .A1(n13191), .A2(n13205), .ZN(P2_U2975) );
  AOI22_X1 U16511 ( .A1(n13208), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n13207), .B2(
        P2_LWORD_REG_9__SCAN_IN), .ZN(n13193) );
  NAND2_X1 U16512 ( .A1(n13193), .A2(n13192), .ZN(P2_U2976) );
  AOI22_X1 U16513 ( .A1(n13208), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13207), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n13194) );
  OAI22_X1 U16514 ( .A1(n13674), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13675), .ZN(n19214) );
  INV_X1 U16515 ( .A(n19214), .ZN(n16172) );
  NAND2_X1 U16516 ( .A1(n13199), .A2(n16172), .ZN(n13203) );
  NAND2_X1 U16517 ( .A1(n13194), .A2(n13203), .ZN(P2_U2973) );
  AOI22_X1 U16518 ( .A1(n13208), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13207), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13196) );
  NAND2_X1 U16519 ( .A1(n13196), .A2(n13195), .ZN(P2_U2980) );
  AOI22_X1 U16520 ( .A1(n13208), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n13207), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13198) );
  NAND2_X1 U16521 ( .A1(n13198), .A2(n13197), .ZN(P2_U2978) );
  AOI22_X1 U16522 ( .A1(n13208), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13207), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n13200) );
  INV_X1 U16523 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16453) );
  INV_X1 U16524 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18173) );
  AOI22_X1 U16525 ( .A1(n13675), .A2(n16453), .B1(n18173), .B2(n13674), .ZN(
        n19096) );
  NAND2_X1 U16526 ( .A1(n13199), .A2(n19096), .ZN(n13201) );
  NAND2_X1 U16527 ( .A1(n13200), .A2(n13201), .ZN(P2_U2971) );
  AOI22_X1 U16528 ( .A1(P2_EAX_REG_20__SCAN_IN), .A2(n13208), .B1(n13207), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13202) );
  NAND2_X1 U16529 ( .A1(n13202), .A2(n13201), .ZN(P2_U2956) );
  AOI22_X1 U16530 ( .A1(P2_EAX_REG_22__SCAN_IN), .A2(n13208), .B1(n13207), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13204) );
  NAND2_X1 U16531 ( .A1(n13204), .A2(n13203), .ZN(P2_U2958) );
  AOI22_X1 U16532 ( .A1(P2_EAX_REG_24__SCAN_IN), .A2(n13208), .B1(n13207), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13206) );
  NAND2_X1 U16533 ( .A1(n13206), .A2(n13205), .ZN(P2_U2960) );
  AOI22_X1 U16534 ( .A1(P2_EAX_REG_18__SCAN_IN), .A2(n13208), .B1(n13207), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13210) );
  NAND2_X1 U16535 ( .A1(n13210), .A2(n13209), .ZN(P2_U2954) );
  OAI22_X1 U16536 ( .A1(n13364), .A2(n13213), .B1(n13212), .B2(n13211), .ZN(
        n19874) );
  INV_X1 U16537 ( .A(n15804), .ZN(n15781) );
  OR2_X2 U16538 ( .A1(n13413), .A2(n20084), .ZN(n13381) );
  NAND3_X1 U16539 ( .A1(n13793), .A2(n15781), .A3(n13381), .ZN(n13214) );
  AND2_X1 U16540 ( .A1(n13214), .A2(n20691), .ZN(n20764) );
  NOR2_X1 U16541 ( .A1(n19874), .A2(n20764), .ZN(n15773) );
  OR2_X1 U16542 ( .A1(n15773), .A2(n19873), .ZN(n13226) );
  INV_X1 U16543 ( .A(n13226), .ZN(n19881) );
  INV_X1 U16544 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13228) );
  NOR2_X1 U16545 ( .A1(n11695), .A2(n20122), .ZN(n13215) );
  NAND4_X1 U16546 ( .A1(n11326), .A2(n13216), .A3(n13215), .A4(n13242), .ZN(
        n13217) );
  AND2_X1 U16547 ( .A1(n13218), .A2(n13217), .ZN(n13224) );
  NAND2_X1 U16548 ( .A1(n13364), .A2(n13342), .ZN(n13223) );
  INV_X1 U16549 ( .A(n13219), .ZN(n13221) );
  NAND2_X1 U16550 ( .A1(n13221), .A2(n13220), .ZN(n13222) );
  OAI211_X1 U16551 ( .C1(n13364), .C2(n13224), .A(n13223), .B(n13222), .ZN(
        n13225) );
  NAND2_X1 U16552 ( .A1(n13225), .A2(n20134), .ZN(n15774) );
  OR2_X1 U16553 ( .A1(n13226), .A2(n15774), .ZN(n13227) );
  OAI21_X1 U16554 ( .B1(n19881), .B2(n13228), .A(n13227), .ZN(P1_U3484) );
  NAND2_X1 U16555 ( .A1(n19196), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13230) );
  AND4_X1 U16556 ( .A1(n13230), .A2(n13229), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n10900), .ZN(n13231) );
  INV_X1 U16557 ( .A(n19830), .ZN(n19231) );
  NAND2_X1 U16558 ( .A1(n19231), .A2(n15018), .ZN(n13233) );
  NAND2_X1 U16559 ( .A1(n15022), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n13232) );
  OAI211_X1 U16560 ( .C1(n15022), .C2(n10260), .A(n13233), .B(n13232), .ZN(
        P2_U2887) );
  MUX2_X1 U16561 ( .A(n10214), .B(n13911), .S(n15027), .Z(n13238) );
  OAI21_X1 U16562 ( .B1(n19183), .B2(n15030), .A(n13238), .ZN(P2_U2886) );
  INV_X1 U16563 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13244) );
  NAND2_X1 U16564 ( .A1(n15804), .A2(n13239), .ZN(n13240) );
  AOI21_X1 U16565 ( .B1(n15760), .B2(n15782), .A(n13240), .ZN(n13241) );
  NAND2_X1 U16566 ( .A1(n20925), .A2(n13242), .ZN(n13483) );
  NAND2_X1 U16567 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16154) );
  INV_X1 U16568 ( .A(n16154), .ZN(n13592) );
  NAND2_X1 U16569 ( .A1(n20676), .A2(n13592), .ZN(n20761) );
  INV_X2 U16570 ( .A(n20761), .ZN(n20021) );
  AOI22_X1 U16571 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20021), .B1(n20007), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13243) );
  OAI21_X1 U16572 ( .B1(n13244), .B2(n13483), .A(n13243), .ZN(P1_U2920) );
  INV_X1 U16573 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13246) );
  AOI22_X1 U16574 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20021), .B1(n20007), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13245) );
  OAI21_X1 U16575 ( .B1(n13246), .B2(n13483), .A(n13245), .ZN(P1_U2915) );
  INV_X1 U16576 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13248) );
  AOI22_X1 U16577 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20021), .B1(n20007), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13247) );
  OAI21_X1 U16578 ( .B1(n13248), .B2(n13483), .A(n13247), .ZN(P1_U2918) );
  INV_X1 U16579 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13250) );
  AOI22_X1 U16580 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20021), .B1(n20007), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13249) );
  OAI21_X1 U16581 ( .B1(n13250), .B2(n13483), .A(n13249), .ZN(P1_U2916) );
  INV_X1 U16582 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13252) );
  AOI22_X1 U16583 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20021), .B1(n20007), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13251) );
  OAI21_X1 U16584 ( .B1(n13252), .B2(n13483), .A(n13251), .ZN(P1_U2919) );
  INV_X1 U16585 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13254) );
  AOI22_X1 U16586 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20021), .B1(n20007), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13253) );
  OAI21_X1 U16587 ( .B1(n13254), .B2(n13483), .A(n13253), .ZN(P1_U2917) );
  INV_X1 U16588 ( .A(n13703), .ZN(n19049) );
  INV_X1 U16589 ( .A(n19111), .ZN(n19054) );
  INV_X1 U16590 ( .A(n13256), .ZN(n13262) );
  INV_X1 U16591 ( .A(n13257), .ZN(n13260) );
  INV_X1 U16592 ( .A(n13258), .ZN(n13259) );
  NAND2_X1 U16593 ( .A1(n13260), .A2(n13259), .ZN(n13261) );
  NAND2_X1 U16594 ( .A1(n13262), .A2(n13261), .ZN(n19024) );
  OAI22_X1 U16595 ( .A1(n19054), .A2(n19024), .B1(n19083), .B2(n13263), .ZN(
        n13265) );
  NOR2_X1 U16596 ( .A1(n19830), .A2(n19024), .ZN(n19114) );
  AOI211_X1 U16597 ( .C1(n19830), .C2(n19024), .A(n19115), .B(n19114), .ZN(
        n13264) );
  AOI211_X1 U16598 ( .C1(n19049), .C2(n19085), .A(n13265), .B(n13264), .ZN(
        n13266) );
  INV_X1 U16599 ( .A(n13266), .ZN(P2_U2919) );
  INV_X1 U16600 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13276) );
  INV_X1 U16601 ( .A(n13267), .ZN(n13268) );
  NAND2_X1 U16602 ( .A1(n13269), .A2(n13268), .ZN(n13271) );
  NAND2_X1 U16603 ( .A1(n13271), .A2(n13270), .ZN(n13272) );
  INV_X1 U16604 ( .A(n19727), .ZN(n19854) );
  NAND2_X1 U16605 ( .A1(n19144), .A2(n13273), .ZN(n13320) );
  INV_X1 U16606 ( .A(n13274), .ZN(n19834) );
  NAND2_X1 U16607 ( .A1(n18828), .A2(n19834), .ZN(n19864) );
  INV_X2 U16608 ( .A(n19864), .ZN(n19152) );
  AOI22_X1 U16609 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n19151), .B1(n19152), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13275) );
  OAI21_X1 U16610 ( .B1(n13276), .B2(n13320), .A(n13275), .ZN(P2_U2928) );
  INV_X1 U16611 ( .A(n13277), .ZN(n15398) );
  NOR2_X1 U16612 ( .A1(n15400), .A2(n13293), .ZN(n13278) );
  AOI211_X1 U16613 ( .C1(n13293), .C2(n15398), .A(n16296), .B(n13278), .ZN(
        n13298) );
  NAND2_X1 U16614 ( .A1(n13280), .A2(n13279), .ZN(n13282) );
  AND2_X1 U16615 ( .A1(n13282), .A2(n9989), .ZN(n19812) );
  INV_X1 U16616 ( .A(n19812), .ZN(n13556) );
  INV_X1 U16617 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19742) );
  OR2_X1 U16618 ( .A1(n16264), .A2(n19742), .ZN(n19172) );
  AOI21_X1 U16619 ( .B1(n13285), .B2(n13284), .A(n13283), .ZN(n19170) );
  INV_X1 U16620 ( .A(n13286), .ZN(n13287) );
  AOI21_X1 U16621 ( .B1(n13289), .B2(n13288), .A(n13287), .ZN(n19168) );
  AOI22_X1 U16622 ( .A1(n16270), .A2(n19170), .B1(n16301), .B2(n19168), .ZN(
        n13290) );
  NAND2_X1 U16623 ( .A1(n19172), .A2(n13290), .ZN(n13291) );
  AOI211_X1 U16624 ( .C1(n13556), .C2(n16280), .A(n13292), .B(n13291), .ZN(
        n13296) );
  AOI22_X1 U16625 ( .A1(n13294), .A2(n13293), .B1(n14011), .B2(n16283), .ZN(
        n13295) );
  OAI211_X1 U16626 ( .C1(n13298), .C2(n13297), .A(n13296), .B(n13295), .ZN(
        P2_U3044) );
  INV_X1 U16627 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14020) );
  AOI22_X1 U16628 ( .A1(n19152), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13299) );
  OAI21_X1 U16629 ( .B1(n14020), .B2(n13320), .A(n13299), .ZN(P2_U2932) );
  INV_X1 U16630 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13301) );
  AOI22_X1 U16631 ( .A1(n19152), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13300) );
  OAI21_X1 U16632 ( .B1(n13301), .B2(n13320), .A(n13300), .ZN(P2_U2930) );
  INV_X1 U16633 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13303) );
  AOI22_X1 U16634 ( .A1(n19152), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13302) );
  OAI21_X1 U16635 ( .B1(n13303), .B2(n13320), .A(n13302), .ZN(P2_U2929) );
  INV_X1 U16636 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13305) );
  AOI22_X1 U16637 ( .A1(n19152), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13304) );
  OAI21_X1 U16638 ( .B1(n13305), .B2(n13320), .A(n13304), .ZN(P2_U2931) );
  INV_X1 U16639 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13307) );
  AOI22_X1 U16640 ( .A1(n19152), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13306) );
  OAI21_X1 U16641 ( .B1(n13307), .B2(n13320), .A(n13306), .ZN(P2_U2934) );
  INV_X1 U16642 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13309) );
  AOI22_X1 U16643 ( .A1(n19152), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13308) );
  OAI21_X1 U16644 ( .B1(n13309), .B2(n13320), .A(n13308), .ZN(P2_U2933) );
  AOI22_X1 U16645 ( .A1(n19152), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13310) );
  OAI21_X1 U16646 ( .B1(n13311), .B2(n13320), .A(n13310), .ZN(P2_U2935) );
  INV_X1 U16647 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n15058) );
  AOI22_X1 U16648 ( .A1(n19152), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13312) );
  OAI21_X1 U16649 ( .B1(n15058), .B2(n13320), .A(n13312), .ZN(P2_U2926) );
  AOI22_X1 U16650 ( .A1(n19152), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13313) );
  OAI21_X1 U16651 ( .B1(n13314), .B2(n13320), .A(n13313), .ZN(P2_U2925) );
  INV_X1 U16652 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15044) );
  AOI22_X1 U16653 ( .A1(n19152), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13315) );
  OAI21_X1 U16654 ( .B1(n15044), .B2(n13320), .A(n13315), .ZN(P2_U2924) );
  INV_X1 U16655 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n20823) );
  AOI22_X1 U16656 ( .A1(n19152), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13316) );
  OAI21_X1 U16657 ( .B1(n20823), .B2(n13320), .A(n13316), .ZN(P2_U2927) );
  AOI22_X1 U16658 ( .A1(n19152), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13317) );
  OAI21_X1 U16659 ( .B1(n20883), .B2(n13320), .A(n13317), .ZN(P2_U2923) );
  INV_X1 U16660 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n15033) );
  AOI22_X1 U16661 ( .A1(n19152), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13318) );
  OAI21_X1 U16662 ( .B1(n15033), .B2(n13320), .A(n13318), .ZN(P2_U2922) );
  AOI22_X1 U16663 ( .A1(n19152), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13319) );
  OAI21_X1 U16664 ( .B1(n13321), .B2(n13320), .A(n13319), .ZN(P2_U2921) );
  MUX2_X1 U16665 ( .A(n19178), .B(n10240), .S(n15022), .Z(n13327) );
  OAI21_X1 U16666 ( .B1(n19810), .B2(n15030), .A(n13327), .ZN(P2_U2885) );
  INV_X1 U16667 ( .A(n13329), .ZN(n13334) );
  NOR2_X1 U16668 ( .A1(n13074), .A2(n13331), .ZN(n13333) );
  NAND3_X1 U16669 ( .A1(n13334), .A2(n13333), .A3(n13332), .ZN(n14831) );
  NAND2_X1 U16670 ( .A1(n13328), .A2(n14831), .ZN(n13354) );
  NOR2_X1 U16671 ( .A1(n13336), .A2(n13345), .ZN(n13338) );
  AND2_X1 U16672 ( .A1(n13338), .A2(n13337), .ZN(n13355) );
  NAND2_X1 U16673 ( .A1(n11340), .A2(n13355), .ZN(n13351) );
  NAND2_X1 U16674 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13339) );
  MUX2_X1 U16675 ( .A(n13340), .B(n13339), .S(n13579), .Z(n13341) );
  INV_X1 U16676 ( .A(n13341), .ZN(n13349) );
  INV_X1 U16677 ( .A(n13342), .ZN(n13343) );
  NAND2_X1 U16678 ( .A1(n13344), .A2(n13343), .ZN(n13573) );
  NOR2_X1 U16679 ( .A1(n13347), .A2(n13346), .ZN(n13348) );
  AOI22_X1 U16680 ( .A1(n14834), .A2(n13349), .B1(n13573), .B2(n13348), .ZN(
        n13350) );
  OAI21_X1 U16681 ( .B1(n14831), .B2(n13351), .A(n13350), .ZN(n13352) );
  INV_X1 U16682 ( .A(n13352), .ZN(n13353) );
  NAND2_X1 U16683 ( .A1(n13354), .A2(n13353), .ZN(n13578) );
  INV_X1 U16684 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20841) );
  AOI22_X1 U16685 ( .A1(n13578), .A2(n16146), .B1(n13355), .B2(n14137), .ZN(
        n13371) );
  INV_X1 U16686 ( .A(n20112), .ZN(n13375) );
  NOR2_X1 U16687 ( .A1(n13375), .A2(n20084), .ZN(n13356) );
  NAND2_X1 U16688 ( .A1(n13357), .A2(n13356), .ZN(n13377) );
  NAND2_X1 U16689 ( .A1(n13377), .A2(n13358), .ZN(n13360) );
  NAND2_X1 U16690 ( .A1(n13360), .A2(n13359), .ZN(n13370) );
  INV_X1 U16691 ( .A(n13361), .ZN(n13367) );
  OAI211_X1 U16692 ( .C1(n14834), .C2(n13074), .A(n15804), .B(n20691), .ZN(
        n13362) );
  INV_X1 U16693 ( .A(n13362), .ZN(n13363) );
  NAND2_X1 U16694 ( .A1(n13364), .A2(n13363), .ZN(n13366) );
  AND4_X1 U16695 ( .A1(n13368), .A2(n13367), .A3(n13366), .A4(n13365), .ZN(
        n13369) );
  NAND2_X1 U16696 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13592), .ZN(n16158) );
  INV_X1 U16697 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19880) );
  OAI22_X1 U16698 ( .A1(n15765), .A2(n19873), .B1(n16158), .B2(n19880), .ZN(
        n16148) );
  AOI21_X1 U16699 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20676), .A(n16148), 
        .ZN(n14139) );
  INV_X1 U16700 ( .A(n14139), .ZN(n16151) );
  MUX2_X1 U16701 ( .A(n13579), .B(n13371), .S(n16151), .Z(n13372) );
  INV_X1 U16702 ( .A(n13372), .ZN(P1_U3469) );
  OAI21_X1 U16703 ( .B1(n13374), .B2(n13373), .A(n13511), .ZN(n13877) );
  NAND4_X1 U16704 ( .A1(n9680), .A2(n13384), .A3(n13530), .A4(n13375), .ZN(
        n13376) );
  NAND2_X1 U16705 ( .A1(n13377), .A2(n13376), .ZN(n13379) );
  NOR2_X1 U16706 ( .A1(n20107), .A2(n19873), .ZN(n13378) );
  INV_X1 U16707 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14838) );
  XNOR2_X1 U16708 ( .A(n13499), .B(n13382), .ZN(n13500) );
  XNOR2_X1 U16709 ( .A(n13500), .B(n13530), .ZN(n13874) );
  AOI22_X1 U16710 ( .A1(n19989), .A2(n13874), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n14438), .ZN(n13383) );
  OAI21_X1 U16711 ( .B1(n13877), .B2(n14455), .A(n13383), .ZN(P1_U2871) );
  NAND2_X1 U16712 ( .A1(n13384), .A2(n20134), .ZN(n13390) );
  AND2_X1 U16713 ( .A1(n13390), .A2(n13385), .ZN(n13386) );
  INV_X1 U16714 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n13387) );
  OR2_X1 U16715 ( .A1(n20080), .A2(n13387), .ZN(n13389) );
  NAND2_X1 U16716 ( .A1(n20080), .A2(DATAI_1_), .ZN(n13388) );
  AND2_X1 U16717 ( .A1(n13389), .A2(n13388), .ZN(n20104) );
  INV_X1 U16718 ( .A(n13390), .ZN(n13391) );
  INV_X1 U16719 ( .A(n15959), .ZN(n13393) );
  INV_X1 U16720 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20020) );
  OAI222_X1 U16721 ( .A1(n14544), .A2(n13877), .B1(n20104), .B2(n14542), .C1(
        n14540), .C2(n20020), .ZN(P1_U2903) );
  NAND2_X1 U16722 ( .A1(n13395), .A2(n13394), .ZN(n13396) );
  NAND2_X1 U16723 ( .A1(n13397), .A2(n13396), .ZN(n20064) );
  OR2_X1 U16724 ( .A1(n20080), .A2(n16462), .ZN(n13399) );
  NAND2_X1 U16725 ( .A1(n20080), .A2(DATAI_0_), .ZN(n13398) );
  AND2_X1 U16726 ( .A1(n13399), .A2(n13398), .ZN(n20093) );
  INV_X1 U16727 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20024) );
  OAI222_X1 U16728 ( .A1(n14544), .A2(n20064), .B1(n20093), .B2(n14542), .C1(
        n14540), .C2(n20024), .ZN(P1_U2904) );
  OR2_X1 U16729 ( .A1(n13400), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13401) );
  NAND2_X1 U16730 ( .A1(n13402), .A2(n13401), .ZN(n16304) );
  OR2_X1 U16731 ( .A1(n18992), .A2(n18848), .ZN(n16302) );
  AOI21_X1 U16732 ( .B1(n19028), .B2(n13404), .A(n13403), .ZN(n16300) );
  NAND2_X1 U16733 ( .A1(n19167), .A2(n16300), .ZN(n13405) );
  OAI211_X1 U16734 ( .C1(n16245), .C2(n16304), .A(n16302), .B(n13405), .ZN(
        n13406) );
  INV_X1 U16735 ( .A(n13406), .ZN(n13409) );
  OAI21_X1 U16736 ( .B1(n19166), .B2(n13407), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13408) );
  OAI211_X1 U16737 ( .C1(n19179), .C2(n10260), .A(n13409), .B(n13408), .ZN(
        P2_U3014) );
  NOR2_X1 U16738 ( .A1(n13410), .A2(n20691), .ZN(n13411) );
  NOR2_X2 U16739 ( .A1(n20052), .A2(n13413), .ZN(n20038) );
  INV_X1 U16740 ( .A(n20104), .ZN(n14526) );
  NAND2_X1 U16741 ( .A1(n20038), .A2(n14526), .ZN(n13417) );
  AND2_X2 U16742 ( .A1(n13414), .A2(n13413), .ZN(n20053) );
  AOI22_X1 U16743 ( .A1(n20053), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20052), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13415) );
  NAND2_X1 U16744 ( .A1(n13417), .A2(n13415), .ZN(P1_U2938) );
  AOI22_X1 U16745 ( .A1(n20053), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20052), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13416) );
  NAND2_X1 U16746 ( .A1(n13417), .A2(n13416), .ZN(P1_U2953) );
  INV_X1 U16747 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n13418) );
  OR2_X1 U16748 ( .A1(n20080), .A2(n13418), .ZN(n13420) );
  NAND2_X1 U16749 ( .A1(n20080), .A2(DATAI_6_), .ZN(n13419) );
  AND2_X1 U16750 ( .A1(n13420), .A2(n13419), .ZN(n20128) );
  INV_X1 U16751 ( .A(n20128), .ZN(n14495) );
  NAND2_X1 U16752 ( .A1(n20038), .A2(n14495), .ZN(n13448) );
  AOI22_X1 U16753 ( .A1(n20053), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20052), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13421) );
  NAND2_X1 U16754 ( .A1(n13448), .A2(n13421), .ZN(P1_U2943) );
  INV_X1 U16755 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n13422) );
  OR2_X1 U16756 ( .A1(n20080), .A2(n13422), .ZN(n13424) );
  NAND2_X1 U16757 ( .A1(n20080), .A2(DATAI_7_), .ZN(n13423) );
  AND2_X1 U16758 ( .A1(n13424), .A2(n13423), .ZN(n20137) );
  INV_X1 U16759 ( .A(n20137), .ZN(n15958) );
  NAND2_X1 U16760 ( .A1(n20038), .A2(n15958), .ZN(n13450) );
  AOI22_X1 U16761 ( .A1(n20053), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20052), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13425) );
  NAND2_X1 U16762 ( .A1(n13450), .A2(n13425), .ZN(P1_U2944) );
  INV_X1 U16763 ( .A(n20093), .ZN(n14533) );
  NAND2_X1 U16764 ( .A1(n20038), .A2(n14533), .ZN(n13428) );
  AOI22_X1 U16765 ( .A1(n20053), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20052), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13426) );
  NAND2_X1 U16766 ( .A1(n13428), .A2(n13426), .ZN(P1_U2937) );
  AOI22_X1 U16767 ( .A1(n20053), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20052), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13427) );
  NAND2_X1 U16768 ( .A1(n13428), .A2(n13427), .ZN(P1_U2952) );
  INV_X1 U16769 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n13429) );
  OR2_X1 U16770 ( .A1(n20080), .A2(n13429), .ZN(n13431) );
  NAND2_X1 U16771 ( .A1(n20080), .A2(DATAI_3_), .ZN(n13430) );
  AND2_X1 U16772 ( .A1(n13431), .A2(n13430), .ZN(n20114) );
  INV_X1 U16773 ( .A(n20114), .ZN(n14514) );
  NAND2_X1 U16774 ( .A1(n20038), .A2(n14514), .ZN(n13444) );
  AOI22_X1 U16775 ( .A1(n20053), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20052), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13432) );
  NAND2_X1 U16776 ( .A1(n13444), .A2(n13432), .ZN(P1_U2940) );
  OR2_X1 U16777 ( .A1(n20080), .A2(n16453), .ZN(n13434) );
  NAND2_X1 U16778 ( .A1(n20080), .A2(DATAI_4_), .ZN(n13433) );
  AND2_X1 U16779 ( .A1(n13434), .A2(n13433), .ZN(n20119) );
  INV_X1 U16780 ( .A(n20119), .ZN(n14507) );
  NAND2_X1 U16781 ( .A1(n20038), .A2(n14507), .ZN(n13454) );
  AOI22_X1 U16782 ( .A1(n20053), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20052), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13435) );
  NAND2_X1 U16783 ( .A1(n13454), .A2(n13435), .ZN(P1_U2941) );
  INV_X1 U16784 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n13436) );
  OR2_X1 U16785 ( .A1(n20080), .A2(n13436), .ZN(n13438) );
  NAND2_X1 U16786 ( .A1(n20080), .A2(DATAI_2_), .ZN(n13437) );
  AND2_X1 U16787 ( .A1(n13438), .A2(n13437), .ZN(n20109) );
  INV_X1 U16788 ( .A(n20109), .ZN(n14520) );
  NAND2_X1 U16789 ( .A1(n20038), .A2(n14520), .ZN(n13452) );
  AOI22_X1 U16790 ( .A1(n20053), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20052), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13439) );
  NAND2_X1 U16791 ( .A1(n13452), .A2(n13439), .ZN(P1_U2939) );
  OR2_X1 U16792 ( .A1(n20080), .A2(n20825), .ZN(n13441) );
  NAND2_X1 U16793 ( .A1(n20080), .A2(DATAI_5_), .ZN(n13440) );
  AND2_X1 U16794 ( .A1(n13441), .A2(n13440), .ZN(n20124) );
  INV_X1 U16795 ( .A(n20124), .ZN(n14501) );
  NAND2_X1 U16796 ( .A1(n20038), .A2(n14501), .ZN(n13446) );
  AOI22_X1 U16797 ( .A1(n20053), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20052), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13442) );
  NAND2_X1 U16798 ( .A1(n13446), .A2(n13442), .ZN(P1_U2942) );
  AOI22_X1 U16799 ( .A1(n20053), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20052), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13443) );
  NAND2_X1 U16800 ( .A1(n13444), .A2(n13443), .ZN(P1_U2955) );
  AOI22_X1 U16801 ( .A1(n20053), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20052), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13445) );
  NAND2_X1 U16802 ( .A1(n13446), .A2(n13445), .ZN(P1_U2957) );
  AOI22_X1 U16803 ( .A1(n20053), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20052), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13447) );
  NAND2_X1 U16804 ( .A1(n13448), .A2(n13447), .ZN(P1_U2958) );
  AOI22_X1 U16805 ( .A1(n20053), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20052), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13449) );
  NAND2_X1 U16806 ( .A1(n13450), .A2(n13449), .ZN(P1_U2959) );
  AOI22_X1 U16807 ( .A1(n20053), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20052), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13451) );
  NAND2_X1 U16808 ( .A1(n13452), .A2(n13451), .ZN(P1_U2954) );
  AOI22_X1 U16809 ( .A1(n20053), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20052), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13453) );
  NAND2_X1 U16810 ( .A1(n13454), .A2(n13453), .ZN(P1_U2956) );
  XNOR2_X1 U16811 ( .A(n13455), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13490) );
  INV_X1 U16812 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20749) );
  NOR2_X1 U16813 ( .A1(n16041), .A2(n20749), .ZN(n13485) );
  AOI211_X1 U16814 ( .C1(n14837), .C2(n13497), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n14695), .ZN(n13456) );
  AOI211_X1 U16815 ( .C1(n20067), .C2(n13874), .A(n13485), .B(n13456), .ZN(
        n13459) );
  OAI21_X1 U16816 ( .B1(n13457), .B2(n13494), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13458) );
  OAI211_X1 U16817 ( .C1(n13490), .C2(n16070), .A(n13459), .B(n13458), .ZN(
        P1_U3030) );
  MUX2_X1 U16818 ( .A(n10253), .B(n10287), .S(n15027), .Z(n13464) );
  OAI21_X1 U16819 ( .B1(n19235), .B2(n15030), .A(n13464), .ZN(P2_U2884) );
  INV_X1 U16820 ( .A(n13841), .ZN(n13465) );
  OAI222_X1 U16821 ( .A1(n20064), .A2(n14455), .B1(n13109), .B2(n19994), .C1(
        n13465), .C2(n14457), .ZN(P1_U2872) );
  INV_X1 U16822 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13467) );
  AOI22_X1 U16823 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13466) );
  OAI21_X1 U16824 ( .B1(n13467), .B2(n13483), .A(n13466), .ZN(P1_U2907) );
  INV_X1 U16825 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13469) );
  AOI22_X1 U16826 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13468) );
  OAI21_X1 U16827 ( .B1(n13469), .B2(n13483), .A(n13468), .ZN(P1_U2914) );
  INV_X1 U16828 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13471) );
  AOI22_X1 U16829 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13470) );
  OAI21_X1 U16830 ( .B1(n13471), .B2(n13483), .A(n13470), .ZN(P1_U2906) );
  INV_X1 U16831 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13473) );
  AOI22_X1 U16832 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13472) );
  OAI21_X1 U16833 ( .B1(n13473), .B2(n13483), .A(n13472), .ZN(P1_U2912) );
  INV_X1 U16834 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13475) );
  AOI22_X1 U16835 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13474) );
  OAI21_X1 U16836 ( .B1(n13475), .B2(n13483), .A(n13474), .ZN(P1_U2908) );
  INV_X1 U16837 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13477) );
  AOI22_X1 U16838 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13476) );
  OAI21_X1 U16839 ( .B1(n13477), .B2(n13483), .A(n13476), .ZN(P1_U2911) );
  INV_X1 U16840 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13479) );
  AOI22_X1 U16841 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13478) );
  OAI21_X1 U16842 ( .B1(n13479), .B2(n13483), .A(n13478), .ZN(P1_U2910) );
  INV_X1 U16843 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13481) );
  AOI22_X1 U16844 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13480) );
  OAI21_X1 U16845 ( .B1(n13481), .B2(n13483), .A(n13480), .ZN(P1_U2913) );
  INV_X1 U16846 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13484) );
  AOI22_X1 U16847 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13482) );
  OAI21_X1 U16848 ( .B1(n13484), .B2(n13483), .A(n13482), .ZN(P1_U2909) );
  INV_X1 U16849 ( .A(n13877), .ZN(n13488) );
  AOI21_X1 U16850 ( .B1(n20058), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13485), .ZN(n13486) );
  OAI21_X1 U16851 ( .B1(n16034), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13486), .ZN(n13487) );
  AOI21_X1 U16852 ( .B1(n13488), .B2(n16031), .A(n13487), .ZN(n13489) );
  OAI21_X1 U16853 ( .B1(n13490), .B2(n19879), .A(n13489), .ZN(P1_U2998) );
  XNOR2_X1 U16854 ( .A(n13492), .B(n13491), .ZN(n13565) );
  INV_X1 U16855 ( .A(n14805), .ZN(n13495) );
  NOR2_X1 U16856 ( .A1(n13498), .A2(n14838), .ZN(n14033) );
  NOR2_X1 U16857 ( .A1(n13494), .A2(n13493), .ZN(n14788) );
  OAI21_X1 U16858 ( .B1(n13495), .B2(n14033), .A(n14788), .ZN(n13617) );
  NAND2_X1 U16859 ( .A1(n14692), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13496) );
  NAND2_X1 U16860 ( .A1(n13497), .A2(n13496), .ZN(n16117) );
  NAND3_X1 U16861 ( .A1(n16117), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n13498), .ZN(n13508) );
  AOI21_X1 U16862 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13776) );
  OAI221_X1 U16863 ( .B1(n13776), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .C1(
        n13776), .C2(n14033), .A(n14690), .ZN(n13507) );
  AOI21_X1 U16864 ( .B1(n13500), .B2(n13530), .A(n13499), .ZN(n13529) );
  BUF_X2 U16865 ( .A(n13501), .Z(n14179) );
  MUX2_X1 U16866 ( .A(n14179), .B(n14276), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n13503) );
  NOR2_X1 U16867 ( .A1(n14277), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13502) );
  NOR2_X1 U16868 ( .A1(n13503), .A2(n13502), .ZN(n13528) );
  XNOR2_X1 U16869 ( .A(n13529), .B(n13528), .ZN(n14370) );
  INV_X1 U16870 ( .A(n14370), .ZN(n13505) );
  INV_X1 U16871 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13504) );
  NOR2_X1 U16872 ( .A1(n16041), .A2(n13504), .ZN(n13560) );
  AOI21_X1 U16873 ( .B1(n20067), .B2(n13505), .A(n13560), .ZN(n13506) );
  NAND3_X1 U16874 ( .A1(n13508), .A2(n13507), .A3(n13506), .ZN(n13509) );
  AOI21_X1 U16875 ( .B1(n13617), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n13509), .ZN(n13510) );
  OAI21_X1 U16876 ( .B1(n16070), .B2(n13565), .A(n13510), .ZN(P1_U3029) );
  INV_X1 U16877 ( .A(n13511), .ZN(n13513) );
  OAI21_X1 U16878 ( .B1(n9676), .B2(n13513), .A(n13512), .ZN(n14375) );
  INV_X1 U16879 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13514) );
  OAI222_X1 U16880 ( .A1(n14375), .A2(n14455), .B1(n13514), .B2(n19994), .C1(
        n14370), .C2(n14457), .ZN(P1_U2870) );
  INV_X1 U16881 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n13515) );
  OAI222_X1 U16882 ( .A1(n14375), .A2(n14544), .B1(n20109), .B2(n14542), .C1(
        n13515), .C2(n14540), .ZN(P1_U2902) );
  NAND2_X1 U16883 ( .A1(n13516), .A2(n13518), .ZN(n13540) );
  AND2_X1 U16884 ( .A1(n19213), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13517) );
  OR2_X1 U16885 ( .A1(n13518), .A2(n13517), .ZN(n13519) );
  OR2_X1 U16886 ( .A1(n13516), .A2(n13519), .ZN(n13520) );
  NAND2_X1 U16887 ( .A1(n13540), .A2(n13520), .ZN(n19098) );
  OR2_X1 U16888 ( .A1(n13522), .A2(n13521), .ZN(n13523) );
  NAND2_X1 U16889 ( .A1(n13523), .A2(n13541), .ZN(n19160) );
  MUX2_X1 U16890 ( .A(n10774), .B(n19160), .S(n15027), .Z(n13524) );
  OAI21_X1 U16891 ( .B1(n19098), .B2(n15030), .A(n13524), .ZN(P2_U2883) );
  OAI21_X1 U16892 ( .B1(n13527), .B2(n13526), .A(n13525), .ZN(n13818) );
  NAND2_X1 U16893 ( .A1(n13529), .A2(n13528), .ZN(n13536) );
  INV_X1 U16894 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13531) );
  NAND2_X1 U16895 ( .A1(n14273), .A2(n13531), .ZN(n13534) );
  NAND2_X1 U16896 ( .A1(n9581), .A2(n13775), .ZN(n13532) );
  OAI211_X1 U16897 ( .C1(n13381), .C2(P1_EBX_REG_3__SCAN_IN), .A(n13532), .B(
        n14290), .ZN(n13533) );
  AND2_X1 U16898 ( .A1(n13534), .A2(n13533), .ZN(n13535) );
  NAND2_X1 U16899 ( .A1(n13536), .A2(n13535), .ZN(n13537) );
  NAND2_X1 U16900 ( .A1(n13627), .A2(n13537), .ZN(n13616) );
  INV_X1 U16901 ( .A(n13616), .ZN(n13805) );
  AOI22_X1 U16902 ( .A1(n19989), .A2(n13805), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14438), .ZN(n13538) );
  OAI21_X1 U16903 ( .B1(n13818), .B2(n14455), .A(n13538), .ZN(P1_U2869) );
  INV_X1 U16904 ( .A(n13540), .ZN(n13635) );
  OR2_X1 U16905 ( .A1(n13540), .A2(n13539), .ZN(n13602) );
  OAI211_X1 U16906 ( .C1(n13635), .C2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n15018), .B(n13602), .ZN(n13548) );
  NAND2_X1 U16907 ( .A1(n13542), .A2(n13541), .ZN(n13545) );
  INV_X1 U16908 ( .A(n13543), .ZN(n13544) );
  INV_X1 U16909 ( .A(n19001), .ZN(n13546) );
  MUX2_X1 U16910 ( .A(n18994), .B(n13546), .S(n15027), .Z(n13547) );
  NAND2_X1 U16911 ( .A1(n13548), .A2(n13547), .ZN(P2_U2882) );
  XNOR2_X1 U16912 ( .A(n19810), .B(n19812), .ZN(n13555) );
  XNOR2_X1 U16913 ( .A(n13550), .B(n13549), .ZN(n19826) );
  INV_X1 U16914 ( .A(n19826), .ZN(n13551) );
  NAND2_X1 U16915 ( .A1(n19183), .A2(n13551), .ZN(n13552) );
  OAI21_X1 U16916 ( .B1(n19183), .B2(n13551), .A(n13552), .ZN(n19113) );
  NOR2_X1 U16917 ( .A1(n19113), .A2(n19114), .ZN(n19112) );
  INV_X1 U16918 ( .A(n13552), .ZN(n13553) );
  NOR2_X1 U16919 ( .A1(n19112), .A2(n13553), .ZN(n13554) );
  NOR2_X1 U16920 ( .A1(n13554), .A2(n13555), .ZN(n19087) );
  AOI21_X1 U16921 ( .B1(n13555), .B2(n13554), .A(n19087), .ZN(n13559) );
  AOI22_X1 U16922 ( .A1(n19085), .A2(n16184), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19110), .ZN(n13558) );
  NAND2_X1 U16923 ( .A1(n13556), .A2(n19111), .ZN(n13557) );
  OAI211_X1 U16924 ( .C1(n13559), .C2(n19115), .A(n13558), .B(n13557), .ZN(
        P2_U2917) );
  INV_X1 U16925 ( .A(n14375), .ZN(n13563) );
  AOI21_X1 U16926 ( .B1(n20058), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13560), .ZN(n13561) );
  OAI21_X1 U16927 ( .B1(n16034), .B2(n14365), .A(n13561), .ZN(n13562) );
  AOI21_X1 U16928 ( .B1(n13563), .B2(n16031), .A(n13562), .ZN(n13564) );
  OAI21_X1 U16929 ( .B1(n19879), .B2(n13565), .A(n13564), .ZN(P1_U2997) );
  INV_X1 U16930 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13566) );
  OR2_X1 U16931 ( .A1(n20080), .A2(n13566), .ZN(n13568) );
  NAND2_X1 U16932 ( .A1(n20080), .A2(DATAI_15_), .ZN(n13567) );
  NAND2_X1 U16933 ( .A1(n13568), .A2(n13567), .ZN(n14539) );
  AOI222_X1 U16934 ( .A1(n20052), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20053), 
        .B2(P1_EAX_REG_15__SCAN_IN), .C1(n14539), .C2(n20038), .ZN(n13569) );
  INV_X1 U16935 ( .A(n13569), .ZN(P1_U2967) );
  INV_X1 U16936 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20017) );
  OAI222_X1 U16937 ( .A1(n14544), .A2(n13818), .B1(n20114), .B2(n14542), .C1(
        n14540), .C2(n20017), .ZN(P1_U2901) );
  NOR2_X1 U16938 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20677), .ZN(n13582) );
  INV_X1 U16939 ( .A(n14848), .ZN(n13570) );
  NAND2_X1 U16940 ( .A1(n11340), .A2(n13570), .ZN(n13577) );
  INV_X1 U16941 ( .A(n13572), .ZN(n20091) );
  NAND2_X1 U16942 ( .A1(n20091), .A2(n14831), .ZN(n13576) );
  XNOR2_X1 U16943 ( .A(n20888), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13574) );
  AOI22_X1 U16944 ( .A1(n14834), .A2(n13574), .B1(n13573), .B2(n14848), .ZN(
        n13575) );
  OAI211_X1 U16945 ( .C1(n14831), .C2(n13577), .A(n13576), .B(n13575), .ZN(
        n14846) );
  MUX2_X1 U16946 ( .A(n14846), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15765), .Z(n15767) );
  AOI22_X1 U16947 ( .A1(n13582), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n20677), .B2(n15767), .ZN(n13584) );
  OR2_X1 U16948 ( .A1(n15765), .A2(n13578), .ZN(n13581) );
  NAND2_X1 U16949 ( .A1(n15765), .A2(n13579), .ZN(n13580) );
  AND2_X1 U16950 ( .A1(n13581), .A2(n13580), .ZN(n15768) );
  AOI22_X1 U16951 ( .A1(n13582), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n15768), .B2(n20677), .ZN(n13583) );
  NOR2_X1 U16952 ( .A1(n13584), .A2(n13583), .ZN(n15771) );
  INV_X1 U16953 ( .A(n14830), .ZN(n13585) );
  NAND2_X1 U16954 ( .A1(n15771), .A2(n13585), .ZN(n13593) );
  MUX2_X1 U16955 ( .A(n19880), .B(n15765), .S(n20677), .Z(n13590) );
  INV_X1 U16956 ( .A(n20250), .ZN(n20510) );
  OR2_X1 U16957 ( .A1(n11453), .A2(n20510), .ZN(n13587) );
  XNOR2_X1 U16958 ( .A(n13587), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19967) );
  NAND2_X1 U16959 ( .A1(n19967), .A2(n13588), .ZN(n16145) );
  NOR2_X1 U16960 ( .A1(n16145), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13589) );
  AOI21_X1 U16961 ( .B1(n13590), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13589), .ZN(n15777) );
  AND3_X1 U16962 ( .A1(n13593), .A2(n15777), .A3(n19880), .ZN(n13591) );
  NOR2_X1 U16963 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20763) );
  OAI21_X1 U16964 ( .B1(n13591), .B2(n16158), .A(n20257), .ZN(n20077) );
  NAND3_X1 U16965 ( .A1(n13593), .A2(n15777), .A3(n13592), .ZN(n15788) );
  INV_X1 U16966 ( .A(n15788), .ZN(n13595) );
  INV_X1 U16967 ( .A(n11712), .ZN(n13843) );
  AND2_X1 U16968 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20841), .ZN(n14827) );
  OAI22_X1 U16969 ( .A1(n20171), .A2(n20620), .B1(n13843), .B2(n14827), .ZN(
        n13594) );
  OAI21_X1 U16970 ( .B1(n13595), .B2(n13594), .A(n20077), .ZN(n13596) );
  OAI21_X1 U16971 ( .B1(n20077), .B2(n20536), .A(n13596), .ZN(P1_U3478) );
  XOR2_X1 U16972 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B(n13602), .Z(n13600)
         );
  OR2_X1 U16973 ( .A1(n13597), .A2(n13543), .ZN(n13598) );
  NAND2_X1 U16974 ( .A1(n13605), .A2(n13598), .ZN(n18986) );
  MUX2_X1 U16975 ( .A(n10780), .B(n18986), .S(n15027), .Z(n13599) );
  OAI21_X1 U16976 ( .B1(n13600), .B2(n15030), .A(n13599), .ZN(P2_U2881) );
  NOR2_X1 U16977 ( .A1(n13602), .A2(n13601), .ZN(n13603) );
  XNOR2_X1 U16978 ( .A(n13603), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13608) );
  NAND2_X1 U16979 ( .A1(n13605), .A2(n13604), .ZN(n13606) );
  NAND2_X1 U16980 ( .A1(n13631), .A2(n13606), .ZN(n18976) );
  MUX2_X1 U16981 ( .A(n10786), .B(n18976), .S(n15027), .Z(n13607) );
  OAI21_X1 U16982 ( .B1(n13608), .B2(n15030), .A(n13607), .ZN(P2_U2880) );
  XNOR2_X1 U16983 ( .A(n13610), .B(n13609), .ZN(n13621) );
  INV_X1 U16984 ( .A(n13818), .ZN(n13613) );
  NAND2_X1 U16985 ( .A1(n16139), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n13615) );
  NAND2_X1 U16986 ( .A1(n20058), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13611) );
  OAI211_X1 U16987 ( .C1(n16034), .C2(n13806), .A(n13615), .B(n13611), .ZN(
        n13612) );
  AOI21_X1 U16988 ( .B1(n13613), .B2(n16031), .A(n13612), .ZN(n13614) );
  OAI21_X1 U16989 ( .B1(n13621), .B2(n19879), .A(n13614), .ZN(P1_U2996) );
  AOI21_X1 U16990 ( .B1(n14033), .B2(n16117), .A(n14690), .ZN(n16093) );
  OAI21_X1 U16991 ( .B1(n16069), .B2(n13616), .A(n13615), .ZN(n13619) );
  AOI21_X1 U16992 ( .B1(n14690), .B2(n13776), .A(n13617), .ZN(n20069) );
  NOR2_X1 U16993 ( .A1(n20069), .A2(n13775), .ZN(n13618) );
  AOI211_X1 U16994 ( .C1(n20074), .C2(n13775), .A(n13619), .B(n13618), .ZN(
        n13620) );
  OAI21_X1 U16995 ( .B1(n16070), .B2(n13621), .A(n13620), .ZN(P1_U3028) );
  NAND2_X1 U16996 ( .A1(n13525), .A2(n13622), .ZN(n13623) );
  AND2_X1 U16997 ( .A1(n13647), .A2(n13623), .ZN(n19984) );
  INV_X1 U16998 ( .A(n19984), .ZN(n13630) );
  INV_X1 U16999 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13629) );
  NAND2_X1 U17000 ( .A1(n14179), .A2(n13629), .ZN(n13626) );
  NAND2_X1 U17001 ( .A1(n14290), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13624) );
  OAI211_X1 U17002 ( .C1(P1_EBX_REG_4__SCAN_IN), .C2(n13381), .A(n13624), .B(
        n9581), .ZN(n13625) );
  NAND2_X1 U17003 ( .A1(n13626), .A2(n13625), .ZN(n13628) );
  NOR2_X2 U17004 ( .A1(n13627), .A2(n13628), .ZN(n13666) );
  AOI21_X1 U17005 ( .B1(n13628), .B2(n13627), .A(n13666), .ZN(n20066) );
  INV_X1 U17006 ( .A(n20066), .ZN(n19976) );
  OAI222_X1 U17007 ( .A1(n13630), .A2(n14455), .B1(n13629), .B2(n19994), .C1(
        n19976), .C2(n14457), .ZN(P1_U2868) );
  INV_X1 U17008 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20015) );
  OAI222_X1 U17009 ( .A1(n13630), .A2(n14544), .B1(n20119), .B2(n14542), .C1(
        n20015), .C2(n14540), .ZN(P1_U2900) );
  INV_X1 U17010 ( .A(n13631), .ZN(n13633) );
  OAI21_X1 U17011 ( .B1(n13633), .B2(n10043), .A(n13642), .ZN(n16235) );
  AND2_X1 U17012 ( .A1(n13635), .A2(n13634), .ZN(n13711) );
  INV_X1 U17013 ( .A(n13711), .ZN(n13637) );
  OR2_X1 U17014 ( .A1(n13637), .A2(n13636), .ZN(n13653) );
  OAI211_X1 U17015 ( .C1(n13711), .C2(n13638), .A(n15018), .B(n13653), .ZN(
        n13640) );
  NAND2_X1 U17016 ( .A1(n15022), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13639) );
  OAI211_X1 U17017 ( .C1(n16235), .C2(n15022), .A(n13640), .B(n13639), .ZN(
        P2_U2879) );
  XNOR2_X1 U17018 ( .A(n13653), .B(n13652), .ZN(n13645) );
  AND2_X1 U17019 ( .A1(n13642), .A2(n13641), .ZN(n13643) );
  OR2_X1 U17020 ( .A1(n13643), .A2(n13656), .ZN(n18966) );
  MUX2_X1 U17021 ( .A(n10793), .B(n18966), .S(n15027), .Z(n13644) );
  OAI21_X1 U17022 ( .B1(n13645), .B2(n15030), .A(n13644), .ZN(P2_U2878) );
  AND2_X1 U17023 ( .A1(n13647), .A2(n13646), .ZN(n13649) );
  OR2_X1 U17024 ( .A1(n13649), .A2(n13648), .ZN(n19959) );
  INV_X1 U17025 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20013) );
  OAI222_X1 U17026 ( .A1(n14544), .A2(n19959), .B1(n20124), .B2(n14542), .C1(
        n14540), .C2(n20013), .ZN(P1_U2899) );
  OAI21_X1 U17027 ( .B1(n13653), .B2(n13652), .A(n13651), .ZN(n13654) );
  NAND3_X1 U17028 ( .A1(n13714), .A2(n13654), .A3(n15018), .ZN(n13659) );
  OR2_X1 U17029 ( .A1(n13656), .A2(n13655), .ZN(n13657) );
  AND2_X1 U17030 ( .A1(n13657), .A2(n13683), .ZN(n16224) );
  NAND2_X1 U17031 ( .A1(n16224), .A2(n15027), .ZN(n13658) );
  OAI211_X1 U17032 ( .C1(n15027), .C2(n13660), .A(n13659), .B(n13658), .ZN(
        P2_U2877) );
  MUX2_X1 U17033 ( .A(n14176), .B(n9581), .S(P1_EBX_REG_5__SCAN_IN), .Z(n13664) );
  NAND2_X1 U17034 ( .A1(n9874), .A2(n13381), .ZN(n14164) );
  NAND2_X1 U17035 ( .A1(n13381), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13662) );
  AND2_X1 U17036 ( .A1(n14164), .A2(n13662), .ZN(n13663) );
  NAND2_X1 U17037 ( .A1(n13664), .A2(n13663), .ZN(n13665) );
  AND2_X2 U17038 ( .A1(n13666), .A2(n13665), .ZN(n16137) );
  NOR2_X1 U17039 ( .A1(n13666), .A2(n13665), .ZN(n13667) );
  OR2_X1 U17040 ( .A1(n16137), .A2(n13667), .ZN(n19956) );
  INV_X1 U17041 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n19961) );
  OAI222_X1 U17042 ( .A1(n19956), .A2(n14457), .B1(n19994), .B2(n19961), .C1(
        n19959), .C2(n14455), .ZN(P1_U2867) );
  NOR2_X1 U17043 ( .A1(n19235), .A2(n19446), .ZN(n19651) );
  NAND2_X1 U17044 ( .A1(n19651), .A2(n19800), .ZN(n13668) );
  NAND2_X1 U17045 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19819), .ZN(
        n19497) );
  OR2_X1 U17046 ( .A1(n19828), .A2(n19497), .ZN(n13677) );
  NAND2_X1 U17047 ( .A1(n13668), .A2(n13677), .ZN(n13673) );
  NAND2_X1 U17048 ( .A1(n10411), .A2(n10900), .ZN(n13671) );
  INV_X1 U17049 ( .A(n19497), .ZN(n13669) );
  AND2_X1 U17050 ( .A1(n19388), .A2(n13669), .ZN(n19539) );
  NOR2_X1 U17051 ( .A1(n19539), .A2(n19802), .ZN(n13670) );
  AOI21_X1 U17052 ( .B1(n13671), .B2(n13670), .A(n19421), .ZN(n13672) );
  NAND2_X1 U17053 ( .A1(n13673), .A2(n13672), .ZN(n19542) );
  INV_X1 U17054 ( .A(n19542), .ZN(n19527) );
  INV_X1 U17055 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13681) );
  AOI22_X1 U17056 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19222), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19221), .ZN(n19565) );
  INV_X1 U17057 ( .A(n19579), .ZN(n19551) );
  AOI22_X1 U17058 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19222), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19221), .ZN(n19673) );
  INV_X1 U17059 ( .A(n19673), .ZN(n19562) );
  AOI22_X1 U17060 ( .A1(n19541), .A2(n19670), .B1(n19551), .B2(n19562), .ZN(
        n13680) );
  OAI21_X1 U17061 ( .B1(n10411), .B2(n19539), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13676) );
  OAI21_X1 U17062 ( .B1(n13677), .B2(n19609), .A(n13676), .ZN(n19540) );
  NOR2_X2 U17063 ( .A1(n13678), .A2(n19421), .ZN(n19669) );
  NAND2_X1 U17064 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19656), .ZN(n19205) );
  AND2_X1 U17065 ( .A1(n10718), .A2(n19223), .ZN(n19668) );
  AOI22_X1 U17066 ( .A1(n19540), .A2(n19669), .B1(n19539), .B2(n19668), .ZN(
        n13679) );
  OAI211_X1 U17067 ( .C1(n19527), .C2(n13681), .A(n13680), .B(n13679), .ZN(
        P2_U3138) );
  INV_X1 U17068 ( .A(n13682), .ZN(n13713) );
  XNOR2_X1 U17069 ( .A(n13714), .B(n13713), .ZN(n13688) );
  NAND2_X1 U17070 ( .A1(n13684), .A2(n13683), .ZN(n13686) );
  INV_X1 U17071 ( .A(n13707), .ZN(n13685) );
  INV_X1 U17072 ( .A(n16219), .ZN(n18945) );
  MUX2_X1 U17073 ( .A(n18944), .B(n18945), .S(n15027), .Z(n13687) );
  OAI21_X1 U17074 ( .B1(n13688), .B2(n15030), .A(n13687), .ZN(P2_U2876) );
  XOR2_X1 U17075 ( .A(n13690), .B(n13689), .Z(n20072) );
  NAND2_X1 U17076 ( .A1(n19984), .A2(n16031), .ZN(n13692) );
  INV_X1 U17077 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20840) );
  NOR2_X1 U17078 ( .A1(n16041), .A2(n20840), .ZN(n20065) );
  AOI21_X1 U17079 ( .B1(n20058), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20065), .ZN(n13691) );
  OAI211_X1 U17080 ( .C1(n16034), .C2(n19987), .A(n13692), .B(n13691), .ZN(
        n13693) );
  AOI21_X1 U17081 ( .B1(n20072), .B2(n20060), .A(n13693), .ZN(n13694) );
  INV_X1 U17082 ( .A(n13694), .ZN(P1_U2995) );
  NAND3_X1 U17083 ( .A1(n19828), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19547) );
  INV_X1 U17084 ( .A(n19547), .ZN(n13700) );
  AOI21_X1 U17085 ( .B1(n19651), .B2(n19352), .A(n13700), .ZN(n13699) );
  NOR2_X1 U17086 ( .A1(n19837), .A2(n19547), .ZN(n19608) );
  INV_X1 U17087 ( .A(n19608), .ZN(n13696) );
  NAND2_X1 U17088 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13696), .ZN(n13695) );
  NOR2_X1 U17089 ( .A1(n10359), .A2(n13695), .ZN(n13702) );
  NAND2_X1 U17090 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n13696), .ZN(n13697) );
  NAND2_X1 U17091 ( .A1(n19656), .A2(n13697), .ZN(n13698) );
  INV_X1 U17092 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13706) );
  NOR2_X2 U17093 ( .A1(n19604), .A2(n19353), .ZN(n19599) );
  AOI22_X1 U17094 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19221), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19222), .ZN(n19620) );
  AOI22_X1 U17095 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19222), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19221), .ZN(n19661) );
  AOI22_X1 U17096 ( .A1(n19599), .A2(n19658), .B1(n19633), .B2(n19606), .ZN(
        n13705) );
  AOI21_X1 U17097 ( .B1(n10900), .B2(n13700), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13701) );
  NOR2_X1 U17098 ( .A1(n13702), .A2(n13701), .ZN(n19597) );
  NOR2_X2 U17099 ( .A1(n13703), .A2(n19421), .ZN(n19650) );
  AND2_X1 U17100 ( .A1(n19852), .A2(n19223), .ZN(n19649) );
  AOI22_X1 U17101 ( .A1(n19597), .A2(n19650), .B1(n19649), .B2(n19608), .ZN(
        n13704) );
  OAI211_X1 U17102 ( .C1(n19602), .C2(n13706), .A(n13705), .B(n13704), .ZN(
        P2_U3152) );
  OR2_X1 U17103 ( .A1(n13708), .A2(n13707), .ZN(n13709) );
  AND2_X1 U17104 ( .A1(n13709), .A2(n13753), .ZN(n18934) );
  INV_X1 U17105 ( .A(n18934), .ZN(n15437) );
  AND2_X1 U17106 ( .A1(n13711), .A2(n13710), .ZN(n13752) );
  INV_X1 U17107 ( .A(n13752), .ZN(n13716) );
  OAI21_X1 U17108 ( .B1(n13714), .B2(n13713), .A(n13712), .ZN(n13715) );
  NAND3_X1 U17109 ( .A1(n13716), .A2(n15018), .A3(n13715), .ZN(n13718) );
  NAND2_X1 U17110 ( .A1(n15022), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13717) );
  OAI211_X1 U17111 ( .C1(n15437), .C2(n15022), .A(n13718), .B(n13717), .ZN(
        P2_U2875) );
  NAND2_X1 U17112 ( .A1(n13721), .A2(n13722), .ZN(n13723) );
  AND2_X1 U17113 ( .A1(n13720), .A2(n13723), .ZN(n19937) );
  INV_X1 U17114 ( .A(n19937), .ZN(n13749) );
  MUX2_X1 U17115 ( .A(n14176), .B(n9581), .S(P1_EBX_REG_7__SCAN_IN), .Z(n13726) );
  NAND2_X1 U17116 ( .A1(n13381), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13724) );
  AND2_X1 U17117 ( .A1(n14164), .A2(n13724), .ZN(n13725) );
  INV_X1 U17118 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n19993) );
  NAND2_X1 U17119 ( .A1(n14179), .A2(n19993), .ZN(n13729) );
  NAND2_X1 U17120 ( .A1(n14290), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13727) );
  OAI211_X1 U17121 ( .C1(n13381), .C2(P1_EBX_REG_6__SCAN_IN), .A(n13727), .B(
        n9581), .ZN(n13728) );
  AND2_X1 U17122 ( .A1(n13729), .A2(n13728), .ZN(n16136) );
  AOI21_X1 U17123 ( .B1(n13730), .B2(n16135), .A(n9881), .ZN(n19931) );
  AOI22_X1 U17124 ( .A1(n19989), .A2(n19931), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n14438), .ZN(n13731) );
  OAI21_X1 U17125 ( .B1(n13749), .B2(n14455), .A(n13731), .ZN(P1_U2865) );
  NOR3_X2 U17126 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19837), .A3(
        n19497), .ZN(n19498) );
  INV_X1 U17127 ( .A(n19498), .ZN(n13732) );
  OAI21_X1 U17128 ( .B1(n13733), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n13732), 
        .ZN(n13735) );
  NAND2_X1 U17129 ( .A1(n19651), .A2(n19232), .ZN(n13739) );
  OR2_X1 U17130 ( .A1(n19497), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13737) );
  NAND2_X1 U17131 ( .A1(n13739), .A2(n13737), .ZN(n13734) );
  MUX2_X1 U17132 ( .A(n13735), .B(n13734), .S(n19802), .Z(n13736) );
  NAND2_X1 U17133 ( .A1(n13736), .A2(n19656), .ZN(n19491) );
  INV_X1 U17134 ( .A(n19491), .ZN(n13747) );
  INV_X1 U17135 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13746) );
  INV_X1 U17136 ( .A(n13737), .ZN(n13738) );
  NAND3_X1 U17137 ( .A1(n13739), .A2(n19802), .A3(n13738), .ZN(n13742) );
  OAI21_X1 U17138 ( .B1(n13740), .B2(n19498), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13741) );
  NAND2_X1 U17139 ( .A1(n13742), .A2(n13741), .ZN(n19490) );
  AOI22_X1 U17140 ( .A1(n19606), .A2(n19499), .B1(n19649), .B2(n19498), .ZN(
        n13743) );
  OAI21_X1 U17141 ( .B1(n19482), .B2(n19620), .A(n13743), .ZN(n13744) );
  AOI21_X1 U17142 ( .B1(n19650), .B2(n19490), .A(n13744), .ZN(n13745) );
  OAI21_X1 U17143 ( .B1(n13747), .B2(n13746), .A(n13745), .ZN(P2_U3120) );
  OAI222_X1 U17144 ( .A1(n14544), .A2(n13749), .B1(n14542), .B2(n20137), .C1(
        n13748), .C2(n14540), .ZN(P1_U2897) );
  OAI211_X1 U17145 ( .C1(n13752), .C2(n13751), .A(n13750), .B(n15018), .ZN(
        n13756) );
  AOI21_X1 U17146 ( .B1(n13754), .B2(n13753), .A(n13833), .ZN(n18924) );
  NAND2_X1 U17147 ( .A1(n15027), .A2(n18924), .ZN(n13755) );
  OAI211_X1 U17148 ( .C1(n15027), .C2(n10805), .A(n13756), .B(n13755), .ZN(
        P2_U2874) );
  XOR2_X1 U17149 ( .A(n13648), .B(n13757), .Z(n19991) );
  INV_X1 U17150 ( .A(n19991), .ZN(n19947) );
  OAI222_X1 U17151 ( .A1(n14544), .A2(n19947), .B1(n14540), .B2(n11757), .C1(
        n14542), .C2(n20128), .ZN(P1_U2898) );
  AOI21_X1 U17152 ( .B1(n13759), .B2(n13720), .A(n13758), .ZN(n13760) );
  INV_X1 U17153 ( .A(n13760), .ZN(n19920) );
  INV_X1 U17154 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13761) );
  NAND2_X1 U17155 ( .A1(n14179), .A2(n13761), .ZN(n13764) );
  NAND2_X1 U17156 ( .A1(n14290), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13762) );
  OAI211_X1 U17157 ( .C1(n13381), .C2(P1_EBX_REG_8__SCAN_IN), .A(n13762), .B(
        n9581), .ZN(n13763) );
  NAND2_X1 U17158 ( .A1(n13764), .A2(n13763), .ZN(n13765) );
  NAND2_X1 U17159 ( .A1(n13766), .A2(n13765), .ZN(n13767) );
  AND2_X1 U17160 ( .A1(n13903), .A2(n13767), .ZN(n19924) );
  AOI22_X1 U17161 ( .A1(n19989), .A2(n19924), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n14438), .ZN(n13768) );
  OAI21_X1 U17162 ( .B1(n19920), .B2(n14455), .A(n13768), .ZN(P1_U2864) );
  OR2_X1 U17163 ( .A1(n20080), .A2(n13769), .ZN(n13771) );
  NAND2_X1 U17164 ( .A1(n20080), .A2(DATAI_8_), .ZN(n13770) );
  NAND2_X1 U17165 ( .A1(n13771), .A2(n13770), .ZN(n20025) );
  AOI22_X1 U17166 ( .A1(n14095), .A2(n20025), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n15957), .ZN(n13772) );
  OAI21_X1 U17167 ( .B1(n19920), .B2(n14544), .A(n13772), .ZN(P1_U2896) );
  XOR2_X1 U17168 ( .A(n13774), .B(n13773), .Z(n16036) );
  NOR2_X1 U17169 ( .A1(n11573), .A2(n13775), .ZN(n13777) );
  NAND2_X1 U17170 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13777), .ZN(
        n14032) );
  NOR2_X1 U17171 ( .A1(n13776), .A2(n14032), .ZN(n14673) );
  OAI21_X1 U17172 ( .B1(n14810), .B2(n14673), .A(n14788), .ZN(n14804) );
  INV_X1 U17173 ( .A(n14033), .ZN(n13778) );
  INV_X1 U17174 ( .A(n13777), .ZN(n20073) );
  OAI21_X1 U17175 ( .B1(n13778), .B2(n20073), .A(n14805), .ZN(n13779) );
  INV_X1 U17176 ( .A(n13779), .ZN(n13780) );
  NOR2_X1 U17177 ( .A1(n14804), .A2(n13780), .ZN(n16119) );
  INV_X1 U17178 ( .A(n19956), .ZN(n13783) );
  INV_X1 U17179 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n13781) );
  OR2_X1 U17180 ( .A1(n16041), .A2(n13781), .ZN(n16037) );
  INV_X1 U17181 ( .A(n16037), .ZN(n13782) );
  AOI21_X1 U17182 ( .B1(n20067), .B2(n13783), .A(n13782), .ZN(n13785) );
  NOR2_X1 U17183 ( .A1(n20073), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16118) );
  NAND2_X1 U17184 ( .A1(n20074), .A2(n16118), .ZN(n13784) );
  OAI211_X1 U17185 ( .C1(n16119), .C2(n11582), .A(n13785), .B(n13784), .ZN(
        n13786) );
  AOI21_X1 U17186 ( .B1(n16036), .B2(n20071), .A(n13786), .ZN(n13787) );
  INV_X1 U17187 ( .A(n13787), .ZN(P1_U3026) );
  NAND2_X1 U17188 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20763), .ZN(n15787) );
  NAND2_X1 U17189 ( .A1(n12142), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13788) );
  MUX2_X1 U17190 ( .A(n15787), .B(n13788), .S(n20676), .Z(n13789) );
  INV_X1 U17191 ( .A(n13789), .ZN(n13790) );
  NOR2_X1 U17192 ( .A1(n13790), .A2(n16139), .ZN(n13791) );
  NOR2_X1 U17193 ( .A1(n13796), .A2(n13793), .ZN(n13794) );
  INV_X1 U17194 ( .A(n19983), .ZN(n14376) );
  NOR2_X1 U17195 ( .A1(n13795), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13799) );
  NAND2_X1 U17196 ( .A1(n19914), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n19979) );
  NOR2_X1 U17197 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n19979), .ZN(n13816) );
  INV_X1 U17198 ( .A(n13328), .ZN(n14828) );
  INV_X1 U17199 ( .A(n13796), .ZN(n13798) );
  NAND2_X1 U17200 ( .A1(n13798), .A2(n13797), .ZN(n19972) );
  AND2_X1 U17201 ( .A1(n20102), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13802) );
  NOR2_X1 U17202 ( .A1(n13799), .A2(n13802), .ZN(n13800) );
  NAND2_X1 U17203 ( .A1(n20691), .A2(n20777), .ZN(n15780) );
  NAND2_X1 U17204 ( .A1(n13802), .A2(n15780), .ZN(n13803) );
  AOI22_X1 U17205 ( .A1(n19974), .A2(P1_EBX_REG_3__SCAN_IN), .B1(n19942), .B2(
        n13805), .ZN(n13814) );
  INV_X1 U17206 ( .A(n13806), .ZN(n13812) );
  NOR2_X1 U17207 ( .A1(n13807), .A2(n20677), .ZN(n13808) );
  NOR2_X1 U17208 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n19979), .ZN(n14371) );
  OAI21_X1 U17209 ( .B1(n19901), .B2(P1_REIP_REG_1__SCAN_IN), .A(n19898), .ZN(
        n14373) );
  OAI21_X1 U17210 ( .B1(n14371), .B2(n14373), .A(P1_REIP_REG_3__SCAN_IN), .ZN(
        n13809) );
  OAI21_X1 U17211 ( .B1(n15945), .B2(n13810), .A(n13809), .ZN(n13811) );
  AOI21_X1 U17212 ( .B1(n13812), .B2(n19909), .A(n13811), .ZN(n13813) );
  OAI211_X1 U17213 ( .C1(n14828), .C2(n19972), .A(n13814), .B(n13813), .ZN(
        n13815) );
  AOI21_X1 U17214 ( .B1(n13816), .B2(P1_REIP_REG_2__SCAN_IN), .A(n13815), .ZN(
        n13817) );
  OAI21_X1 U17215 ( .B1(n13818), .B2(n14376), .A(n13817), .ZN(P1_U2837) );
  INV_X1 U17216 ( .A(n19039), .ZN(n19012) );
  NAND2_X1 U17217 ( .A1(n13017), .A2(n13819), .ZN(n13820) );
  XNOR2_X1 U17218 ( .A(n16252), .B(n13820), .ZN(n13821) );
  NAND2_X1 U17219 ( .A1(n13821), .A2(n19002), .ZN(n13832) );
  INV_X1 U17220 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19744) );
  OAI22_X1 U17221 ( .A1(n10253), .A2(n19009), .B1(n19744), .B2(n18993), .ZN(
        n13822) );
  AOI21_X1 U17222 ( .B1(n19041), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13822), .ZN(n13823) );
  OAI21_X1 U17223 ( .B1(n19008), .B2(n13824), .A(n13823), .ZN(n13830) );
  OR2_X1 U17224 ( .A1(n13826), .A2(n13825), .ZN(n13828) );
  NAND2_X1 U17225 ( .A1(n13828), .A2(n13827), .ZN(n19088) );
  NOR2_X1 U17226 ( .A1(n19088), .A2(n19006), .ZN(n13829) );
  AOI211_X1 U17227 ( .C1(n19022), .C2(n15599), .A(n13830), .B(n13829), .ZN(
        n13831) );
  OAI211_X1 U17228 ( .C1(n19012), .C2(n19235), .A(n13832), .B(n13831), .ZN(
        P2_U2852) );
  OR2_X1 U17229 ( .A1(n13834), .A2(n13833), .ZN(n13835) );
  AND2_X1 U17230 ( .A1(n13958), .A2(n13835), .ZN(n16282) );
  INV_X1 U17231 ( .A(n16282), .ZN(n13980) );
  INV_X1 U17232 ( .A(n13750), .ZN(n13838) );
  OAI211_X1 U17233 ( .C1(n13838), .C2(n12280), .A(n15018), .B(n13837), .ZN(
        n13840) );
  NAND2_X1 U17234 ( .A1(n15022), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13839) );
  OAI211_X1 U17235 ( .C1(n13980), .C2(n15022), .A(n13840), .B(n13839), .ZN(
        P2_U2873) );
  NAND2_X1 U17236 ( .A1(n19901), .A2(n19898), .ZN(n19955) );
  INV_X1 U17237 ( .A(n19955), .ZN(n13849) );
  AOI22_X1 U17238 ( .A1(n19974), .A2(P1_EBX_REG_0__SCAN_IN), .B1(n19923), .B2(
        n13841), .ZN(n13847) );
  INV_X1 U17239 ( .A(n20064), .ZN(n13845) );
  OAI21_X1 U17240 ( .B1(n19969), .B2(n19909), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13842) );
  OAI21_X1 U17241 ( .B1(n19972), .B2(n13843), .A(n13842), .ZN(n13844) );
  AOI21_X1 U17242 ( .B1(n13845), .B2(n19983), .A(n13844), .ZN(n13846) );
  OAI211_X1 U17243 ( .C1(n13849), .C2(n13848), .A(n13847), .B(n13846), .ZN(
        P1_U2840) );
  NOR2_X1 U17244 ( .A1(n13016), .A2(n13850), .ZN(n13851) );
  XNOR2_X1 U17245 ( .A(n13851), .B(n16242), .ZN(n13852) );
  NAND2_X1 U17246 ( .A1(n13852), .A2(n19002), .ZN(n13859) );
  AOI21_X1 U17247 ( .B1(n13853), .B2(n15518), .A(n15481), .ZN(n19079) );
  AOI22_X1 U17248 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19041), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19031), .ZN(n13854) );
  OAI211_X1 U17249 ( .C1(n19009), .C2(n13855), .A(n13854), .B(n16264), .ZN(
        n13857) );
  NOR2_X1 U17250 ( .A1(n16235), .A2(n19011), .ZN(n13856) );
  AOI211_X1 U17251 ( .C1(n19079), .C2(n19027), .A(n13857), .B(n13856), .ZN(
        n13858) );
  OAI211_X1 U17252 ( .C1(n19008), .C2(n13860), .A(n13859), .B(n13858), .ZN(
        P2_U2847) );
  NOR2_X1 U17253 ( .A1(n13016), .A2(n13861), .ZN(n13912) );
  XNOR2_X1 U17254 ( .A(n13912), .B(n19171), .ZN(n13862) );
  NAND2_X1 U17255 ( .A1(n13862), .A2(n19002), .ZN(n13869) );
  OAI22_X1 U17256 ( .A1(n10240), .A2(n19009), .B1(n19742), .B2(n18993), .ZN(
        n13863) );
  AOI21_X1 U17257 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19041), .A(
        n13863), .ZN(n13864) );
  OAI21_X1 U17258 ( .B1(n19008), .B2(n13865), .A(n13864), .ZN(n13867) );
  NOR2_X1 U17259 ( .A1(n19812), .A2(n19006), .ZN(n13866) );
  AOI211_X1 U17260 ( .C1(n19022), .C2(n14011), .A(n13867), .B(n13866), .ZN(
        n13868) );
  OAI211_X1 U17261 ( .C1(n19012), .C2(n19810), .A(n13869), .B(n13868), .ZN(
        P2_U2853) );
  NOR2_X1 U17262 ( .A1(n19972), .A2(n20372), .ZN(n13873) );
  INV_X1 U17263 ( .A(n19898), .ZN(n15929) );
  AOI22_X1 U17264 ( .A1(n19969), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n15929), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13871) );
  OAI21_X1 U17265 ( .B1(n19986), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13871), .ZN(n13872) );
  AOI211_X1 U17266 ( .C1(n13874), .C2(n19942), .A(n13873), .B(n13872), .ZN(
        n13876) );
  AOI22_X1 U17267 ( .A1(n19914), .A2(n20749), .B1(n19974), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13875) );
  OAI211_X1 U17268 ( .C1(n14376), .C2(n13877), .A(n13876), .B(n13875), .ZN(
        P1_U2839) );
  NAND2_X1 U17269 ( .A1(n13879), .A2(n13878), .ZN(n13881) );
  XNOR2_X1 U17270 ( .A(n13881), .B(n13880), .ZN(n16256) );
  INV_X1 U17271 ( .A(n16256), .ZN(n13891) );
  INV_X1 U17272 ( .A(n19088), .ZN(n19804) );
  OAI22_X1 U17273 ( .A1(n10287), .A2(n16295), .B1(n19744), .B2(n16264), .ZN(
        n13886) );
  INV_X1 U17274 ( .A(n13882), .ZN(n13883) );
  MUX2_X1 U17275 ( .A(n13884), .B(n13883), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n13885) );
  AOI211_X1 U17276 ( .C1(n16280), .C2(n19804), .A(n13886), .B(n13885), .ZN(
        n13890) );
  NAND3_X1 U17277 ( .A1(n16253), .A2(n16270), .A3(n13888), .ZN(n13889) );
  OAI211_X1 U17278 ( .C1(n13891), .C2(n16274), .A(n13890), .B(n13889), .ZN(
        P2_U3043) );
  NOR2_X1 U17279 ( .A1(n13758), .A2(n13893), .ZN(n13894) );
  OR2_X1 U17280 ( .A1(n13892), .A2(n13894), .ZN(n19907) );
  OR2_X1 U17281 ( .A1(n20080), .A2(n13895), .ZN(n13897) );
  NAND2_X1 U17282 ( .A1(n20080), .A2(DATAI_9_), .ZN(n13896) );
  NAND2_X1 U17283 ( .A1(n13897), .A2(n13896), .ZN(n20027) );
  AOI22_X1 U17284 ( .A1(n14095), .A2(n20027), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15957), .ZN(n13898) );
  OAI21_X1 U17285 ( .B1(n19907), .B2(n14544), .A(n13898), .ZN(P1_U2895) );
  INV_X1 U17286 ( .A(n13903), .ZN(n13905) );
  MUX2_X1 U17287 ( .A(n14176), .B(n9581), .S(P1_EBX_REG_9__SCAN_IN), .Z(n13901) );
  NAND2_X1 U17288 ( .A1(n13381), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13899) );
  AND2_X1 U17289 ( .A1(n14164), .A2(n13899), .ZN(n13900) );
  NAND2_X1 U17290 ( .A1(n13901), .A2(n13900), .ZN(n13904) );
  INV_X1 U17291 ( .A(n13904), .ZN(n13902) );
  INV_X1 U17292 ( .A(n13925), .ZN(n13927) );
  OAI21_X1 U17293 ( .B1(n13905), .B2(n13904), .A(n13927), .ZN(n19903) );
  INV_X1 U17294 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n13906) );
  OAI222_X1 U17295 ( .A1(n19903), .A2(n14457), .B1(n13906), .B2(n19994), .C1(
        n19907), .C2(n14455), .ZN(P1_U2863) );
  NOR2_X1 U17296 ( .A1(n19008), .A2(n15244), .ZN(n13908) );
  OAI22_X1 U17297 ( .A1(n19009), .A2(n10214), .B1(n18991), .B2(n15241), .ZN(
        n13907) );
  AOI211_X1 U17298 ( .C1(n19031), .C2(P2_REIP_REG_1__SCAN_IN), .A(n13908), .B(
        n13907), .ZN(n13910) );
  NAND2_X1 U17299 ( .A1(n19826), .A2(n19027), .ZN(n13909) );
  OAI211_X1 U17300 ( .C1(n13911), .C2(n19011), .A(n13910), .B(n13909), .ZN(
        n13915) );
  NAND2_X1 U17301 ( .A1(n13016), .A2(n19002), .ZN(n18881) );
  OAI21_X1 U17302 ( .B1(n13931), .B2(n13913), .A(n13912), .ZN(n13930) );
  OAI22_X1 U17303 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18881), .B1(
        n13930), .B2(n19720), .ZN(n13914) );
  AOI211_X1 U17304 ( .C1(n19039), .C2(n19822), .A(n13915), .B(n13914), .ZN(
        n13916) );
  INV_X1 U17305 ( .A(n13916), .ZN(P2_U2854) );
  OAI21_X1 U17306 ( .B1(n13892), .B2(n13918), .A(n13917), .ZN(n15946) );
  OR2_X1 U17307 ( .A1(n20080), .A2(n16445), .ZN(n13920) );
  NAND2_X1 U17308 ( .A1(n20080), .A2(DATAI_10_), .ZN(n13919) );
  NAND2_X1 U17309 ( .A1(n13920), .A2(n13919), .ZN(n20029) );
  AOI22_X1 U17310 ( .A1(n14095), .A2(n20029), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15957), .ZN(n13921) );
  OAI21_X1 U17311 ( .B1(n15946), .B2(n14544), .A(n13921), .ZN(P1_U2894) );
  MUX2_X1 U17312 ( .A(n14179), .B(n14276), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n13923) );
  NOR2_X1 U17313 ( .A1(n14277), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13922) );
  NOR2_X1 U17314 ( .A1(n13923), .A2(n13922), .ZN(n13924) );
  INV_X1 U17315 ( .A(n13924), .ZN(n13928) );
  INV_X1 U17316 ( .A(n15931), .ZN(n13926) );
  AOI21_X1 U17317 ( .B1(n13928), .B2(n13927), .A(n13926), .ZN(n16109) );
  AOI22_X1 U17318 ( .A1(n19989), .A2(n16109), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14438), .ZN(n13929) );
  OAI21_X1 U17319 ( .B1(n15946), .B2(n14455), .A(n13929), .ZN(P1_U2862) );
  OAI21_X1 U17320 ( .B1(n13017), .B2(n15248), .A(n13930), .ZN(n14014) );
  INV_X1 U17321 ( .A(n14014), .ZN(n13941) );
  INV_X1 U17322 ( .A(n13931), .ZN(n19038) );
  AOI22_X1 U17323 ( .A1(n13016), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19038), .B2(n13017), .ZN(n15576) );
  NOR2_X1 U17324 ( .A1(n15576), .A2(n19712), .ZN(n14013) );
  INV_X1 U17325 ( .A(n13932), .ZN(n15598) );
  INV_X1 U17326 ( .A(n13933), .ZN(n13935) );
  NOR2_X1 U17327 ( .A1(n13935), .A2(n13934), .ZN(n15578) );
  NOR2_X1 U17328 ( .A1(n13937), .A2(n13936), .ZN(n13938) );
  INV_X1 U17329 ( .A(n10868), .ZN(n15579) );
  OAI22_X1 U17330 ( .A1(n15578), .A2(n13938), .B1(n15579), .B2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13939) );
  AOI21_X1 U17331 ( .B1(n15568), .B2(n15598), .A(n13939), .ZN(n16325) );
  OAI22_X1 U17332 ( .A1(n19183), .A2(n15601), .B1(n15600), .B2(n16325), .ZN(
        n13940) );
  AOI21_X1 U17333 ( .B1(n13941), .B2(n14013), .A(n13940), .ZN(n13944) );
  NAND2_X1 U17334 ( .A1(n15602), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13943) );
  OAI21_X1 U17335 ( .B1(n13944), .B2(n15602), .A(n13943), .ZN(P2_U3600) );
  XNOR2_X1 U17336 ( .A(n13945), .B(n13948), .ZN(n19156) );
  INV_X1 U17337 ( .A(n19156), .ZN(n13955) );
  XNOR2_X1 U17338 ( .A(n13946), .B(n9674), .ZN(n19157) );
  NAND2_X1 U17339 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19155), .ZN(n13947) );
  OAI221_X1 U17340 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15557), .C1(
        n13948), .C2(n15559), .A(n13947), .ZN(n13953) );
  NAND2_X1 U17341 ( .A1(n13949), .A2(n13827), .ZN(n13951) );
  INV_X1 U17342 ( .A(n15556), .ZN(n13950) );
  AND2_X1 U17343 ( .A1(n13951), .A2(n13950), .ZN(n19097) );
  INV_X1 U17344 ( .A(n19097), .ZN(n19089) );
  OAI22_X1 U17345 ( .A1(n19160), .A2(n16295), .B1(n16294), .B2(n19089), .ZN(
        n13952) );
  AOI211_X1 U17346 ( .C1(n19157), .C2(n16301), .A(n13953), .B(n13952), .ZN(
        n13954) );
  OAI21_X1 U17347 ( .B1(n13955), .B2(n16305), .A(n13954), .ZN(P2_U3042) );
  XNOR2_X1 U17348 ( .A(n13837), .B(n13956), .ZN(n13961) );
  NAND2_X1 U17349 ( .A1(n13958), .A2(n13957), .ZN(n13959) );
  AND2_X1 U17350 ( .A1(n13998), .A2(n13959), .ZN(n16269) );
  MUX2_X1 U17351 ( .A(n10814), .B(n18912), .S(n15027), .Z(n13960) );
  OAI21_X1 U17352 ( .B1(n13961), .B2(n15030), .A(n13960), .ZN(P2_U2872) );
  INV_X1 U17353 ( .A(n13962), .ZN(n13964) );
  OAI21_X1 U17354 ( .B1(n13964), .B2(n9688), .A(n13963), .ZN(n15031) );
  OAI21_X1 U17355 ( .B1(n15412), .B2(n13966), .A(n13965), .ZN(n15405) );
  INV_X1 U17356 ( .A(n15405), .ZN(n18885) );
  NAND2_X1 U17357 ( .A1(n19051), .A2(BUF1_REG_17__SCAN_IN), .ZN(n13970) );
  NAND2_X1 U17358 ( .A1(n19052), .A2(BUF2_REG_17__SCAN_IN), .ZN(n13969) );
  AOI22_X1 U17359 ( .A1(n19050), .A2(n13967), .B1(n19110), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n13968) );
  NAND3_X1 U17360 ( .A1(n13970), .A2(n13969), .A3(n13968), .ZN(n13971) );
  AOI21_X1 U17361 ( .B1(n18885), .B2(n19111), .A(n13971), .ZN(n13972) );
  OAI21_X1 U17362 ( .B1(n19115), .B2(n15031), .A(n13972), .ZN(P2_U2902) );
  NOR2_X1 U17363 ( .A1(n13016), .A2(n13973), .ZN(n13974) );
  XNOR2_X1 U17364 ( .A(n13974), .B(n16208), .ZN(n13975) );
  NAND2_X1 U17365 ( .A1(n13975), .A2(n19002), .ZN(n13986) );
  AND2_X1 U17366 ( .A1(n13977), .A2(n13976), .ZN(n16263) );
  AOI21_X1 U17367 ( .B1(n13978), .B2(n15423), .A(n16263), .ZN(n19062) );
  OAI22_X1 U17368 ( .A1(n19011), .A2(n13980), .B1(n19009), .B2(n13979), .ZN(
        n13984) );
  INV_X1 U17369 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19763) );
  AOI22_X1 U17370 ( .A1(n13981), .A2(n19030), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19041), .ZN(n13982) );
  OAI211_X1 U17371 ( .C1(n19763), .C2(n18993), .A(n13982), .B(n18992), .ZN(
        n13983) );
  AOI211_X1 U17372 ( .C1(n19027), .C2(n19062), .A(n13984), .B(n13983), .ZN(
        n13985) );
  NAND2_X1 U17373 ( .A1(n13986), .A2(n13985), .ZN(P2_U2841) );
  XOR2_X1 U17374 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n13987), .Z(
        n13988) );
  XNOR2_X1 U17375 ( .A(n13989), .B(n13988), .ZN(n16125) );
  NAND2_X1 U17376 ( .A1(n16125), .A2(n20060), .ZN(n13993) );
  INV_X1 U17377 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n13990) );
  NOR2_X1 U17378 ( .A1(n16041), .A2(n13990), .ZN(n16122) );
  NOR2_X1 U17379 ( .A1(n16034), .A2(n19917), .ZN(n13991) );
  AOI211_X1 U17380 ( .C1(n20058), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16122), .B(n13991), .ZN(n13992) );
  OAI211_X1 U17381 ( .C1(n20081), .C2(n19920), .A(n13993), .B(n13992), .ZN(
        P1_U2991) );
  OR2_X1 U17382 ( .A1(n13995), .A2(n13994), .ZN(n13996) );
  NAND2_X1 U17383 ( .A1(n13962), .A2(n13996), .ZN(n19053) );
  OR2_X1 U17384 ( .A1(n15027), .A2(n18899), .ZN(n14001) );
  NAND2_X1 U17385 ( .A1(n13998), .A2(n13997), .ZN(n13999) );
  AND2_X1 U17386 ( .A1(n15024), .A2(n13999), .ZN(n18901) );
  NAND2_X1 U17387 ( .A1(n15027), .A2(n18901), .ZN(n14000) );
  OAI211_X1 U17388 ( .C1(n19053), .C2(n15030), .A(n14001), .B(n14000), .ZN(
        P2_U2871) );
  OR2_X1 U17389 ( .A1(n14003), .A2(n14002), .ZN(n15588) );
  NOR2_X1 U17390 ( .A1(n15589), .A2(n10308), .ZN(n14006) );
  NOR2_X1 U17391 ( .A1(n14004), .A2(n10739), .ZN(n14005) );
  AOI22_X1 U17392 ( .A1(n15588), .A2(n14006), .B1(n14005), .B2(n10868), .ZN(
        n14009) );
  OR2_X1 U17393 ( .A1(n16311), .A2(n16309), .ZN(n15587) );
  INV_X1 U17394 ( .A(n14006), .ZN(n14007) );
  NAND2_X1 U17395 ( .A1(n15587), .A2(n14007), .ZN(n14008) );
  NAND2_X1 U17396 ( .A1(n14009), .A2(n14008), .ZN(n14010) );
  AOI21_X1 U17397 ( .B1(n14011), .B2(n15598), .A(n14010), .ZN(n16307) );
  OAI22_X1 U17398 ( .A1(n19810), .A2(n15601), .B1(n15600), .B2(n16307), .ZN(
        n14012) );
  AOI21_X1 U17399 ( .B1(n14014), .B2(n14013), .A(n14012), .ZN(n14015) );
  MUX2_X1 U17400 ( .A(n14015), .B(n10458), .S(n15602), .Z(n14016) );
  INV_X1 U17401 ( .A(n14016), .ZN(P2_U3599) );
  XNOR2_X1 U17402 ( .A(n14932), .B(n14017), .ZN(n18875) );
  AOI21_X1 U17403 ( .B1(n9686), .B2(n10029), .A(n15006), .ZN(n15014) );
  INV_X1 U17404 ( .A(n19051), .ZN(n14023) );
  INV_X1 U17405 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n14515) );
  INV_X1 U17406 ( .A(n19050), .ZN(n15065) );
  OAI22_X1 U17407 ( .A1(n15065), .A2(n19202), .B1(n19083), .B2(n14020), .ZN(
        n14021) );
  AOI21_X1 U17408 ( .B1(n19052), .B2(BUF2_REG_19__SCAN_IN), .A(n14021), .ZN(
        n14022) );
  OAI21_X1 U17409 ( .B1(n14023), .B2(n14515), .A(n14022), .ZN(n14024) );
  AOI21_X1 U17410 ( .B1(n15014), .B2(n19100), .A(n14024), .ZN(n14025) );
  OAI21_X1 U17411 ( .B1(n18875), .B2(n19054), .A(n14025), .ZN(P2_U2900) );
  MUX2_X1 U17412 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n11614), .S(
        n15965), .Z(n14027) );
  XOR2_X1 U17413 ( .A(n14027), .B(n14026), .Z(n14039) );
  INV_X1 U17414 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n14028) );
  OAI22_X1 U17415 ( .A1(n16039), .A2(n11806), .B1(n16041), .B2(n14028), .ZN(
        n14030) );
  NOR2_X1 U17416 ( .A1(n19907), .A2(n20081), .ZN(n14029) );
  AOI211_X1 U17417 ( .C1(n16007), .C2(n19908), .A(n14030), .B(n14029), .ZN(
        n14031) );
  OAI21_X1 U17418 ( .B1(n14039), .B2(n19879), .A(n14031), .ZN(P1_U2990) );
  NAND2_X1 U17419 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16123) );
  NOR2_X1 U17420 ( .A1(n16129), .A2(n16123), .ZN(n14671) );
  INV_X1 U17421 ( .A(n14032), .ZN(n14036) );
  NAND2_X1 U17422 ( .A1(n14033), .A2(n14036), .ZN(n14807) );
  AOI21_X1 U17423 ( .B1(n14805), .B2(n14807), .A(n14804), .ZN(n14034) );
  AND2_X1 U17424 ( .A1(n14695), .A2(n14788), .ZN(n14687) );
  AOI21_X1 U17425 ( .B1(n14671), .B2(n14034), .A(n14687), .ZN(n16110) );
  OAI22_X1 U17426 ( .A1(n16069), .A2(n19903), .B1(n14028), .B2(n16041), .ZN(
        n14035) );
  AOI21_X1 U17427 ( .B1(n16110), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n14035), .ZN(n14038) );
  NAND2_X1 U17428 ( .A1(n14036), .A2(n20074), .ZN(n16144) );
  NOR3_X1 U17429 ( .A1(n16129), .A2(n16123), .A3(n16144), .ZN(n16112) );
  NAND2_X1 U17430 ( .A1(n16112), .A2(n11614), .ZN(n14037) );
  OAI211_X1 U17431 ( .C1(n14039), .C2(n16070), .A(n14038), .B(n14037), .ZN(
        P1_U3022) );
  INV_X1 U17432 ( .A(n14040), .ZN(n14100) );
  OAI21_X1 U17433 ( .B1(n14048), .B2(n14041), .A(n14100), .ZN(n15915) );
  OR2_X1 U17434 ( .A1(n20080), .A2(n14042), .ZN(n14044) );
  NAND2_X1 U17435 ( .A1(n20080), .A2(DATAI_14_), .ZN(n14043) );
  NAND2_X1 U17436 ( .A1(n14044), .A2(n14043), .ZN(n20037) );
  AOI22_X1 U17437 ( .A1(n14095), .A2(n20037), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15957), .ZN(n14045) );
  OAI21_X1 U17438 ( .B1(n15915), .B2(n14544), .A(n14045), .ZN(P1_U2890) );
  OAI21_X1 U17439 ( .B1(n11818), .B2(n11817), .A(n14047), .ZN(n14081) );
  OAI21_X1 U17440 ( .B1(n14081), .B2(n14082), .A(n14047), .ZN(n14088) );
  INV_X1 U17441 ( .A(n14048), .ZN(n14049) );
  OR2_X1 U17442 ( .A1(n20080), .A2(n14051), .ZN(n14053) );
  NAND2_X1 U17443 ( .A1(n20080), .A2(DATAI_13_), .ZN(n14052) );
  NAND2_X1 U17444 ( .A1(n14053), .A2(n14052), .ZN(n20035) );
  AOI22_X1 U17445 ( .A1(n14095), .A2(n20035), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15957), .ZN(n14054) );
  OAI21_X1 U17446 ( .B1(n14663), .B2(n14544), .A(n14054), .ZN(P1_U2891) );
  INV_X1 U17447 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15954) );
  NAND2_X1 U17448 ( .A1(n14179), .A2(n15954), .ZN(n14057) );
  NAND2_X1 U17449 ( .A1(n14290), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14055) );
  OAI211_X1 U17450 ( .C1(n13381), .C2(P1_EBX_REG_12__SCAN_IN), .A(n14055), .B(
        n9581), .ZN(n14056) );
  AND2_X1 U17451 ( .A1(n14057), .A2(n14056), .ZN(n14797) );
  INV_X1 U17452 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15956) );
  NAND2_X1 U17453 ( .A1(n14273), .A2(n15956), .ZN(n14061) );
  INV_X1 U17454 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14058) );
  NAND2_X1 U17455 ( .A1(n9581), .A2(n14058), .ZN(n14059) );
  OAI211_X1 U17456 ( .C1(n13381), .C2(P1_EBX_REG_11__SCAN_IN), .A(n14059), .B(
        n14290), .ZN(n14060) );
  NAND2_X1 U17457 ( .A1(n14061), .A2(n14060), .ZN(n15930) );
  NAND2_X1 U17458 ( .A1(n14797), .A2(n15930), .ZN(n14062) );
  MUX2_X1 U17459 ( .A(n14176), .B(n9581), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n14065) );
  NAND2_X1 U17460 ( .A1(n13381), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14063) );
  AND2_X1 U17461 ( .A1(n14164), .A2(n14063), .ZN(n14064) );
  NAND2_X1 U17462 ( .A1(n14065), .A2(n14064), .ZN(n14077) );
  XNOR2_X1 U17463 ( .A(n14800), .B(n14077), .ZN(n16095) );
  AOI22_X1 U17464 ( .A1(n19989), .A2(n16095), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14438), .ZN(n14066) );
  OAI21_X1 U17465 ( .B1(n14663), .B2(n14455), .A(n14066), .ZN(P1_U2859) );
  INV_X1 U17466 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n14802) );
  INV_X1 U17467 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15937) );
  NAND2_X1 U17468 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n19980) );
  NOR3_X1 U17469 ( .A1(n20840), .A2(n20749), .A3(n19980), .ZN(n19913) );
  NAND3_X1 U17470 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n19915) );
  NOR2_X1 U17471 ( .A1(n13990), .A2(n19915), .ZN(n19897) );
  NAND2_X1 U17472 ( .A1(n19913), .A2(n19897), .ZN(n19900) );
  NOR2_X1 U17473 ( .A1(n14028), .A2(n19900), .ZN(n15940) );
  NAND2_X1 U17474 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n15940), .ZN(n15938) );
  NOR3_X1 U17475 ( .A1(n14802), .A2(n15937), .A3(n15938), .ZN(n14355) );
  OAI21_X1 U17476 ( .B1(n19901), .B2(n14355), .A(n19898), .ZN(n15892) );
  AOI22_X1 U17477 ( .A1(n14658), .A2(n19909), .B1(n19942), .B2(n16095), .ZN(
        n14068) );
  NAND2_X1 U17478 ( .A1(n19898), .A2(n14067), .ZN(n19944) );
  OAI211_X1 U17479 ( .C1(n15945), .C2(n14069), .A(n14068), .B(n19944), .ZN(
        n14070) );
  AOI21_X1 U17480 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15892), .A(n14070), 
        .ZN(n14073) );
  INV_X1 U17481 ( .A(n14355), .ZN(n14071) );
  NOR2_X1 U17482 ( .A1(n19901), .A2(n14071), .ZN(n15908) );
  INV_X1 U17483 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20712) );
  AOI22_X1 U17484 ( .A1(n15908), .A2(n20712), .B1(n19974), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14072) );
  OAI211_X1 U17485 ( .C1(n14663), .C2(n19946), .A(n14073), .B(n14072), .ZN(
        P1_U2827) );
  INV_X1 U17486 ( .A(n14800), .ZN(n14076) );
  MUX2_X1 U17487 ( .A(n14179), .B(n14276), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n14075) );
  NOR2_X1 U17488 ( .A1(n14277), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14074) );
  NOR2_X1 U17489 ( .A1(n14075), .A2(n14074), .ZN(n14078) );
  AOI21_X1 U17490 ( .B1(n14076), .B2(n14077), .A(n14078), .ZN(n14080) );
  NAND2_X1 U17491 ( .A1(n14078), .A2(n14077), .ZN(n14079) );
  OR2_X1 U17492 ( .A1(n14080), .A2(n14106), .ZN(n15909) );
  INV_X1 U17493 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15913) );
  OAI222_X1 U17494 ( .A1(n15909), .A2(n14457), .B1(n15913), .B2(n19994), .C1(
        n15915), .C2(n14455), .ZN(P1_U2858) );
  XOR2_X1 U17495 ( .A(n14082), .B(n14081), .Z(n16017) );
  INV_X1 U17496 ( .A(n16017), .ZN(n14087) );
  OR2_X1 U17497 ( .A1(n20080), .A2(n14083), .ZN(n14085) );
  NAND2_X1 U17498 ( .A1(n20080), .A2(DATAI_11_), .ZN(n14084) );
  NAND2_X1 U17499 ( .A1(n14085), .A2(n14084), .ZN(n20031) );
  AOI22_X1 U17500 ( .A1(n14095), .A2(n20031), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n15957), .ZN(n14086) );
  OAI21_X1 U17501 ( .B1(n14087), .B2(n14544), .A(n14086), .ZN(P1_U2893) );
  INV_X1 U17502 ( .A(n14088), .ZN(n14092) );
  INV_X1 U17503 ( .A(n14089), .ZN(n14091) );
  INV_X1 U17504 ( .A(n16005), .ZN(n14097) );
  OR2_X1 U17505 ( .A1(n20080), .A2(n16442), .ZN(n14094) );
  NAND2_X1 U17506 ( .A1(n20080), .A2(DATAI_12_), .ZN(n14093) );
  NAND2_X1 U17507 ( .A1(n14094), .A2(n14093), .ZN(n20033) );
  AOI22_X1 U17508 ( .A1(n14095), .A2(n20033), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n15957), .ZN(n14096) );
  OAI21_X1 U17509 ( .B1(n14097), .B2(n14544), .A(n14096), .ZN(P1_U2892) );
  INV_X1 U17510 ( .A(n14098), .ZN(n14101) );
  INV_X1 U17511 ( .A(n14099), .ZN(n14454) );
  AOI21_X1 U17512 ( .B1(n14101), .B2(n14100), .A(n14454), .ZN(n16001) );
  NAND2_X1 U17513 ( .A1(n9581), .A2(n16077), .ZN(n14102) );
  OAI211_X1 U17514 ( .C1(n13381), .C2(P1_EBX_REG_15__SCAN_IN), .A(n14102), .B(
        n14290), .ZN(n14103) );
  OAI21_X1 U17515 ( .B1(n14176), .B2(P1_EBX_REG_15__SCAN_IN), .A(n14103), .ZN(
        n14105) );
  INV_X1 U17516 ( .A(n14450), .ZN(n14104) );
  OAI21_X1 U17517 ( .B1(n14106), .B2(n14105), .A(n14104), .ZN(n15904) );
  INV_X1 U17518 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14107) );
  OAI22_X1 U17519 ( .A1(n15904), .A2(n14457), .B1(n14107), .B2(n19994), .ZN(
        n14108) );
  AOI21_X1 U17520 ( .B1(n16001), .B2(n19990), .A(n14108), .ZN(n14109) );
  INV_X1 U17521 ( .A(n14109), .ZN(P1_U2857) );
  AOI22_X1 U17522 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14110) );
  OAI21_X1 U17523 ( .B1(n12721), .B2(n14111), .A(n14110), .ZN(n14120) );
  AOI22_X1 U17524 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14118) );
  OAI22_X1 U17525 ( .A1(n17113), .A2(n18160), .B1(n17146), .B2(n17128), .ZN(
        n14116) );
  AOI22_X1 U17526 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15648), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14114) );
  AOI22_X1 U17527 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17056), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14113) );
  AOI22_X1 U17528 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14112) );
  NAND3_X1 U17529 ( .A1(n14114), .A2(n14113), .A3(n14112), .ZN(n14115) );
  AOI211_X1 U17530 ( .C1(n17156), .C2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n14116), .B(n14115), .ZN(n14117) );
  OAI211_X1 U17531 ( .C1(n17004), .C2(n17134), .A(n14118), .B(n14117), .ZN(
        n14119) );
  AOI211_X1 U17532 ( .C1(n17032), .C2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n14120), .B(n14119), .ZN(n17272) );
  INV_X1 U17533 ( .A(n17272), .ZN(n14129) );
  INV_X1 U17534 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17038) );
  INV_X1 U17535 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n14126) );
  INV_X1 U17536 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n14125) );
  INV_X1 U17537 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17159) );
  INV_X1 U17538 ( .A(n18601), .ZN(n14122) );
  NAND3_X1 U17539 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17180) );
  INV_X1 U17540 ( .A(n17180), .ZN(n17176) );
  AND2_X1 U17541 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17176), .ZN(n17173) );
  NAND2_X1 U17542 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17173), .ZN(n17172) );
  NOR2_X1 U17543 ( .A1(n17240), .A2(n17022), .ZN(n17036) );
  AOI21_X1 U17544 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17036), .A(
        P3_EBX_REG_17__SCAN_IN), .ZN(n14127) );
  NOR2_X1 U17545 ( .A1(n17008), .A2(n14127), .ZN(n14128) );
  INV_X2 U17546 ( .A(n17188), .ZN(n17186) );
  MUX2_X1 U17547 ( .A(n14129), .B(n14128), .S(n17186), .Z(P3_U2686) );
  INV_X1 U17548 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16923) );
  INV_X1 U17549 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16948) );
  NOR3_X1 U17550 ( .A1(n16584), .A2(n16605), .A3(n16948), .ZN(n14130) );
  NAND3_X1 U17551 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(n14130), .ZN(n16920) );
  NAND2_X1 U17552 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16919) );
  OR2_X1 U17553 ( .A1(n16920), .A2(n16919), .ZN(n14131) );
  NOR4_X1 U17554 ( .A1(n16923), .A2(n16977), .A3(n16963), .A4(n14131), .ZN(
        n16888) );
  NAND2_X1 U17555 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16888), .ZN(n14132) );
  NOR2_X1 U17556 ( .A1(n17240), .A2(n14132), .ZN(n14134) );
  NAND2_X1 U17557 ( .A1(n17186), .A2(n14132), .ZN(n16913) );
  INV_X1 U17558 ( .A(n16913), .ZN(n14133) );
  MUX2_X1 U17559 ( .A(n14134), .B(n14133), .S(P3_EBX_REG_31__SCAN_IN), .Z(
        P3_U2672) );
  AOI22_X1 U17560 ( .A1(n11712), .A2(n14831), .B1(n14832), .B2(n11345), .ZN(
        n15759) );
  INV_X1 U17561 ( .A(n16146), .ZN(n14135) );
  OAI22_X1 U17562 ( .A1(n15759), .A2(n14135), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n20677), .ZN(n14136) );
  AOI21_X1 U17563 ( .B1(n14137), .B2(n11345), .A(n14136), .ZN(n14140) );
  AOI21_X1 U17564 ( .B1(n14834), .B2(n16146), .A(n14139), .ZN(n14138) );
  OAI22_X1 U17565 ( .A1(n14140), .A2(n14139), .B1(n14138), .B2(n11345), .ZN(
        P1_U3474) );
  INV_X1 U17566 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14191) );
  MUX2_X1 U17567 ( .A(n14179), .B(n14276), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n14144) );
  NOR2_X1 U17568 ( .A1(n14277), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14143) );
  NOR2_X1 U17569 ( .A1(n14144), .A2(n14143), .ZN(n14449) );
  MUX2_X1 U17570 ( .A(n14176), .B(n9581), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n14147) );
  NAND2_X1 U17571 ( .A1(n13381), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14145) );
  AND2_X1 U17572 ( .A1(n14164), .A2(n14145), .ZN(n14146) );
  MUX2_X1 U17573 ( .A(n14179), .B(n14276), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n14148) );
  INV_X1 U17574 ( .A(n14148), .ZN(n14150) );
  NAND2_X1 U17575 ( .A1(n14168), .A2(n16067), .ZN(n14149) );
  NAND2_X1 U17576 ( .A1(n14150), .A2(n14149), .ZN(n14362) );
  NOR2_X2 U17577 ( .A1(n14447), .A2(n14362), .ZN(n14433) );
  NAND2_X1 U17578 ( .A1(n9581), .A2(n15806), .ZN(n14151) );
  OAI211_X1 U17579 ( .C1(n13381), .C2(P1_EBX_REG_19__SCAN_IN), .A(n14151), .B(
        n14290), .ZN(n14152) );
  OAI21_X1 U17580 ( .B1(n14176), .B2(P1_EBX_REG_19__SCAN_IN), .A(n14152), .ZN(
        n14432) );
  NAND2_X1 U17581 ( .A1(n14433), .A2(n14432), .ZN(n14435) );
  INV_X1 U17582 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14153) );
  NAND2_X1 U17583 ( .A1(n14179), .A2(n14153), .ZN(n14156) );
  NAND2_X1 U17584 ( .A1(n14290), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14154) );
  OAI211_X1 U17585 ( .C1(n13381), .C2(P1_EBX_REG_20__SCAN_IN), .A(n14154), .B(
        n9581), .ZN(n14155) );
  NAND2_X1 U17586 ( .A1(n14156), .A2(n14155), .ZN(n14428) );
  INV_X1 U17587 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14421) );
  NAND2_X1 U17588 ( .A1(n14273), .A2(n14421), .ZN(n14159) );
  NAND2_X1 U17589 ( .A1(n9581), .A2(n14772), .ZN(n14157) );
  OAI211_X1 U17590 ( .C1(n13381), .C2(P1_EBX_REG_21__SCAN_IN), .A(n14157), .B(
        n14290), .ZN(n14158) );
  AND2_X1 U17591 ( .A1(n14159), .A2(n14158), .ZN(n14418) );
  MUX2_X1 U17592 ( .A(n14179), .B(n14276), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n14160) );
  INV_X1 U17593 ( .A(n14160), .ZN(n14162) );
  INV_X1 U17594 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14619) );
  NAND2_X1 U17595 ( .A1(n14168), .A2(n14619), .ZN(n14161) );
  NAND2_X1 U17596 ( .A1(n14162), .A2(n14161), .ZN(n14410) );
  MUX2_X1 U17597 ( .A(n14176), .B(n9581), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n14166) );
  NAND2_X1 U17598 ( .A1(n13381), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14163) );
  AND2_X1 U17599 ( .A1(n14164), .A2(n14163), .ZN(n14165) );
  NAND2_X1 U17600 ( .A1(n14166), .A2(n14165), .ZN(n14404) );
  MUX2_X1 U17601 ( .A(n14179), .B(n14276), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n14167) );
  INV_X1 U17602 ( .A(n14167), .ZN(n14170) );
  NAND2_X1 U17603 ( .A1(n14168), .A2(n14609), .ZN(n14169) );
  NAND2_X1 U17604 ( .A1(n14170), .A2(n14169), .ZN(n14345) );
  OR2_X2 U17605 ( .A1(n14403), .A2(n14345), .ZN(n14392) );
  INV_X1 U17606 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14395) );
  NAND2_X1 U17607 ( .A1(n14273), .A2(n14395), .ZN(n14173) );
  NAND2_X1 U17608 ( .A1(n9581), .A2(n14741), .ZN(n14171) );
  OAI211_X1 U17609 ( .C1(n13381), .C2(P1_EBX_REG_25__SCAN_IN), .A(n14171), .B(
        n14290), .ZN(n14172) );
  AND2_X1 U17610 ( .A1(n14173), .A2(n14172), .ZN(n14391) );
  MUX2_X1 U17611 ( .A(n14179), .B(n14276), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n14175) );
  NOR2_X1 U17612 ( .A1(n14277), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14174) );
  NOR2_X1 U17613 ( .A1(n14175), .A2(n14174), .ZN(n14331) );
  MUX2_X1 U17614 ( .A(n14176), .B(n9581), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n14178) );
  NAND2_X1 U17615 ( .A1(n13381), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14177) );
  NAND2_X1 U17616 ( .A1(n14178), .A2(n14177), .ZN(n14319) );
  MUX2_X1 U17617 ( .A(n14179), .B(n14276), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n14181) );
  NOR2_X1 U17618 ( .A1(n14277), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14180) );
  NOR2_X1 U17619 ( .A1(n14181), .A2(n14180), .ZN(n14182) );
  AOI21_X1 U17620 ( .B1(n14333), .B2(n14319), .A(n14182), .ZN(n14183) );
  OR2_X1 U17621 ( .A1(n14304), .A2(n14183), .ZN(n14184) );
  INV_X1 U17622 ( .A(n14184), .ZN(n14723) );
  INV_X1 U17623 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20726) );
  INV_X1 U17624 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20723) );
  NAND2_X1 U17625 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .ZN(n15893) );
  NAND3_X1 U17626 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14356) );
  NOR2_X1 U17627 ( .A1(n15893), .A2(n14356), .ZN(n14357) );
  INV_X1 U17628 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20720) );
  INV_X1 U17629 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n15873) );
  NOR2_X1 U17630 ( .A1(n20720), .A2(n15873), .ZN(n15872) );
  NAND4_X1 U17631 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n14355), .A3(n14357), 
        .A4(n15872), .ZN(n15849) );
  NOR2_X1 U17632 ( .A1(n20723), .A2(n15849), .ZN(n15846) );
  NAND2_X1 U17633 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n15846), .ZN(n15840) );
  NOR2_X1 U17634 ( .A1(n20726), .A2(n15840), .ZN(n14347) );
  NAND2_X1 U17635 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n14347), .ZN(n15829) );
  INV_X1 U17636 ( .A(n15829), .ZN(n14185) );
  AND2_X1 U17637 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n14185), .ZN(n14334) );
  AND2_X1 U17638 ( .A1(n14334), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14324) );
  NAND2_X1 U17639 ( .A1(n14324), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14186) );
  NOR2_X1 U17640 ( .A1(n19901), .A2(n14186), .ZN(n14307) );
  AND2_X1 U17641 ( .A1(n19898), .A2(n14324), .ZN(n14320) );
  NAND3_X1 U17642 ( .A1(n14320), .A2(P1_REIP_REG_27__SCAN_IN), .A3(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14187) );
  NAND2_X1 U17643 ( .A1(n19955), .A2(n14187), .ZN(n14313) );
  INV_X1 U17644 ( .A(n14313), .ZN(n14188) );
  OAI21_X1 U17645 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n14307), .A(n14188), 
        .ZN(n14190) );
  AOI22_X1 U17646 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19969), .B1(
        n19909), .B2(n14578), .ZN(n14189) );
  OAI211_X1 U17647 ( .C1(n19960), .C2(n14191), .A(n14190), .B(n14189), .ZN(
        n14192) );
  AOI21_X1 U17648 ( .B1(n14723), .B2(n19923), .A(n14192), .ZN(n14193) );
  OAI21_X1 U17649 ( .B1(n14575), .B2(n19946), .A(n14193), .ZN(P1_U2812) );
  XOR2_X1 U17650 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n9677), .Z(n15087) );
  AOI21_X1 U17651 ( .B1(n15100), .B2(n14194), .A(n9677), .ZN(n15102) );
  OAI21_X1 U17652 ( .B1(n14195), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14194), .ZN(n15115) );
  INV_X1 U17653 ( .A(n15115), .ZN(n14883) );
  NOR2_X1 U17654 ( .A1(n14883), .A2(n14882), .ZN(n14881) );
  NOR2_X1 U17655 ( .A1(n13016), .A2(n14881), .ZN(n14865) );
  NAND2_X1 U17656 ( .A1(n14857), .A2(n14198), .ZN(n14207) );
  NAND2_X1 U17657 ( .A1(n19031), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n14200) );
  NAND2_X1 U17658 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19041), .ZN(
        n14199) );
  OAI211_X1 U17659 ( .C1(n14201), .C2(n19009), .A(n14200), .B(n14199), .ZN(
        n14204) );
  NOR2_X1 U17660 ( .A1(n14202), .A2(n19011), .ZN(n14203) );
  AOI211_X1 U17661 ( .C1(n14205), .C2(n19027), .A(n14204), .B(n14203), .ZN(
        n14206) );
  OAI211_X1 U17662 ( .C1(n14208), .C2(n19008), .A(n14207), .B(n14206), .ZN(
        P2_U2825) );
  NAND2_X1 U17663 ( .A1(n10673), .A2(n15128), .ZN(n14210) );
  XNOR2_X1 U17664 ( .A(n15129), .B(n14210), .ZN(n14230) );
  INV_X1 U17665 ( .A(n14211), .ZN(n15299) );
  AND2_X1 U17666 ( .A1(n14899), .A2(n14212), .ZN(n14213) );
  OR2_X1 U17667 ( .A1(n14213), .A2(n14965), .ZN(n14977) );
  OR2_X1 U17668 ( .A1(n14905), .A2(n14214), .ZN(n14215) );
  AND2_X1 U17669 ( .A1(n15052), .A2(n14215), .ZN(n15060) );
  NAND2_X1 U17670 ( .A1(n15288), .A2(n15291), .ZN(n14216) );
  INV_X1 U17671 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19781) );
  OR2_X1 U17672 ( .A1(n16264), .A2(n19781), .ZN(n14224) );
  NAND2_X1 U17673 ( .A1(n14216), .A2(n14224), .ZN(n14217) );
  AOI21_X1 U17674 ( .B1(n16280), .B2(n15060), .A(n14217), .ZN(n14218) );
  OAI21_X1 U17675 ( .B1(n14977), .B2(n16295), .A(n14218), .ZN(n14222) );
  INV_X1 U17676 ( .A(n14219), .ZN(n14220) );
  NOR2_X1 U17677 ( .A1(n14220), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14226) );
  NOR2_X1 U17678 ( .A1(n14219), .A2(n15291), .ZN(n15135) );
  NOR3_X1 U17679 ( .A1(n14226), .A2(n15135), .A3(n16305), .ZN(n14221) );
  AOI211_X1 U17680 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n15299), .A(
        n14222), .B(n14221), .ZN(n14223) );
  OAI21_X1 U17681 ( .B1(n14230), .B2(n16274), .A(n14223), .ZN(P2_U3021) );
  INV_X1 U17682 ( .A(n19179), .ZN(n16248) );
  INV_X1 U17683 ( .A(n14977), .ZN(n14895) );
  NAND2_X1 U17684 ( .A1(n19175), .A2(n14888), .ZN(n14225) );
  OAI211_X1 U17685 ( .C1(n16259), .C2(n14893), .A(n14225), .B(n14224), .ZN(
        n14228) );
  NOR3_X1 U17686 ( .A1(n14226), .A2(n15135), .A3(n16245), .ZN(n14227) );
  AOI211_X1 U17687 ( .C1(n16248), .C2(n14895), .A(n14228), .B(n14227), .ZN(
        n14229) );
  OAI21_X1 U17688 ( .B1(n14230), .B2(n16243), .A(n14229), .ZN(P2_U2989) );
  INV_X1 U17689 ( .A(n14234), .ZN(n14238) );
  NOR2_X1 U17690 ( .A1(n14235), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14237) );
  MUX2_X1 U17691 ( .A(n14238), .B(n14237), .S(n14236), .Z(n14854) );
  NAND2_X1 U17692 ( .A1(n14854), .A2(n14239), .ZN(n14240) );
  NAND2_X1 U17693 ( .A1(n15098), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14241) );
  INV_X1 U17694 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n14245) );
  NAND2_X1 U17695 ( .A1(n10771), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14244) );
  AOI22_X1 U17696 ( .A1(n14242), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14243) );
  OAI211_X1 U17697 ( .C1(n10856), .C2(n14245), .A(n14244), .B(n14243), .ZN(
        n14246) );
  INV_X1 U17698 ( .A(n14262), .ZN(n14259) );
  AOI222_X1 U17699 ( .A1(n10910), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n14248), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n10944), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14249) );
  OAI21_X1 U17700 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15384), .A(
        n14252), .ZN(n14257) );
  INV_X1 U17701 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n14255) );
  OR2_X1 U17702 ( .A1(n16264), .A2(n14255), .ZN(n14264) );
  AOI21_X2 U17703 ( .B1(n14267), .B2(n16270), .A(n14260), .ZN(n14261) );
  OAI21_X1 U17704 ( .B1(n14270), .B2(n16274), .A(n14261), .ZN(P2_U3015) );
  NAND2_X1 U17705 ( .A1(n19166), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14263) );
  OAI211_X1 U17706 ( .C1(n19165), .C2(n14265), .A(n14264), .B(n14263), .ZN(
        n14266) );
  AOI21_X1 U17707 ( .B1(n14262), .B2(n16248), .A(n14266), .ZN(n14269) );
  NAND2_X1 U17708 ( .A1(n14267), .A2(n19169), .ZN(n14268) );
  OAI211_X1 U17709 ( .C1(n14270), .C2(n16243), .A(n14269), .B(n14268), .ZN(
        P2_U2983) );
  NAND2_X1 U17710 ( .A1(n14277), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n14272) );
  NAND2_X1 U17711 ( .A1(n13381), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14271) );
  NAND2_X1 U17712 ( .A1(n14272), .A2(n14271), .ZN(n14291) );
  OAI22_X1 U17713 ( .A1(n14277), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(n13381), .ZN(n14288) );
  OR2_X1 U17714 ( .A1(n14288), .A2(n14276), .ZN(n14275) );
  INV_X1 U17715 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14382) );
  NAND2_X1 U17716 ( .A1(n14273), .A2(n14382), .ZN(n14274) );
  NAND2_X1 U17717 ( .A1(n14275), .A2(n14274), .ZN(n14303) );
  MUX2_X1 U17718 ( .A(n14276), .B(n14291), .S(n14306), .Z(n14280) );
  NAND2_X1 U17719 ( .A1(n14306), .A2(n14291), .ZN(n14279) );
  AOI22_X1 U17720 ( .A1(n14277), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13381), .ZN(n14278) );
  MUX2_X1 U17721 ( .A(n14280), .B(n14279), .S(n14278), .Z(n14669) );
  NAND2_X1 U17722 ( .A1(n14281), .A2(n19936), .ZN(n14286) );
  INV_X1 U17723 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20736) );
  INV_X1 U17724 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14550) );
  OAI21_X1 U17725 ( .B1(n20736), .B2(n14550), .A(n19955), .ZN(n14282) );
  NAND2_X1 U17726 ( .A1(n14282), .A2(n14313), .ZN(n14294) );
  INV_X1 U17727 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14377) );
  OAI22_X1 U17728 ( .A1(n19960), .A2(n14377), .B1(n20885), .B2(n15945), .ZN(
        n14284) );
  NAND3_X1 U17729 ( .A1(n14307), .A2(P1_REIP_REG_28__SCAN_IN), .A3(
        P1_REIP_REG_29__SCAN_IN), .ZN(n14293) );
  NOR3_X1 U17730 ( .A1(n14293), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14550), 
        .ZN(n14283) );
  AOI211_X1 U17731 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14294), .A(n14284), 
        .B(n14283), .ZN(n14285) );
  OAI211_X1 U17732 ( .C1(n14669), .C2(n19977), .A(n14286), .B(n14285), .ZN(
        P1_U2809) );
  INV_X1 U17733 ( .A(n14304), .ZN(n14289) );
  OAI22_X1 U17734 ( .A1(n14306), .A2(n14290), .B1(n14289), .B2(n14288), .ZN(
        n14292) );
  XNOR2_X1 U17735 ( .A(n14292), .B(n14291), .ZN(n14378) );
  INV_X1 U17736 ( .A(n14378), .ZN(n14704) );
  INV_X1 U17737 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14379) );
  INV_X1 U17738 ( .A(n14293), .ZN(n14295) );
  OAI21_X1 U17739 ( .B1(n14295), .B2(P1_REIP_REG_30__SCAN_IN), .A(n14294), 
        .ZN(n14297) );
  AOI22_X1 U17740 ( .A1(n14549), .A2(n19909), .B1(n19969), .B2(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14296) );
  OAI211_X1 U17741 ( .C1(n19960), .C2(n14379), .A(n14297), .B(n14296), .ZN(
        n14298) );
  AOI21_X1 U17742 ( .B1(n14704), .B2(n19942), .A(n14298), .ZN(n14299) );
  OAI21_X1 U17743 ( .B1(n14380), .B2(n19946), .A(n14299), .ZN(P1_U2810) );
  AOI21_X1 U17744 ( .B1(n14302), .B2(n14301), .A(n14300), .ZN(n14563) );
  INV_X1 U17745 ( .A(n14563), .ZN(n14383) );
  NOR2_X1 U17746 ( .A1(n14304), .A2(n14303), .ZN(n14305) );
  INV_X1 U17747 ( .A(n14381), .ZN(n14715) );
  NAND3_X1 U17748 ( .A1(n14307), .A2(P1_REIP_REG_28__SCAN_IN), .A3(n20736), 
        .ZN(n14312) );
  INV_X1 U17749 ( .A(n14561), .ZN(n14308) );
  AOI22_X1 U17750 ( .A1(n14308), .A2(n19909), .B1(n19969), .B2(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14309) );
  OAI21_X1 U17751 ( .B1(n19960), .B2(n14382), .A(n14309), .ZN(n14310) );
  INV_X1 U17752 ( .A(n14310), .ZN(n14311) );
  OAI211_X1 U17753 ( .C1(n14313), .C2(n20736), .A(n14312), .B(n14311), .ZN(
        n14314) );
  AOI21_X1 U17754 ( .B1(n14715), .B2(n19923), .A(n14314), .ZN(n14315) );
  OAI21_X1 U17755 ( .B1(n14383), .B2(n19946), .A(n14315), .ZN(P1_U2811) );
  INV_X1 U17756 ( .A(n14316), .ZN(n14317) );
  AOI21_X1 U17757 ( .B1(n14318), .B2(n14317), .A(n14141), .ZN(n14587) );
  INV_X1 U17758 ( .A(n14587), .ZN(n14385) );
  XOR2_X1 U17759 ( .A(n14319), .B(n14333), .Z(n14730) );
  INV_X1 U17760 ( .A(n14320), .ZN(n14321) );
  NAND2_X1 U17761 ( .A1(n19955), .A2(n14321), .ZN(n14337) );
  INV_X1 U17762 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20733) );
  OAI22_X1 U17763 ( .A1(n14322), .A2(n15945), .B1(n19986), .B2(n14585), .ZN(
        n14323) );
  AOI21_X1 U17764 ( .B1(n19974), .B2(P1_EBX_REG_27__SCAN_IN), .A(n14323), .ZN(
        n14326) );
  NAND3_X1 U17765 ( .A1(n19914), .A2(n14324), .A3(n20733), .ZN(n14325) );
  OAI211_X1 U17766 ( .C1(n14337), .C2(n20733), .A(n14326), .B(n14325), .ZN(
        n14327) );
  AOI21_X1 U17767 ( .B1(n14730), .B2(n19923), .A(n14327), .ZN(n14328) );
  OAI21_X1 U17768 ( .B1(n14385), .B2(n19946), .A(n14328), .ZN(P1_U2813) );
  AOI21_X1 U17769 ( .B1(n14330), .B2(n14329), .A(n14316), .ZN(n14596) );
  INV_X1 U17770 ( .A(n14596), .ZN(n14388) );
  NOR2_X1 U17771 ( .A1(n14393), .A2(n14331), .ZN(n14332) );
  OR2_X1 U17772 ( .A1(n14333), .A2(n14332), .ZN(n14386) );
  INV_X1 U17773 ( .A(n14386), .ZN(n14739) );
  AOI21_X1 U17774 ( .B1(n19914), .B2(n14334), .A(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14338) );
  AOI22_X1 U17775 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19969), .B1(
        n19909), .B2(n14592), .ZN(n14336) );
  NAND2_X1 U17776 ( .A1(n19974), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14335) );
  OAI211_X1 U17777 ( .C1(n14338), .C2(n14337), .A(n14336), .B(n14335), .ZN(
        n14339) );
  AOI21_X1 U17778 ( .B1(n14739), .B2(n19923), .A(n14339), .ZN(n14340) );
  OAI21_X1 U17779 ( .B1(n14388), .B2(n19946), .A(n14340), .ZN(P1_U2814) );
  INV_X1 U17780 ( .A(n14342), .ZN(n14343) );
  OAI21_X1 U17781 ( .B1(n14344), .B2(n14341), .A(n14343), .ZN(n14612) );
  NAND2_X1 U17782 ( .A1(n14403), .A2(n14345), .ZN(n14346) );
  AND2_X1 U17783 ( .A1(n14392), .A2(n14346), .ZN(n14755) );
  OAI21_X1 U17784 ( .B1(n19901), .B2(n14347), .A(n19898), .ZN(n15842) );
  AOI22_X1 U17785 ( .A1(n14615), .A2(n19909), .B1(P1_REIP_REG_24__SCAN_IN), 
        .B2(n15842), .ZN(n14349) );
  NOR2_X1 U17786 ( .A1(n19901), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15835) );
  AOI22_X1 U17787 ( .A1(n15835), .A2(n14347), .B1(n19974), .B2(
        P1_EBX_REG_24__SCAN_IN), .ZN(n14348) );
  OAI211_X1 U17788 ( .C1(n14611), .C2(n15945), .A(n14349), .B(n14348), .ZN(
        n14350) );
  AOI21_X1 U17789 ( .B1(n14755), .B2(n19923), .A(n14350), .ZN(n14351) );
  OAI21_X1 U17790 ( .B1(n14612), .B2(n19946), .A(n14351), .ZN(P1_U2816) );
  INV_X1 U17791 ( .A(n14352), .ZN(n14443) );
  AOI21_X1 U17792 ( .B1(n14354), .B2(n14443), .A(n14353), .ZN(n14631) );
  INV_X1 U17793 ( .A(n14631), .ZN(n14440) );
  NAND4_X1 U17794 ( .A1(n19914), .A2(n14355), .A3(P1_REIP_REG_14__SCAN_IN), 
        .A4(P1_REIP_REG_13__SCAN_IN), .ZN(n15907) );
  NOR2_X1 U17795 ( .A1(n14356), .A2(n15907), .ZN(n15874) );
  INV_X1 U17796 ( .A(n15892), .ZN(n15928) );
  OAI21_X1 U17797 ( .B1(n19901), .B2(n14357), .A(n15928), .ZN(n15884) );
  INV_X1 U17798 ( .A(n14629), .ZN(n14358) );
  AOI22_X1 U17799 ( .A1(n19974), .A2(P1_EBX_REG_18__SCAN_IN), .B1(n19909), 
        .B2(n14358), .ZN(n14359) );
  OAI211_X1 U17800 ( .C1(n15945), .C2(n14360), .A(n14359), .B(n19944), .ZN(
        n14361) );
  AOI221_X1 U17801 ( .B1(n15874), .B2(n15873), .C1(n15884), .C2(
        P1_REIP_REG_18__SCAN_IN), .A(n14361), .ZN(n14364) );
  AOI21_X1 U17802 ( .B1(n14362), .B2(n14447), .A(n14433), .ZN(n16063) );
  NAND2_X1 U17803 ( .A1(n16063), .A2(n19923), .ZN(n14363) );
  OAI211_X1 U17804 ( .C1(n14440), .C2(n19946), .A(n14364), .B(n14363), .ZN(
        P1_U2822) );
  INV_X1 U17805 ( .A(n14365), .ZN(n14366) );
  AOI22_X1 U17806 ( .A1(n14366), .A2(n19909), .B1(n19969), .B2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14367) );
  OAI21_X1 U17807 ( .B1(n13572), .B2(n19972), .A(n14367), .ZN(n14368) );
  AOI21_X1 U17808 ( .B1(n19974), .B2(P1_EBX_REG_2__SCAN_IN), .A(n14368), .ZN(
        n14369) );
  OAI21_X1 U17809 ( .B1(n19977), .B2(n14370), .A(n14369), .ZN(n14372) );
  AOI211_X1 U17810 ( .C1(P1_REIP_REG_2__SCAN_IN), .C2(n14373), .A(n14372), .B(
        n14371), .ZN(n14374) );
  OAI21_X1 U17811 ( .B1(n14376), .B2(n14375), .A(n14374), .ZN(P1_U2838) );
  OAI22_X1 U17812 ( .A1(n14669), .A2(n14457), .B1(n19994), .B2(n14377), .ZN(
        P1_U2841) );
  OAI222_X1 U17813 ( .A1(n14455), .A2(n14380), .B1(n14379), .B2(n19994), .C1(
        n14378), .C2(n14457), .ZN(P1_U2842) );
  OAI222_X1 U17814 ( .A1(n14455), .A2(n14383), .B1(n14382), .B2(n19994), .C1(
        n14381), .C2(n14457), .ZN(P1_U2843) );
  AOI22_X1 U17815 ( .A1(n14730), .A2(n19989), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n14438), .ZN(n14384) );
  OAI21_X1 U17816 ( .B1(n14385), .B2(n14455), .A(n14384), .ZN(P1_U2845) );
  INV_X1 U17817 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14387) );
  OAI222_X1 U17818 ( .A1(n14455), .A2(n14388), .B1(n19994), .B2(n14387), .C1(
        n14386), .C2(n14457), .ZN(P1_U2846) );
  OR2_X1 U17819 ( .A1(n14342), .A2(n14389), .ZN(n14390) );
  AND2_X1 U17820 ( .A1(n14329), .A2(n14390), .ZN(n15834) );
  AND2_X1 U17821 ( .A1(n14392), .A2(n14391), .ZN(n14394) );
  OR2_X1 U17822 ( .A1(n14394), .A2(n14393), .ZN(n15838) );
  OAI22_X1 U17823 ( .A1(n15838), .A2(n14457), .B1(n14395), .B2(n19994), .ZN(
        n14396) );
  AOI21_X1 U17824 ( .B1(n15834), .B2(n19990), .A(n14396), .ZN(n14397) );
  INV_X1 U17825 ( .A(n14397), .ZN(P1_U2847) );
  AOI22_X1 U17826 ( .A1(n14755), .A2(n19989), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n14438), .ZN(n14398) );
  OAI21_X1 U17827 ( .B1(n14612), .B2(n14455), .A(n14398), .ZN(P1_U2848) );
  INV_X1 U17828 ( .A(n14399), .ZN(n14400) );
  AND2_X1 U17829 ( .A1(n14400), .A2(n14401), .ZN(n14402) );
  NOR2_X1 U17830 ( .A1(n14341), .A2(n14402), .ZN(n15968) );
  INV_X1 U17831 ( .A(n15968), .ZN(n14406) );
  INV_X1 U17832 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14405) );
  OAI21_X1 U17833 ( .B1(n14412), .B2(n14404), .A(n14403), .ZN(n16042) );
  OAI222_X1 U17834 ( .A1(n14406), .A2(n14455), .B1(n14405), .B2(n19994), .C1(
        n16042), .C2(n14457), .ZN(P1_U2849) );
  NAND2_X1 U17835 ( .A1(n14407), .A2(n14408), .ZN(n14409) );
  INV_X1 U17836 ( .A(n15848), .ZN(n14414) );
  AND2_X1 U17837 ( .A1(n14420), .A2(n14410), .ZN(n14411) );
  NOR2_X1 U17838 ( .A1(n14412), .A2(n14411), .ZN(n16052) );
  AOI22_X1 U17839 ( .A1(n16052), .A2(n19989), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n14438), .ZN(n14413) );
  OAI21_X1 U17840 ( .B1(n14414), .B2(n14455), .A(n14413), .ZN(P1_U2850) );
  OAI21_X1 U17841 ( .B1(n14415), .B2(n14416), .A(n14407), .ZN(n14417) );
  NAND2_X1 U17842 ( .A1(n14427), .A2(n14418), .ZN(n14419) );
  NAND2_X1 U17843 ( .A1(n14420), .A2(n14419), .ZN(n15861) );
  OAI22_X1 U17844 ( .A1(n15861), .A2(n14457), .B1(n14421), .B2(n19994), .ZN(
        n14422) );
  AOI21_X1 U17845 ( .B1(n15973), .B2(n19990), .A(n14422), .ZN(n14423) );
  INV_X1 U17846 ( .A(n14423), .ZN(P1_U2851) );
  INV_X1 U17847 ( .A(n14415), .ZN(n14425) );
  OAI21_X1 U17848 ( .B1(n14426), .B2(n14424), .A(n14425), .ZN(n15978) );
  AOI21_X1 U17849 ( .B1(n14428), .B2(n14435), .A(n9879), .ZN(n15865) );
  AOI22_X1 U17850 ( .A1(n15865), .A2(n19989), .B1(P1_EBX_REG_20__SCAN_IN), 
        .B2(n14438), .ZN(n14429) );
  OAI21_X1 U17851 ( .B1(n15978), .B2(n14455), .A(n14429), .ZN(P1_U2852) );
  NOR2_X1 U17852 ( .A1(n14353), .A2(n14430), .ZN(n14431) );
  OR2_X1 U17853 ( .A1(n14424), .A2(n14431), .ZN(n15985) );
  OR2_X1 U17854 ( .A1(n14433), .A2(n14432), .ZN(n14434) );
  NAND2_X1 U17855 ( .A1(n14435), .A2(n14434), .ZN(n15879) );
  INV_X1 U17856 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15869) );
  OAI22_X1 U17857 ( .A1(n15879), .A2(n14457), .B1(n15869), .B2(n19994), .ZN(
        n14436) );
  AOI21_X1 U17858 ( .B1(n15876), .B2(n19990), .A(n14436), .ZN(n14437) );
  INV_X1 U17859 ( .A(n14437), .ZN(P1_U2853) );
  AOI22_X1 U17860 ( .A1(n16063), .A2(n19989), .B1(P1_EBX_REG_18__SCAN_IN), 
        .B2(n14438), .ZN(n14439) );
  OAI21_X1 U17861 ( .B1(n14440), .B2(n14455), .A(n14439), .ZN(P1_U2854) );
  AOI21_X1 U17862 ( .B1(n14444), .B2(n14452), .A(n14352), .ZN(n15997) );
  INV_X1 U17863 ( .A(n15997), .ZN(n14448) );
  INV_X1 U17864 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15881) );
  NAND2_X1 U17865 ( .A1(n9658), .A2(n14445), .ZN(n14446) );
  NAND2_X1 U17866 ( .A1(n14447), .A2(n14446), .ZN(n16068) );
  OAI222_X1 U17867 ( .A1(n14448), .A2(n14455), .B1(n19994), .B2(n15881), .C1(
        n16068), .C2(n14457), .ZN(P1_U2855) );
  OAI21_X1 U17868 ( .B1(n14450), .B2(n14449), .A(n9658), .ZN(n15889) );
  INV_X1 U17869 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14456) );
  INV_X1 U17870 ( .A(n14451), .ZN(n14453) );
  OAI21_X1 U17871 ( .B1(n14454), .B2(n14453), .A(n14452), .ZN(n15894) );
  OAI222_X1 U17872 ( .A1(n15889), .A2(n14457), .B1(n14456), .B2(n19994), .C1(
        n15894), .C2(n14455), .ZN(P1_U2856) );
  NAND2_X1 U17873 ( .A1(n14554), .A2(n15961), .ZN(n14463) );
  AOI22_X1 U17874 ( .A1(n15959), .A2(n20037), .B1(n15957), .B2(
        P1_EAX_REG_30__SCAN_IN), .ZN(n14462) );
  NAND2_X1 U17875 ( .A1(n15960), .A2(DATAI_30_), .ZN(n14461) );
  INV_X1 U17876 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n14459) );
  OR2_X1 U17877 ( .A1(n15964), .A2(n14459), .ZN(n14460) );
  NAND4_X1 U17878 ( .A1(n14463), .A2(n14462), .A3(n14461), .A4(n14460), .ZN(
        P1_U2874) );
  NAND2_X1 U17879 ( .A1(n14563), .A2(n15961), .ZN(n14468) );
  AOI22_X1 U17880 ( .A1(n15959), .A2(n20035), .B1(n15957), .B2(
        P1_EAX_REG_29__SCAN_IN), .ZN(n14467) );
  NAND2_X1 U17881 ( .A1(n15960), .A2(DATAI_29_), .ZN(n14466) );
  INV_X1 U17882 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n14464) );
  OR2_X1 U17883 ( .A1(n15964), .A2(n14464), .ZN(n14465) );
  NAND4_X1 U17884 ( .A1(n14468), .A2(n14467), .A3(n14466), .A4(n14465), .ZN(
        P1_U2875) );
  INV_X1 U17885 ( .A(n14575), .ZN(n14469) );
  NAND2_X1 U17886 ( .A1(n14469), .A2(n15961), .ZN(n14474) );
  AOI22_X1 U17887 ( .A1(n15959), .A2(n20033), .B1(n15957), .B2(
        P1_EAX_REG_28__SCAN_IN), .ZN(n14473) );
  NAND2_X1 U17888 ( .A1(n15960), .A2(DATAI_28_), .ZN(n14472) );
  INV_X1 U17889 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n14470) );
  OR2_X1 U17890 ( .A1(n15964), .A2(n14470), .ZN(n14471) );
  NAND4_X1 U17891 ( .A1(n14474), .A2(n14473), .A3(n14472), .A4(n14471), .ZN(
        P1_U2876) );
  NAND2_X1 U17892 ( .A1(n14587), .A2(n15961), .ZN(n14478) );
  AOI22_X1 U17893 ( .A1(n15959), .A2(n20031), .B1(n15957), .B2(
        P1_EAX_REG_27__SCAN_IN), .ZN(n14477) );
  NAND2_X1 U17894 ( .A1(n15960), .A2(DATAI_27_), .ZN(n14476) );
  INV_X1 U17895 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16426) );
  OR2_X1 U17896 ( .A1(n15964), .A2(n16426), .ZN(n14475) );
  NAND4_X1 U17897 ( .A1(n14478), .A2(n14477), .A3(n14476), .A4(n14475), .ZN(
        P1_U2877) );
  NAND2_X1 U17898 ( .A1(n14596), .A2(n15961), .ZN(n14483) );
  AOI22_X1 U17899 ( .A1(n15959), .A2(n20029), .B1(n15957), .B2(
        P1_EAX_REG_26__SCAN_IN), .ZN(n14482) );
  NAND2_X1 U17900 ( .A1(n15960), .A2(DATAI_26_), .ZN(n14481) );
  INV_X1 U17901 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n14479) );
  OR2_X1 U17902 ( .A1(n15964), .A2(n14479), .ZN(n14480) );
  NAND4_X1 U17903 ( .A1(n14483), .A2(n14482), .A3(n14481), .A4(n14480), .ZN(
        P1_U2878) );
  INV_X1 U17904 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n14486) );
  NAND2_X1 U17905 ( .A1(n15960), .A2(DATAI_25_), .ZN(n14485) );
  AOI22_X1 U17906 ( .A1(n15959), .A2(n20027), .B1(n15957), .B2(
        P1_EAX_REG_25__SCAN_IN), .ZN(n14484) );
  OAI211_X1 U17907 ( .C1(n14486), .C2(n15964), .A(n14485), .B(n14484), .ZN(
        n14487) );
  AOI21_X1 U17908 ( .B1(n15834), .B2(n15961), .A(n14487), .ZN(n14488) );
  INV_X1 U17909 ( .A(n14488), .ZN(P1_U2879) );
  INV_X1 U17910 ( .A(n14612), .ZN(n14493) );
  INV_X1 U17911 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n14491) );
  NAND2_X1 U17912 ( .A1(n15960), .A2(DATAI_24_), .ZN(n14490) );
  AOI22_X1 U17913 ( .A1(n15959), .A2(n20025), .B1(n15957), .B2(
        P1_EAX_REG_24__SCAN_IN), .ZN(n14489) );
  OAI211_X1 U17914 ( .C1(n14491), .C2(n15964), .A(n14490), .B(n14489), .ZN(
        n14492) );
  AOI21_X1 U17915 ( .B1(n14493), .B2(n15961), .A(n14492), .ZN(n14494) );
  INV_X1 U17916 ( .A(n14494), .ZN(P1_U2880) );
  INV_X1 U17917 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n14498) );
  NAND2_X1 U17918 ( .A1(n15960), .A2(DATAI_22_), .ZN(n14497) );
  AOI22_X1 U17919 ( .A1(n15959), .A2(n14495), .B1(n15957), .B2(
        P1_EAX_REG_22__SCAN_IN), .ZN(n14496) );
  OAI211_X1 U17920 ( .C1(n15964), .C2(n14498), .A(n14497), .B(n14496), .ZN(
        n14499) );
  AOI21_X1 U17921 ( .B1(n15848), .B2(n15961), .A(n14499), .ZN(n14500) );
  INV_X1 U17922 ( .A(n14500), .ZN(P1_U2882) );
  NAND2_X1 U17923 ( .A1(n15973), .A2(n15961), .ZN(n14506) );
  AOI22_X1 U17924 ( .A1(n15959), .A2(n14501), .B1(n15957), .B2(
        P1_EAX_REG_21__SCAN_IN), .ZN(n14505) );
  NAND2_X1 U17925 ( .A1(n15960), .A2(DATAI_21_), .ZN(n14504) );
  INV_X1 U17926 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n14502) );
  OR2_X1 U17927 ( .A1(n15964), .A2(n14502), .ZN(n14503) );
  NAND4_X1 U17928 ( .A1(n14506), .A2(n14505), .A3(n14504), .A4(n14503), .ZN(
        P1_U2883) );
  INV_X1 U17929 ( .A(n15978), .ZN(n14512) );
  INV_X1 U17930 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n14510) );
  NAND2_X1 U17931 ( .A1(n15960), .A2(DATAI_20_), .ZN(n14509) );
  AOI22_X1 U17932 ( .A1(n15959), .A2(n14507), .B1(n15957), .B2(
        P1_EAX_REG_20__SCAN_IN), .ZN(n14508) );
  OAI211_X1 U17933 ( .C1(n15964), .C2(n14510), .A(n14509), .B(n14508), .ZN(
        n14511) );
  AOI21_X1 U17934 ( .B1(n14512), .B2(n15961), .A(n14511), .ZN(n14513) );
  INV_X1 U17935 ( .A(n14513), .ZN(P1_U2884) );
  NAND2_X1 U17936 ( .A1(n15876), .A2(n15961), .ZN(n14519) );
  AOI22_X1 U17937 ( .A1(n15959), .A2(n14514), .B1(n15957), .B2(
        P1_EAX_REG_19__SCAN_IN), .ZN(n14518) );
  NAND2_X1 U17938 ( .A1(n15960), .A2(DATAI_19_), .ZN(n14517) );
  OR2_X1 U17939 ( .A1(n15964), .A2(n14515), .ZN(n14516) );
  NAND4_X1 U17940 ( .A1(n14519), .A2(n14518), .A3(n14517), .A4(n14516), .ZN(
        P1_U2885) );
  NAND2_X1 U17941 ( .A1(n14631), .A2(n15961), .ZN(n14525) );
  AOI22_X1 U17942 ( .A1(n15959), .A2(n14520), .B1(n15957), .B2(
        P1_EAX_REG_18__SCAN_IN), .ZN(n14524) );
  NAND2_X1 U17943 ( .A1(n15960), .A2(DATAI_18_), .ZN(n14523) );
  INV_X1 U17944 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n14521) );
  OR2_X1 U17945 ( .A1(n15964), .A2(n14521), .ZN(n14522) );
  NAND4_X1 U17946 ( .A1(n14525), .A2(n14524), .A3(n14523), .A4(n14522), .ZN(
        P1_U2886) );
  NAND2_X1 U17947 ( .A1(n15997), .A2(n15961), .ZN(n14531) );
  AOI22_X1 U17948 ( .A1(n15959), .A2(n14526), .B1(n15957), .B2(
        P1_EAX_REG_17__SCAN_IN), .ZN(n14530) );
  NAND2_X1 U17949 ( .A1(n15960), .A2(DATAI_17_), .ZN(n14529) );
  INV_X1 U17950 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n14527) );
  OR2_X1 U17951 ( .A1(n15964), .A2(n14527), .ZN(n14528) );
  NAND4_X1 U17952 ( .A1(n14531), .A2(n14530), .A3(n14529), .A4(n14528), .ZN(
        P1_U2887) );
  INV_X1 U17953 ( .A(n15894), .ZN(n14532) );
  NAND2_X1 U17954 ( .A1(n14532), .A2(n15961), .ZN(n14538) );
  AOI22_X1 U17955 ( .A1(n15959), .A2(n14533), .B1(n15957), .B2(
        P1_EAX_REG_16__SCAN_IN), .ZN(n14537) );
  NAND2_X1 U17956 ( .A1(n15960), .A2(DATAI_16_), .ZN(n14536) );
  INV_X1 U17957 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n14534) );
  OR2_X1 U17958 ( .A1(n15964), .A2(n14534), .ZN(n14535) );
  NAND4_X1 U17959 ( .A1(n14538), .A2(n14537), .A3(n14536), .A4(n14535), .ZN(
        P1_U2888) );
  INV_X1 U17960 ( .A(n16001), .ZN(n14543) );
  INV_X1 U17961 ( .A(n14539), .ZN(n14541) );
  INV_X1 U17962 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n19996) );
  OAI222_X1 U17963 ( .A1(n14544), .A2(n14543), .B1(n14542), .B2(n14541), .C1(
        n14540), .C2(n19996), .ZN(P1_U2889) );
  INV_X1 U17964 ( .A(n14545), .ZN(n14546) );
  OAI21_X1 U17965 ( .B1(n14557), .B2(n14547), .A(n14546), .ZN(n14548) );
  XNOR2_X1 U17966 ( .A(n14548), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14710) );
  INV_X1 U17967 ( .A(n14549), .ZN(n14552) );
  NOR2_X1 U17968 ( .A1(n16041), .A2(n14550), .ZN(n14703) );
  AOI21_X1 U17969 ( .B1(n20058), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14703), .ZN(n14551) );
  OAI21_X1 U17970 ( .B1(n16034), .B2(n14552), .A(n14551), .ZN(n14553) );
  OAI21_X1 U17971 ( .B1(n14710), .B2(n19879), .A(n14555), .ZN(P1_U2969) );
  NAND2_X1 U17972 ( .A1(n14557), .A2(n14556), .ZN(n14559) );
  XOR2_X1 U17973 ( .A(n14559), .B(n14558), .Z(n14717) );
  NOR2_X1 U17974 ( .A1(n16041), .A2(n20736), .ZN(n14714) );
  AOI21_X1 U17975 ( .B1(n20058), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14714), .ZN(n14560) );
  OAI21_X1 U17976 ( .B1(n16034), .B2(n14561), .A(n14560), .ZN(n14562) );
  AOI21_X1 U17977 ( .B1(n14563), .B2(n16031), .A(n14562), .ZN(n14564) );
  OAI21_X1 U17978 ( .B1(n19879), .B2(n14717), .A(n14564), .ZN(P1_U2970) );
  NAND2_X1 U17979 ( .A1(n15965), .A2(n14736), .ZN(n14565) );
  NAND2_X1 U17980 ( .A1(n15967), .A2(n14565), .ZN(n14570) );
  NAND2_X1 U17981 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14566) );
  NOR2_X1 U17982 ( .A1(n14570), .A2(n14566), .ZN(n14572) );
  INV_X1 U17983 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14582) );
  INV_X1 U17984 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14580) );
  NAND2_X1 U17985 ( .A1(n14582), .A2(n14580), .ZN(n14567) );
  NOR2_X1 U17986 ( .A1(n14568), .A2(n14567), .ZN(n14569) );
  AND2_X1 U17987 ( .A1(n14570), .A2(n14569), .ZN(n14571) );
  MUX2_X1 U17988 ( .A(n14572), .B(n14571), .S(n16013), .Z(n14573) );
  XNOR2_X1 U17989 ( .A(n14573), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14726) );
  INV_X1 U17990 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14574) );
  NAND2_X1 U17991 ( .A1(n16139), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14718) );
  OAI21_X1 U17992 ( .B1(n16039), .B2(n14574), .A(n14718), .ZN(n14577) );
  NOR2_X1 U17993 ( .A1(n14575), .A2(n20081), .ZN(n14576) );
  OAI21_X1 U17994 ( .B1(n19879), .B2(n14726), .A(n14579), .ZN(P1_U2971) );
  NAND2_X1 U17995 ( .A1(n14590), .A2(n14580), .ZN(n14581) );
  MUX2_X1 U17996 ( .A(n9645), .B(n14581), .S(n16013), .Z(n14583) );
  XNOR2_X1 U17997 ( .A(n14583), .B(n14582), .ZN(n14734) );
  NOR2_X1 U17998 ( .A1(n16041), .A2(n20733), .ZN(n14729) );
  AOI21_X1 U17999 ( .B1(n20058), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14729), .ZN(n14584) );
  OAI21_X1 U18000 ( .B1(n16034), .B2(n14585), .A(n14584), .ZN(n14586) );
  AOI21_X1 U18001 ( .B1(n14587), .B2(n16031), .A(n14586), .ZN(n14588) );
  OAI21_X1 U18002 ( .B1(n19879), .B2(n14734), .A(n14588), .ZN(P1_U2972) );
  INV_X1 U18003 ( .A(n15967), .ZN(n14606) );
  NOR2_X1 U18004 ( .A1(n14606), .A2(n14736), .ZN(n14589) );
  MUX2_X1 U18005 ( .A(n14590), .B(n14589), .S(n15965), .Z(n14591) );
  XNOR2_X1 U18006 ( .A(n14591), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14746) );
  INV_X1 U18007 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14594) );
  NAND2_X1 U18008 ( .A1(n16007), .A2(n14592), .ZN(n14593) );
  NAND2_X1 U18009 ( .A1(n16139), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14735) );
  OAI211_X1 U18010 ( .C1(n16039), .C2(n14594), .A(n14593), .B(n14735), .ZN(
        n14595) );
  AOI21_X1 U18011 ( .B1(n14596), .B2(n16031), .A(n14595), .ZN(n14597) );
  OAI21_X1 U18012 ( .B1(n19879), .B2(n14746), .A(n14597), .ZN(P1_U2973) );
  NAND2_X1 U18013 ( .A1(n14598), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14607) );
  NAND2_X1 U18014 ( .A1(n14606), .A2(n16047), .ZN(n14599) );
  MUX2_X1 U18015 ( .A(n14599), .B(n14609), .S(n15965), .Z(n14600) );
  AOI21_X1 U18016 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14607), .A(
        n14600), .ZN(n14601) );
  XNOR2_X1 U18017 ( .A(n14601), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14752) );
  NAND2_X1 U18018 ( .A1(n16007), .A2(n15830), .ZN(n14602) );
  NAND2_X1 U18019 ( .A1(n16139), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14747) );
  OAI211_X1 U18020 ( .C1(n16039), .C2(n14603), .A(n14602), .B(n14747), .ZN(
        n14604) );
  AOI21_X1 U18021 ( .B1(n15834), .B2(n16031), .A(n14604), .ZN(n14605) );
  OAI21_X1 U18022 ( .B1(n19879), .B2(n14752), .A(n14605), .ZN(P1_U2974) );
  NAND2_X1 U18023 ( .A1(n14607), .A2(n14606), .ZN(n14608) );
  MUX2_X1 U18024 ( .A(n14608), .B(n14607), .S(n15965), .Z(n14610) );
  XNOR2_X1 U18025 ( .A(n14610), .B(n14609), .ZN(n14762) );
  NAND2_X1 U18026 ( .A1(n16139), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14756) );
  OAI21_X1 U18027 ( .B1(n16039), .B2(n14611), .A(n14756), .ZN(n14614) );
  NOR2_X1 U18028 ( .A1(n14612), .A2(n20081), .ZN(n14613) );
  AOI211_X1 U18029 ( .C1(n16007), .C2(n14615), .A(n14614), .B(n14613), .ZN(
        n14616) );
  OAI21_X1 U18030 ( .B1(n19879), .B2(n14762), .A(n14616), .ZN(P1_U2975) );
  NAND2_X1 U18031 ( .A1(n14618), .A2(n14617), .ZN(n14620) );
  XNOR2_X1 U18032 ( .A(n14620), .B(n14619), .ZN(n16049) );
  NAND2_X1 U18033 ( .A1(n15848), .A2(n16031), .ZN(n14625) );
  INV_X1 U18034 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n14621) );
  OAI22_X1 U18035 ( .A1(n16039), .A2(n14622), .B1(n16041), .B2(n14621), .ZN(
        n14623) );
  AOI21_X1 U18036 ( .B1(n16007), .B2(n15847), .A(n14623), .ZN(n14624) );
  OAI211_X1 U18037 ( .C1(n16049), .C2(n19879), .A(n14625), .B(n14624), .ZN(
        P1_U2977) );
  OAI21_X1 U18038 ( .B1(n14627), .B2(n14626), .A(n15809), .ZN(n16062) );
  AOI22_X1 U18039 ( .A1(n20058), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n16139), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14628) );
  OAI21_X1 U18040 ( .B1(n16034), .B2(n14629), .A(n14628), .ZN(n14630) );
  AOI21_X1 U18041 ( .B1(n14631), .B2(n16031), .A(n14630), .ZN(n14632) );
  OAI21_X1 U18042 ( .B1(n19879), .B2(n16062), .A(n14632), .ZN(P1_U2981) );
  INV_X1 U18043 ( .A(n14635), .ZN(n14636) );
  OAI21_X1 U18044 ( .B1(n14781), .B2(n14637), .A(n14782), .ZN(n15992) );
  XNOR2_X1 U18045 ( .A(n15992), .B(n15990), .ZN(n16080) );
  NAND2_X1 U18046 ( .A1(n16080), .A2(n20060), .ZN(n14641) );
  INV_X1 U18047 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14638) );
  NOR2_X1 U18048 ( .A1(n16041), .A2(n14638), .ZN(n16074) );
  NOR2_X1 U18049 ( .A1(n16039), .A2(n15891), .ZN(n14639) );
  AOI211_X1 U18050 ( .C1(n16007), .C2(n15897), .A(n16074), .B(n14639), .ZN(
        n14640) );
  OAI211_X1 U18051 ( .C1(n20081), .C2(n15894), .A(n14641), .B(n14640), .ZN(
        P1_U2983) );
  OAI21_X1 U18052 ( .B1(n14643), .B2(n15965), .A(n14642), .ZN(n14645) );
  XNOR2_X1 U18053 ( .A(n15965), .B(n16085), .ZN(n14644) );
  XNOR2_X1 U18054 ( .A(n14645), .B(n14644), .ZN(n16089) );
  NAND2_X1 U18055 ( .A1(n16089), .A2(n20060), .ZN(n14649) );
  INV_X1 U18056 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n14646) );
  NOR2_X1 U18057 ( .A1(n16041), .A2(n14646), .ZN(n16087) );
  NOR2_X1 U18058 ( .A1(n16034), .A2(n15916), .ZN(n14647) );
  AOI211_X1 U18059 ( .C1(n20058), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16087), .B(n14647), .ZN(n14648) );
  OAI211_X1 U18060 ( .C1(n20081), .C2(n15915), .A(n14649), .B(n14648), .ZN(
        P1_U2985) );
  INV_X1 U18061 ( .A(n14650), .ZN(n14651) );
  AOI22_X1 U18062 ( .A1(n14653), .A2(n14652), .B1(n16013), .B2(n14651), .ZN(
        n14795) );
  INV_X1 U18063 ( .A(n14655), .ZN(n14654) );
  AOI21_X1 U18064 ( .B1(n16013), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n14654), .ZN(n14794) );
  NAND2_X1 U18065 ( .A1(n14795), .A2(n14794), .ZN(n14793) );
  NAND2_X1 U18066 ( .A1(n14793), .A2(n14655), .ZN(n14657) );
  XNOR2_X1 U18067 ( .A(n14657), .B(n14656), .ZN(n16097) );
  NAND2_X1 U18068 ( .A1(n16097), .A2(n20060), .ZN(n14662) );
  NOR2_X1 U18069 ( .A1(n16041), .A2(n20712), .ZN(n16094) );
  INV_X1 U18070 ( .A(n14658), .ZN(n14659) );
  NOR2_X1 U18071 ( .A1(n16034), .A2(n14659), .ZN(n14660) );
  AOI211_X1 U18072 ( .C1(n20058), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16094), .B(n14660), .ZN(n14661) );
  OAI211_X1 U18073 ( .C1(n20081), .C2(n14663), .A(n14662), .B(n14661), .ZN(
        P1_U2986) );
  MUX2_X1 U18074 ( .A(n16011), .B(n16012), .S(n16013), .Z(n14664) );
  XNOR2_X1 U18075 ( .A(n14664), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16111) );
  NAND2_X1 U18076 ( .A1(n16111), .A2(n20060), .ZN(n14668) );
  INV_X1 U18077 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14665) );
  NOR2_X1 U18078 ( .A1(n16041), .A2(n14665), .ZN(n16108) );
  NOR2_X1 U18079 ( .A1(n16034), .A2(n15941), .ZN(n14666) );
  AOI211_X1 U18080 ( .C1(n20058), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16108), .B(n14666), .ZN(n14667) );
  OAI211_X1 U18081 ( .C1(n20081), .C2(n15946), .A(n14668), .B(n14667), .ZN(
        P1_U2989) );
  INV_X1 U18082 ( .A(n14669), .ZN(n14682) );
  INV_X1 U18083 ( .A(n14670), .ZN(n14681) );
  NAND3_X1 U18084 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n14671), .ZN(n14806) );
  NOR2_X1 U18085 ( .A1(n14058), .A2(n14806), .ZN(n14811) );
  NAND2_X1 U18086 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14811), .ZN(
        n14672) );
  NOR2_X1 U18087 ( .A1(n14807), .A2(n14672), .ZN(n14683) );
  INV_X1 U18088 ( .A(n14672), .ZN(n14674) );
  NAND2_X1 U18089 ( .A1(n14674), .A2(n14673), .ZN(n14684) );
  NAND3_X1 U18090 ( .A1(n14692), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n14683), .ZN(n14675) );
  OAI21_X1 U18091 ( .B1(n14684), .B2(n14810), .A(n14675), .ZN(n15807) );
  AOI21_X1 U18092 ( .B1(n15808), .B2(n14683), .A(n15807), .ZN(n16100) );
  NOR2_X1 U18093 ( .A1(n16100), .A2(n14643), .ZN(n16061) );
  INV_X1 U18094 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16083) );
  NOR2_X1 U18095 ( .A1(n16077), .A2(n16083), .ZN(n16076) );
  NAND3_X1 U18096 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n16076), .ZN(n16059) );
  NOR2_X1 U18097 ( .A1(n16067), .A2(n16059), .ZN(n14685) );
  AND4_X1 U18098 ( .A1(n14685), .A2(n14688), .A3(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14676) );
  NAND2_X1 U18099 ( .A1(n16061), .A2(n14676), .ZN(n16048) );
  INV_X1 U18100 ( .A(n14736), .ZN(n14677) );
  NAND2_X1 U18101 ( .A1(n14677), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14678) );
  NOR2_X1 U18102 ( .A1(n16048), .A2(n14678), .ZN(n14719) );
  NAND3_X1 U18103 ( .A1(n14719), .A2(n11633), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14705) );
  INV_X1 U18104 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14679) );
  NOR3_X1 U18105 ( .A1(n14705), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14679), .ZN(n14680) );
  AOI211_X1 U18106 ( .C1(n14682), .C2(n20067), .A(n14681), .B(n14680), .ZN(
        n14702) );
  INV_X1 U18107 ( .A(n14695), .ZN(n16121) );
  NAND2_X1 U18108 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16053) );
  INV_X1 U18109 ( .A(n14683), .ZN(n14786) );
  NAND2_X1 U18110 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14685), .ZN(
        n14775) );
  NOR2_X1 U18111 ( .A1(n14643), .A2(n14684), .ZN(n16086) );
  OAI221_X1 U18112 ( .B1(n14810), .B2(n14685), .C1(n14810), .C2(n16086), .A(
        n14788), .ZN(n14686) );
  AOI221_X1 U18113 ( .B1(n14786), .B2(n14805), .C1(n14775), .C2(n14805), .A(
        n14686), .ZN(n15821) );
  AOI21_X1 U18114 ( .B1(n15821), .B2(n14688), .A(n14687), .ZN(n16050) );
  AOI21_X1 U18115 ( .B1(n16121), .B2(n16053), .A(n16050), .ZN(n16046) );
  OR2_X1 U18116 ( .A1(n14810), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14689) );
  AND2_X1 U18117 ( .A1(n16046), .A2(n14689), .ZN(n14753) );
  OR2_X1 U18118 ( .A1(n15808), .A2(n14690), .ZN(n14693) );
  INV_X1 U18119 ( .A(n14742), .ZN(n14691) );
  AOI22_X1 U18120 ( .A1(n14693), .A2(n14736), .B1(n14692), .B2(n14691), .ZN(
        n14694) );
  NAND2_X1 U18121 ( .A1(n14740), .A2(n14695), .ZN(n14700) );
  NAND3_X1 U18122 ( .A1(n14740), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14696) );
  AOI211_X1 U18123 ( .C1(n14698), .C2(n14700), .A(n14697), .B(n14731), .ZN(
        n14712) );
  INV_X1 U18124 ( .A(n14700), .ZN(n14699) );
  OAI21_X1 U18125 ( .B1(n14712), .B2(n14699), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14706) );
  NAND3_X1 U18126 ( .A1(n14706), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14700), .ZN(n14701) );
  OAI211_X1 U18127 ( .C1(n9563), .C2(n16070), .A(n14702), .B(n14701), .ZN(
        P1_U3000) );
  AOI21_X1 U18128 ( .B1(n14704), .B2(n20067), .A(n14703), .ZN(n14709) );
  INV_X1 U18129 ( .A(n14705), .ZN(n14707) );
  OAI21_X1 U18130 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14707), .A(
        n14706), .ZN(n14708) );
  OAI211_X1 U18131 ( .C1(n14710), .C2(n16070), .A(n14709), .B(n14708), .ZN(
        P1_U3001) );
  AOI21_X1 U18132 ( .B1(n14719), .B2(n11633), .A(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14711) );
  NOR2_X1 U18133 ( .A1(n14712), .A2(n14711), .ZN(n14713) );
  AOI211_X1 U18134 ( .C1(n20067), .C2(n14715), .A(n14714), .B(n14713), .ZN(
        n14716) );
  OAI21_X1 U18135 ( .B1(n14717), .B2(n16070), .A(n14716), .ZN(P1_U3002) );
  INV_X1 U18136 ( .A(n14718), .ZN(n14722) );
  INV_X1 U18137 ( .A(n14719), .ZN(n14727) );
  NOR3_X1 U18138 ( .A1(n14727), .A2(n11633), .A3(n14720), .ZN(n14721) );
  AOI211_X1 U18139 ( .C1(n14723), .C2(n20067), .A(n14722), .B(n14721), .ZN(
        n14725) );
  NAND2_X1 U18140 ( .A1(n14731), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14724) );
  OAI211_X1 U18141 ( .C1(n14726), .C2(n16070), .A(n14725), .B(n14724), .ZN(
        P1_U3003) );
  NOR2_X1 U18142 ( .A1(n14727), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14728) );
  AOI211_X1 U18143 ( .C1(n14730), .C2(n20067), .A(n14729), .B(n14728), .ZN(
        n14733) );
  NAND2_X1 U18144 ( .A1(n14731), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14732) );
  OAI211_X1 U18145 ( .C1(n14734), .C2(n16070), .A(n14733), .B(n14732), .ZN(
        P1_U3004) );
  INV_X1 U18146 ( .A(n14735), .ZN(n14738) );
  NOR3_X1 U18147 ( .A1(n16048), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14736), .ZN(n14737) );
  AOI211_X1 U18148 ( .C1(n14739), .C2(n20067), .A(n14738), .B(n14737), .ZN(
        n14745) );
  INV_X1 U18149 ( .A(n14740), .ZN(n14750) );
  NAND2_X1 U18150 ( .A1(n14742), .A2(n14741), .ZN(n14743) );
  NOR2_X1 U18151 ( .A1(n16048), .A2(n14743), .ZN(n14749) );
  OAI21_X1 U18152 ( .B1(n14750), .B2(n14749), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14744) );
  OAI211_X1 U18153 ( .C1(n14746), .C2(n16070), .A(n14745), .B(n14744), .ZN(
        P1_U3005) );
  OAI21_X1 U18154 ( .B1(n15838), .B2(n16069), .A(n14747), .ZN(n14748) );
  AOI211_X1 U18155 ( .C1(n14750), .C2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n14749), .B(n14748), .ZN(n14751) );
  OAI21_X1 U18156 ( .B1(n14752), .B2(n16070), .A(n14751), .ZN(P1_U3006) );
  INV_X1 U18157 ( .A(n16117), .ZN(n14754) );
  OAI21_X1 U18158 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14754), .A(
        n14753), .ZN(n14760) );
  NOR3_X1 U18159 ( .A1(n16048), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n16047), .ZN(n14759) );
  INV_X1 U18160 ( .A(n14755), .ZN(n14757) );
  OAI21_X1 U18161 ( .B1(n14757), .B2(n16069), .A(n14756), .ZN(n14758) );
  AOI211_X1 U18162 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n14760), .A(
        n14759), .B(n14758), .ZN(n14761) );
  OAI21_X1 U18163 ( .B1(n14762), .B2(n16070), .A(n14761), .ZN(P1_U3007) );
  INV_X1 U18164 ( .A(n16050), .ZN(n14771) );
  NOR2_X1 U18165 ( .A1(n15809), .A2(n14767), .ZN(n14765) );
  NAND2_X1 U18166 ( .A1(n16013), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14763) );
  NAND2_X1 U18167 ( .A1(n15809), .A2(n14763), .ZN(n14774) );
  NOR3_X1 U18168 ( .A1(n14774), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14764) );
  MUX2_X1 U18169 ( .A(n14765), .B(n14764), .S(n16013), .Z(n14766) );
  XNOR2_X1 U18170 ( .A(n14766), .B(n14772), .ZN(n15972) );
  NAND2_X1 U18171 ( .A1(n15972), .A2(n20071), .ZN(n14770) );
  NOR3_X1 U18172 ( .A1(n16100), .A2(n14775), .A3(n14767), .ZN(n16054) );
  OAI22_X1 U18173 ( .A1(n15861), .A2(n16069), .B1(n16041), .B2(n20723), .ZN(
        n14768) );
  AOI21_X1 U18174 ( .B1(n16054), .B2(n14772), .A(n14768), .ZN(n14769) );
  OAI211_X1 U18175 ( .C1(n14772), .C2(n14771), .A(n14770), .B(n14769), .ZN(
        P1_U3010) );
  XNOR2_X1 U18176 ( .A(n15965), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14773) );
  XNOR2_X1 U18177 ( .A(n14774), .B(n14773), .ZN(n15984) );
  NOR2_X1 U18178 ( .A1(n16100), .A2(n14775), .ZN(n15814) );
  OAI22_X1 U18179 ( .A1(n15879), .A2(n16069), .B1(n20720), .B2(n16041), .ZN(
        n14776) );
  AOI21_X1 U18180 ( .B1(n15814), .B2(n15806), .A(n14776), .ZN(n14778) );
  OR2_X1 U18181 ( .A1(n15821), .A2(n15806), .ZN(n14777) );
  OAI211_X1 U18182 ( .C1(n15984), .C2(n16070), .A(n14778), .B(n14777), .ZN(
        P1_U3012) );
  INV_X1 U18183 ( .A(n14779), .ZN(n14780) );
  NOR2_X1 U18184 ( .A1(n14781), .A2(n14780), .ZN(n14785) );
  NAND2_X1 U18185 ( .A1(n14783), .A2(n14782), .ZN(n14784) );
  XNOR2_X1 U18186 ( .A(n14785), .B(n14784), .ZN(n16004) );
  OAI21_X1 U18187 ( .B1(n14643), .B2(n14786), .A(n14805), .ZN(n14787) );
  OAI211_X1 U18188 ( .C1(n16086), .C2(n14810), .A(n14788), .B(n14787), .ZN(
        n16096) );
  AOI21_X1 U18189 ( .B1(n16085), .B2(n16121), .A(n16096), .ZN(n16084) );
  AND2_X1 U18190 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16061), .ZN(
        n16078) );
  NAND2_X1 U18191 ( .A1(n16077), .A2(n16078), .ZN(n14789) );
  OAI21_X1 U18192 ( .B1(n16077), .B2(n16084), .A(n14789), .ZN(n14791) );
  NOR2_X1 U18193 ( .A1(n15904), .A2(n16069), .ZN(n14790) );
  AOI211_X1 U18194 ( .C1(n16139), .C2(P1_REIP_REG_15__SCAN_IN), .A(n14791), 
        .B(n14790), .ZN(n14792) );
  OAI21_X1 U18195 ( .B1(n16004), .B2(n16070), .A(n14792), .ZN(P1_U3016) );
  OAI21_X1 U18196 ( .B1(n14795), .B2(n14794), .A(n14793), .ZN(n14796) );
  INV_X1 U18197 ( .A(n14796), .ZN(n16010) );
  INV_X1 U18198 ( .A(n15930), .ZN(n14799) );
  INV_X1 U18199 ( .A(n14797), .ZN(n14798) );
  OAI21_X1 U18200 ( .B1(n15931), .B2(n14799), .A(n14798), .ZN(n14801) );
  AND2_X1 U18201 ( .A1(n14801), .A2(n14800), .ZN(n15952) );
  NOR2_X1 U18202 ( .A1(n16041), .A2(n14802), .ZN(n14816) );
  INV_X1 U18203 ( .A(n14811), .ZN(n14803) );
  NOR2_X1 U18204 ( .A1(n14803), .A2(n16144), .ZN(n14814) );
  NOR2_X1 U18205 ( .A1(n14806), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16101) );
  INV_X1 U18206 ( .A(n14804), .ZN(n14809) );
  OAI21_X1 U18207 ( .B1(n14807), .B2(n14806), .A(n14805), .ZN(n14808) );
  OAI211_X1 U18208 ( .C1(n14811), .C2(n14810), .A(n14809), .B(n14808), .ZN(
        n16103) );
  AOI21_X1 U18209 ( .B1(n16117), .B2(n16101), .A(n16103), .ZN(n14812) );
  INV_X1 U18210 ( .A(n14812), .ZN(n14813) );
  MUX2_X1 U18211 ( .A(n14814), .B(n14813), .S(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n14815) );
  AOI211_X1 U18212 ( .C1(n20067), .C2(n15952), .A(n14816), .B(n14815), .ZN(
        n14817) );
  OAI21_X1 U18213 ( .B1(n16010), .B2(n16070), .A(n14817), .ZN(P1_U3019) );
  NAND2_X1 U18214 ( .A1(n20172), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20477) );
  OAI211_X1 U18215 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20172), .A(n20477), 
        .B(n20481), .ZN(n14818) );
  OAI21_X1 U18216 ( .B1(n14827), .B2(n20372), .A(n14818), .ZN(n14819) );
  MUX2_X1 U18217 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14819), .S(
        n20077), .Z(P1_U3477) );
  XOR2_X1 U18218 ( .A(n20477), .B(n9587), .Z(n14820) );
  OAI22_X1 U18219 ( .A1(n14820), .A2(n20620), .B1(n13572), .B2(n14827), .ZN(
        n14821) );
  MUX2_X1 U18220 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14821), .S(
        n20077), .Z(P1_U3476) );
  NOR2_X1 U18221 ( .A1(n20483), .A2(n20777), .ZN(n14823) );
  OAI22_X1 U18222 ( .A1(n14823), .A2(n11720), .B1(n20477), .B2(n20348), .ZN(
        n14824) );
  NAND2_X1 U18223 ( .A1(n14824), .A2(n20481), .ZN(n14826) );
  NOR3_X1 U18224 ( .A1(n20172), .A2(n20620), .A3(n20777), .ZN(n20146) );
  NAND2_X1 U18225 ( .A1(n20564), .A2(n20146), .ZN(n20540) );
  OAI211_X1 U18226 ( .C1(n14828), .C2(n14827), .A(n14826), .B(n20540), .ZN(
        n14829) );
  MUX2_X1 U18227 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n14829), .S(
        n20077), .Z(P1_U3475) );
  INV_X1 U18228 ( .A(n14833), .ZN(n14841) );
  INV_X1 U18229 ( .A(n14831), .ZN(n14836) );
  AOI22_X1 U18230 ( .A1(n14834), .A2(n11357), .B1(n14833), .B2(n14832), .ZN(
        n14835) );
  OAI21_X1 U18231 ( .B1(n20372), .B2(n14836), .A(n14835), .ZN(n15761) );
  NOR2_X1 U18232 ( .A1(n20677), .A2(n14837), .ZN(n14845) );
  INV_X1 U18233 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14839) );
  OAI22_X1 U18234 ( .A1(n14839), .A2(n14838), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14843) );
  AOI22_X1 U18235 ( .A1(n15761), .A2(n16146), .B1(n14845), .B2(n14843), .ZN(
        n14840) );
  OAI21_X1 U18236 ( .B1(n14849), .B2(n14841), .A(n14840), .ZN(n14842) );
  MUX2_X1 U18237 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14842), .S(
        n16151), .Z(P1_U3473) );
  INV_X1 U18238 ( .A(n14843), .ZN(n14844) );
  AOI22_X1 U18239 ( .A1(n14846), .A2(n16146), .B1(n14845), .B2(n14844), .ZN(
        n14847) );
  OAI21_X1 U18240 ( .B1(n14849), .B2(n14848), .A(n14847), .ZN(n14850) );
  MUX2_X1 U18241 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14850), .S(
        n16151), .Z(P1_U3472) );
  NAND2_X1 U18242 ( .A1(n13017), .A2(n19002), .ZN(n19036) );
  AOI22_X1 U18243 ( .A1(n19025), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19041), .ZN(n14852) );
  NAND2_X1 U18244 ( .A1(n19031), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14851) );
  OAI211_X1 U18245 ( .C1(n19045), .C2(n19006), .A(n14852), .B(n14851), .ZN(
        n14853) );
  AOI21_X1 U18246 ( .B1(n14854), .B2(n19030), .A(n14853), .ZN(n14856) );
  NAND2_X1 U18247 ( .A1(n14262), .A2(n19022), .ZN(n14855) );
  OAI211_X1 U18248 ( .C1(n14857), .C2(n19036), .A(n14856), .B(n14855), .ZN(
        P2_U2824) );
  XNOR2_X1 U18249 ( .A(n14869), .B(n14858), .ZN(n15259) );
  OR2_X1 U18250 ( .A1(n14872), .A2(n14859), .ZN(n14860) );
  NAND2_X1 U18251 ( .A1(n11113), .A2(n14860), .ZN(n15258) );
  AOI22_X1 U18252 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n19025), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19031), .ZN(n14863) );
  AOI22_X1 U18253 ( .A1(n14861), .A2(n19030), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19041), .ZN(n14862) );
  OAI211_X1 U18254 ( .C1(n15258), .C2(n19006), .A(n14863), .B(n14862), .ZN(
        n14867) );
  AOI211_X1 U18255 ( .C1(n15102), .C2(n14865), .A(n14864), .B(n19720), .ZN(
        n14866) );
  NOR2_X1 U18256 ( .A1(n14867), .A2(n14866), .ZN(n14868) );
  OAI21_X1 U18257 ( .B1(n15259), .B2(n19011), .A(n14868), .ZN(P2_U2826) );
  AOI21_X1 U18258 ( .B1(n14871), .B2(n14870), .A(n14869), .ZN(n15266) );
  AOI21_X1 U18259 ( .B1(n14874), .B2(n14873), .A(n14872), .ZN(n15270) );
  NAND2_X1 U18260 ( .A1(n19031), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n14876) );
  NAND2_X1 U18261 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19041), .ZN(
        n14875) );
  OAI211_X1 U18262 ( .C1(n19009), .C2(n14877), .A(n14876), .B(n14875), .ZN(
        n14878) );
  AOI21_X1 U18263 ( .B1(n15270), .B2(n19027), .A(n14878), .ZN(n14879) );
  OAI21_X1 U18264 ( .B1(n14880), .B2(n19008), .A(n14879), .ZN(n14885) );
  AOI211_X1 U18265 ( .C1(n14883), .C2(n14882), .A(n14881), .B(n19720), .ZN(
        n14884) );
  AOI211_X1 U18266 ( .C1(n19022), .C2(n15266), .A(n14885), .B(n14884), .ZN(
        n14886) );
  INV_X1 U18267 ( .A(n14886), .ZN(P2_U2827) );
  AOI211_X1 U18268 ( .C1(n14889), .C2(n14888), .A(n14887), .B(n19720), .ZN(
        n14890) );
  INV_X1 U18269 ( .A(n14890), .ZN(n14897) );
  NAND2_X1 U18270 ( .A1(n19027), .A2(n15060), .ZN(n14892) );
  AOI22_X1 U18271 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n19025), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19031), .ZN(n14891) );
  OAI211_X1 U18272 ( .C1(n18991), .C2(n14893), .A(n14892), .B(n14891), .ZN(
        n14894) );
  AOI21_X1 U18273 ( .B1(n14895), .B2(n19022), .A(n14894), .ZN(n14896) );
  OAI211_X1 U18274 ( .C1(n19008), .C2(n14898), .A(n14897), .B(n14896), .ZN(
        P2_U2830) );
  INV_X1 U18275 ( .A(n14899), .ZN(n14900) );
  AOI21_X1 U18276 ( .B1(n14902), .B2(n14901), .A(n14900), .ZN(n15148) );
  INV_X1 U18277 ( .A(n15148), .ZN(n15306) );
  NOR2_X1 U18278 ( .A1(n13039), .A2(n14903), .ZN(n14904) );
  OR2_X1 U18279 ( .A1(n14905), .A2(n14904), .ZN(n15064) );
  AOI22_X1 U18280 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n19025), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19031), .ZN(n14909) );
  OAI22_X1 U18281 ( .A1(n14906), .A2(n19008), .B1(n18991), .B2(n9966), .ZN(
        n14907) );
  INV_X1 U18282 ( .A(n14907), .ZN(n14908) );
  OAI211_X1 U18283 ( .C1(n15064), .C2(n19006), .A(n14909), .B(n14908), .ZN(
        n14913) );
  AOI211_X1 U18284 ( .C1(n14911), .C2(n9971), .A(n14910), .B(n19720), .ZN(
        n14912) );
  NOR2_X1 U18285 ( .A1(n14913), .A2(n14912), .ZN(n14914) );
  OAI21_X1 U18286 ( .B1(n15306), .B2(n19011), .A(n14914), .ZN(P2_U2831) );
  NOR2_X1 U18287 ( .A1(n14916), .A2(n14915), .ZN(n14917) );
  OR2_X1 U18288 ( .A1(n15079), .A2(n14917), .ZN(n16179) );
  INV_X1 U18289 ( .A(n16179), .ZN(n14918) );
  NAND2_X1 U18290 ( .A1(n14918), .A2(n19027), .ZN(n14931) );
  INV_X1 U18291 ( .A(n15164), .ZN(n14919) );
  INV_X1 U18292 ( .A(n18881), .ZN(n19040) );
  AOI22_X1 U18293 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19041), .B1(
        n14919), .B2(n19040), .ZN(n14930) );
  OAI211_X1 U18294 ( .C1(n14920), .C2(n15164), .A(n19002), .B(n18855), .ZN(
        n14929) );
  AND2_X1 U18295 ( .A1(n15013), .A2(n14921), .ZN(n14923) );
  OR2_X1 U18296 ( .A1(n14923), .A2(n14922), .ZN(n15361) );
  NAND2_X1 U18297 ( .A1(n19031), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n14925) );
  NAND2_X1 U18298 ( .A1(n19025), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n14924) );
  OAI211_X1 U18299 ( .C1(n15361), .C2(n19011), .A(n14925), .B(n14924), .ZN(
        n14926) );
  AOI21_X1 U18300 ( .B1(n14927), .B2(n19030), .A(n14926), .ZN(n14928) );
  NAND4_X1 U18301 ( .A1(n14931), .A2(n14930), .A3(n14929), .A4(n14928), .ZN(
        P2_U2835) );
  INV_X1 U18302 ( .A(n14932), .ZN(n14933) );
  AOI21_X1 U18303 ( .B1(n14934), .B2(n13965), .A(n14933), .ZN(n16186) );
  INV_X1 U18304 ( .A(n16186), .ZN(n14948) );
  INV_X1 U18305 ( .A(n14935), .ZN(n14946) );
  OR2_X1 U18306 ( .A1(n15026), .A2(n14936), .ZN(n14937) );
  AND2_X1 U18307 ( .A1(n15011), .A2(n14937), .ZN(n15389) );
  INV_X1 U18308 ( .A(n15389), .ZN(n15021) );
  INV_X1 U18309 ( .A(n15185), .ZN(n14938) );
  OAI211_X1 U18310 ( .C1(n14939), .C2(n13016), .A(n14938), .B(n19002), .ZN(
        n14944) );
  NOR2_X1 U18311 ( .A1(n14939), .A2(n19036), .ZN(n18886) );
  AOI22_X1 U18312 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19041), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19031), .ZN(n14940) );
  OAI211_X1 U18313 ( .C1(n19009), .C2(n14941), .A(n14940), .B(n16264), .ZN(
        n14942) );
  AOI21_X1 U18314 ( .B1(n15185), .B2(n18886), .A(n14942), .ZN(n14943) );
  OAI211_X1 U18315 ( .C1(n19011), .C2(n15021), .A(n14944), .B(n14943), .ZN(
        n14945) );
  AOI21_X1 U18316 ( .B1(n14946), .B2(n19030), .A(n14945), .ZN(n14947) );
  OAI21_X1 U18317 ( .B1(n14948), .B2(n19006), .A(n14947), .ZN(P2_U2837) );
  MUX2_X1 U18318 ( .A(n14262), .B(P2_EBX_REG_31__SCAN_IN), .S(n15022), .Z(
        P2_U2856) );
  OR2_X1 U18319 ( .A1(n14950), .A2(n14949), .ZN(n15032) );
  NAND3_X1 U18320 ( .A1(n15032), .A2(n14951), .A3(n15018), .ZN(n14953) );
  NAND2_X1 U18321 ( .A1(n15022), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14952) );
  OAI211_X1 U18322 ( .C1(n15259), .C2(n15022), .A(n14953), .B(n14952), .ZN(
        P2_U2858) );
  NAND2_X1 U18323 ( .A1(n10017), .A2(n14954), .ZN(n14956) );
  XNOR2_X1 U18324 ( .A(n14956), .B(n14955), .ZN(n15043) );
  NAND2_X1 U18325 ( .A1(n15022), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n14958) );
  NAND2_X1 U18326 ( .A1(n15266), .A2(n15027), .ZN(n14957) );
  OAI211_X1 U18327 ( .C1(n15043), .C2(n15030), .A(n14958), .B(n14957), .ZN(
        P2_U2859) );
  OAI21_X1 U18328 ( .B1(n14961), .B2(n14960), .A(n14959), .ZN(n15048) );
  NOR2_X1 U18329 ( .A1(n15283), .A2(n15022), .ZN(n14962) );
  AOI21_X1 U18330 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n15022), .A(n14962), .ZN(
        n14963) );
  OAI21_X1 U18331 ( .B1(n15048), .B2(n15030), .A(n14963), .ZN(P2_U2860) );
  OR2_X1 U18332 ( .A1(n14965), .A2(n14964), .ZN(n14966) );
  NAND2_X1 U18333 ( .A1(n14967), .A2(n14966), .ZN(n16167) );
  AOI21_X1 U18334 ( .B1(n14970), .B2(n14969), .A(n14968), .ZN(n15049) );
  NAND2_X1 U18335 ( .A1(n15049), .A2(n15018), .ZN(n14972) );
  NAND2_X1 U18336 ( .A1(n15022), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14971) );
  OAI211_X1 U18337 ( .C1(n16167), .C2(n15022), .A(n14972), .B(n14971), .ZN(
        P2_U2861) );
  OAI21_X1 U18338 ( .B1(n14975), .B2(n14974), .A(n14973), .ZN(n15063) );
  MUX2_X1 U18339 ( .A(n14977), .B(n14976), .S(n15022), .Z(n14978) );
  OAI21_X1 U18340 ( .B1(n15063), .B2(n15030), .A(n14978), .ZN(P2_U2862) );
  AOI21_X1 U18341 ( .B1(n9668), .B2(n14980), .A(n14979), .ZN(n14981) );
  XOR2_X1 U18342 ( .A(n14982), .B(n14981), .Z(n15069) );
  NOR2_X1 U18343 ( .A1(n15027), .A2(n14983), .ZN(n14984) );
  AOI21_X1 U18344 ( .B1(n15148), .B2(n15027), .A(n14984), .ZN(n14985) );
  OAI21_X1 U18345 ( .B1(n15069), .B2(n15030), .A(n14985), .ZN(P2_U2863) );
  AOI21_X1 U18346 ( .B1(n14988), .B2(n14987), .A(n14986), .ZN(n15070) );
  NAND2_X1 U18347 ( .A1(n15070), .A2(n15018), .ZN(n14991) );
  INV_X1 U18348 ( .A(n15321), .ZN(n14989) );
  NAND2_X1 U18349 ( .A1(n14989), .A2(n15027), .ZN(n14990) );
  OAI211_X1 U18350 ( .C1(n15027), .C2(n10839), .A(n14991), .B(n14990), .ZN(
        P2_U2864) );
  OR2_X1 U18351 ( .A1(n12633), .A2(n14992), .ZN(n14993) );
  AND2_X1 U18352 ( .A1(n14994), .A2(n14993), .ZN(n16191) );
  INV_X1 U18353 ( .A(n16191), .ZN(n14999) );
  AOI21_X1 U18354 ( .B1(n14996), .B2(n15003), .A(n14995), .ZN(n16174) );
  NAND2_X1 U18355 ( .A1(n16174), .A2(n15018), .ZN(n14998) );
  NAND2_X1 U18356 ( .A1(n15022), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14997) );
  OAI211_X1 U18357 ( .C1(n14999), .C2(n15022), .A(n14998), .B(n14997), .ZN(
        P2_U2865) );
  NAND2_X1 U18358 ( .A1(n15000), .A2(n15001), .ZN(n15002) );
  NAND2_X1 U18359 ( .A1(n15003), .A2(n15002), .ZN(n15085) );
  MUX2_X1 U18360 ( .A(n18862), .B(n18859), .S(n15022), .Z(n15004) );
  OAI21_X1 U18361 ( .B1(n15085), .B2(n15030), .A(n15004), .ZN(P2_U2866) );
  OR2_X1 U18362 ( .A1(n15006), .A2(n15005), .ZN(n15007) );
  NAND2_X1 U18363 ( .A1(n15000), .A2(n15007), .ZN(n16178) );
  NOR2_X1 U18364 ( .A1(n15361), .A2(n15022), .ZN(n15008) );
  AOI21_X1 U18365 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(n15022), .A(n15008), .ZN(
        n15009) );
  OAI21_X1 U18366 ( .B1(n16178), .B2(n15030), .A(n15009), .ZN(P2_U2867) );
  NAND2_X1 U18367 ( .A1(n15011), .A2(n15010), .ZN(n15012) );
  NAND2_X1 U18368 ( .A1(n15013), .A2(n15012), .ZN(n18874) );
  NAND2_X1 U18369 ( .A1(n15014), .A2(n15018), .ZN(n15016) );
  NAND2_X1 U18370 ( .A1(n15022), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15015) );
  OAI211_X1 U18371 ( .C1(n18874), .C2(n15022), .A(n15016), .B(n15015), .ZN(
        P2_U2868) );
  AOI21_X1 U18372 ( .B1(n15017), .B2(n13963), .A(n14018), .ZN(n16185) );
  NAND2_X1 U18373 ( .A1(n16185), .A2(n15018), .ZN(n15020) );
  NAND2_X1 U18374 ( .A1(n15022), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n15019) );
  OAI211_X1 U18375 ( .C1(n15021), .C2(n15022), .A(n15020), .B(n15019), .ZN(
        P2_U2869) );
  NAND2_X1 U18376 ( .A1(n15022), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15029) );
  AND2_X1 U18377 ( .A1(n15024), .A2(n15023), .ZN(n15025) );
  NOR2_X1 U18378 ( .A1(n15026), .A2(n15025), .ZN(n18884) );
  NAND2_X1 U18379 ( .A1(n18884), .A2(n15027), .ZN(n15028) );
  OAI211_X1 U18380 ( .C1(n15031), .C2(n15030), .A(n15029), .B(n15028), .ZN(
        P2_U2870) );
  NAND3_X1 U18381 ( .A1(n15032), .A2(n14951), .A3(n19100), .ZN(n15038) );
  INV_X1 U18382 ( .A(n15258), .ZN(n15035) );
  OAI22_X1 U18383 ( .A1(n15065), .A2(n19066), .B1(n19083), .B2(n15033), .ZN(
        n15034) );
  AOI21_X1 U18384 ( .B1(n19111), .B2(n15035), .A(n15034), .ZN(n15037) );
  AOI22_X1 U18385 ( .A1(n19052), .A2(BUF2_REG_29__SCAN_IN), .B1(n19051), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n15036) );
  NAND3_X1 U18386 ( .A1(n15038), .A2(n15037), .A3(n15036), .ZN(P2_U2890) );
  INV_X1 U18387 ( .A(n19069), .ZN(n15039) );
  OAI22_X1 U18388 ( .A1(n15065), .A2(n15039), .B1(n19083), .B2(n20883), .ZN(
        n15040) );
  AOI21_X1 U18389 ( .B1(n19111), .B2(n15270), .A(n15040), .ZN(n15042) );
  AOI22_X1 U18390 ( .A1(n19052), .A2(BUF2_REG_28__SCAN_IN), .B1(n19051), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15041) );
  OAI211_X1 U18391 ( .C1(n15043), .C2(n19115), .A(n15042), .B(n15041), .ZN(
        P2_U2891) );
  OAI22_X1 U18392 ( .A1(n15065), .A2(n19072), .B1(n19083), .B2(n15044), .ZN(
        n15045) );
  AOI21_X1 U18393 ( .B1(n19111), .B2(n15280), .A(n15045), .ZN(n15047) );
  AOI22_X1 U18394 ( .A1(n19052), .A2(BUF2_REG_27__SCAN_IN), .B1(n19051), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15046) );
  OAI211_X1 U18395 ( .C1(n15048), .C2(n19115), .A(n15047), .B(n15046), .ZN(
        P2_U2892) );
  NAND2_X1 U18396 ( .A1(n15049), .A2(n19100), .ZN(n15057) );
  AOI22_X1 U18397 ( .A1(n19050), .A2(n19074), .B1(n19110), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15056) );
  AOI22_X1 U18398 ( .A1(n19052), .A2(BUF2_REG_26__SCAN_IN), .B1(n19051), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15055) );
  INV_X1 U18399 ( .A(n15050), .ZN(n15051) );
  AOI21_X1 U18400 ( .B1(n15053), .B2(n15052), .A(n15051), .ZN(n16170) );
  NAND2_X1 U18401 ( .A1(n19111), .A2(n16170), .ZN(n15054) );
  NAND4_X1 U18402 ( .A1(n15057), .A2(n15056), .A3(n15055), .A4(n15054), .ZN(
        P2_U2893) );
  OAI22_X1 U18403 ( .A1(n15065), .A2(n19077), .B1(n19083), .B2(n15058), .ZN(
        n15059) );
  AOI21_X1 U18404 ( .B1(n19111), .B2(n15060), .A(n15059), .ZN(n15062) );
  AOI22_X1 U18405 ( .A1(n19052), .A2(BUF2_REG_25__SCAN_IN), .B1(n19051), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15061) );
  OAI211_X1 U18406 ( .C1(n15063), .C2(n19115), .A(n15062), .B(n15061), .ZN(
        P2_U2894) );
  INV_X1 U18407 ( .A(n15064), .ZN(n15304) );
  OAI22_X1 U18408 ( .A1(n15065), .A2(n19080), .B1(n19083), .B2(n20823), .ZN(
        n15066) );
  AOI21_X1 U18409 ( .B1(n19111), .B2(n15304), .A(n15066), .ZN(n15068) );
  AOI22_X1 U18410 ( .A1(n19052), .A2(BUF2_REG_24__SCAN_IN), .B1(n19051), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15067) );
  OAI211_X1 U18411 ( .C1(n15069), .C2(n19115), .A(n15068), .B(n15067), .ZN(
        P2_U2895) );
  NAND2_X1 U18412 ( .A1(n15070), .A2(n19100), .ZN(n15075) );
  AOI22_X1 U18413 ( .A1(n19050), .A2(n15071), .B1(n19110), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n15074) );
  AOI22_X1 U18414 ( .A1(n19052), .A2(BUF2_REG_23__SCAN_IN), .B1(n19051), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n15073) );
  NAND2_X1 U18415 ( .A1(n19111), .A2(n15318), .ZN(n15072) );
  NAND4_X1 U18416 ( .A1(n15075), .A2(n15074), .A3(n15073), .A4(n15072), .ZN(
        P2_U2896) );
  NAND2_X1 U18417 ( .A1(n19052), .A2(BUF2_REG_21__SCAN_IN), .ZN(n15077) );
  AOI22_X1 U18418 ( .A1(n19050), .A2(n19086), .B1(n19110), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15076) );
  NAND2_X1 U18419 ( .A1(n15077), .A2(n15076), .ZN(n15083) );
  OR2_X1 U18420 ( .A1(n15079), .A2(n15078), .ZN(n15081) );
  INV_X1 U18421 ( .A(n15334), .ZN(n15080) );
  NAND2_X1 U18422 ( .A1(n15081), .A2(n15080), .ZN(n18863) );
  NOR2_X1 U18423 ( .A1(n18863), .A2(n19054), .ZN(n15082) );
  AOI211_X1 U18424 ( .C1(BUF1_REG_21__SCAN_IN), .C2(n19051), .A(n15083), .B(
        n15082), .ZN(n15084) );
  OAI21_X1 U18425 ( .B1(n19115), .B2(n15085), .A(n15084), .ZN(P2_U2898) );
  AOI21_X1 U18426 ( .B1(n19166), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15086), .ZN(n15089) );
  NAND2_X1 U18427 ( .A1(n19175), .A2(n15087), .ZN(n15088) );
  OAI211_X1 U18428 ( .C1(n14202), .C2(n19179), .A(n15089), .B(n15088), .ZN(
        n15090) );
  AOI21_X1 U18429 ( .B1(n15091), .B2(n19169), .A(n15090), .ZN(n15092) );
  OAI21_X1 U18430 ( .B1(n15093), .B2(n16243), .A(n15092), .ZN(P2_U2984) );
  NOR2_X1 U18431 ( .A1(n15095), .A2(n15094), .ZN(n15097) );
  XOR2_X1 U18432 ( .A(n15097), .B(n15096), .Z(n15265) );
  AOI21_X1 U18433 ( .B1(n15099), .B2(n15116), .A(n15098), .ZN(n15262) );
  NAND2_X1 U18434 ( .A1(n19155), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15257) );
  OAI21_X1 U18435 ( .B1(n16259), .B2(n15100), .A(n15257), .ZN(n15101) );
  AOI21_X1 U18436 ( .B1(n19175), .B2(n15102), .A(n15101), .ZN(n15103) );
  OAI21_X1 U18437 ( .B1(n15259), .B2(n19179), .A(n15103), .ZN(n15104) );
  AOI21_X1 U18438 ( .B1(n15262), .B2(n19169), .A(n15104), .ZN(n15105) );
  OAI21_X1 U18439 ( .B1(n15265), .B2(n16243), .A(n15105), .ZN(P2_U2985) );
  NOR2_X1 U18440 ( .A1(n15107), .A2(n15106), .ZN(n15108) );
  XNOR2_X1 U18441 ( .A(n15108), .B(n15110), .ZN(n15120) );
  INV_X1 U18442 ( .A(n15108), .ZN(n15109) );
  AOI22_X1 U18443 ( .A1(n15120), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n15110), .B2(n15109), .ZN(n15113) );
  XNOR2_X1 U18444 ( .A(n15111), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15112) );
  XNOR2_X1 U18445 ( .A(n15113), .B(n15112), .ZN(n15276) );
  NAND2_X1 U18446 ( .A1(n19155), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15267) );
  NAND2_X1 U18447 ( .A1(n19166), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15114) );
  OAI211_X1 U18448 ( .C1(n19165), .C2(n15115), .A(n15267), .B(n15114), .ZN(
        n15118) );
  NOR2_X1 U18449 ( .A1(n15273), .A2(n16245), .ZN(n15117) );
  OAI21_X1 U18450 ( .B1(n15276), .B2(n16243), .A(n15119), .ZN(P2_U2986) );
  XNOR2_X1 U18451 ( .A(n15120), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15287) );
  AOI21_X1 U18452 ( .B1(n15253), .B2(n15134), .A(n15121), .ZN(n15285) );
  INV_X1 U18453 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19786) );
  NOR2_X1 U18454 ( .A1(n16264), .A2(n19786), .ZN(n15278) );
  AOI21_X1 U18455 ( .B1(n19166), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15278), .ZN(n15124) );
  NAND2_X1 U18456 ( .A1(n19175), .A2(n15122), .ZN(n15123) );
  OAI211_X1 U18457 ( .C1(n15283), .C2(n19179), .A(n15124), .B(n15123), .ZN(
        n15125) );
  AOI21_X1 U18458 ( .B1(n15285), .B2(n19169), .A(n15125), .ZN(n15126) );
  OAI21_X1 U18459 ( .B1(n15287), .B2(n16243), .A(n15126), .ZN(P2_U2987) );
  AOI21_X1 U18460 ( .B1(n15129), .B2(n15128), .A(n15127), .ZN(n15130) );
  XOR2_X1 U18461 ( .A(n15131), .B(n15130), .Z(n15301) );
  INV_X1 U18462 ( .A(n16167), .ZN(n15138) );
  INV_X1 U18463 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19783) );
  NOR2_X1 U18464 ( .A1(n16264), .A2(n19783), .ZN(n15294) );
  AOI21_X1 U18465 ( .B1(n19166), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15294), .ZN(n15132) );
  OAI21_X1 U18466 ( .B1(n19165), .B2(n15133), .A(n15132), .ZN(n15137) );
  OAI21_X1 U18467 ( .B1(n15135), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15134), .ZN(n15296) );
  NOR2_X1 U18468 ( .A1(n15296), .A2(n16245), .ZN(n15136) );
  AOI211_X1 U18469 ( .C1(n16248), .C2(n15138), .A(n15137), .B(n15136), .ZN(
        n15139) );
  OAI21_X1 U18470 ( .B1(n15301), .B2(n16243), .A(n15139), .ZN(P2_U2988) );
  XNOR2_X1 U18471 ( .A(n15140), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15141) );
  XNOR2_X1 U18472 ( .A(n15142), .B(n15141), .ZN(n15312) );
  INV_X1 U18473 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19779) );
  NOR2_X1 U18474 ( .A1(n16264), .A2(n19779), .ZN(n15302) );
  AOI21_X1 U18475 ( .B1(n19166), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15302), .ZN(n15143) );
  OAI21_X1 U18476 ( .B1(n19165), .B2(n15144), .A(n15143), .ZN(n15147) );
  OR2_X1 U18477 ( .A1(n15152), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15145) );
  NAND2_X1 U18478 ( .A1(n14219), .A2(n15145), .ZN(n15307) );
  NOR2_X1 U18479 ( .A1(n15307), .A2(n16245), .ZN(n15146) );
  AOI211_X1 U18480 ( .C1(n16248), .C2(n15148), .A(n15147), .B(n15146), .ZN(
        n15149) );
  OAI21_X1 U18481 ( .B1(n15312), .B2(n16243), .A(n15149), .ZN(P2_U2990) );
  XNOR2_X1 U18482 ( .A(n15151), .B(n15150), .ZN(n15325) );
  AOI21_X1 U18483 ( .B1(n15315), .B2(n15331), .A(n15152), .ZN(n15323) );
  NOR2_X1 U18484 ( .A1(n16264), .A2(n19777), .ZN(n15317) );
  AOI21_X1 U18485 ( .B1(n19166), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15317), .ZN(n15155) );
  NAND2_X1 U18486 ( .A1(n19175), .A2(n15153), .ZN(n15154) );
  OAI211_X1 U18487 ( .C1(n15321), .C2(n19179), .A(n15155), .B(n15154), .ZN(
        n15156) );
  AOI21_X1 U18488 ( .B1(n15323), .B2(n19169), .A(n15156), .ZN(n15157) );
  OAI21_X1 U18489 ( .B1(n15325), .B2(n16243), .A(n15157), .ZN(P2_U2991) );
  INV_X1 U18490 ( .A(n15158), .ZN(n15159) );
  NOR2_X1 U18491 ( .A1(n15160), .A2(n15159), .ZN(n15161) );
  XNOR2_X1 U18492 ( .A(n15162), .B(n15161), .ZN(n15373) );
  AOI21_X1 U18493 ( .B1(n15364), .B2(n15169), .A(n15163), .ZN(n15371) );
  INV_X1 U18494 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19772) );
  NOR2_X1 U18495 ( .A1(n16264), .A2(n19772), .ZN(n15363) );
  NOR2_X1 U18496 ( .A1(n19165), .A2(n15164), .ZN(n15165) );
  AOI211_X1 U18497 ( .C1(n19166), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15363), .B(n15165), .ZN(n15166) );
  OAI21_X1 U18498 ( .B1(n19179), .B2(n15361), .A(n15166), .ZN(n15167) );
  AOI21_X1 U18499 ( .B1(n15371), .B2(n19169), .A(n15167), .ZN(n15168) );
  OAI21_X1 U18500 ( .B1(n15373), .B2(n16243), .A(n15168), .ZN(P2_U2994) );
  OAI21_X1 U18501 ( .B1(n15181), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15169), .ZN(n15383) );
  NAND2_X1 U18502 ( .A1(n19155), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15376) );
  OAI21_X1 U18503 ( .B1(n16259), .B2(n15172), .A(n15376), .ZN(n15174) );
  NOR2_X1 U18504 ( .A1(n19179), .A2(n18874), .ZN(n15173) );
  AOI211_X1 U18505 ( .C1(n19175), .C2(n18870), .A(n15174), .B(n15173), .ZN(
        n15175) );
  OAI211_X1 U18506 ( .C1(n16245), .C2(n15383), .A(n15176), .B(n15175), .ZN(
        P2_U2995) );
  NAND2_X1 U18507 ( .A1(n9767), .A2(n15178), .ZN(n15179) );
  XNOR2_X1 U18508 ( .A(n15180), .B(n15179), .ZN(n15397) );
  NAND2_X1 U18509 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15402) );
  AOI21_X1 U18510 ( .B1(n15201), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15182) );
  NOR2_X1 U18511 ( .A1(n15182), .A2(n15181), .ZN(n15395) );
  INV_X1 U18512 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19769) );
  NOR2_X1 U18513 ( .A1(n16264), .A2(n19769), .ZN(n15388) );
  AOI21_X1 U18514 ( .B1(n19166), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15388), .ZN(n15184) );
  NAND2_X1 U18515 ( .A1(n16248), .A2(n15389), .ZN(n15183) );
  OAI211_X1 U18516 ( .C1(n19165), .C2(n15185), .A(n15184), .B(n15183), .ZN(
        n15186) );
  AOI21_X1 U18517 ( .B1(n15395), .B2(n19169), .A(n15186), .ZN(n15187) );
  OAI21_X1 U18518 ( .B1(n15397), .B2(n16243), .A(n15187), .ZN(P2_U2996) );
  XNOR2_X1 U18519 ( .A(n15201), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15195) );
  XNOR2_X1 U18520 ( .A(n15189), .B(n15188), .ZN(n15401) );
  NAND2_X1 U18521 ( .A1(n15401), .A2(n19167), .ZN(n15194) );
  INV_X1 U18522 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19767) );
  NOR2_X1 U18523 ( .A1(n19767), .A2(n16264), .ZN(n15192) );
  OAI22_X1 U18524 ( .A1(n16259), .A2(n15190), .B1(n19165), .B2(n18887), .ZN(
        n15191) );
  AOI211_X1 U18525 ( .C1(n16248), .C2(n18884), .A(n15192), .B(n15191), .ZN(
        n15193) );
  OAI211_X1 U18526 ( .C1(n16245), .C2(n15195), .A(n15194), .B(n15193), .ZN(
        P2_U2997) );
  XNOR2_X1 U18527 ( .A(n15197), .B(n15196), .ZN(n15420) );
  INV_X1 U18528 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19765) );
  NOR2_X1 U18529 ( .A1(n19765), .A2(n16264), .ZN(n15200) );
  INV_X1 U18530 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15198) );
  OAI22_X1 U18531 ( .A1(n16259), .A2(n15198), .B1(n19165), .B2(n18894), .ZN(
        n15199) );
  AOI211_X1 U18532 ( .C1(n16248), .C2(n18901), .A(n15200), .B(n15199), .ZN(
        n15204) );
  INV_X1 U18533 ( .A(n15201), .ZN(n15403) );
  OAI21_X1 U18534 ( .B1(n16198), .B2(n16267), .A(n20859), .ZN(n15202) );
  NAND3_X1 U18535 ( .A1(n15403), .A2(n19169), .A3(n15202), .ZN(n15203) );
  OAI211_X1 U18536 ( .C1(n15420), .C2(n16243), .A(n15204), .B(n15203), .ZN(
        P2_U2998) );
  NAND2_X1 U18537 ( .A1(n15206), .A2(n15205), .ZN(n15208) );
  XOR2_X1 U18538 ( .A(n15208), .B(n15207), .Z(n16275) );
  XNOR2_X1 U18539 ( .A(n16198), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16271) );
  INV_X1 U18540 ( .A(n15209), .ZN(n18908) );
  OAI22_X1 U18541 ( .A1(n16259), .A2(n15210), .B1(n19165), .B2(n18908), .ZN(
        n15213) );
  INV_X1 U18542 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n15211) );
  OAI22_X1 U18543 ( .A1(n19179), .A2(n18912), .B1(n15211), .B2(n18992), .ZN(
        n15212) );
  AOI211_X1 U18544 ( .C1(n16271), .C2(n19169), .A(n15213), .B(n15212), .ZN(
        n15214) );
  OAI21_X1 U18545 ( .B1(n16275), .B2(n16243), .A(n15214), .ZN(P2_U2999) );
  OAI21_X1 U18546 ( .B1(n15433), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n16196), .ZN(n15431) );
  NAND2_X1 U18547 ( .A1(n15216), .A2(n15215), .ZN(n15218) );
  XOR2_X1 U18548 ( .A(n15218), .B(n15217), .Z(n15421) );
  NAND2_X1 U18549 ( .A1(n15421), .A2(n19167), .ZN(n15223) );
  INV_X1 U18550 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n20796) );
  OAI22_X1 U18551 ( .A1(n16259), .A2(n18917), .B1(n20796), .B2(n18992), .ZN(
        n15221) );
  INV_X1 U18552 ( .A(n18923), .ZN(n15219) );
  NOR2_X1 U18553 ( .A1(n19165), .A2(n15219), .ZN(n15220) );
  AOI211_X1 U18554 ( .C1(n18924), .C2(n16248), .A(n15221), .B(n15220), .ZN(
        n15222) );
  OAI211_X1 U18555 ( .C1(n16245), .C2(n15431), .A(n15223), .B(n15222), .ZN(
        P2_U3001) );
  XNOR2_X1 U18556 ( .A(n15225), .B(n15224), .ZN(n15530) );
  NAND2_X1 U18557 ( .A1(n15227), .A2(n15226), .ZN(n15511) );
  NAND2_X1 U18558 ( .A1(n15508), .A2(n15510), .ZN(n15228) );
  XNOR2_X1 U18559 ( .A(n15511), .B(n15228), .ZN(n15528) );
  INV_X1 U18560 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19751) );
  OAI22_X1 U18561 ( .A1(n16259), .A2(n15229), .B1(n19751), .B2(n16264), .ZN(
        n15230) );
  AOI21_X1 U18562 ( .B1(n19175), .B2(n18972), .A(n15230), .ZN(n15231) );
  OAI21_X1 U18563 ( .B1(n19179), .B2(n18976), .A(n15231), .ZN(n15232) );
  AOI21_X1 U18564 ( .B1(n15528), .B2(n19167), .A(n15232), .ZN(n15233) );
  OAI21_X1 U18565 ( .B1(n15530), .B2(n16245), .A(n15233), .ZN(P2_U3007) );
  XNOR2_X1 U18566 ( .A(n15234), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15546) );
  INV_X1 U18567 ( .A(n15235), .ZN(n15236) );
  XNOR2_X1 U18568 ( .A(n15237), .B(n15236), .ZN(n15544) );
  INV_X1 U18569 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19749) );
  OAI22_X1 U18570 ( .A1(n19749), .A2(n18992), .B1(n19165), .B2(n18985), .ZN(
        n15239) );
  OAI22_X1 U18571 ( .A1(n19179), .A2(n18986), .B1(n16259), .B2(n9963), .ZN(
        n15238) );
  AOI211_X1 U18572 ( .C1(n15544), .C2(n19167), .A(n15239), .B(n15238), .ZN(
        n15240) );
  OAI21_X1 U18573 ( .B1(n15546), .B2(n16245), .A(n15240), .ZN(P2_U3008) );
  AOI22_X1 U18574 ( .A1(n15241), .A2(n19175), .B1(n16248), .B2(n15568), .ZN(
        n15251) );
  OAI21_X1 U18575 ( .B1(n15244), .B2(n15243), .A(n15242), .ZN(n15245) );
  XOR2_X1 U18576 ( .A(n15245), .B(n15248), .Z(n15570) );
  NOR2_X1 U18577 ( .A1(n18992), .A2(n19740), .ZN(n15567) );
  AOI21_X1 U18578 ( .B1(n19167), .B2(n15570), .A(n15567), .ZN(n15250) );
  AOI21_X1 U18579 ( .B1(n15248), .B2(n15247), .A(n15246), .ZN(n15569) );
  AOI22_X1 U18580 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19166), .B1(
        n19169), .B2(n15569), .ZN(n15249) );
  NAND3_X1 U18581 ( .A1(n15251), .A2(n15250), .A3(n15249), .ZN(P2_U3013) );
  NOR2_X1 U18582 ( .A1(n15252), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15279) );
  OR2_X1 U18583 ( .A1(n15277), .A2(n15279), .ZN(n15275) );
  INV_X1 U18584 ( .A(n15252), .ZN(n15255) );
  OAI21_X1 U18585 ( .B1(n15253), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15254) );
  OAI211_X1 U18586 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(n15255), .B(n15254), .ZN(
        n15256) );
  OAI211_X1 U18587 ( .C1(n16294), .C2(n15258), .A(n15257), .B(n15256), .ZN(
        n15261) );
  NOR2_X1 U18588 ( .A1(n15259), .A2(n16295), .ZN(n15260) );
  AOI211_X1 U18589 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15275), .A(
        n15261), .B(n15260), .ZN(n15264) );
  NAND2_X1 U18590 ( .A1(n15262), .A2(n16270), .ZN(n15263) );
  OAI211_X1 U18591 ( .C1(n15265), .C2(n16274), .A(n15264), .B(n15263), .ZN(
        P2_U3017) );
  INV_X1 U18592 ( .A(n15266), .ZN(n15272) );
  OAI21_X1 U18593 ( .B1(n15268), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15267), .ZN(n15269) );
  AOI21_X1 U18594 ( .B1(n16280), .B2(n15270), .A(n15269), .ZN(n15271) );
  OAI21_X1 U18595 ( .B1(n15272), .B2(n16295), .A(n15271), .ZN(n15274) );
  NAND2_X1 U18596 ( .A1(n15277), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15282) );
  AOI211_X1 U18597 ( .C1(n16280), .C2(n15280), .A(n15279), .B(n15278), .ZN(
        n15281) );
  OAI211_X1 U18598 ( .C1(n15283), .C2(n16295), .A(n15282), .B(n15281), .ZN(
        n15284) );
  AOI21_X1 U18599 ( .B1(n15285), .B2(n16270), .A(n15284), .ZN(n15286) );
  OAI21_X1 U18600 ( .B1(n15287), .B2(n16274), .A(n15286), .ZN(P2_U3019) );
  INV_X1 U18601 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15292) );
  INV_X1 U18602 ( .A(n15288), .ZN(n15289) );
  AOI211_X1 U18603 ( .C1(n15292), .C2(n15291), .A(n15290), .B(n15289), .ZN(
        n15293) );
  AOI211_X1 U18604 ( .C1(n16280), .C2(n16170), .A(n15294), .B(n15293), .ZN(
        n15295) );
  OAI21_X1 U18605 ( .B1(n16167), .B2(n16295), .A(n15295), .ZN(n15298) );
  NOR2_X1 U18606 ( .A1(n15296), .A2(n16305), .ZN(n15297) );
  AOI211_X1 U18607 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n15299), .A(
        n15298), .B(n15297), .ZN(n15300) );
  OAI21_X1 U18608 ( .B1(n15301), .B2(n16274), .A(n15300), .ZN(P2_U3020) );
  AOI211_X1 U18609 ( .C1(n16280), .C2(n15304), .A(n15303), .B(n15302), .ZN(
        n15305) );
  OAI21_X1 U18610 ( .B1(n15306), .B2(n16295), .A(n15305), .ZN(n15309) );
  NOR2_X1 U18611 ( .A1(n15307), .A2(n16305), .ZN(n15308) );
  AOI211_X1 U18612 ( .C1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n15310), .A(
        n15309), .B(n15308), .ZN(n15311) );
  OAI21_X1 U18613 ( .B1(n15312), .B2(n16274), .A(n15311), .ZN(P2_U3022) );
  INV_X1 U18614 ( .A(n15337), .ZN(n15313) );
  AOI211_X1 U18615 ( .C1(n15315), .C2(n15342), .A(n15314), .B(n15313), .ZN(
        n15316) );
  AOI211_X1 U18616 ( .C1(n16280), .C2(n15318), .A(n15317), .B(n15316), .ZN(
        n15320) );
  NAND2_X1 U18617 ( .A1(n15357), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15319) );
  OAI211_X1 U18618 ( .C1(n15321), .C2(n16295), .A(n15320), .B(n15319), .ZN(
        n15322) );
  AOI21_X1 U18619 ( .B1(n15323), .B2(n16270), .A(n15322), .ZN(n15324) );
  OAI21_X1 U18620 ( .B1(n15325), .B2(n16274), .A(n15324), .ZN(P2_U3023) );
  INV_X1 U18621 ( .A(n15326), .ZN(n15327) );
  NOR2_X1 U18622 ( .A1(n15328), .A2(n15327), .ZN(n15329) );
  XNOR2_X1 U18623 ( .A(n15330), .B(n15329), .ZN(n16192) );
  INV_X1 U18624 ( .A(n16192), .ZN(n15346) );
  INV_X1 U18625 ( .A(n15331), .ZN(n15332) );
  AOI21_X1 U18626 ( .B1(n15342), .B2(n15333), .A(n15332), .ZN(n16190) );
  INV_X1 U18627 ( .A(n15357), .ZN(n15343) );
  OR2_X1 U18628 ( .A1(n15335), .A2(n15334), .ZN(n15336) );
  NAND2_X1 U18629 ( .A1(n15336), .A2(n9614), .ZN(n15746) );
  NAND2_X1 U18630 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19155), .ZN(n15339) );
  NAND2_X1 U18631 ( .A1(n15337), .A2(n15342), .ZN(n15338) );
  OAI211_X1 U18632 ( .C1(n16294), .C2(n15746), .A(n15339), .B(n15338), .ZN(
        n15340) );
  AOI21_X1 U18633 ( .B1(n16191), .B2(n16283), .A(n15340), .ZN(n15341) );
  OAI21_X1 U18634 ( .B1(n15343), .B2(n15342), .A(n15341), .ZN(n15344) );
  AOI21_X1 U18635 ( .B1(n16190), .B2(n16270), .A(n15344), .ZN(n15345) );
  OAI21_X1 U18636 ( .B1(n15346), .B2(n16274), .A(n15345), .ZN(P2_U3024) );
  NAND2_X1 U18637 ( .A1(n15347), .A2(n16301), .ZN(n15359) );
  INV_X1 U18638 ( .A(n15449), .ZN(n15348) );
  NOR2_X1 U18639 ( .A1(n15486), .A2(n15482), .ZN(n15466) );
  NAND2_X1 U18640 ( .A1(n15348), .A2(n15466), .ZN(n16276) );
  NAND2_X1 U18641 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15349), .ZN(
        n15350) );
  INV_X1 U18642 ( .A(n15351), .ZN(n15367) );
  NOR3_X1 U18643 ( .A1(n16261), .A2(n20881), .A3(n15367), .ZN(n15365) );
  NAND3_X1 U18644 ( .A1(n15365), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n15352), .ZN(n15353) );
  OAI211_X1 U18645 ( .C1(n18862), .C2(n16295), .A(n15354), .B(n15353), .ZN(
        n15356) );
  NOR2_X1 U18646 ( .A1(n18863), .A2(n16294), .ZN(n15355) );
  AOI211_X1 U18647 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15357), .A(
        n15356), .B(n15355), .ZN(n15358) );
  OAI211_X1 U18648 ( .C1(n15360), .C2(n16305), .A(n15359), .B(n15358), .ZN(
        P2_U3025) );
  NOR2_X1 U18649 ( .A1(n15361), .A2(n16295), .ZN(n15362) );
  AOI211_X1 U18650 ( .C1(n15365), .C2(n15364), .A(n15363), .B(n15362), .ZN(
        n15369) );
  OAI21_X1 U18651 ( .B1(n15366), .B2(n15384), .A(n15487), .ZN(n15380) );
  NOR3_X1 U18652 ( .A1(n16261), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n15367), .ZN(n15375) );
  OAI21_X1 U18653 ( .B1(n15380), .B2(n15375), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15368) );
  OAI211_X1 U18654 ( .C1(n16179), .C2(n16294), .A(n15369), .B(n15368), .ZN(
        n15370) );
  AOI21_X1 U18655 ( .B1(n15371), .B2(n16270), .A(n15370), .ZN(n15372) );
  OAI21_X1 U18656 ( .B1(n15373), .B2(n16274), .A(n15372), .ZN(P2_U3026) );
  NAND2_X1 U18657 ( .A1(n15374), .A2(n16301), .ZN(n15382) );
  INV_X1 U18658 ( .A(n15375), .ZN(n15377) );
  OAI211_X1 U18659 ( .C1(n16295), .C2(n18874), .A(n15377), .B(n15376), .ZN(
        n15379) );
  NOR2_X1 U18660 ( .A1(n18875), .A2(n16294), .ZN(n15378) );
  AOI211_X1 U18661 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15380), .A(
        n15379), .B(n15378), .ZN(n15381) );
  OAI211_X1 U18662 ( .C1(n15383), .C2(n16305), .A(n15382), .B(n15381), .ZN(
        P2_U3027) );
  OAI21_X1 U18663 ( .B1(n15385), .B2(n15384), .A(n15487), .ZN(n16266) );
  AOI21_X1 U18664 ( .B1(n15386), .B2(n16297), .A(n16266), .ZN(n15393) );
  NAND2_X1 U18665 ( .A1(n16186), .A2(n16280), .ZN(n15391) );
  NOR3_X1 U18666 ( .A1(n16261), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15386), .ZN(n15387) );
  AOI211_X1 U18667 ( .C1(n16283), .C2(n15389), .A(n15388), .B(n15387), .ZN(
        n15390) );
  OAI211_X1 U18668 ( .C1(n15393), .C2(n15392), .A(n15391), .B(n15390), .ZN(
        n15394) );
  AOI21_X1 U18669 ( .B1(n15395), .B2(n16270), .A(n15394), .ZN(n15396) );
  OAI21_X1 U18670 ( .B1(n15397), .B2(n16274), .A(n15396), .ZN(P2_U3028) );
  INV_X1 U18671 ( .A(n16266), .ZN(n15399) );
  NAND2_X1 U18672 ( .A1(n15401), .A2(n16301), .ZN(n15409) );
  OAI22_X1 U18673 ( .A1(n15403), .A2(n16305), .B1(n16261), .B2(n15402), .ZN(
        n15407) );
  AOI22_X1 U18674 ( .A1(n16283), .A2(n18884), .B1(P2_REIP_REG_17__SCAN_IN), 
        .B2(n19155), .ZN(n15404) );
  OAI21_X1 U18675 ( .B1(n15405), .B2(n16294), .A(n15404), .ZN(n15406) );
  AOI21_X1 U18676 ( .B1(n15407), .B2(n15410), .A(n15406), .ZN(n15408) );
  AND2_X1 U18677 ( .A1(n9662), .A2(n15411), .ZN(n15413) );
  OR2_X1 U18678 ( .A1(n15413), .A2(n15412), .ZN(n19055) );
  OAI21_X1 U18679 ( .B1(n16198), .B2(n16305), .A(n16261), .ZN(n15414) );
  NAND3_X1 U18680 ( .A1(n15414), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n20859), .ZN(n15416) );
  AOI22_X1 U18681 ( .A1(n16283), .A2(n18901), .B1(P2_REIP_REG_16__SCAN_IN), 
        .B2(n19155), .ZN(n15415) );
  OAI211_X1 U18682 ( .C1(n16294), .C2(n19055), .A(n15416), .B(n15415), .ZN(
        n15417) );
  AOI21_X1 U18683 ( .B1(n15418), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15417), .ZN(n15419) );
  OAI21_X1 U18684 ( .B1(n15420), .B2(n16274), .A(n15419), .ZN(P2_U3030) );
  NAND2_X1 U18685 ( .A1(n15421), .A2(n16301), .ZN(n15430) );
  OAI21_X1 U18686 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15482), .A(
        n15487), .ZN(n15465) );
  AOI21_X1 U18687 ( .B1(n15449), .B2(n16297), .A(n15465), .ZN(n15439) );
  OAI21_X1 U18688 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16276), .A(
        n15439), .ZN(n16288) );
  OR2_X1 U18689 ( .A1(n15422), .A2(n15435), .ZN(n15424) );
  NAND2_X1 U18690 ( .A1(n15424), .A2(n15423), .ZN(n19067) );
  NAND2_X1 U18691 ( .A1(n16283), .A2(n18924), .ZN(n15427) );
  NOR2_X1 U18692 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16276), .ZN(
        n16289) );
  NOR2_X1 U18693 ( .A1(n20796), .A2(n16264), .ZN(n15425) );
  AOI21_X1 U18694 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16289), .A(
        n15425), .ZN(n15426) );
  OAI211_X1 U18695 ( .C1(n19067), .C2(n16294), .A(n15427), .B(n15426), .ZN(
        n15428) );
  AOI21_X1 U18696 ( .B1(n16288), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15428), .ZN(n15429) );
  OAI211_X1 U18697 ( .C1(n15431), .C2(n16305), .A(n15430), .B(n15429), .ZN(
        P2_U3033) );
  AND2_X1 U18698 ( .A1(n15448), .A2(n15432), .ZN(n15434) );
  OR2_X1 U18699 ( .A1(n15434), .A2(n15433), .ZN(n16212) );
  AOI21_X1 U18700 ( .B1(n15453), .B2(n15436), .A(n15435), .ZN(n19068) );
  NOR2_X1 U18701 ( .A1(n16295), .A2(n15437), .ZN(n15441) );
  NAND2_X1 U18702 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19155), .ZN(n15438) );
  OAI221_X1 U18703 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16276), 
        .C1(n15432), .C2(n15439), .A(n15438), .ZN(n15440) );
  AOI211_X1 U18704 ( .C1(n16280), .C2(n19068), .A(n15441), .B(n15440), .ZN(
        n15447) );
  AND2_X1 U18705 ( .A1(n15443), .A2(n15442), .ZN(n15444) );
  XNOR2_X1 U18706 ( .A(n15445), .B(n15444), .ZN(n16209) );
  NAND2_X1 U18707 ( .A1(n16209), .A2(n16301), .ZN(n15446) );
  OAI211_X1 U18708 ( .C1(n16212), .C2(n16305), .A(n15447), .B(n15446), .ZN(
        P2_U3034) );
  NOR2_X1 U18709 ( .A1(n15478), .A2(n20795), .ZN(n15463) );
  OAI21_X1 U18710 ( .B1(n15463), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15448), .ZN(n16217) );
  INV_X1 U18711 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n15452) );
  NAND2_X1 U18712 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15465), .ZN(
        n15451) );
  OAI211_X1 U18713 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n15449), .B(n15466), .ZN(
        n15450) );
  OAI211_X1 U18714 ( .C1(n16264), .C2(n15452), .A(n15451), .B(n15450), .ZN(
        n15457) );
  OAI21_X1 U18715 ( .B1(n15455), .B2(n15454), .A(n15453), .ZN(n19073) );
  NOR2_X1 U18716 ( .A1(n19073), .A2(n16294), .ZN(n15456) );
  AOI211_X1 U18717 ( .C1(n16283), .C2(n16219), .A(n15457), .B(n15456), .ZN(
        n15462) );
  XNOR2_X1 U18718 ( .A(n15459), .B(n9843), .ZN(n15460) );
  XNOR2_X1 U18719 ( .A(n15458), .B(n15460), .ZN(n16216) );
  OR2_X1 U18720 ( .A1(n16216), .A2(n16274), .ZN(n15461) );
  OAI211_X1 U18721 ( .C1(n16217), .C2(n16305), .A(n15462), .B(n15461), .ZN(
        P2_U3035) );
  AOI21_X1 U18722 ( .B1(n20795), .B2(n15478), .A(n15463), .ZN(n16223) );
  NAND2_X1 U18723 ( .A1(n16223), .A2(n16270), .ZN(n15477) );
  INV_X1 U18724 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19757) );
  NOR2_X1 U18725 ( .A1(n19757), .A2(n16264), .ZN(n15464) );
  AOI221_X1 U18726 ( .B1(n15466), .B2(n20795), .C1(n15465), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n15464), .ZN(n15476) );
  XNOR2_X1 U18727 ( .A(n15479), .B(n15467), .ZN(n19076) );
  INV_X1 U18728 ( .A(n16224), .ZN(n18955) );
  OAI22_X1 U18729 ( .A1(n19076), .A2(n16294), .B1(n16295), .B2(n18955), .ZN(
        n15468) );
  INV_X1 U18730 ( .A(n15468), .ZN(n15475) );
  INV_X1 U18731 ( .A(n15488), .ZN(n15492) );
  OR2_X1 U18732 ( .A1(n15469), .A2(n15492), .ZN(n15473) );
  NAND2_X1 U18733 ( .A1(n15471), .A2(n15470), .ZN(n15472) );
  XNOR2_X1 U18734 ( .A(n15473), .B(n15472), .ZN(n16225) );
  NAND2_X1 U18735 ( .A1(n16225), .A2(n16301), .ZN(n15474) );
  NAND4_X1 U18736 ( .A1(n15477), .A2(n15476), .A3(n15475), .A4(n15474), .ZN(
        P2_U3036) );
  OAI21_X1 U18737 ( .B1(n12640), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15478), .ZN(n16229) );
  OAI21_X1 U18738 ( .B1(n15481), .B2(n15480), .A(n15479), .ZN(n19078) );
  INV_X1 U18739 ( .A(n19078), .ZN(n15498) );
  INV_X1 U18740 ( .A(n18966), .ZN(n16231) );
  NOR2_X1 U18741 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15482), .ZN(
        n15484) );
  INV_X1 U18742 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19755) );
  NOR2_X1 U18743 ( .A1(n19755), .A2(n16264), .ZN(n15483) );
  AOI211_X1 U18744 ( .C1(n16283), .C2(n16231), .A(n15484), .B(n15483), .ZN(
        n15485) );
  OAI21_X1 U18745 ( .B1(n15487), .B2(n15486), .A(n15485), .ZN(n15497) );
  NAND2_X1 U18746 ( .A1(n15469), .A2(n15488), .ZN(n15495) );
  NAND2_X1 U18747 ( .A1(n15490), .A2(n15489), .ZN(n15491) );
  OAI21_X1 U18748 ( .B1(n15493), .B2(n15492), .A(n15491), .ZN(n15494) );
  NAND2_X1 U18749 ( .A1(n15495), .A2(n15494), .ZN(n16228) );
  NOR2_X1 U18750 ( .A1(n16228), .A2(n16274), .ZN(n15496) );
  AOI211_X1 U18751 ( .C1(n16280), .C2(n15498), .A(n15497), .B(n15496), .ZN(
        n15499) );
  OAI21_X1 U18752 ( .B1(n16305), .B2(n16229), .A(n15499), .ZN(P2_U3037) );
  XNOR2_X1 U18753 ( .A(n15501), .B(n15500), .ZN(n16236) );
  INV_X1 U18754 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19753) );
  OAI22_X1 U18755 ( .A1(n16295), .A2(n16235), .B1(n19753), .B2(n18992), .ZN(
        n15505) );
  OAI21_X1 U18756 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n15521), .ZN(n15502) );
  OAI22_X1 U18757 ( .A1(n15538), .A2(n11174), .B1(n15503), .B2(n15502), .ZN(
        n15504) );
  AOI211_X1 U18758 ( .C1(n16280), .C2(n19079), .A(n15505), .B(n15504), .ZN(
        n15515) );
  NAND2_X1 U18759 ( .A1(n15507), .A2(n15506), .ZN(n15513) );
  INV_X1 U18760 ( .A(n15508), .ZN(n15509) );
  AOI21_X1 U18761 ( .B1(n15511), .B2(n15510), .A(n15509), .ZN(n15512) );
  XOR2_X1 U18762 ( .A(n15513), .B(n15512), .Z(n16239) );
  NAND2_X1 U18763 ( .A1(n16239), .A2(n16301), .ZN(n15514) );
  OAI211_X1 U18764 ( .C1(n16236), .C2(n16305), .A(n15515), .B(n15514), .ZN(
        P2_U3038) );
  OR2_X1 U18765 ( .A1(n15517), .A2(n15516), .ZN(n15519) );
  NAND2_X1 U18766 ( .A1(n15519), .A2(n15518), .ZN(n19082) );
  NAND2_X1 U18767 ( .A1(n15521), .A2(n15520), .ZN(n15526) );
  INV_X1 U18768 ( .A(n15538), .ZN(n15524) );
  NOR2_X1 U18769 ( .A1(n19751), .A2(n16264), .ZN(n15523) );
  NOR2_X1 U18770 ( .A1(n16295), .A2(n18976), .ZN(n15522) );
  AOI211_X1 U18771 ( .C1(n15524), .C2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n15523), .B(n15522), .ZN(n15525) );
  OAI211_X1 U18772 ( .C1(n16294), .C2(n19082), .A(n15526), .B(n15525), .ZN(
        n15527) );
  AOI21_X1 U18773 ( .B1(n15528), .B2(n16301), .A(n15527), .ZN(n15529) );
  OAI21_X1 U18774 ( .B1(n15530), .B2(n16305), .A(n15529), .ZN(P2_U3039) );
  NOR3_X1 U18775 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15531), .A3(
        n15557), .ZN(n15542) );
  XNOR2_X1 U18776 ( .A(n15533), .B(n15532), .ZN(n19084) );
  INV_X1 U18777 ( .A(n18986), .ZN(n15535) );
  NOR2_X1 U18778 ( .A1(n19749), .A2(n16264), .ZN(n15534) );
  AOI21_X1 U18779 ( .B1(n16283), .B2(n15535), .A(n15534), .ZN(n15536) );
  OAI21_X1 U18780 ( .B1(n15538), .B2(n15537), .A(n15536), .ZN(n15539) );
  INV_X1 U18781 ( .A(n15539), .ZN(n15540) );
  OAI21_X1 U18782 ( .B1(n19084), .B2(n16294), .A(n15540), .ZN(n15541) );
  OR2_X1 U18783 ( .A1(n15542), .A2(n15541), .ZN(n15543) );
  AOI21_X1 U18784 ( .B1(n15544), .B2(n16301), .A(n15543), .ZN(n15545) );
  OAI21_X1 U18785 ( .B1(n15546), .B2(n16305), .A(n15545), .ZN(P2_U3040) );
  XNOR2_X1 U18786 ( .A(n15547), .B(n15548), .ZN(n16244) );
  OAI21_X1 U18787 ( .B1(n10034), .B2(n15551), .A(n15550), .ZN(n15552) );
  OAI21_X1 U18788 ( .B1(n15553), .B2(n10034), .A(n15552), .ZN(n16246) );
  INV_X1 U18789 ( .A(n16246), .ZN(n15565) );
  OAI21_X1 U18790 ( .B1(n15556), .B2(n15555), .A(n15554), .ZN(n19094) );
  OAI22_X1 U18791 ( .A1(n15559), .A2(n20886), .B1(n15558), .B2(n15557), .ZN(
        n15561) );
  INV_X1 U18792 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19748) );
  NOR2_X1 U18793 ( .A1(n19748), .A2(n16264), .ZN(n15560) );
  AOI221_X1 U18794 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n15561), .C1(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n15561), .A(n15560), .ZN(
        n15563) );
  NAND2_X1 U18795 ( .A1(n16283), .A2(n19001), .ZN(n15562) );
  OAI211_X1 U18796 ( .C1(n19094), .C2(n16294), .A(n15563), .B(n15562), .ZN(
        n15564) );
  AOI21_X1 U18797 ( .B1(n15565), .B2(n16270), .A(n15564), .ZN(n15566) );
  OAI21_X1 U18798 ( .B1(n16274), .B2(n16244), .A(n15566), .ZN(P2_U3041) );
  AOI22_X1 U18799 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n16296), .B1(
        n16280), .B2(n19826), .ZN(n15575) );
  AOI21_X1 U18800 ( .B1(n16283), .B2(n15568), .A(n15567), .ZN(n15574) );
  AOI22_X1 U18801 ( .A1(n16301), .A2(n15570), .B1(n16270), .B2(n15569), .ZN(
        n15573) );
  OAI211_X1 U18802 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n16297), .B(n15571), .ZN(n15572) );
  NAND4_X1 U18803 ( .A1(n15575), .A2(n15574), .A3(n15573), .A4(n15572), .ZN(
        P2_U3045) );
  NAND2_X1 U18804 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15576), .ZN(n15583) );
  NAND2_X1 U18805 ( .A1(n19023), .A2(n15598), .ZN(n15581) );
  MUX2_X1 U18806 ( .A(n15579), .B(n15578), .S(n15577), .Z(n15580) );
  NAND2_X1 U18807 ( .A1(n15581), .A2(n15580), .ZN(n16328) );
  NAND2_X1 U18808 ( .A1(n16328), .A2(n19801), .ZN(n15582) );
  OAI211_X1 U18809 ( .C1(n15584), .C2(n15601), .A(n15583), .B(n15582), .ZN(
        n15585) );
  MUX2_X1 U18810 ( .A(n15585), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n15602), .Z(P2_U3601) );
  INV_X1 U18811 ( .A(n15589), .ZN(n15586) );
  AOI22_X1 U18812 ( .A1(n15587), .A2(n15586), .B1(n10739), .B2(n10868), .ZN(
        n15594) );
  NAND2_X1 U18813 ( .A1(n15588), .A2(n12399), .ZN(n15592) );
  INV_X1 U18814 ( .A(n10739), .ZN(n15590) );
  AOI21_X1 U18815 ( .B1(n10868), .B2(n15590), .A(n15589), .ZN(n15591) );
  AND2_X1 U18816 ( .A1(n15592), .A2(n15591), .ZN(n15593) );
  MUX2_X1 U18817 ( .A(n15594), .B(n15593), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15596) );
  NAND2_X1 U18818 ( .A1(n15596), .A2(n15595), .ZN(n15597) );
  AOI21_X1 U18819 ( .B1(n15599), .B2(n15598), .A(n15597), .ZN(n16334) );
  OAI22_X1 U18820 ( .A1(n19235), .A2(n15601), .B1(n15600), .B2(n16334), .ZN(
        n15603) );
  MUX2_X1 U18821 ( .A(n15603), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15602), .Z(P2_U3596) );
  NOR2_X1 U18822 ( .A1(n17240), .A2(n17184), .ZN(n17187) );
  NOR2_X1 U18823 ( .A1(n17188), .A2(n16928), .ZN(n16932) );
  AOI21_X1 U18824 ( .B1(n17187), .B2(n16919), .A(n16932), .ZN(n16924) );
  INV_X1 U18825 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n15683) );
  AOI22_X1 U18826 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12691), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15604) );
  OAI21_X1 U18827 ( .B1(n12721), .B2(n18160), .A(n15604), .ZN(n15614) );
  AOI22_X1 U18828 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15684), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15612) );
  AOI22_X1 U18829 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15605) );
  OAI21_X1 U18830 ( .B1(n17004), .B2(n17124), .A(n15605), .ZN(n15610) );
  AOI22_X1 U18831 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15607) );
  AOI22_X1 U18832 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15648), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15606) );
  OAI211_X1 U18833 ( .C1(n17090), .C2(n15608), .A(n15607), .B(n15606), .ZN(
        n15609) );
  AOI211_X1 U18834 ( .C1(n17131), .C2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n15610), .B(n15609), .ZN(n15611) );
  OAI211_X1 U18835 ( .C1(n17113), .C2(n17128), .A(n15612), .B(n15611), .ZN(
        n15613) );
  AOI211_X1 U18836 ( .C1(n17141), .C2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n15614), .B(n15613), .ZN(n16939) );
  AOI22_X1 U18837 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15625) );
  AOI22_X1 U18838 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15624) );
  OAI22_X1 U18839 ( .A1(n17113), .A2(n15615), .B1(n17146), .B2(n20773), .ZN(
        n15622) );
  AOI22_X1 U18840 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15684), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15620) );
  AOI22_X1 U18841 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15617) );
  AOI22_X1 U18842 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15648), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15616) );
  OAI211_X1 U18843 ( .C1(n17090), .C2(n17035), .A(n15617), .B(n15616), .ZN(
        n15618) );
  AOI21_X1 U18844 ( .B1(n17131), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n15618), .ZN(n15619) );
  OAI211_X1 U18845 ( .C1(n17004), .C2(n17024), .A(n15620), .B(n15619), .ZN(
        n15621) );
  AOI211_X1 U18846 ( .C1(n17156), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n15622), .B(n15621), .ZN(n15623) );
  NAND3_X1 U18847 ( .A1(n15625), .A2(n15624), .A3(n15623), .ZN(n16943) );
  AOI22_X1 U18848 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17105), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17149), .ZN(n15635) );
  AOI22_X1 U18849 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15627) );
  AOI22_X1 U18850 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n15684), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17143), .ZN(n15626) );
  OAI211_X1 U18851 ( .C1(n9565), .C2(n18244), .A(n15627), .B(n15626), .ZN(
        n15633) );
  AOI22_X1 U18852 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n16899), .ZN(n15631) );
  AOI22_X1 U18853 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n9568), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n17122), .ZN(n15630) );
  AOI22_X1 U18854 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n15648), .ZN(n15629) );
  NAND2_X1 U18855 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n9574), .ZN(
        n15628) );
  NAND4_X1 U18856 ( .A1(n15631), .A2(n15630), .A3(n15629), .A4(n15628), .ZN(
        n15632) );
  AOI211_X1 U18857 ( .C1(n17131), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n15633), .B(n15632), .ZN(n15634) );
  OAI211_X1 U18858 ( .C1(n15636), .C2(n17090), .A(n15635), .B(n15634), .ZN(
        n16944) );
  NAND2_X1 U18859 ( .A1(n16943), .A2(n16944), .ZN(n16942) );
  NOR2_X1 U18860 ( .A1(n16939), .A2(n16942), .ZN(n16936) );
  AOI22_X1 U18861 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9574), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15647) );
  AOI22_X1 U18862 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15684), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15637) );
  OAI21_X1 U18863 ( .B1(n10053), .B2(n17118), .A(n15637), .ZN(n15645) );
  AOI22_X1 U18864 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15642) );
  AOI22_X1 U18865 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15648), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15639) );
  AOI22_X1 U18866 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12691), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15638) );
  OAI211_X1 U18867 ( .C1(n17146), .C2(n18228), .A(n15639), .B(n15638), .ZN(
        n15640) );
  AOI21_X1 U18868 ( .B1(n17156), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n15640), .ZN(n15641) );
  OAI211_X1 U18869 ( .C1(n17108), .C2(n15643), .A(n15642), .B(n15641), .ZN(
        n15644) );
  AOI211_X1 U18870 ( .C1(n17148), .C2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n15645), .B(n15644), .ZN(n15646) );
  OAI211_X1 U18871 ( .C1(n9616), .C2(n17112), .A(n15647), .B(n15646), .ZN(
        n16935) );
  NAND2_X1 U18872 ( .A1(n16936), .A2(n16935), .ZN(n16934) );
  INV_X1 U18873 ( .A(n16934), .ZN(n16931) );
  AOI22_X1 U18874 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15658) );
  INV_X1 U18875 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18232) );
  AOI22_X1 U18876 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15650) );
  AOI22_X1 U18877 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15648), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15649) );
  OAI211_X1 U18878 ( .C1(n17146), .C2(n18232), .A(n15650), .B(n15649), .ZN(
        n15656) );
  AOI22_X1 U18879 ( .A1(n17122), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15684), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15654) );
  AOI22_X1 U18880 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15653) );
  AOI22_X1 U18881 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15652) );
  NAND2_X1 U18882 ( .A1(n12701), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n15651) );
  NAND4_X1 U18883 ( .A1(n15654), .A2(n15653), .A3(n15652), .A4(n15651), .ZN(
        n15655) );
  AOI211_X1 U18884 ( .C1(n17131), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n15656), .B(n15655), .ZN(n15657) );
  OAI211_X1 U18885 ( .C1(n17004), .C2(n20809), .A(n15658), .B(n15657), .ZN(
        n16930) );
  AOI22_X1 U18886 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15669) );
  INV_X1 U18887 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15661) );
  AOI22_X1 U18888 ( .A1(n9568), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15660) );
  AOI22_X1 U18889 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15659) );
  OAI211_X1 U18890 ( .C1(n9565), .C2(n15661), .A(n15660), .B(n15659), .ZN(
        n15667) );
  AOI22_X1 U18891 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15665) );
  AOI22_X1 U18892 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15664) );
  AOI22_X1 U18893 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15684), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15663) );
  NAND2_X1 U18894 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n15662) );
  NAND4_X1 U18895 ( .A1(n15665), .A2(n15664), .A3(n15663), .A4(n15662), .ZN(
        n15666) );
  AOI211_X1 U18896 ( .C1(n17131), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n15667), .B(n15666), .ZN(n15668) );
  OAI211_X1 U18897 ( .C1(n17113), .C2(n17083), .A(n15669), .B(n15668), .ZN(
        n16926) );
  NAND3_X1 U18898 ( .A1(n16931), .A2(n16930), .A3(n16926), .ZN(n16925) );
  INV_X1 U18899 ( .A(n16925), .ZN(n16915) );
  AOI22_X1 U18900 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15680) );
  AOI22_X1 U18901 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15670) );
  OAI21_X1 U18902 ( .B1(n12661), .B2(n15671), .A(n15670), .ZN(n15678) );
  OAI22_X1 U18903 ( .A1(n9564), .A2(n15686), .B1(n12721), .B2(n18184), .ZN(
        n15672) );
  AOI21_X1 U18904 ( .B1(n9574), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A(n15672), .ZN(n15676) );
  AOI22_X1 U18905 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15675) );
  AOI22_X1 U18906 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15684), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15674) );
  AOI22_X1 U18907 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15673) );
  NAND4_X1 U18908 ( .A1(n15676), .A2(n15675), .A3(n15674), .A4(n15673), .ZN(
        n15677) );
  AOI211_X1 U18909 ( .C1(n16899), .C2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n15678), .B(n15677), .ZN(n15679) );
  OAI211_X1 U18910 ( .C1(n17113), .C2(n16966), .A(n15680), .B(n15679), .ZN(
        n16916) );
  XOR2_X1 U18911 ( .A(n16915), .B(n16916), .Z(n17211) );
  INV_X1 U18912 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16927) );
  NOR2_X1 U18913 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16927), .ZN(n15681) );
  AOI22_X1 U18914 ( .A1(n17188), .A2(n17211), .B1(n16928), .B2(n15681), .ZN(
        n15682) );
  OAI21_X1 U18915 ( .B1(n16924), .B2(n15683), .A(n15682), .ZN(P3_U2675) );
  AOI22_X1 U18916 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15684), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15685) );
  OAI21_X1 U18917 ( .B1(n17088), .B2(n15686), .A(n15685), .ZN(n15696) );
  INV_X1 U18918 ( .A(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15694) );
  AOI22_X1 U18919 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15693) );
  AOI22_X1 U18920 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15687) );
  OAI21_X1 U18921 ( .B1(n17146), .B2(n18184), .A(n15687), .ZN(n15691) );
  AOI22_X1 U18922 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15689) );
  AOI22_X1 U18923 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15688) );
  OAI211_X1 U18924 ( .C1(n9565), .C2(n16966), .A(n15689), .B(n15688), .ZN(
        n15690) );
  AOI211_X1 U18925 ( .C1(n12701), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n15691), .B(n15690), .ZN(n15692) );
  OAI211_X1 U18926 ( .C1(n17004), .C2(n15694), .A(n15693), .B(n15692), .ZN(
        n15695) );
  AOI211_X1 U18927 ( .C1(n17032), .C2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n15696), .B(n15695), .ZN(n17289) );
  AND2_X1 U18928 ( .A1(n18193), .A2(n17055), .ZN(n17085) );
  OAI21_X1 U18929 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17085), .A(n15697), .ZN(
        n15698) );
  AOI22_X1 U18930 ( .A1(n17188), .A2(n17289), .B1(n15698), .B2(n17186), .ZN(
        P3_U2690) );
  NOR2_X1 U18931 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18759), .ZN(
        n18199) );
  NOR3_X1 U18932 ( .A1(n18809), .A2(n18770), .A3(n18805), .ZN(n18663) );
  NAND3_X1 U18933 ( .A1(n17113), .A2(n15717), .A3(n18607), .ZN(n18139) );
  AOI221_X1 U18934 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n18663), .C1(n18139), .C2(
        n18663), .A(n18508), .ZN(n15699) );
  NOR2_X1 U18935 ( .A1(n18199), .A2(n15699), .ZN(n15701) );
  INV_X1 U18936 ( .A(n15699), .ZN(n18145) );
  INV_X1 U18937 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18407) );
  OAI22_X1 U18938 ( .A1(n17788), .A2(n18811), .B1(n18407), .B2(n18759), .ZN(
        n15704) );
  NAND3_X1 U18939 ( .A1(n18635), .A2(n18145), .A3(n15704), .ZN(n15700) );
  OAI221_X1 U18940 ( .B1(n18635), .B2(n15701), .C1(n18635), .C2(n18505), .A(
        n15700), .ZN(P3_U2864) );
  NAND2_X1 U18941 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18384) );
  NOR2_X1 U18942 ( .A1(n17788), .A2(n18811), .ZN(n15703) );
  INV_X1 U18943 ( .A(n15701), .ZN(n15702) );
  AOI221_X1 U18944 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18384), .C1(n15703), 
        .C2(n18384), .A(n15702), .ZN(n18144) );
  INV_X1 U18945 ( .A(n18505), .ZN(n18246) );
  OAI221_X1 U18946 ( .B1(n18246), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18246), .C2(n15704), .A(n18145), .ZN(n18142) );
  AOI22_X1 U18947 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18144), .B1(
        n18142), .B2(n18640), .ZN(P3_U2865) );
  AOI21_X1 U18948 ( .B1(n17408), .B2(n18804), .A(n15705), .ZN(n15825) );
  NOR2_X1 U18949 ( .A1(n15707), .A2(n15706), .ZN(n18651) );
  INV_X1 U18950 ( .A(n18675), .ZN(n18803) );
  OAI21_X1 U18951 ( .B1(n15708), .B2(n18651), .A(n18803), .ZN(n17348) );
  INV_X1 U18952 ( .A(n18599), .ZN(n16504) );
  AOI211_X1 U18953 ( .C1(n15825), .C2(n17348), .A(n16504), .B(n18806), .ZN(
        n15713) );
  INV_X1 U18954 ( .A(n15709), .ZN(n15712) );
  OAI211_X1 U18955 ( .C1(n16496), .C2(n15712), .A(n15711), .B(n15710), .ZN(
        n15728) );
  NOR3_X1 U18956 ( .A1(n15714), .A2(n15713), .A3(n15728), .ZN(n18638) );
  INV_X1 U18957 ( .A(n18638), .ZN(n18627) );
  INV_X1 U18958 ( .A(n18663), .ZN(n18758) );
  INV_X1 U18959 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18140) );
  OAI22_X1 U18960 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18759), .B1(n18758), 
        .B2(n18140), .ZN(n15715) );
  AOI21_X1 U18961 ( .B1(n15717), .B2(n18607), .A(n15716), .ZN(n18650) );
  NAND3_X1 U18962 ( .A1(n18788), .A2(n18786), .A3(n18650), .ZN(n15718) );
  OAI21_X1 U18963 ( .B1(n18788), .B2(n18607), .A(n15718), .ZN(P3_U3284) );
  INV_X1 U18964 ( .A(n17596), .ZN(n17933) );
  NAND3_X1 U18965 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15720) );
  INV_X1 U18966 ( .A(n15720), .ZN(n17935) );
  AOI21_X1 U18967 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18079) );
  INV_X1 U18968 ( .A(n18079), .ZN(n18098) );
  NAND2_X1 U18969 ( .A1(n17935), .A2(n18098), .ZN(n18047) );
  NAND3_X1 U18970 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15719) );
  NOR2_X1 U18971 ( .A1(n18047), .A2(n15719), .ZN(n18011) );
  NAND3_X1 U18972 ( .A1(n17933), .A2(n17888), .A3(n18011), .ZN(n15735) );
  INV_X1 U18973 ( .A(n15735), .ZN(n17928) );
  AOI21_X1 U18974 ( .B1(n18628), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18608), .ZN(n17934) );
  INV_X1 U18975 ( .A(n17934), .ZN(n18104) );
  INV_X1 U18976 ( .A(n15719), .ZN(n15721) );
  NAND2_X1 U18977 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18077) );
  NOR2_X1 U18978 ( .A1(n15720), .A2(n18077), .ZN(n18045) );
  NAND2_X1 U18979 ( .A1(n15721), .A2(n18045), .ZN(n17949) );
  NOR2_X1 U18980 ( .A1(n9944), .A2(n17949), .ZN(n17889) );
  AND2_X1 U18981 ( .A1(n17933), .A2(n17889), .ZN(n15722) );
  AOI22_X1 U18982 ( .A1(n18609), .A2(n17928), .B1(n18104), .B2(n15722), .ZN(
        n17852) );
  NOR2_X1 U18983 ( .A1(n17852), .A2(n16410), .ZN(n16389) );
  NAND2_X1 U18984 ( .A1(n17316), .A2(n18111), .ZN(n18041) );
  OAI22_X1 U18985 ( .A1(n18107), .A2(n17836), .B1(n16374), .B2(n18041), .ZN(
        n15734) );
  INV_X1 U18986 ( .A(n18602), .ZN(n15733) );
  OAI21_X1 U18987 ( .B1(n15724), .B2(n15723), .A(n18175), .ZN(n15730) );
  OAI21_X1 U18988 ( .B1(n18163), .B2(n18804), .A(n18675), .ZN(n15725) );
  OAI21_X1 U18989 ( .B1(n15726), .B2(n15725), .A(n18814), .ZN(n16501) );
  AOI211_X1 U18990 ( .C1(n18163), .C2(n15727), .A(n16504), .B(n16501), .ZN(
        n15729) );
  AOI211_X1 U18991 ( .C1(n18601), .C2(n15730), .A(n15729), .B(n15728), .ZN(
        n15732) );
  AOI221_X4 U18992 ( .B1(n15733), .B2(n15732), .C1(n15731), .C2(n15732), .A(
        n18657), .ZN(n18129) );
  OAI211_X1 U18993 ( .C1(n16389), .C2(n15734), .A(n18129), .B(n16375), .ZN(
        n15799) );
  NOR2_X1 U18994 ( .A1(n9586), .A2(n18116), .ZN(n18124) );
  NOR2_X1 U18995 ( .A1(n18608), .A2(n18609), .ZN(n18022) );
  INV_X1 U18996 ( .A(n18022), .ZN(n17988) );
  INV_X1 U18997 ( .A(n15736), .ZN(n17880) );
  NOR2_X1 U18998 ( .A1(n17880), .A2(n15735), .ZN(n17869) );
  AOI21_X1 U18999 ( .B1(n16361), .B2(n17869), .A(n18626), .ZN(n15738) );
  NAND2_X1 U19000 ( .A1(n18029), .A2(n18630), .ZN(n18078) );
  INV_X1 U19001 ( .A(n18078), .ZN(n18099) );
  NAND2_X1 U19002 ( .A1(n18628), .A2(n18787), .ZN(n18100) );
  NAND2_X1 U19003 ( .A1(n17889), .A2(n18100), .ZN(n17930) );
  NAND2_X1 U19004 ( .A1(n17933), .A2(n15736), .ZN(n16360) );
  OAI21_X1 U19005 ( .B1(n17930), .B2(n16360), .A(n18078), .ZN(n17866) );
  OAI21_X1 U19006 ( .B1(n16361), .B2(n18099), .A(n17866), .ZN(n15737) );
  NOR2_X1 U19007 ( .A1(n15738), .A2(n15737), .ZN(n17833) );
  OAI211_X1 U19008 ( .C1(n18029), .C2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n18129), .B(n17833), .ZN(n15796) );
  AOI21_X1 U19009 ( .B1(n17484), .B2(n17988), .A(n15796), .ZN(n16405) );
  NAND2_X1 U19010 ( .A1(n18597), .A2(n18129), .ZN(n18127) );
  INV_X1 U19011 ( .A(n18127), .ZN(n18134) );
  NAND2_X1 U19012 ( .A1(n16390), .A2(n17461), .ZN(n16358) );
  INV_X1 U19013 ( .A(n18111), .ZN(n18603) );
  INV_X1 U19014 ( .A(n18132), .ZN(n18076) );
  NOR3_X1 U19015 ( .A1(n16359), .A2(n16403), .A3(n18076), .ZN(n15739) );
  AOI21_X1 U19016 ( .B1(n18134), .B2(n16358), .A(n15739), .ZN(n15802) );
  OAI21_X1 U19017 ( .B1(n9577), .B2(n16405), .A(n15802), .ZN(n15740) );
  AOI21_X1 U19018 ( .B1(n18124), .B2(n20916), .A(n15740), .ZN(n15745) );
  INV_X1 U19019 ( .A(n18137), .ZN(n18044) );
  NAND2_X1 U19020 ( .A1(n15742), .A2(n15741), .ZN(n15743) );
  XOR2_X1 U19021 ( .A(n15743), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n16380) );
  AOI22_X1 U19022 ( .A1(n18044), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n18033), 
        .B2(n16380), .ZN(n15744) );
  OAI221_X1 U19023 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15799), 
        .C1(n16377), .C2(n15745), .A(n15744), .ZN(P3_U2833) );
  INV_X1 U19024 ( .A(n15746), .ZN(n16173) );
  AOI22_X1 U19025 ( .A1(n16191), .A2(n19022), .B1(n19027), .B2(n16173), .ZN(
        n15757) );
  AOI211_X1 U19026 ( .C1(n15749), .C2(n15748), .A(n15747), .B(n19720), .ZN(
        n15755) );
  INV_X1 U19027 ( .A(n15750), .ZN(n15753) );
  INV_X1 U19028 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n15751) );
  OAI222_X1 U19029 ( .A1(n19008), .A2(n15753), .B1(n19009), .B2(n15752), .C1(
        n18993), .C2(n15751), .ZN(n15754) );
  AOI211_X1 U19030 ( .C1(n19041), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15755), .B(n15754), .ZN(n15756) );
  NAND2_X1 U19031 ( .A1(n15757), .A2(n15756), .ZN(P2_U2833) );
  NOR2_X1 U19032 ( .A1(n15758), .A2(n15787), .ZN(n15795) );
  INV_X1 U19033 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20078) );
  OAI211_X1 U19034 ( .C1(n11345), .C2(n15760), .A(n15759), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n15762) );
  OAI21_X1 U19035 ( .B1(n15762), .B2(n20615), .A(n15761), .ZN(n15764) );
  NAND2_X1 U19036 ( .A1(n15762), .A2(n20615), .ZN(n15763) );
  OAI21_X1 U19037 ( .B1(n15765), .B2(n15764), .A(n15763), .ZN(n15766) );
  AOI222_X1 U19038 ( .A1(n20371), .A2(n15767), .B1(n20371), .B2(n15766), .C1(
        n15767), .C2(n15766), .ZN(n15770) );
  INV_X1 U19039 ( .A(n15768), .ZN(n15769) );
  AOI222_X1 U19040 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15770), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15769), .C1(n15770), 
        .C2(n15769), .ZN(n15772) );
  AOI21_X1 U19041 ( .B1(n20078), .B2(n15772), .A(n15771), .ZN(n15779) );
  OAI21_X1 U19042 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15773), .ZN(n15775) );
  AND4_X1 U19043 ( .A1(n15777), .A2(n15776), .A3(n15775), .A4(n15774), .ZN(
        n15778) );
  NOR3_X1 U19044 ( .A1(n15782), .A2(n15781), .A3(n15780), .ZN(n15783) );
  AOI221_X1 U19045 ( .B1(n15785), .B2(n15784), .C1(n20691), .C2(n15784), .A(
        n15783), .ZN(n16153) );
  OAI221_X1 U19046 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n15786), 
        .A(n16153), .ZN(n16159) );
  NAND2_X1 U19047 ( .A1(n16159), .A2(n20676), .ZN(n15794) );
  INV_X1 U19048 ( .A(n15786), .ZN(n15790) );
  OAI211_X1 U19049 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20691), .A(n15788), 
        .B(n15787), .ZN(n15789) );
  AOI21_X1 U19050 ( .B1(n15791), .B2(n15790), .A(n15789), .ZN(n15792) );
  AND2_X1 U19051 ( .A1(n16159), .A2(n15792), .ZN(n15793) );
  OAI22_X1 U19052 ( .A1(n15795), .A2(n15794), .B1(n15793), .B2(n20676), .ZN(
        P1_U3161) );
  INV_X1 U19053 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16370) );
  INV_X1 U19054 ( .A(n9586), .ZN(n17874) );
  OAI221_X1 U19055 ( .B1(n15796), .B2(n17874), .C1(n15796), .C2(n16362), .A(
        n18137), .ZN(n16398) );
  INV_X1 U19056 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18746) );
  NOR2_X1 U19057 ( .A1(n18137), .A2(n18746), .ZN(n16363) );
  NOR3_X1 U19058 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16377), .A3(
        n15799), .ZN(n15800) );
  OAI221_X1 U19059 ( .B1(n16370), .B2(n15802), .C1(n16370), .C2(n16398), .A(
        n15801), .ZN(P3_U2832) );
  INV_X1 U19060 ( .A(HOLD), .ZN(n20684) );
  INV_X1 U19061 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20692) );
  NOR2_X1 U19062 ( .A1(n20692), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n19878) );
  INV_X1 U19063 ( .A(n19878), .ZN(n20689) );
  INV_X1 U19064 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20769) );
  AOI211_X1 U19065 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(HOLD), .A(n20695), .B(
        n20769), .ZN(n15803) );
  AOI211_X1 U19066 ( .C1(n20762), .C2(P1_STATE_REG_1__SCAN_IN), .A(n15804), 
        .B(n15803), .ZN(n15805) );
  OAI21_X1 U19067 ( .B1(n20684), .B2(n20689), .A(n15805), .ZN(P1_U3195) );
  AND2_X1 U19068 ( .A1(n20924), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  OAI21_X1 U19069 ( .B1(n15808), .B2(n15807), .A(n15806), .ZN(n15820) );
  INV_X1 U19070 ( .A(n15809), .ZN(n15810) );
  NAND2_X1 U19071 ( .A1(n15810), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15811) );
  MUX2_X1 U19072 ( .A(n15812), .B(n15811), .S(n15965), .Z(n15813) );
  XNOR2_X1 U19073 ( .A(n15813), .B(n15822), .ZN(n15977) );
  INV_X1 U19074 ( .A(n15977), .ZN(n15818) );
  INV_X1 U19075 ( .A(n15865), .ZN(n15816) );
  NAND3_X1 U19076 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15814), .A3(
        n15822), .ZN(n15815) );
  NAND2_X1 U19077 ( .A1(n16139), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15981) );
  OAI211_X1 U19078 ( .C1(n15816), .C2(n16069), .A(n15815), .B(n15981), .ZN(
        n15817) );
  AOI21_X1 U19079 ( .B1(n15818), .B2(n20071), .A(n15817), .ZN(n15819) );
  OAI221_X1 U19080 ( .B1(n15822), .B2(n15821), .C1(n15822), .C2(n15820), .A(
        n15819), .ZN(P1_U3011) );
  NAND2_X1 U19081 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19860), .ZN(n19716) );
  NOR2_X1 U19082 ( .A1(n19711), .A2(n19716), .ZN(n16344) );
  NOR3_X1 U19083 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15823) );
  NOR4_X1 U19084 ( .A1(n19857), .A2(n16344), .A3(n16345), .A4(n15823), .ZN(
        P2_U3178) );
  INV_X1 U19085 ( .A(n16346), .ZN(n19843) );
  AOI221_X1 U19086 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16345), .C1(n19843), .C2(
        n16345), .A(n19656), .ZN(n19838) );
  INV_X1 U19087 ( .A(n19838), .ZN(n19835) );
  NOR2_X1 U19088 ( .A1(n15824), .A2(n19835), .ZN(P2_U3047) );
  OAI33_X1 U19089 ( .A1(n16820), .A2(n18804), .A3(n15826), .B1(n15825), .B2(
        n17409), .B3(n18806), .ZN(n17192) );
  INV_X1 U19090 ( .A(n9585), .ZN(n17340) );
  NOR2_X1 U19091 ( .A1(n17240), .A2(n17340), .ZN(n17343) );
  INV_X1 U19092 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17407) );
  NOR2_X1 U19093 ( .A1(n15827), .A2(n17340), .ZN(n17311) );
  AOI22_X1 U19094 ( .A1(n17341), .A2(BUF2_REG_0__SCAN_IN), .B1(n17311), .B2(
        n17826), .ZN(n15828) );
  OAI221_X1 U19095 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17326), .C1(n17407), 
        .C2(n9585), .A(n15828), .ZN(P3_U2735) );
  NOR3_X1 U19096 ( .A1(n19901), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n15829), 
        .ZN(n15833) );
  AOI22_X1 U19097 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19969), .B1(
        n19909), .B2(n15830), .ZN(n15831) );
  OAI21_X1 U19098 ( .B1(n19960), .B2(n14395), .A(n15831), .ZN(n15832) );
  AOI211_X1 U19099 ( .C1(n15834), .C2(n19936), .A(n15833), .B(n15832), .ZN(
        n15837) );
  OAI21_X1 U19100 ( .B1(n15835), .B2(n15842), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n15836) );
  OAI211_X1 U19101 ( .C1(n19977), .C2(n15838), .A(n15837), .B(n15836), .ZN(
        P1_U2815) );
  INV_X1 U19102 ( .A(n15971), .ZN(n15839) );
  AOI222_X1 U19103 ( .A1(n19974), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19969), .C1(n15839), .C2(
        n19909), .ZN(n15844) );
  OAI21_X1 U19104 ( .B1(n19901), .B2(n15840), .A(n20726), .ZN(n15841) );
  AOI22_X1 U19105 ( .A1(n15968), .A2(n19936), .B1(n15842), .B2(n15841), .ZN(
        n15843) );
  OAI211_X1 U19106 ( .C1(n19977), .C2(n16042), .A(n15844), .B(n15843), .ZN(
        P1_U2817) );
  AOI22_X1 U19107 ( .A1(n19974), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19969), .ZN(n15854) );
  NOR2_X1 U19108 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n19901), .ZN(n15845) );
  AOI22_X1 U19109 ( .A1(n15847), .A2(n19909), .B1(n15846), .B2(n15845), .ZN(
        n15853) );
  AOI22_X1 U19110 ( .A1(n15848), .A2(n19936), .B1(n19942), .B2(n16052), .ZN(
        n15852) );
  OAI21_X1 U19111 ( .B1(n15929), .B2(n15849), .A(n19955), .ZN(n15862) );
  INV_X1 U19112 ( .A(n15862), .ZN(n15850) );
  NOR3_X1 U19113 ( .A1(n19901), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n15849), 
        .ZN(n15858) );
  OAI21_X1 U19114 ( .B1(n15850), .B2(n15858), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15851) );
  NAND4_X1 U19115 ( .A1(n15854), .A2(n15853), .A3(n15852), .A4(n15851), .ZN(
        P1_U2818) );
  OAI22_X1 U19116 ( .A1(n15976), .A2(n19986), .B1(n20723), .B2(n15862), .ZN(
        n15855) );
  INV_X1 U19117 ( .A(n15855), .ZN(n15860) );
  AOI22_X1 U19118 ( .A1(n19974), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n19969), .ZN(n15856) );
  INV_X1 U19119 ( .A(n15856), .ZN(n15857) );
  AOI211_X1 U19120 ( .C1(n15973), .C2(n19936), .A(n15858), .B(n15857), .ZN(
        n15859) );
  OAI211_X1 U19121 ( .C1(n19977), .C2(n15861), .A(n15860), .B(n15859), .ZN(
        P1_U2819) );
  AOI22_X1 U19122 ( .A1(n19974), .A2(P1_EBX_REG_20__SCAN_IN), .B1(n19909), 
        .B2(n15980), .ZN(n15867) );
  AOI21_X1 U19123 ( .B1(n15872), .B2(n15874), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15863) );
  OAI22_X1 U19124 ( .A1(n15978), .A2(n19946), .B1(n15863), .B2(n15862), .ZN(
        n15864) );
  AOI21_X1 U19125 ( .B1(n19942), .B2(n15865), .A(n15864), .ZN(n15866) );
  OAI211_X1 U19126 ( .C1(n15983), .C2(n15945), .A(n15867), .B(n15866), .ZN(
        P1_U2820) );
  AOI21_X1 U19127 ( .B1(n19969), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n19968), .ZN(n15868) );
  INV_X1 U19128 ( .A(n15868), .ZN(n15871) );
  OAI22_X1 U19129 ( .A1(n19960), .A2(n15869), .B1(n19986), .B2(n15989), .ZN(
        n15870) );
  AOI211_X1 U19130 ( .C1(P1_REIP_REG_19__SCAN_IN), .C2(n15884), .A(n15871), 
        .B(n15870), .ZN(n15878) );
  AOI21_X1 U19131 ( .B1(n20720), .B2(n15873), .A(n15872), .ZN(n15875) );
  AOI22_X1 U19132 ( .A1(n15876), .A2(n19936), .B1(n15875), .B2(n15874), .ZN(
        n15877) );
  OAI211_X1 U19133 ( .C1(n19977), .C2(n15879), .A(n15878), .B(n15877), .ZN(
        P1_U2821) );
  OAI22_X1 U19134 ( .A1(n19960), .A2(n15881), .B1(n15880), .B2(n15945), .ZN(
        n15882) );
  AOI211_X1 U19135 ( .C1(n19909), .C2(n15996), .A(n19968), .B(n15882), .ZN(
        n15887) );
  NAND2_X1 U19136 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15888) );
  INV_X1 U19137 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n15883) );
  OAI21_X1 U19138 ( .B1(n15888), .B2(n15907), .A(n15883), .ZN(n15885) );
  AOI22_X1 U19139 ( .A1(n15997), .A2(n19936), .B1(n15885), .B2(n15884), .ZN(
        n15886) );
  OAI211_X1 U19140 ( .C1(n19977), .C2(n16068), .A(n15887), .B(n15886), .ZN(
        P1_U2823) );
  OAI21_X1 U19141 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n15888), .ZN(n15899) );
  INV_X1 U19142 ( .A(n15889), .ZN(n16075) );
  AOI22_X1 U19143 ( .A1(n16075), .A2(n19942), .B1(n19974), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n15890) );
  OAI211_X1 U19144 ( .C1(n15945), .C2(n15891), .A(n15890), .B(n19944), .ZN(
        n15896) );
  AOI21_X1 U19145 ( .B1(n19914), .B2(n15893), .A(n15892), .ZN(n15922) );
  OAI22_X1 U19146 ( .A1(n15894), .A2(n19946), .B1(n14638), .B2(n15922), .ZN(
        n15895) );
  AOI211_X1 U19147 ( .C1(n15897), .C2(n19909), .A(n15896), .B(n15895), .ZN(
        n15898) );
  OAI21_X1 U19148 ( .B1(n15907), .B2(n15899), .A(n15898), .ZN(P1_U2824) );
  INV_X1 U19149 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20714) );
  INV_X1 U19150 ( .A(n16000), .ZN(n15901) );
  AOI21_X1 U19151 ( .B1(n19969), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n19968), .ZN(n15900) );
  OAI21_X1 U19152 ( .B1(n19986), .B2(n15901), .A(n15900), .ZN(n15902) );
  AOI21_X1 U19153 ( .B1(n19974), .B2(P1_EBX_REG_15__SCAN_IN), .A(n15902), .ZN(
        n15903) );
  OAI21_X1 U19154 ( .B1(n19977), .B2(n15904), .A(n15903), .ZN(n15905) );
  AOI21_X1 U19155 ( .B1(n16001), .B2(n19936), .A(n15905), .ZN(n15906) );
  OAI221_X1 U19156 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n15907), .C1(n20714), 
        .C2(n15922), .A(n15906), .ZN(P1_U2825) );
  AOI21_X1 U19157 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15908), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n15921) );
  INV_X1 U19158 ( .A(n15909), .ZN(n16088) );
  NAND2_X1 U19159 ( .A1(n19923), .A2(n16088), .ZN(n15912) );
  NAND2_X1 U19160 ( .A1(n19969), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15910) );
  AND2_X1 U19161 ( .A1(n15910), .A2(n19944), .ZN(n15911) );
  OAI211_X1 U19162 ( .C1(n15913), .C2(n19960), .A(n15912), .B(n15911), .ZN(
        n15914) );
  INV_X1 U19163 ( .A(n15914), .ZN(n15920) );
  INV_X1 U19164 ( .A(n15915), .ZN(n15918) );
  INV_X1 U19165 ( .A(n15916), .ZN(n15917) );
  AOI22_X1 U19166 ( .A1(n15918), .A2(n19936), .B1(n15917), .B2(n19909), .ZN(
        n15919) );
  OAI211_X1 U19167 ( .C1(n15922), .C2(n15921), .A(n15920), .B(n15919), .ZN(
        P1_U2826) );
  NOR2_X1 U19168 ( .A1(n19901), .A2(n15938), .ZN(n15932) );
  AOI21_X1 U19169 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15932), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15927) );
  OAI22_X1 U19170 ( .A1(n19960), .A2(n15954), .B1(n15923), .B2(n15945), .ZN(
        n15924) );
  AOI211_X1 U19171 ( .C1(n15952), .C2(n19923), .A(n19968), .B(n15924), .ZN(
        n15926) );
  AOI22_X1 U19172 ( .A1(n16006), .A2(n19909), .B1(n19936), .B2(n16005), .ZN(
        n15925) );
  OAI211_X1 U19173 ( .C1(n15928), .C2(n15927), .A(n15926), .B(n15925), .ZN(
        P1_U2828) );
  AOI21_X1 U19174 ( .B1(n19914), .B2(n15938), .A(n15929), .ZN(n15951) );
  XNOR2_X1 U19175 ( .A(n15931), .B(n15930), .ZN(n16102) );
  AOI22_X1 U19176 ( .A1(n19942), .A2(n16102), .B1(n15932), .B2(n15937), .ZN(
        n15936) );
  AOI22_X1 U19177 ( .A1(n19974), .A2(P1_EBX_REG_11__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19969), .ZN(n15933) );
  OAI211_X1 U19178 ( .C1(n19986), .C2(n16020), .A(n15933), .B(n19944), .ZN(
        n15934) );
  AOI21_X1 U19179 ( .B1(n19936), .B2(n16017), .A(n15934), .ZN(n15935) );
  OAI211_X1 U19180 ( .C1(n15951), .C2(n15937), .A(n15936), .B(n15935), .ZN(
        P1_U2829) );
  AND2_X1 U19181 ( .A1(n15938), .A2(n19914), .ZN(n15939) );
  AOI22_X1 U19182 ( .A1(n19942), .A2(n16109), .B1(n15940), .B2(n15939), .ZN(
        n15950) );
  INV_X1 U19183 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15944) );
  INV_X1 U19184 ( .A(n15941), .ZN(n15942) );
  NAND2_X1 U19185 ( .A1(n19909), .A2(n15942), .ZN(n15943) );
  OAI211_X1 U19186 ( .C1(n15945), .C2(n15944), .A(n19944), .B(n15943), .ZN(
        n15948) );
  NOR2_X1 U19187 ( .A1(n15946), .A2(n19946), .ZN(n15947) );
  AOI211_X1 U19188 ( .C1(n19974), .C2(P1_EBX_REG_10__SCAN_IN), .A(n15948), .B(
        n15947), .ZN(n15949) );
  OAI211_X1 U19189 ( .C1(n15951), .C2(n14665), .A(n15950), .B(n15949), .ZN(
        P1_U2830) );
  AOI22_X1 U19190 ( .A1(n16005), .A2(n19990), .B1(n19989), .B2(n15952), .ZN(
        n15953) );
  OAI21_X1 U19191 ( .B1(n19994), .B2(n15954), .A(n15953), .ZN(P1_U2860) );
  AOI22_X1 U19192 ( .A1(n16017), .A2(n19990), .B1(n19989), .B2(n16102), .ZN(
        n15955) );
  OAI21_X1 U19193 ( .B1(n19994), .B2(n15956), .A(n15955), .ZN(P1_U2861) );
  INV_X1 U19194 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n19220) );
  AOI22_X1 U19195 ( .A1(n15959), .A2(n15958), .B1(n15957), .B2(
        P1_EAX_REG_23__SCAN_IN), .ZN(n15963) );
  AOI22_X1 U19196 ( .A1(n15968), .A2(n15961), .B1(n15960), .B2(DATAI_23_), 
        .ZN(n15962) );
  OAI211_X1 U19197 ( .C1(n15964), .C2(n19220), .A(n15963), .B(n15962), .ZN(
        P1_U2881) );
  AOI22_X1 U19198 ( .A1(n20058), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n16139), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n15970) );
  XNOR2_X1 U19199 ( .A(n15965), .B(n16047), .ZN(n15966) );
  XNOR2_X1 U19200 ( .A(n15967), .B(n15966), .ZN(n16044) );
  AOI22_X1 U19201 ( .A1(n15968), .A2(n16031), .B1(n20060), .B2(n16044), .ZN(
        n15969) );
  OAI211_X1 U19202 ( .C1(n16034), .C2(n15971), .A(n15970), .B(n15969), .ZN(
        P1_U2976) );
  AOI22_X1 U19203 ( .A1(n20058), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n16139), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15975) );
  AOI22_X1 U19204 ( .A1(n15973), .A2(n16031), .B1(n15972), .B2(n20060), .ZN(
        n15974) );
  OAI211_X1 U19205 ( .C1(n16034), .C2(n15976), .A(n15975), .B(n15974), .ZN(
        P1_U2978) );
  OAI22_X1 U19206 ( .A1(n15978), .A2(n20081), .B1(n15977), .B2(n19879), .ZN(
        n15979) );
  AOI21_X1 U19207 ( .B1(n16007), .B2(n15980), .A(n15979), .ZN(n15982) );
  OAI211_X1 U19208 ( .C1(n15983), .C2(n16039), .A(n15982), .B(n15981), .ZN(
        P1_U2979) );
  AOI22_X1 U19209 ( .A1(n20058), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n16139), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15988) );
  OAI22_X1 U19210 ( .A1(n15985), .A2(n20081), .B1(n15984), .B2(n19879), .ZN(
        n15986) );
  INV_X1 U19211 ( .A(n15986), .ZN(n15987) );
  OAI211_X1 U19212 ( .C1(n16034), .C2(n15989), .A(n15988), .B(n15987), .ZN(
        P1_U2980) );
  INV_X1 U19213 ( .A(n15990), .ZN(n15991) );
  NOR2_X1 U19214 ( .A1(n15992), .A2(n15991), .ZN(n15994) );
  NOR2_X1 U19215 ( .A1(n15994), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15993) );
  MUX2_X1 U19216 ( .A(n15994), .B(n15993), .S(n16013), .Z(n15995) );
  AOI22_X1 U19217 ( .A1(n20058), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n16139), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15999) );
  AOI22_X1 U19218 ( .A1(n15997), .A2(n16031), .B1(n15996), .B2(n16007), .ZN(
        n15998) );
  OAI211_X1 U19219 ( .C1(n19879), .C2(n16071), .A(n15999), .B(n15998), .ZN(
        P1_U2982) );
  AOI22_X1 U19220 ( .A1(n20058), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n16139), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16003) );
  AOI22_X1 U19221 ( .A1(n16001), .A2(n16031), .B1(n16007), .B2(n16000), .ZN(
        n16002) );
  OAI211_X1 U19222 ( .C1(n16004), .C2(n19879), .A(n16003), .B(n16002), .ZN(
        P1_U2984) );
  AOI22_X1 U19223 ( .A1(n20058), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n16139), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16009) );
  AOI22_X1 U19224 ( .A1(n16007), .A2(n16006), .B1(n16031), .B2(n16005), .ZN(
        n16008) );
  OAI211_X1 U19225 ( .C1(n16010), .C2(n19879), .A(n16009), .B(n16008), .ZN(
        P1_U2987) );
  AOI22_X1 U19226 ( .A1(n20058), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16139), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16019) );
  INV_X1 U19227 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16113) );
  NOR2_X1 U19228 ( .A1(n16011), .A2(n16113), .ZN(n16015) );
  NOR2_X1 U19229 ( .A1(n16012), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16014) );
  MUX2_X1 U19230 ( .A(n16015), .B(n16014), .S(n16013), .Z(n16016) );
  XNOR2_X1 U19231 ( .A(n16016), .B(n14058), .ZN(n16104) );
  AOI22_X1 U19232 ( .A1(n20060), .A2(n16104), .B1(n16031), .B2(n16017), .ZN(
        n16018) );
  OAI211_X1 U19233 ( .C1(n16034), .C2(n16020), .A(n16019), .B(n16018), .ZN(
        P1_U2988) );
  AOI22_X1 U19234 ( .A1(n20058), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16139), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16026) );
  NAND2_X1 U19235 ( .A1(n16022), .A2(n16021), .ZN(n16023) );
  NAND2_X1 U19236 ( .A1(n16024), .A2(n16023), .ZN(n16130) );
  AOI22_X1 U19237 ( .A1(n16130), .A2(n20060), .B1(n16031), .B2(n19937), .ZN(
        n16025) );
  OAI211_X1 U19238 ( .C1(n16034), .C2(n19934), .A(n16026), .B(n16025), .ZN(
        P1_U2992) );
  AOI22_X1 U19239 ( .A1(n20058), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n16139), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16033) );
  NAND2_X1 U19240 ( .A1(n16028), .A2(n16027), .ZN(n16029) );
  XNOR2_X1 U19241 ( .A(n16030), .B(n16029), .ZN(n16141) );
  AOI22_X1 U19242 ( .A1(n16141), .A2(n20060), .B1(n16031), .B2(n19991), .ZN(
        n16032) );
  OAI211_X1 U19243 ( .C1(n16034), .C2(n19945), .A(n16033), .B(n16032), .ZN(
        P1_U2993) );
  OAI22_X1 U19244 ( .A1(n19959), .A2(n20081), .B1(n19957), .B2(n16034), .ZN(
        n16035) );
  AOI21_X1 U19245 ( .B1(n16036), .B2(n20060), .A(n16035), .ZN(n16038) );
  OAI211_X1 U19246 ( .C1(n16040), .C2(n16039), .A(n16038), .B(n16037), .ZN(
        P1_U2994) );
  OAI22_X1 U19247 ( .A1(n16042), .A2(n16069), .B1(n20726), .B2(n16041), .ZN(
        n16043) );
  AOI21_X1 U19248 ( .B1(n16044), .B2(n20071), .A(n16043), .ZN(n16045) );
  OAI221_X1 U19249 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16048), 
        .C1(n16047), .C2(n16046), .A(n16045), .ZN(P1_U3008) );
  INV_X1 U19250 ( .A(n16049), .ZN(n16051) );
  AOI22_X1 U19251 ( .A1(n16051), .A2(n20071), .B1(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n16050), .ZN(n16058) );
  NAND2_X1 U19252 ( .A1(n16139), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n16057) );
  NAND2_X1 U19253 ( .A1(n16052), .A2(n20067), .ZN(n16056) );
  OAI211_X1 U19254 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16054), .B(n16053), .ZN(
        n16055) );
  NAND4_X1 U19255 ( .A1(n16058), .A2(n16057), .A3(n16056), .A4(n16055), .ZN(
        P1_U3009) );
  AOI21_X1 U19256 ( .B1(n16121), .B2(n16059), .A(n16096), .ZN(n16073) );
  NOR2_X1 U19257 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16059), .ZN(
        n16060) );
  AOI22_X1 U19258 ( .A1(n16139), .A2(P1_REIP_REG_18__SCAN_IN), .B1(n16061), 
        .B2(n16060), .ZN(n16066) );
  INV_X1 U19259 ( .A(n16062), .ZN(n16064) );
  AOI22_X1 U19260 ( .A1(n16064), .A2(n20071), .B1(n20067), .B2(n16063), .ZN(
        n16065) );
  OAI211_X1 U19261 ( .C1(n16073), .C2(n16067), .A(n16066), .B(n16065), .ZN(
        P1_U3013) );
  AOI21_X1 U19262 ( .B1(n16076), .B2(n16078), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16072) );
  AOI21_X1 U19263 ( .B1(n16075), .B2(n20067), .A(n16074), .ZN(n16082) );
  AOI21_X1 U19264 ( .B1(n16077), .B2(n16083), .A(n16076), .ZN(n16079) );
  AOI22_X1 U19265 ( .A1(n16080), .A2(n20071), .B1(n16079), .B2(n16078), .ZN(
        n16081) );
  OAI211_X1 U19266 ( .C1(n16084), .C2(n16083), .A(n16082), .B(n16081), .ZN(
        P1_U3015) );
  NAND2_X1 U19267 ( .A1(n16086), .A2(n16085), .ZN(n16092) );
  AOI21_X1 U19268 ( .B1(n16088), .B2(n20067), .A(n16087), .ZN(n16091) );
  AOI22_X1 U19269 ( .A1(n16089), .A2(n20071), .B1(n16096), .B2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16090) );
  OAI211_X1 U19270 ( .C1(n16093), .C2(n16092), .A(n16091), .B(n16090), .ZN(
        P1_U3017) );
  AOI21_X1 U19271 ( .B1(n20067), .B2(n16095), .A(n16094), .ZN(n16099) );
  AOI22_X1 U19272 ( .A1(n16097), .A2(n20071), .B1(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16096), .ZN(n16098) );
  OAI211_X1 U19273 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n16100), .A(
        n16099), .B(n16098), .ZN(P1_U3018) );
  INV_X1 U19274 ( .A(n16101), .ZN(n16107) );
  AOI22_X1 U19275 ( .A1(n20067), .A2(n16102), .B1(n16139), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16106) );
  AOI22_X1 U19276 ( .A1(n16104), .A2(n20071), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16103), .ZN(n16105) );
  OAI211_X1 U19277 ( .C1(n16144), .C2(n16107), .A(n16106), .B(n16105), .ZN(
        P1_U3020) );
  AOI21_X1 U19278 ( .B1(n20067), .B2(n16109), .A(n16108), .ZN(n16116) );
  AOI22_X1 U19279 ( .A1(n16111), .A2(n20071), .B1(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16110), .ZN(n16115) );
  OAI221_X1 U19280 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n16113), .C2(n11614), .A(
        n16112), .ZN(n16114) );
  NAND3_X1 U19281 ( .A1(n16116), .A2(n16115), .A3(n16114), .ZN(P1_U3021) );
  INV_X1 U19282 ( .A(n16118), .ZN(n16120) );
  OAI21_X1 U19283 ( .B1(n14754), .B2(n16120), .A(n16119), .ZN(n16140) );
  AOI21_X1 U19284 ( .B1(n16129), .B2(n16121), .A(n16140), .ZN(n16132) );
  INV_X1 U19285 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16128) );
  AOI21_X1 U19286 ( .B1(n20067), .B2(n19924), .A(n16122), .ZN(n16127) );
  INV_X1 U19287 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16133) );
  AOI211_X1 U19288 ( .C1(n16128), .C2(n16133), .A(n16129), .B(n16144), .ZN(
        n16124) );
  AOI22_X1 U19289 ( .A1(n16125), .A2(n20071), .B1(n16124), .B2(n16123), .ZN(
        n16126) );
  OAI211_X1 U19290 ( .C1(n16132), .C2(n16128), .A(n16127), .B(n16126), .ZN(
        P1_U3023) );
  OR2_X1 U19291 ( .A1(n16129), .A2(n16144), .ZN(n16134) );
  AOI222_X1 U19292 ( .A1(n16130), .A2(n20071), .B1(n20067), .B2(n19931), .C1(
        P1_REIP_REG_7__SCAN_IN), .C2(n16139), .ZN(n16131) );
  OAI221_X1 U19293 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16134), .C1(
        n16133), .C2(n16132), .A(n16131), .ZN(P1_U3024) );
  OAI21_X1 U19294 ( .B1(n16137), .B2(n16136), .A(n16135), .ZN(n16138) );
  INV_X1 U19295 ( .A(n16138), .ZN(n19988) );
  AOI22_X1 U19296 ( .A1(n20067), .A2(n19988), .B1(n16139), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16143) );
  AOI22_X1 U19297 ( .A1(n16141), .A2(n20071), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16140), .ZN(n16142) );
  OAI211_X1 U19298 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16144), .A(
        n16143), .B(n16142), .ZN(P1_U3025) );
  INV_X1 U19299 ( .A(n16145), .ZN(n16147) );
  NAND3_X1 U19300 ( .A1(n16148), .A2(n16147), .A3(n16146), .ZN(n16149) );
  OAI21_X1 U19301 ( .B1(n16151), .B2(n16150), .A(n16149), .ZN(P1_U3468) );
  NAND2_X1 U19302 ( .A1(n20841), .A2(n20691), .ZN(n16157) );
  NOR2_X1 U19303 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20762), .ZN(n16152) );
  OAI221_X1 U19304 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n20676), .C2(n16152), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n20678) );
  AOI21_X1 U19305 ( .B1(n20678), .B2(n16154), .A(n16153), .ZN(n16156) );
  AOI21_X1 U19306 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n16159), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16155) );
  AOI211_X1 U19307 ( .C1(n20763), .C2(n16157), .A(n16156), .B(n16155), .ZN(
        P1_U3162) );
  OAI221_X1 U19308 ( .B1(n20841), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n20841), 
        .C2(n16159), .A(n16158), .ZN(P1_U3466) );
  AOI211_X1 U19309 ( .C1(n16162), .C2(n16161), .A(n16160), .B(n19720), .ZN(
        n16169) );
  AOI22_X1 U19310 ( .A1(n19025), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19041), .ZN(n16163) );
  OAI21_X1 U19311 ( .B1(n18993), .B2(n19783), .A(n16163), .ZN(n16164) );
  AOI21_X1 U19312 ( .B1(n16165), .B2(n19030), .A(n16164), .ZN(n16166) );
  OAI21_X1 U19313 ( .B1(n16167), .B2(n19011), .A(n16166), .ZN(n16168) );
  AOI211_X1 U19314 ( .C1(n19027), .C2(n16170), .A(n16169), .B(n16168), .ZN(
        n16171) );
  INV_X1 U19315 ( .A(n16171), .ZN(P2_U2829) );
  AOI22_X1 U19316 ( .A1(n19050), .A2(n16172), .B1(n19110), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16177) );
  AOI22_X1 U19317 ( .A1(n19052), .A2(BUF2_REG_22__SCAN_IN), .B1(n19051), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n16176) );
  AOI22_X1 U19318 ( .A1(n16174), .A2(n19100), .B1(n19111), .B2(n16173), .ZN(
        n16175) );
  NAND3_X1 U19319 ( .A1(n16177), .A2(n16176), .A3(n16175), .ZN(P2_U2897) );
  AOI22_X1 U19320 ( .A1(n19050), .A2(n19096), .B1(n19110), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16183) );
  AOI22_X1 U19321 ( .A1(n19052), .A2(BUF2_REG_20__SCAN_IN), .B1(n19051), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16182) );
  OAI22_X1 U19322 ( .A1(n16179), .A2(n19054), .B1(n19115), .B2(n16178), .ZN(
        n16180) );
  INV_X1 U19323 ( .A(n16180), .ZN(n16181) );
  NAND3_X1 U19324 ( .A1(n16183), .A2(n16182), .A3(n16181), .ZN(P2_U2899) );
  AOI22_X1 U19325 ( .A1(n19050), .A2(n16184), .B1(n19110), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16189) );
  AOI22_X1 U19326 ( .A1(n19052), .A2(BUF2_REG_18__SCAN_IN), .B1(n19051), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16188) );
  AOI22_X1 U19327 ( .A1(n16186), .A2(n19111), .B1(n19100), .B2(n16185), .ZN(
        n16187) );
  NAND3_X1 U19328 ( .A1(n16189), .A2(n16188), .A3(n16187), .ZN(P2_U2901) );
  AOI22_X1 U19329 ( .A1(n19166), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19155), .ZN(n16194) );
  AOI222_X1 U19330 ( .A1(n16192), .A2(n19167), .B1(n16248), .B2(n16191), .C1(
        n19169), .C2(n16190), .ZN(n16193) );
  OAI211_X1 U19331 ( .C1(n19165), .C2(n16195), .A(n16194), .B(n16193), .ZN(
        P2_U2992) );
  AOI22_X1 U19332 ( .A1(n19166), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19155), .ZN(n16207) );
  NAND2_X1 U19333 ( .A1(n16196), .A2(n16278), .ZN(n16197) );
  NAND2_X1 U19334 ( .A1(n16198), .A2(n16197), .ZN(n16286) );
  AND2_X1 U19335 ( .A1(n16200), .A2(n16199), .ZN(n16201) );
  XNOR2_X1 U19336 ( .A(n16202), .B(n16201), .ZN(n16281) );
  NAND2_X1 U19337 ( .A1(n16281), .A2(n19167), .ZN(n16204) );
  NAND2_X1 U19338 ( .A1(n16248), .A2(n16282), .ZN(n16203) );
  OAI211_X1 U19339 ( .C1(n16245), .C2(n16286), .A(n16204), .B(n16203), .ZN(
        n16205) );
  INV_X1 U19340 ( .A(n16205), .ZN(n16206) );
  OAI211_X1 U19341 ( .C1(n19165), .C2(n16208), .A(n16207), .B(n16206), .ZN(
        P2_U3000) );
  AOI22_X1 U19342 ( .A1(n19166), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19155), .ZN(n16215) );
  NAND2_X1 U19343 ( .A1(n16248), .A2(n18934), .ZN(n16211) );
  NAND2_X1 U19344 ( .A1(n16209), .A2(n19167), .ZN(n16210) );
  OAI211_X1 U19345 ( .C1(n16212), .C2(n16245), .A(n16211), .B(n16210), .ZN(
        n16213) );
  INV_X1 U19346 ( .A(n16213), .ZN(n16214) );
  OAI211_X1 U19347 ( .C1(n19165), .C2(n18929), .A(n16215), .B(n16214), .ZN(
        P2_U3002) );
  AOI22_X1 U19348 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19155), .B1(n19175), 
        .B2(n18939), .ZN(n16221) );
  OAI22_X1 U19349 ( .A1(n16217), .A2(n16245), .B1(n16216), .B2(n16243), .ZN(
        n16218) );
  AOI21_X1 U19350 ( .B1(n16248), .B2(n16219), .A(n16218), .ZN(n16220) );
  OAI211_X1 U19351 ( .C1(n16259), .C2(n16222), .A(n16221), .B(n16220), .ZN(
        P2_U3003) );
  AOI22_X1 U19352 ( .A1(n19166), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19155), .ZN(n16227) );
  AOI222_X1 U19353 ( .A1(n16225), .A2(n19167), .B1(n16248), .B2(n16224), .C1(
        n19169), .C2(n16223), .ZN(n16226) );
  OAI211_X1 U19354 ( .C1(n19165), .C2(n18954), .A(n16227), .B(n16226), .ZN(
        P2_U3004) );
  AOI22_X1 U19355 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19155), .B1(n19175), 
        .B2(n18962), .ZN(n16233) );
  OAI22_X1 U19356 ( .A1(n16229), .A2(n16245), .B1(n16243), .B2(n16228), .ZN(
        n16230) );
  AOI21_X1 U19357 ( .B1(n16248), .B2(n16231), .A(n16230), .ZN(n16232) );
  OAI211_X1 U19358 ( .C1(n16259), .C2(n16234), .A(n16233), .B(n16232), .ZN(
        P2_U3005) );
  AOI22_X1 U19359 ( .A1(n19166), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19155), .ZN(n16241) );
  INV_X1 U19360 ( .A(n16235), .ZN(n16238) );
  INV_X1 U19361 ( .A(n16236), .ZN(n16237) );
  AOI222_X1 U19362 ( .A1(n16239), .A2(n19167), .B1(n16248), .B2(n16238), .C1(
        n16237), .C2(n19169), .ZN(n16240) );
  OAI211_X1 U19363 ( .C1(n19165), .C2(n16242), .A(n16241), .B(n16240), .ZN(
        P2_U3006) );
  AOI22_X1 U19364 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19155), .B1(n19175), 
        .B2(n19000), .ZN(n16250) );
  OAI22_X1 U19365 ( .A1(n16246), .A2(n16245), .B1(n16244), .B2(n16243), .ZN(
        n16247) );
  AOI21_X1 U19366 ( .B1(n16248), .B2(n19001), .A(n16247), .ZN(n16249) );
  OAI211_X1 U19367 ( .C1(n16259), .C2(n16251), .A(n16250), .B(n16249), .ZN(
        P2_U3009) );
  AOI22_X1 U19368 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19155), .B1(n19175), 
        .B2(n16252), .ZN(n16258) );
  NAND3_X1 U19369 ( .A1(n16253), .A2(n19169), .A3(n13888), .ZN(n16254) );
  OAI21_X1 U19370 ( .B1(n19179), .B2(n10287), .A(n16254), .ZN(n16255) );
  AOI21_X1 U19371 ( .B1(n16256), .B2(n19167), .A(n16255), .ZN(n16257) );
  OAI211_X1 U19372 ( .C1(n16260), .C2(n16259), .A(n16258), .B(n16257), .ZN(
        P2_U3011) );
  INV_X1 U19373 ( .A(n16261), .ZN(n16268) );
  OAI21_X1 U19374 ( .B1(n16263), .B2(n16262), .A(n9662), .ZN(n19061) );
  OAI22_X1 U19375 ( .A1(n19061), .A2(n16294), .B1(n15211), .B2(n16264), .ZN(
        n16265) );
  AOI221_X1 U19376 ( .B1(n16268), .B2(n16267), .C1(n16266), .C2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(n16265), .ZN(n16273) );
  AOI22_X1 U19377 ( .A1(n16271), .A2(n16270), .B1(n16283), .B2(n16269), .ZN(
        n16272) );
  OAI211_X1 U19378 ( .C1(n16275), .C2(n16274), .A(n16273), .B(n16272), .ZN(
        P2_U3031) );
  NOR2_X1 U19379 ( .A1(n16277), .A2(n16276), .ZN(n16279) );
  AOI22_X1 U19380 ( .A1(n16280), .A2(n19062), .B1(n16279), .B2(n16278), .ZN(
        n16293) );
  NAND2_X1 U19381 ( .A1(n16281), .A2(n16301), .ZN(n16285) );
  NAND2_X1 U19382 ( .A1(n16283), .A2(n16282), .ZN(n16284) );
  OAI211_X1 U19383 ( .C1(n16286), .C2(n16305), .A(n16285), .B(n16284), .ZN(
        n16287) );
  INV_X1 U19384 ( .A(n16287), .ZN(n16292) );
  NAND2_X1 U19385 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19155), .ZN(n16291) );
  OAI21_X1 U19386 ( .B1(n16289), .B2(n16288), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16290) );
  NAND4_X1 U19387 ( .A1(n16293), .A2(n16292), .A3(n16291), .A4(n16290), .ZN(
        P2_U3032) );
  OAI22_X1 U19388 ( .A1(n10260), .A2(n16295), .B1(n16294), .B2(n19024), .ZN(
        n16299) );
  MUX2_X1 U19389 ( .A(n16297), .B(n16296), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n16298) );
  AOI211_X1 U19390 ( .C1(n16301), .C2(n16300), .A(n16299), .B(n16298), .ZN(
        n16303) );
  OAI211_X1 U19391 ( .C1(n16305), .C2(n16304), .A(n16303), .B(n16302), .ZN(
        P2_U3046) );
  INV_X1 U19392 ( .A(n16306), .ZN(n16342) );
  MUX2_X1 U19393 ( .A(n10458), .B(n16307), .S(n16306), .Z(n16330) );
  OAI21_X1 U19394 ( .B1(n16330), .B2(n10115), .A(n16308), .ZN(n16341) );
  NOR3_X1 U19395 ( .A1(n16330), .A2(n16334), .A3(n16342), .ZN(n16324) );
  INV_X1 U19396 ( .A(n16309), .ZN(n16313) );
  AOI22_X1 U19397 ( .A1(n16314), .A2(n16311), .B1(n11117), .B2(n16310), .ZN(
        n16312) );
  OAI21_X1 U19398 ( .B1(n16314), .B2(n16313), .A(n16312), .ZN(n19846) );
  INV_X1 U19399 ( .A(n16315), .ZN(n16317) );
  NOR3_X1 U19400 ( .A1(n16318), .A2(n16317), .A3(n16316), .ZN(n18831) );
  OAI21_X1 U19401 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n18831), .ZN(n16320) );
  OAI211_X1 U19402 ( .C1(n16322), .C2(n16321), .A(n16320), .B(n16319), .ZN(
        n16323) );
  OR3_X1 U19403 ( .A1(n16324), .A2(n19846), .A3(n16323), .ZN(n16340) );
  AOI21_X1 U19404 ( .B1(n16325), .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n19388), .ZN(n16329) );
  NAND2_X1 U19405 ( .A1(n16334), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16327) );
  AOI21_X1 U19406 ( .B1(n16325), .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16342), .ZN(n16326) );
  OAI211_X1 U19407 ( .C1(n16329), .C2(n16328), .A(n16327), .B(n16326), .ZN(
        n16331) );
  NAND2_X1 U19408 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16331), .ZN(
        n16333) );
  OAI22_X1 U19409 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16331), .B1(
        n16330), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n16332) );
  NAND2_X1 U19410 ( .A1(n16333), .A2(n16332), .ZN(n16338) );
  INV_X1 U19411 ( .A(n16334), .ZN(n16336) );
  NAND2_X1 U19412 ( .A1(n16336), .A2(n16335), .ZN(n16337) );
  AOI21_X1 U19413 ( .B1(n16338), .B2(n16337), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16339) );
  AOI211_X1 U19414 ( .C1(n16342), .C2(n16341), .A(n16340), .B(n16339), .ZN(
        n16356) );
  AOI211_X1 U19415 ( .C1(n16346), .C2(n16345), .A(n16344), .B(n16343), .ZN(
        n16355) );
  NOR3_X1 U19416 ( .A1(n16348), .A2(n16347), .A3(n19851), .ZN(n16349) );
  NOR3_X1 U19417 ( .A1(n16349), .A2(n19861), .A3(n19860), .ZN(n16351) );
  OAI221_X1 U19418 ( .B1(n18828), .B2(n16356), .C1(n18828), .C2(n19712), .A(
        n16351), .ZN(n19719) );
  INV_X1 U19419 ( .A(n19719), .ZN(n16353) );
  AOI22_X1 U19420 ( .A1(n19865), .A2(n16351), .B1(n19857), .B2(n16350), .ZN(
        n16352) );
  AOI22_X1 U19421 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16353), .B1(n16352), 
        .B2(n18828), .ZN(n16354) );
  OAI211_X1 U19422 ( .C1(n16356), .C2(n19714), .A(n16355), .B(n16354), .ZN(
        P2_U3176) );
  OAI21_X1 U19423 ( .B1(n10900), .B2(n19719), .A(n16357), .ZN(P2_U3593) );
  NAND2_X1 U19424 ( .A1(n17816), .A2(n16358), .ZN(n16373) );
  OR2_X1 U19425 ( .A1(n9615), .A2(n16359), .ZN(n16376) );
  INV_X1 U19426 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16538) );
  XNOR2_X1 U19427 ( .A(n16538), .B(n16381), .ZN(n16537) );
  AOI21_X1 U19428 ( .B1(n17682), .B2(n16537), .A(n16363), .ZN(n16364) );
  OAI221_X1 U19429 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16366), .C1(
        n16538), .C2(n16365), .A(n16364), .ZN(n16367) );
  OAI221_X1 U19430 ( .B1(n16370), .B2(n16373), .C1(n16370), .C2(n16376), .A(
        n16369), .ZN(P3_U2800) );
  AOI22_X1 U19431 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16372), .B1(
        n9689), .B2(n16371), .ZN(n16386) );
  NAND2_X1 U19432 ( .A1(n16375), .A2(n17461), .ZN(n16407) );
  AOI21_X1 U19433 ( .B1(n16377), .B2(n16407), .A(n16373), .ZN(n16379) );
  INV_X1 U19434 ( .A(n16374), .ZN(n17834) );
  NAND2_X1 U19435 ( .A1(n17834), .A2(n16375), .ZN(n16399) );
  AOI21_X1 U19436 ( .B1(n16377), .B2(n16399), .A(n16376), .ZN(n16378) );
  AOI211_X1 U19437 ( .C1(n17722), .C2(n16380), .A(n16379), .B(n16378), .ZN(
        n16385) );
  NAND2_X1 U19438 ( .A1(n18044), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16384) );
  AOI21_X1 U19439 ( .B1(n9753), .B2(n16522), .A(n16381), .ZN(n16546) );
  OAI21_X1 U19440 ( .B1(n16382), .B2(n17682), .A(n16546), .ZN(n16383) );
  NAND4_X1 U19441 ( .A1(n16386), .A2(n16385), .A3(n16384), .A4(n16383), .ZN(
        P3_U2801) );
  INV_X1 U19442 ( .A(n18041), .ZN(n18008) );
  AOI22_X1 U19443 ( .A1(n18008), .A2(n16388), .B1(n16387), .B2(n17874), .ZN(
        n16392) );
  NAND4_X1 U19444 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16390), .A3(
        n16389), .A4(n18772), .ZN(n16391) );
  OAI211_X1 U19445 ( .C1(n16393), .C2(n18107), .A(n16392), .B(n16391), .ZN(
        n16394) );
  AOI22_X1 U19446 ( .A1(n16395), .A2(n18033), .B1(n18129), .B2(n16394), .ZN(
        n16397) );
  INV_X1 U19447 ( .A(n16399), .ZN(n16406) );
  OAI22_X1 U19448 ( .A1(n17734), .A2(n20916), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17632), .ZN(n16413) );
  INV_X1 U19449 ( .A(n16413), .ZN(n17471) );
  OAI21_X1 U19450 ( .B1(n17475), .B2(n17734), .A(n16401), .ZN(n17470) );
  NAND2_X1 U19451 ( .A1(n17471), .A2(n17470), .ZN(n17469) );
  NAND2_X1 U19452 ( .A1(n16402), .A2(n17475), .ZN(n16412) );
  NAND4_X1 U19453 ( .A1(n18111), .A2(n16403), .A3(n17469), .A4(n16412), .ZN(
        n16404) );
  OAI211_X1 U19454 ( .C1(n16406), .C2(n18041), .A(n16405), .B(n16404), .ZN(
        n16408) );
  OAI221_X1 U19455 ( .B1(n16408), .B2(n18597), .C1(n16408), .C2(n16407), .A(
        n18137), .ZN(n16417) );
  AOI22_X1 U19456 ( .A1(n18597), .A2(n17698), .B1(n17699), .B2(n18008), .ZN(
        n17936) );
  NAND2_X1 U19457 ( .A1(n17933), .A2(n17888), .ZN(n16409) );
  OAI21_X1 U19458 ( .B1(n17936), .B2(n16409), .A(n17852), .ZN(n17882) );
  NAND2_X1 U19459 ( .A1(n18129), .A2(n17882), .ZN(n17903) );
  NOR2_X1 U19460 ( .A1(n16410), .A2(n17903), .ZN(n17837) );
  NAND2_X1 U19461 ( .A1(n20916), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17474) );
  INV_X1 U19462 ( .A(n17474), .ZN(n16411) );
  AOI22_X1 U19463 ( .A1(n18044), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n17837), 
        .B2(n16411), .ZN(n16416) );
  NOR2_X1 U19464 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16412), .ZN(
        n16414) );
  OAI221_X1 U19465 ( .B1(n16414), .B2(n16400), .C1(n16414), .C2(n16413), .A(
        n18033), .ZN(n16415) );
  OAI211_X1 U19466 ( .C1(n20916), .C2(n16417), .A(n16416), .B(n16415), .ZN(
        P3_U2834) );
  NOR3_X1 U19467 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16419) );
  NOR4_X1 U19468 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16418) );
  NAND4_X1 U19469 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16419), .A3(n16418), .A4(
        U215), .ZN(U213) );
  INV_X1 U19470 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19120) );
  INV_X2 U19471 ( .A(U214), .ZN(n16459) );
  NOR2_X1 U19472 ( .A1(n16459), .A2(n16420), .ZN(n16456) );
  INV_X1 U19473 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16421) );
  INV_X1 U19474 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16491) );
  OAI222_X1 U19475 ( .A1(U212), .A2(n19120), .B1(n16461), .B2(n16421), .C1(
        U214), .C2(n16491), .ZN(U216) );
  AOI22_X1 U19476 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16458), .ZN(n16422) );
  OAI21_X1 U19477 ( .B1(n14459), .B2(n16461), .A(n16422), .ZN(U217) );
  AOI22_X1 U19478 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16458), .ZN(n16423) );
  OAI21_X1 U19479 ( .B1(n14464), .B2(n16461), .A(n16423), .ZN(U218) );
  AOI22_X1 U19480 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16458), .ZN(n16424) );
  OAI21_X1 U19481 ( .B1(n14470), .B2(n16461), .A(n16424), .ZN(U219) );
  AOI22_X1 U19482 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16458), .ZN(n16425) );
  OAI21_X1 U19483 ( .B1(n16426), .B2(n16461), .A(n16425), .ZN(U220) );
  AOI22_X1 U19484 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16458), .ZN(n16427) );
  OAI21_X1 U19485 ( .B1(n14479), .B2(n16461), .A(n16427), .ZN(U221) );
  AOI22_X1 U19486 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16458), .ZN(n16428) );
  OAI21_X1 U19487 ( .B1(n14486), .B2(n16461), .A(n16428), .ZN(U222) );
  AOI22_X1 U19488 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16458), .ZN(n16429) );
  OAI21_X1 U19489 ( .B1(n14491), .B2(n16461), .A(n16429), .ZN(U223) );
  AOI222_X1 U19490 ( .A1(n16459), .A2(P1_DATAO_REG_23__SCAN_IN), .B1(n16456), 
        .B2(BUF1_REG_23__SCAN_IN), .C1(n16458), .C2(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n16430) );
  INV_X1 U19491 ( .A(n16430), .ZN(U224) );
  AOI22_X1 U19492 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16458), .ZN(n16431) );
  OAI21_X1 U19493 ( .B1(n14498), .B2(n16461), .A(n16431), .ZN(U225) );
  AOI22_X1 U19494 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16458), .ZN(n16432) );
  OAI21_X1 U19495 ( .B1(n14502), .B2(n16461), .A(n16432), .ZN(U226) );
  AOI22_X1 U19496 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16458), .ZN(n16433) );
  OAI21_X1 U19497 ( .B1(n14510), .B2(n16461), .A(n16433), .ZN(U227) );
  AOI22_X1 U19498 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16458), .ZN(n16434) );
  OAI21_X1 U19499 ( .B1(n14515), .B2(n16461), .A(n16434), .ZN(U228) );
  AOI22_X1 U19500 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16458), .ZN(n16435) );
  OAI21_X1 U19501 ( .B1(n14521), .B2(n16461), .A(n16435), .ZN(U229) );
  AOI22_X1 U19502 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16458), .ZN(n16436) );
  OAI21_X1 U19503 ( .B1(n14527), .B2(n16461), .A(n16436), .ZN(U230) );
  AOI22_X1 U19504 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16458), .ZN(n16437) );
  OAI21_X1 U19505 ( .B1(n14534), .B2(n16461), .A(n16437), .ZN(U231) );
  AOI22_X1 U19506 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16458), .ZN(n16438) );
  OAI21_X1 U19507 ( .B1(n13566), .B2(n16461), .A(n16438), .ZN(U232) );
  AOI22_X1 U19508 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16458), .ZN(n16439) );
  OAI21_X1 U19509 ( .B1(n14042), .B2(n16461), .A(n16439), .ZN(U233) );
  AOI22_X1 U19510 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16458), .ZN(n16440) );
  OAI21_X1 U19511 ( .B1(n14051), .B2(n16461), .A(n16440), .ZN(U234) );
  AOI22_X1 U19512 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16458), .ZN(n16441) );
  OAI21_X1 U19513 ( .B1(n16442), .B2(n16461), .A(n16441), .ZN(U235) );
  AOI22_X1 U19514 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16458), .ZN(n16443) );
  OAI21_X1 U19515 ( .B1(n14083), .B2(n16461), .A(n16443), .ZN(U236) );
  AOI22_X1 U19516 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16458), .ZN(n16444) );
  OAI21_X1 U19517 ( .B1(n16445), .B2(n16461), .A(n16444), .ZN(U237) );
  INV_X1 U19518 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n20776) );
  AOI22_X1 U19519 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16456), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16459), .ZN(n16446) );
  OAI21_X1 U19520 ( .B1(n20776), .B2(U212), .A(n16446), .ZN(U238) );
  INV_X1 U19521 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16448) );
  AOI22_X1 U19522 ( .A1(BUF1_REG_8__SCAN_IN), .A2(n16456), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16459), .ZN(n16447) );
  OAI21_X1 U19523 ( .B1(n16448), .B2(U212), .A(n16447), .ZN(U239) );
  INV_X1 U19524 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16467) );
  AOI22_X1 U19525 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16456), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16459), .ZN(n16449) );
  OAI21_X1 U19526 ( .B1(n16467), .B2(U212), .A(n16449), .ZN(U240) );
  AOI222_X1 U19527 ( .A1(n16459), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n16456), 
        .B2(BUF1_REG_6__SCAN_IN), .C1(n16458), .C2(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n16450) );
  INV_X1 U19528 ( .A(n16450), .ZN(U241) );
  INV_X1 U19529 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n20825) );
  AOI22_X1 U19530 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16458), .ZN(n16451) );
  OAI21_X1 U19531 ( .B1(n20825), .B2(n16461), .A(n16451), .ZN(U242) );
  AOI22_X1 U19532 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16458), .ZN(n16452) );
  OAI21_X1 U19533 ( .B1(n16453), .B2(n16461), .A(n16452), .ZN(U243) );
  INV_X1 U19534 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n20838) );
  AOI22_X1 U19535 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16456), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16459), .ZN(n16454) );
  OAI21_X1 U19536 ( .B1(n20838), .B2(U212), .A(n16454), .ZN(U244) );
  AOI222_X1 U19537 ( .A1(n16458), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n16456), 
        .B2(BUF1_REG_2__SCAN_IN), .C1(n16459), .C2(P1_DATAO_REG_2__SCAN_IN), 
        .ZN(n16455) );
  INV_X1 U19538 ( .A(n16455), .ZN(U245) );
  INV_X1 U19539 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16464) );
  AOI22_X1 U19540 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16456), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16459), .ZN(n16457) );
  OAI21_X1 U19541 ( .B1(n16464), .B2(U212), .A(n16457), .ZN(U246) );
  INV_X1 U19542 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16462) );
  AOI22_X1 U19543 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16458), .ZN(n16460) );
  OAI21_X1 U19544 ( .B1(n16462), .B2(n16461), .A(n16460), .ZN(U247) );
  OAI22_X1 U19545 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16488), .ZN(n16463) );
  INV_X1 U19546 ( .A(n16463), .ZN(U251) );
  INV_X1 U19547 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18156) );
  AOI22_X1 U19548 ( .A1(n16490), .A2(n16464), .B1(n18156), .B2(U215), .ZN(U252) );
  INV_X1 U19549 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n19146) );
  INV_X1 U19550 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18162) );
  AOI22_X1 U19551 ( .A1(n16490), .A2(n19146), .B1(n18162), .B2(U215), .ZN(U253) );
  INV_X1 U19552 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18167) );
  AOI22_X1 U19553 ( .A1(n16490), .A2(n20838), .B1(n18167), .B2(U215), .ZN(U254) );
  OAI22_X1 U19554 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16490), .ZN(n16465) );
  INV_X1 U19555 ( .A(n16465), .ZN(U255) );
  OAI22_X1 U19556 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16490), .ZN(n16466) );
  INV_X1 U19557 ( .A(n16466), .ZN(U256) );
  INV_X1 U19558 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n20858) );
  INV_X1 U19559 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18186) );
  AOI22_X1 U19560 ( .A1(n16490), .A2(n20858), .B1(n18186), .B2(U215), .ZN(U257) );
  INV_X1 U19561 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18191) );
  AOI22_X1 U19562 ( .A1(n16490), .A2(n16467), .B1(n18191), .B2(U215), .ZN(U258) );
  OAI22_X1 U19563 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16490), .ZN(n16468) );
  INV_X1 U19564 ( .A(n16468), .ZN(U259) );
  INV_X1 U19565 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17441) );
  AOI22_X1 U19566 ( .A1(n16490), .A2(n20776), .B1(n17441), .B2(U215), .ZN(U260) );
  OAI22_X1 U19567 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16490), .ZN(n16469) );
  INV_X1 U19568 ( .A(n16469), .ZN(U261) );
  OAI22_X1 U19569 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16490), .ZN(n16470) );
  INV_X1 U19570 ( .A(n16470), .ZN(U262) );
  OAI22_X1 U19571 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16490), .ZN(n16471) );
  INV_X1 U19572 ( .A(n16471), .ZN(U263) );
  OAI22_X1 U19573 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16490), .ZN(n16472) );
  INV_X1 U19574 ( .A(n16472), .ZN(U264) );
  OAI22_X1 U19575 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16490), .ZN(n16473) );
  INV_X1 U19576 ( .A(n16473), .ZN(U265) );
  OAI22_X1 U19577 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16490), .ZN(n16474) );
  INV_X1 U19578 ( .A(n16474), .ZN(U266) );
  OAI22_X1 U19579 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16490), .ZN(n16475) );
  INV_X1 U19580 ( .A(n16475), .ZN(U267) );
  OAI22_X1 U19581 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16488), .ZN(n16476) );
  INV_X1 U19582 ( .A(n16476), .ZN(U268) );
  OAI22_X1 U19583 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16490), .ZN(n16477) );
  INV_X1 U19584 ( .A(n16477), .ZN(U269) );
  OAI22_X1 U19585 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16488), .ZN(n16478) );
  INV_X1 U19586 ( .A(n16478), .ZN(U270) );
  OAI22_X1 U19587 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16490), .ZN(n16479) );
  INV_X1 U19588 ( .A(n16479), .ZN(U271) );
  OAI22_X1 U19589 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16488), .ZN(n16480) );
  INV_X1 U19590 ( .A(n16480), .ZN(U272) );
  OAI22_X1 U19591 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16490), .ZN(n16481) );
  INV_X1 U19592 ( .A(n16481), .ZN(U273) );
  INV_X1 U19593 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n20790) );
  INV_X1 U19594 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n19218) );
  AOI22_X1 U19595 ( .A1(n16490), .A2(n20790), .B1(n19218), .B2(U215), .ZN(U274) );
  OAI22_X1 U19596 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16490), .ZN(n16482) );
  INV_X1 U19597 ( .A(n16482), .ZN(U275) );
  OAI22_X1 U19598 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16488), .ZN(n16483) );
  INV_X1 U19599 ( .A(n16483), .ZN(U276) );
  OAI22_X1 U19600 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16488), .ZN(n16484) );
  INV_X1 U19601 ( .A(n16484), .ZN(U277) );
  OAI22_X1 U19602 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16488), .ZN(n16485) );
  INV_X1 U19603 ( .A(n16485), .ZN(U278) );
  OAI22_X1 U19604 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16488), .ZN(n16486) );
  INV_X1 U19605 ( .A(n16486), .ZN(U279) );
  OAI22_X1 U19606 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16488), .ZN(n16487) );
  INV_X1 U19607 ( .A(n16487), .ZN(U280) );
  OAI22_X1 U19608 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16488), .ZN(n16489) );
  INV_X1 U19609 ( .A(n16489), .ZN(U281) );
  INV_X1 U19610 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n20856) );
  AOI22_X1 U19611 ( .A1(n16490), .A2(n19120), .B1(n20856), .B2(U215), .ZN(U282) );
  INV_X1 U19612 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17349) );
  AOI222_X1 U19613 ( .A1(n16491), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19120), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n17349), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16492) );
  INV_X2 U19614 ( .A(n16494), .ZN(n16493) );
  INV_X1 U19615 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18704) );
  INV_X1 U19616 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19758) );
  AOI22_X1 U19617 ( .A1(n16493), .A2(n18704), .B1(n19758), .B2(n16494), .ZN(
        U347) );
  INV_X1 U19618 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18702) );
  INV_X1 U19619 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19756) );
  AOI22_X1 U19620 ( .A1(n16493), .A2(n18702), .B1(n19756), .B2(n16494), .ZN(
        U348) );
  INV_X1 U19621 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18699) );
  INV_X1 U19622 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19754) );
  AOI22_X1 U19623 ( .A1(n16493), .A2(n18699), .B1(n19754), .B2(n16494), .ZN(
        U349) );
  INV_X1 U19624 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18698) );
  INV_X1 U19625 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19752) );
  AOI22_X1 U19626 ( .A1(n16493), .A2(n18698), .B1(n19752), .B2(n16494), .ZN(
        U350) );
  INV_X1 U19627 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18696) );
  INV_X1 U19628 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19750) );
  AOI22_X1 U19629 ( .A1(n16493), .A2(n18696), .B1(n19750), .B2(n16494), .ZN(
        U351) );
  INV_X1 U19630 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18693) );
  INV_X1 U19631 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20810) );
  AOI22_X1 U19632 ( .A1(n16493), .A2(n18693), .B1(n20810), .B2(n16494), .ZN(
        U352) );
  INV_X1 U19633 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18692) );
  INV_X1 U19634 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19747) );
  AOI22_X1 U19635 ( .A1(n16493), .A2(n18692), .B1(n19747), .B2(n16494), .ZN(
        U353) );
  INV_X1 U19636 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18690) );
  AOI22_X1 U19637 ( .A1(n16493), .A2(n18690), .B1(n19745), .B2(n16494), .ZN(
        U354) );
  INV_X1 U19638 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18745) );
  INV_X1 U19639 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19791) );
  AOI22_X1 U19640 ( .A1(n16493), .A2(n18745), .B1(n19791), .B2(n16494), .ZN(
        U355) );
  INV_X1 U19641 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18742) );
  INV_X1 U19642 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20865) );
  AOI22_X1 U19643 ( .A1(n16493), .A2(n18742), .B1(n20865), .B2(n16494), .ZN(
        U356) );
  INV_X1 U19644 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18738) );
  INV_X1 U19645 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19788) );
  AOI22_X1 U19646 ( .A1(n16493), .A2(n18738), .B1(n19788), .B2(n16494), .ZN(
        U357) );
  INV_X1 U19647 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18737) );
  INV_X1 U19648 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19785) );
  AOI22_X1 U19649 ( .A1(n16493), .A2(n18737), .B1(n19785), .B2(n16494), .ZN(
        U358) );
  INV_X1 U19650 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20868) );
  INV_X1 U19651 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19784) );
  AOI22_X1 U19652 ( .A1(n16493), .A2(n20868), .B1(n19784), .B2(n16494), .ZN(
        U359) );
  INV_X1 U19653 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18734) );
  INV_X1 U19654 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19782) );
  AOI22_X1 U19655 ( .A1(n16493), .A2(n18734), .B1(n19782), .B2(n16494), .ZN(
        U360) );
  INV_X1 U19656 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18732) );
  INV_X1 U19657 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19780) );
  AOI22_X1 U19658 ( .A1(n16493), .A2(n18732), .B1(n19780), .B2(n16494), .ZN(
        U361) );
  INV_X1 U19659 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18729) );
  INV_X1 U19660 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19778) );
  AOI22_X1 U19661 ( .A1(n16493), .A2(n18729), .B1(n19778), .B2(n16494), .ZN(
        U362) );
  INV_X1 U19662 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18728) );
  INV_X1 U19663 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19776) );
  AOI22_X1 U19664 ( .A1(n16493), .A2(n18728), .B1(n19776), .B2(n16494), .ZN(
        U363) );
  INV_X1 U19665 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18725) );
  INV_X1 U19666 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19775) );
  AOI22_X1 U19667 ( .A1(n16493), .A2(n18725), .B1(n19775), .B2(n16494), .ZN(
        U364) );
  INV_X1 U19668 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18688) );
  INV_X1 U19669 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19743) );
  AOI22_X1 U19670 ( .A1(n16493), .A2(n18688), .B1(n19743), .B2(n16494), .ZN(
        U365) );
  INV_X1 U19671 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18724) );
  INV_X1 U19672 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19773) );
  AOI22_X1 U19673 ( .A1(n16493), .A2(n18724), .B1(n19773), .B2(n16494), .ZN(
        U366) );
  INV_X1 U19674 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18721) );
  INV_X1 U19675 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20783) );
  AOI22_X1 U19676 ( .A1(n16493), .A2(n18721), .B1(n20783), .B2(n16494), .ZN(
        U367) );
  INV_X1 U19677 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18720) );
  INV_X1 U19678 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19770) );
  AOI22_X1 U19679 ( .A1(n16493), .A2(n18720), .B1(n19770), .B2(n16494), .ZN(
        U368) );
  INV_X1 U19680 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18717) );
  INV_X1 U19681 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19768) );
  AOI22_X1 U19682 ( .A1(n16493), .A2(n18717), .B1(n19768), .B2(n16494), .ZN(
        U369) );
  INV_X1 U19683 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18716) );
  INV_X1 U19684 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19766) );
  AOI22_X1 U19685 ( .A1(n16493), .A2(n18716), .B1(n19766), .B2(n16494), .ZN(
        U370) );
  INV_X1 U19686 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18714) );
  INV_X1 U19687 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20873) );
  AOI22_X1 U19688 ( .A1(n16493), .A2(n18714), .B1(n20873), .B2(n16494), .ZN(
        U371) );
  INV_X1 U19689 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18711) );
  INV_X1 U19690 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19764) );
  AOI22_X1 U19691 ( .A1(n16493), .A2(n18711), .B1(n19764), .B2(n16494), .ZN(
        U372) );
  INV_X1 U19692 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18710) );
  INV_X1 U19693 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19762) );
  AOI22_X1 U19694 ( .A1(n16493), .A2(n18710), .B1(n19762), .B2(n16494), .ZN(
        U373) );
  INV_X1 U19695 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18708) );
  INV_X1 U19696 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19761) );
  AOI22_X1 U19697 ( .A1(n16493), .A2(n18708), .B1(n19761), .B2(n16494), .ZN(
        U374) );
  INV_X1 U19698 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18706) );
  INV_X1 U19699 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19759) );
  AOI22_X1 U19700 ( .A1(n16493), .A2(n18706), .B1(n19759), .B2(n16494), .ZN(
        U375) );
  INV_X1 U19701 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18686) );
  INV_X1 U19702 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19741) );
  AOI22_X1 U19703 ( .A1(n16493), .A2(n18686), .B1(n19741), .B2(n16494), .ZN(
        U376) );
  INV_X1 U19704 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18685) );
  NAND2_X1 U19705 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18685), .ZN(n18677) );
  NOR2_X1 U19706 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n16498) );
  INV_X1 U19707 ( .A(n16498), .ZN(n18669) );
  OAI21_X1 U19708 ( .B1(n18682), .B2(n18677), .A(n18669), .ZN(n18757) );
  AOI21_X1 U19709 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18757), .ZN(n16495) );
  INV_X1 U19710 ( .A(n16495), .ZN(P3_U2633) );
  NOR2_X1 U19711 ( .A1(n17408), .A2(n16496), .ZN(n16502) );
  OAI21_X1 U19712 ( .B1(n16502), .B2(n17409), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16497) );
  OAI21_X1 U19713 ( .B1(n18818), .B2(n18809), .A(n16497), .ZN(P3_U2634) );
  AOI22_X1 U19714 ( .A1(n16498), .A2(n18685), .B1(P3_D_C_N_REG_SCAN_IN), .B2(
        n18817), .ZN(n16499) );
  OAI21_X1 U19715 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n18817), .A(n16499), 
        .ZN(P3_U2635) );
  NOR2_X1 U19716 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18667) );
  OAI21_X1 U19717 ( .B1(n18667), .B2(BS16), .A(n18757), .ZN(n18755) );
  OAI21_X1 U19718 ( .B1(n18757), .B2(n16500), .A(n18755), .ZN(P3_U2636) );
  INV_X1 U19719 ( .A(n16501), .ZN(n16503) );
  NOR3_X1 U19720 ( .A1(n16504), .A2(n16503), .A3(n16502), .ZN(n18604) );
  NOR2_X1 U19721 ( .A1(n18604), .A2(n18657), .ZN(n18801) );
  OAI21_X1 U19722 ( .B1(n18801), .B2(n18140), .A(n9617), .ZN(P3_U2637) );
  NOR4_X1 U19723 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16508) );
  NOR4_X1 U19724 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16507) );
  NOR4_X1 U19725 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16506) );
  NOR4_X1 U19726 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16505) );
  NAND4_X1 U19727 ( .A1(n16508), .A2(n16507), .A3(n16506), .A4(n16505), .ZN(
        n16514) );
  NOR4_X1 U19728 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16512) );
  AOI211_X1 U19729 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16511) );
  NOR4_X1 U19730 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16510) );
  NOR4_X1 U19731 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16509) );
  NAND4_X1 U19732 ( .A1(n16512), .A2(n16511), .A3(n16510), .A4(n16509), .ZN(
        n16513) );
  NOR2_X1 U19733 ( .A1(n16514), .A2(n16513), .ZN(n18794) );
  INV_X1 U19734 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16516) );
  NOR3_X1 U19735 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16517) );
  OAI21_X1 U19736 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16517), .A(n18794), .ZN(
        n16515) );
  OAI21_X1 U19737 ( .B1(n18794), .B2(n16516), .A(n16515), .ZN(P3_U2638) );
  INV_X1 U19738 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n20843) );
  INV_X1 U19739 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18756) );
  AOI21_X1 U19740 ( .B1(n20843), .B2(n18756), .A(n16517), .ZN(n16519) );
  INV_X1 U19741 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16518) );
  INV_X1 U19742 ( .A(n18794), .ZN(n18797) );
  AOI22_X1 U19743 ( .A1(n18794), .A2(n16519), .B1(n16518), .B2(n18797), .ZN(
        P3_U2639) );
  NAND4_X1 U19744 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16555), .ZN(n16527) );
  NOR3_X1 U19745 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18746), .A3(n16527), 
        .ZN(n16521) );
  AOI21_X1 U19746 ( .B1(n16881), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16521), .ZN(
        n16533) );
  NAND2_X1 U19747 ( .A1(n16572), .A2(n16927), .ZN(n16571) );
  NOR2_X1 U19748 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16571), .ZN(n16556) );
  NAND2_X1 U19749 ( .A1(n16556), .A2(n16923), .ZN(n16535) );
  NOR2_X1 U19750 ( .A1(n16849), .A2(n16535), .ZN(n16542) );
  INV_X1 U19751 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16531) );
  INV_X1 U19752 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17481) );
  NOR2_X1 U19753 ( .A1(n16524), .A2(n17481), .ZN(n16523) );
  OAI21_X1 U19754 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16523), .A(
        n16522), .ZN(n17466) );
  INV_X1 U19755 ( .A(n17466), .ZN(n16559) );
  AOI21_X1 U19756 ( .B1(n16524), .B2(n17481), .A(n16523), .ZN(n17477) );
  NOR2_X1 U19757 ( .A1(n9636), .A2(n9590), .ZN(n16567) );
  NOR2_X1 U19758 ( .A1(n17477), .A2(n16567), .ZN(n16566) );
  NOR2_X1 U19759 ( .A1(n9637), .A2(n9590), .ZN(n16536) );
  NOR2_X1 U19760 ( .A1(n9590), .A2(n16824), .ZN(n16856) );
  INV_X1 U19761 ( .A(n16856), .ZN(n16702) );
  NOR3_X1 U19762 ( .A1(n16537), .A2(n16536), .A3(n16702), .ZN(n16530) );
  NAND3_X1 U19763 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16526) );
  NOR2_X1 U19764 ( .A1(n16872), .A2(n16869), .ZN(n16691) );
  INV_X1 U19765 ( .A(n16691), .ZN(n16883) );
  AOI21_X1 U19766 ( .B1(n16526), .B2(n16883), .A(n16525), .ZN(n16554) );
  NOR2_X1 U19767 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16527), .ZN(n16540) );
  INV_X1 U19768 ( .A(n16540), .ZN(n16528) );
  INV_X1 U19769 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18744) );
  AOI21_X1 U19770 ( .B1(n16554), .B2(n16528), .A(n18744), .ZN(n16529) );
  AOI211_X1 U19771 ( .C1(n16542), .C2(n16531), .A(n16530), .B(n16529), .ZN(
        n16532) );
  OAI211_X1 U19772 ( .C1(n16534), .C2(n16866), .A(n16533), .B(n16532), .ZN(
        P3_U2640) );
  NAND2_X1 U19773 ( .A1(n16880), .A2(n16535), .ZN(n16550) );
  XOR2_X1 U19774 ( .A(n16537), .B(n16536), .Z(n16541) );
  OAI22_X1 U19775 ( .A1(n16554), .A2(n18746), .B1(n16538), .B2(n16866), .ZN(
        n16539) );
  AOI211_X1 U19776 ( .C1(n16541), .C2(n18660), .A(n16540), .B(n16539), .ZN(
        n16544) );
  OAI21_X1 U19777 ( .B1(n16881), .B2(n16542), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16543) );
  OAI211_X1 U19778 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16550), .A(n16544), .B(
        n16543), .ZN(P3_U2641) );
  INV_X1 U19779 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18741) );
  AOI211_X1 U19780 ( .C1(n16546), .C2(n16545), .A(n9637), .B(n16824), .ZN(
        n16549) );
  NAND3_X1 U19781 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16555), .ZN(n16547) );
  OAI22_X1 U19782 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16547), .B1(n9753), 
        .B2(n16866), .ZN(n16548) );
  AOI211_X1 U19783 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16863), .A(n16549), .B(
        n16548), .ZN(n16553) );
  INV_X1 U19784 ( .A(n16550), .ZN(n16551) );
  OAI21_X1 U19785 ( .B1(n16556), .B2(n16923), .A(n16551), .ZN(n16552) );
  OAI211_X1 U19786 ( .C1(n16554), .C2(n18741), .A(n16553), .B(n16552), .ZN(
        P3_U2642) );
  NAND2_X1 U19787 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16555), .ZN(n16565) );
  AOI22_X1 U19788 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16875), .B1(
        n16881), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16564) );
  INV_X1 U19789 ( .A(n16555), .ZN(n16568) );
  OAI21_X1 U19790 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16568), .A(n16575), 
        .ZN(n16562) );
  AOI211_X1 U19791 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16571), .A(n16556), .B(
        n16849), .ZN(n16561) );
  AOI211_X1 U19792 ( .C1(n16559), .C2(n16558), .A(n16557), .B(n16824), .ZN(
        n16560) );
  AOI211_X1 U19793 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16562), .A(n16561), 
        .B(n16560), .ZN(n16563) );
  OAI211_X1 U19794 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16565), .A(n16564), 
        .B(n16563), .ZN(P3_U2643) );
  INV_X1 U19795 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18736) );
  AOI211_X1 U19796 ( .C1(n17477), .C2(n16567), .A(n16566), .B(n16824), .ZN(
        n16570) );
  OAI22_X1 U19797 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16568), .B1(n17481), 
        .B2(n16866), .ZN(n16569) );
  AOI211_X1 U19798 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16863), .A(n16570), .B(
        n16569), .ZN(n16574) );
  OAI211_X1 U19799 ( .C1(n16572), .C2(n16927), .A(n16880), .B(n16571), .ZN(
        n16573) );
  OAI211_X1 U19800 ( .C1(n16575), .C2(n18736), .A(n16574), .B(n16573), .ZN(
        P3_U2644) );
  INV_X1 U19801 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18731) );
  OAI21_X1 U19802 ( .B1(n16599), .B2(n16830), .A(n16884), .ZN(n16596) );
  AOI21_X1 U19803 ( .B1(n16872), .B2(n18731), .A(n16596), .ZN(n16587) );
  AOI211_X1 U19804 ( .C1(n16578), .C2(n16577), .A(n16576), .B(n16843), .ZN(
        n16582) );
  NAND2_X1 U19805 ( .A1(n16872), .A2(n18733), .ZN(n16579) );
  OAI22_X1 U19806 ( .A1(n16833), .A2(n16584), .B1(n16580), .B2(n16579), .ZN(
        n16581) );
  AOI211_X1 U19807 ( .C1(n16875), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16582), .B(n16581), .ZN(n16586) );
  OAI211_X1 U19808 ( .C1(n16589), .C2(n16584), .A(n16880), .B(n16583), .ZN(
        n16585) );
  OAI211_X1 U19809 ( .C1(n16587), .C2(n18733), .A(n16586), .B(n16585), .ZN(
        P3_U2646) );
  NOR2_X1 U19810 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16830), .ZN(n16588) );
  AOI22_X1 U19811 ( .A1(n16881), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16599), 
        .B2(n16588), .ZN(n16595) );
  AOI211_X1 U19812 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16604), .A(n16589), .B(
        n16849), .ZN(n16593) );
  AOI211_X1 U19813 ( .C1(n17513), .C2(n16591), .A(n16590), .B(n16824), .ZN(
        n16592) );
  AOI211_X1 U19814 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16596), .A(n16593), 
        .B(n16592), .ZN(n16594) );
  OAI211_X1 U19815 ( .C1(n17517), .C2(n16866), .A(n16595), .B(n16594), .ZN(
        P3_U2647) );
  INV_X1 U19816 ( .A(n16596), .ZN(n16608) );
  AOI211_X1 U19817 ( .C1(n17528), .C2(n16598), .A(n16597), .B(n16824), .ZN(
        n16603) );
  OR2_X1 U19818 ( .A1(n16830), .A2(n16599), .ZN(n16600) );
  OAI22_X1 U19819 ( .A1(n16833), .A2(n16605), .B1(n16601), .B2(n16600), .ZN(
        n16602) );
  AOI211_X1 U19820 ( .C1(n16875), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16603), .B(n16602), .ZN(n16607) );
  OAI211_X1 U19821 ( .C1(n16611), .C2(n16605), .A(n16880), .B(n16604), .ZN(
        n16606) );
  OAI211_X1 U19822 ( .C1(n16608), .C2(n18730), .A(n16607), .B(n16606), .ZN(
        P3_U2648) );
  NOR2_X1 U19823 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16830), .ZN(n16609) );
  AOI22_X1 U19824 ( .A1(n16881), .A2(P3_EBX_REG_22__SCAN_IN), .B1(n16610), 
        .B2(n16609), .ZN(n16617) );
  OAI21_X1 U19825 ( .B1(n16610), .B2(n16830), .A(n16884), .ZN(n16625) );
  AOI211_X1 U19826 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16626), .A(n16611), .B(
        n16849), .ZN(n16615) );
  AOI211_X1 U19827 ( .C1(n17545), .C2(n16613), .A(n16612), .B(n16824), .ZN(
        n16614) );
  AOI211_X1 U19828 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16625), .A(n16615), 
        .B(n16614), .ZN(n16616) );
  OAI211_X1 U19829 ( .C1(n16618), .C2(n16866), .A(n16617), .B(n16616), .ZN(
        P3_U2649) );
  AOI22_X1 U19830 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16875), .B1(
        n16881), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n16629) );
  OAI21_X1 U19831 ( .B1(n16830), .B2(n16619), .A(n18726), .ZN(n16624) );
  AOI211_X1 U19832 ( .C1(n16622), .C2(n16621), .A(n16620), .B(n16843), .ZN(
        n16623) );
  AOI21_X1 U19833 ( .B1(n16625), .B2(n16624), .A(n16623), .ZN(n16628) );
  OAI211_X1 U19834 ( .C1(n16630), .C2(n16977), .A(n16880), .B(n16626), .ZN(
        n16627) );
  NAND3_X1 U19835 ( .A1(n16629), .A2(n16628), .A3(n16627), .ZN(P3_U2650) );
  AOI22_X1 U19836 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16875), .B1(
        n16881), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n16640) );
  NOR2_X1 U19837 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16830), .ZN(n16635) );
  AOI211_X1 U19838 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16650), .A(n16630), .B(
        n16849), .ZN(n16634) );
  AOI211_X1 U19839 ( .C1(n17570), .C2(n16632), .A(n16631), .B(n16843), .ZN(
        n16633) );
  AOI211_X1 U19840 ( .C1(n16636), .C2(n16635), .A(n16634), .B(n16633), .ZN(
        n16639) );
  NOR2_X1 U19841 ( .A1(n16869), .A2(n16677), .ZN(n16690) );
  INV_X1 U19842 ( .A(n16690), .ZN(n16678) );
  OAI211_X1 U19843 ( .C1(n16637), .C2(n16678), .A(P3_REIP_REG_20__SCAN_IN), 
        .B(n16883), .ZN(n16638) );
  NAND3_X1 U19844 ( .A1(n16640), .A2(n16639), .A3(n16638), .ZN(P3_U2651) );
  AOI22_X1 U19845 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n16875), .B1(
        n16881), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n16653) );
  AOI21_X1 U19846 ( .B1(n16641), .B2(n16690), .A(n16691), .ZN(n16671) );
  INV_X1 U19847 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18722) );
  INV_X1 U19848 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18719) );
  NOR3_X1 U19849 ( .A1(n16830), .A2(n16677), .A3(n16679), .ZN(n16670) );
  NAND2_X1 U19850 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16670), .ZN(n16664) );
  AOI221_X1 U19851 ( .B1(P3_REIP_REG_19__SCAN_IN), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n18722), .C2(n18719), .A(n16664), .ZN(n16649) );
  INV_X1 U19852 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17591) );
  NAND2_X1 U19853 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16642), .ZN(
        n16656) );
  NOR2_X1 U19854 ( .A1(n17591), .A2(n16656), .ZN(n16645) );
  INV_X1 U19855 ( .A(n16645), .ZN(n16655) );
  NOR2_X1 U19856 ( .A1(n16643), .A2(n9590), .ZN(n16694) );
  AOI21_X1 U19857 ( .B1(n16838), .B2(n16655), .A(n16694), .ZN(n16647) );
  OAI21_X1 U19858 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16645), .A(
        n16644), .ZN(n17582) );
  OAI21_X1 U19859 ( .B1(n16647), .B2(n17582), .A(n18660), .ZN(n16646) );
  AOI21_X1 U19860 ( .B1(n16647), .B2(n17582), .A(n16646), .ZN(n16648) );
  AOI211_X1 U19861 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n16671), .A(n16649), 
        .B(n16648), .ZN(n16652) );
  OAI211_X1 U19862 ( .C1(n16654), .C2(n16993), .A(n16880), .B(n16650), .ZN(
        n16651) );
  NAND4_X1 U19863 ( .A1(n16653), .A2(n16652), .A3(n18137), .A4(n16651), .ZN(
        P3_U2652) );
  INV_X1 U19864 ( .A(n16671), .ZN(n16663) );
  AOI211_X1 U19865 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16672), .A(n16654), .B(
        n16849), .ZN(n16661) );
  INV_X1 U19866 ( .A(n16656), .ZN(n17576) );
  OAI21_X1 U19867 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17576), .A(
        n16655), .ZN(n17588) );
  OAI21_X1 U19868 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16656), .A(
        n16838), .ZN(n16658) );
  AOI21_X1 U19869 ( .B1(n17588), .B2(n16658), .A(n16843), .ZN(n16657) );
  OAI21_X1 U19870 ( .B1(n17588), .B2(n16658), .A(n16657), .ZN(n16659) );
  OAI211_X1 U19871 ( .C1(n16833), .C2(n9734), .A(n18137), .B(n16659), .ZN(
        n16660) );
  AOI211_X1 U19872 ( .C1(n16875), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16661), .B(n16660), .ZN(n16662) );
  OAI221_X1 U19873 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16664), .C1(n18719), 
        .C2(n16663), .A(n16662), .ZN(P3_U2653) );
  INV_X1 U19874 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17601) );
  NAND3_X1 U19875 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A3(n17616), .ZN(n16680) );
  AOI21_X1 U19876 ( .B1(n17601), .B2(n16680), .A(n17576), .ZN(n17606) );
  NOR2_X1 U19877 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17823), .ZN(
        n16857) );
  AOI21_X1 U19878 ( .B1(n16665), .B2(n16857), .A(n9590), .ZN(n16667) );
  AOI21_X1 U19879 ( .B1(n17606), .B2(n16667), .A(n16843), .ZN(n16666) );
  OAI21_X1 U19880 ( .B1(n17606), .B2(n16667), .A(n16666), .ZN(n16668) );
  OAI211_X1 U19881 ( .C1(n17601), .C2(n16866), .A(n18137), .B(n16668), .ZN(
        n16669) );
  AOI221_X1 U19882 ( .B1(n16671), .B2(P3_REIP_REG_17__SCAN_IN), .C1(n16670), 
        .C2(n18718), .A(n16669), .ZN(n16674) );
  OAI211_X1 U19883 ( .C1(n16676), .C2(n16675), .A(n16880), .B(n16672), .ZN(
        n16673) );
  OAI211_X1 U19884 ( .C1(n16675), .C2(n16833), .A(n16674), .B(n16673), .ZN(
        P3_U2654) );
  AOI211_X1 U19885 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16695), .A(n16676), .B(
        n16849), .ZN(n16686) );
  NOR2_X1 U19886 ( .A1(n16830), .A2(n16677), .ZN(n16693) );
  AOI21_X1 U19887 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16693), .A(
        P3_REIP_REG_16__SCAN_IN), .ZN(n16684) );
  OAI21_X1 U19888 ( .B1(n16679), .B2(n16678), .A(n16883), .ZN(n16683) );
  OAI21_X1 U19889 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16681), .A(
        n16680), .ZN(n17621) );
  XOR2_X1 U19890 ( .A(n16694), .B(n17621), .Z(n16682) );
  OAI22_X1 U19891 ( .A1(n16684), .A2(n16683), .B1(n16824), .B2(n16682), .ZN(
        n16685) );
  AOI211_X1 U19892 ( .C1(n16875), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16686), .B(n16685), .ZN(n16687) );
  OAI211_X1 U19893 ( .C1(n16833), .C2(n17038), .A(n16687), .B(n18137), .ZN(
        P3_U2655) );
  OAI21_X1 U19894 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17616), .A(
        n16688), .ZN(n17627) );
  AOI21_X1 U19895 ( .B1(n16838), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16843), .ZN(n16870) );
  INV_X1 U19896 ( .A(n16870), .ZN(n16799) );
  AOI211_X1 U19897 ( .C1(n16838), .C2(n16703), .A(n17627), .B(n16799), .ZN(
        n16689) );
  NOR2_X1 U19898 ( .A1(n9577), .A2(n16689), .ZN(n16700) );
  NOR2_X1 U19899 ( .A1(n16691), .A2(n16690), .ZN(n16709) );
  INV_X1 U19900 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18713) );
  OAI22_X1 U19901 ( .A1(n17630), .A2(n16866), .B1(n16833), .B2(n16696), .ZN(
        n16692) );
  AOI221_X1 U19902 ( .B1(n16709), .B2(P3_REIP_REG_15__SCAN_IN), .C1(n16693), 
        .C2(n18713), .A(n16692), .ZN(n16699) );
  NAND3_X1 U19903 ( .A1(n18660), .A2(n16694), .A3(n17627), .ZN(n16698) );
  OAI211_X1 U19904 ( .C1(n16706), .C2(n16696), .A(n16880), .B(n16695), .ZN(
        n16697) );
  NAND4_X1 U19905 ( .A1(n16700), .A2(n16699), .A3(n16698), .A4(n16697), .ZN(
        P3_U2656) );
  NOR2_X1 U19906 ( .A1(n16701), .A2(n17663), .ZN(n16714) );
  INV_X1 U19907 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20887) );
  AOI21_X1 U19908 ( .B1(n16714), .B2(n20887), .A(n16702), .ZN(n16719) );
  OAI21_X1 U19909 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16714), .A(
        n16703), .ZN(n17649) );
  AOI21_X1 U19910 ( .B1(n16719), .B2(n17649), .A(n9577), .ZN(n16713) );
  NAND2_X1 U19911 ( .A1(n16714), .A2(n20887), .ZN(n16704) );
  AOI211_X1 U19912 ( .C1(n16838), .C2(n16704), .A(n16843), .B(n17649), .ZN(
        n16705) );
  AOI21_X1 U19913 ( .B1(n16875), .B2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16705), .ZN(n16712) );
  AOI211_X1 U19914 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16724), .A(n16706), .B(
        n16849), .ZN(n16707) );
  AOI21_X1 U19915 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n16881), .A(n16707), .ZN(
        n16711) );
  AND2_X1 U19916 ( .A1(n16872), .A2(n16708), .ZN(n16718) );
  OAI221_X1 U19917 ( .B1(P3_REIP_REG_14__SCAN_IN), .B2(P3_REIP_REG_13__SCAN_IN), .C1(P3_REIP_REG_14__SCAN_IN), .C2(n16718), .A(n16709), .ZN(n16710) );
  NAND4_X1 U19918 ( .A1(n16713), .A2(n16712), .A3(n16711), .A4(n16710), .ZN(
        P3_U2657) );
  INV_X1 U19919 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17667) );
  INV_X1 U19920 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17677) );
  NOR2_X1 U19921 ( .A1(n17677), .A2(n17663), .ZN(n16729) );
  INV_X1 U19922 ( .A(n16729), .ZN(n16716) );
  AOI21_X1 U19923 ( .B1(n17667), .B2(n16716), .A(n16714), .ZN(n16715) );
  INV_X1 U19924 ( .A(n16715), .ZN(n17665) );
  AOI211_X1 U19925 ( .C1(n16838), .C2(n16716), .A(n17665), .B(n16799), .ZN(
        n16723) );
  AOI21_X1 U19926 ( .B1(n16872), .B2(n16732), .A(n16869), .ZN(n16741) );
  OAI21_X1 U19927 ( .B1(n16830), .B2(P3_REIP_REG_12__SCAN_IN), .A(n16741), 
        .ZN(n16717) );
  INV_X1 U19928 ( .A(n16717), .ZN(n16721) );
  INV_X1 U19929 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18709) );
  AOI22_X1 U19930 ( .A1(n16719), .A2(n17665), .B1(n16718), .B2(n18709), .ZN(
        n16720) );
  OAI211_X1 U19931 ( .C1(n16721), .C2(n18709), .A(n16720), .B(n18137), .ZN(
        n16722) );
  AOI211_X1 U19932 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n16881), .A(n16723), .B(
        n16722), .ZN(n16727) );
  OAI211_X1 U19933 ( .C1(n16728), .C2(n16725), .A(n16880), .B(n16724), .ZN(
        n16726) );
  OAI211_X1 U19934 ( .C1(n16866), .C2(n17667), .A(n16727), .B(n16726), .ZN(
        P3_U2658) );
  AOI21_X1 U19935 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n16875), .A(
        n9577), .ZN(n16737) );
  AOI211_X1 U19936 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16744), .A(n16728), .B(
        n16849), .ZN(n16735) );
  AOI21_X1 U19937 ( .B1(n17677), .B2(n17663), .A(n16729), .ZN(n17681) );
  OAI21_X1 U19938 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17663), .A(
        n16838), .ZN(n16730) );
  XOR2_X1 U19939 ( .A(n17681), .B(n16730), .Z(n16733) );
  NAND2_X1 U19940 ( .A1(n16872), .A2(n18707), .ZN(n16731) );
  OAI22_X1 U19941 ( .A1(n16843), .A2(n16733), .B1(n16732), .B2(n16731), .ZN(
        n16734) );
  AOI211_X1 U19942 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16863), .A(n16735), .B(
        n16734), .ZN(n16736) );
  OAI211_X1 U19943 ( .C1(n18707), .C2(n16741), .A(n16737), .B(n16736), .ZN(
        P3_U2659) );
  INV_X1 U19944 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18703) );
  INV_X1 U19945 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18701) );
  NOR2_X1 U19946 ( .A1(n18703), .A2(n18701), .ZN(n16756) );
  NOR4_X1 U19947 ( .A1(n16830), .A2(n18700), .A3(n16787), .A4(n16788), .ZN(
        n16765) );
  AOI21_X1 U19948 ( .B1(n16756), .B2(n16765), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16742) );
  INV_X1 U19949 ( .A(n16808), .ZN(n17770) );
  NOR2_X1 U19950 ( .A1(n17823), .A2(n17770), .ZN(n16821) );
  NAND2_X1 U19951 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n16821), .ZN(
        n16809) );
  INV_X1 U19952 ( .A(n16809), .ZN(n16798) );
  NAND2_X1 U19953 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16798), .ZN(
        n16797) );
  OAI21_X1 U19954 ( .B1(n16797), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16838), .ZN(n16785) );
  INV_X1 U19955 ( .A(n16785), .ZN(n16800) );
  AOI21_X1 U19956 ( .B1(n16838), .B2(n16738), .A(n16800), .ZN(n16739) );
  NAND2_X1 U19957 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17691) );
  NAND2_X1 U19958 ( .A1(n9684), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17729) );
  NOR2_X1 U19959 ( .A1(n17823), .A2(n17729), .ZN(n16784) );
  NAND2_X1 U19960 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16784), .ZN(
        n16773) );
  NOR2_X1 U19961 ( .A1(n17691), .A2(n16773), .ZN(n16752) );
  OAI21_X1 U19962 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16752), .A(
        n17663), .ZN(n17692) );
  XNOR2_X1 U19963 ( .A(n16739), .B(n17692), .ZN(n16740) );
  OAI22_X1 U19964 ( .A1(n16742), .A2(n16741), .B1(n16824), .B2(n16740), .ZN(
        n16743) );
  AOI211_X1 U19965 ( .C1(n16881), .C2(P3_EBX_REG_11__SCAN_IN), .A(n9577), .B(
        n16743), .ZN(n16747) );
  OAI211_X1 U19966 ( .C1(n16749), .C2(n16745), .A(n16880), .B(n16744), .ZN(
        n16746) );
  OAI211_X1 U19967 ( .C1(n16866), .C2(n16748), .A(n16747), .B(n16746), .ZN(
        P3_U2660) );
  AOI211_X1 U19968 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16750), .A(n16749), .B(
        n16849), .ZN(n16751) );
  AOI21_X1 U19969 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n16881), .A(n16751), .ZN(
        n16760) );
  INV_X1 U19970 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17714) );
  NOR2_X1 U19971 ( .A1(n17714), .A2(n16773), .ZN(n16766) );
  AOI21_X1 U19972 ( .B1(n16766), .B2(n20887), .A(n9590), .ZN(n16769) );
  INV_X1 U19973 ( .A(n16752), .ZN(n16753) );
  OAI21_X1 U19974 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16766), .A(
        n16753), .ZN(n17704) );
  XNOR2_X1 U19975 ( .A(n16769), .B(n17704), .ZN(n16754) );
  AOI22_X1 U19976 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16875), .B1(
        n18660), .B2(n16754), .ZN(n16759) );
  OAI21_X1 U19977 ( .B1(n16755), .B2(n16830), .A(n16884), .ZN(n16779) );
  AOI21_X1 U19978 ( .B1(n18703), .B2(n18701), .A(n16756), .ZN(n16757) );
  AOI22_X1 U19979 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n16779), .B1(n16765), 
        .B2(n16757), .ZN(n16758) );
  NAND4_X1 U19980 ( .A1(n16760), .A2(n16759), .A3(n16758), .A4(n18137), .ZN(
        P3_U2661) );
  NOR2_X1 U19981 ( .A1(n16761), .A2(n16849), .ZN(n16777) );
  AOI22_X1 U19982 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16875), .B1(
        n16777), .B2(n16762), .ZN(n16772) );
  INV_X1 U19983 ( .A(n16761), .ZN(n16763) );
  AOI221_X1 U19984 ( .B1(n16849), .B2(n16833), .C1(n16763), .C2(n16833), .A(
        n16762), .ZN(n16764) );
  AOI221_X1 U19985 ( .B1(n16779), .B2(P3_REIP_REG_9__SCAN_IN), .C1(n16765), 
        .C2(n18701), .A(n16764), .ZN(n16771) );
  AOI21_X1 U19986 ( .B1(n17714), .B2(n16773), .A(n16766), .ZN(n17718) );
  NAND2_X1 U19987 ( .A1(n9590), .A2(n18660), .ZN(n16860) );
  INV_X1 U19988 ( .A(n16860), .ZN(n16768) );
  AOI221_X1 U19989 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17718), .C1(
        n16773), .C2(n17718), .A(n16843), .ZN(n16767) );
  OAI22_X1 U19990 ( .A1(n17718), .A2(n16769), .B1(n16768), .B2(n16767), .ZN(
        n16770) );
  NAND4_X1 U19991 ( .A1(n16772), .A2(n16771), .A3(n18137), .A4(n16770), .ZN(
        P3_U2662) );
  AOI21_X1 U19992 ( .B1(n16784), .B2(n20887), .A(n9590), .ZN(n16774) );
  OAI21_X1 U19993 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16784), .A(
        n16773), .ZN(n17742) );
  XOR2_X1 U19994 ( .A(n16774), .B(n17742), .Z(n16775) );
  OAI22_X1 U19995 ( .A1(n16833), .A2(n17159), .B1(n16824), .B2(n16775), .ZN(
        n16776) );
  AOI211_X1 U19996 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n16875), .A(
        n9577), .B(n16776), .ZN(n16783) );
  INV_X1 U19997 ( .A(n16792), .ZN(n16778) );
  OAI21_X1 U19998 ( .B1(n16778), .B2(n17159), .A(n16777), .ZN(n16782) );
  NOR3_X1 U19999 ( .A1(n16830), .A2(n16787), .A3(n16788), .ZN(n16780) );
  OAI21_X1 U20000 ( .B1(P3_REIP_REG_8__SCAN_IN), .B2(n16780), .A(n16779), .ZN(
        n16781) );
  NAND3_X1 U20001 ( .A1(n16783), .A2(n16782), .A3(n16781), .ZN(P3_U2663) );
  INV_X1 U20002 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17748) );
  AOI21_X1 U20003 ( .B1(n16872), .B2(n16787), .A(n16869), .ZN(n16811) );
  INV_X1 U20004 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18697) );
  AOI21_X1 U20005 ( .B1(n17748), .B2(n16797), .A(n16784), .ZN(n17752) );
  INV_X1 U20006 ( .A(n17752), .ZN(n16786) );
  OAI221_X1 U20007 ( .B1(n17752), .B2(n16800), .C1(n16786), .C2(n16785), .A(
        n18660), .ZN(n16790) );
  NOR2_X1 U20008 ( .A1(n16830), .A2(n16787), .ZN(n16804) );
  OAI211_X1 U20009 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(P3_REIP_REG_6__SCAN_IN), 
        .A(n16804), .B(n16788), .ZN(n16789) );
  OAI211_X1 U20010 ( .C1(n16811), .C2(n18697), .A(n16790), .B(n16789), .ZN(
        n16791) );
  AOI211_X1 U20011 ( .C1(n16881), .C2(P3_EBX_REG_7__SCAN_IN), .A(n9577), .B(
        n16791), .ZN(n16794) );
  OAI211_X1 U20012 ( .C1(n16795), .C2(n17163), .A(n16880), .B(n16792), .ZN(
        n16793) );
  OAI211_X1 U20013 ( .C1(n16866), .C2(n17748), .A(n16794), .B(n16793), .ZN(
        P3_U2664) );
  INV_X1 U20014 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18695) );
  AOI211_X1 U20015 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16814), .A(n16795), .B(
        n16849), .ZN(n16796) );
  AOI21_X1 U20016 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n16863), .A(n16796), .ZN(
        n16806) );
  OAI21_X1 U20017 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16798), .A(
        n16797), .ZN(n17763) );
  AOI211_X1 U20018 ( .C1(n16838), .C2(n16809), .A(n17763), .B(n16799), .ZN(
        n16803) );
  NAND3_X1 U20019 ( .A1(n18660), .A2(n16800), .A3(n17763), .ZN(n16801) );
  OAI211_X1 U20020 ( .C1(n17759), .C2(n16866), .A(n18137), .B(n16801), .ZN(
        n16802) );
  AOI211_X1 U20021 ( .C1(n16804), .C2(n18695), .A(n16803), .B(n16802), .ZN(
        n16805) );
  OAI211_X1 U20022 ( .C1(n18695), .C2(n16811), .A(n16806), .B(n16805), .ZN(
        P3_U2665) );
  AOI21_X1 U20023 ( .B1(n16872), .B2(n16807), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n16812) );
  AOI21_X1 U20024 ( .B1(n16808), .B2(n16857), .A(n9590), .ZN(n16823) );
  OAI21_X1 U20025 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16821), .A(
        n16809), .ZN(n17775) );
  XOR2_X1 U20026 ( .A(n16823), .B(n17775), .Z(n16810) );
  OAI22_X1 U20027 ( .A1(n16812), .A2(n16811), .B1(n16824), .B2(n16810), .ZN(
        n16813) );
  AOI211_X1 U20028 ( .C1(n16881), .C2(P3_EBX_REG_5__SCAN_IN), .A(n9577), .B(
        n16813), .ZN(n16817) );
  OAI211_X1 U20029 ( .C1(n16818), .C2(n16815), .A(n16880), .B(n16814), .ZN(
        n16816) );
  OAI211_X1 U20030 ( .C1(n16866), .C2(n9757), .A(n16817), .B(n16816), .ZN(
        P3_U2666) );
  INV_X1 U20031 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n16834) );
  AOI211_X1 U20032 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16819), .A(n16818), .B(
        n16849), .ZN(n16829) );
  AOI21_X1 U20033 ( .B1(n16872), .B2(n16840), .A(n16869), .ZN(n16848) );
  NOR2_X1 U20034 ( .A1(n16820), .A2(n18821), .ZN(n16882) );
  NOR2_X1 U20035 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17787), .ZN(
        n17782) );
  OR2_X1 U20036 ( .A1(n17823), .A2(n17787), .ZN(n16837) );
  AOI21_X1 U20037 ( .B1(n17789), .B2(n16837), .A(n16821), .ZN(n16822) );
  INV_X1 U20038 ( .A(n16822), .ZN(n17790) );
  AOI22_X1 U20039 ( .A1(n16857), .A2(n17782), .B1(n16823), .B2(n17790), .ZN(
        n16825) );
  OAI22_X1 U20040 ( .A1(n16825), .A2(n16824), .B1(n17790), .B2(n16860), .ZN(
        n16826) );
  AOI221_X1 U20041 ( .B1(n17156), .B2(n16882), .C1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n16882), .A(n16826), .ZN(
        n16827) );
  OAI211_X1 U20042 ( .C1(n16848), .C2(n18691), .A(n16827), .B(n18137), .ZN(
        n16828) );
  AOI211_X1 U20043 ( .C1(n16875), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16829), .B(n16828), .ZN(n16832) );
  OR3_X1 U20044 ( .A1(n16830), .A2(n16840), .A3(P3_REIP_REG_4__SCAN_IN), .ZN(
        n16831) );
  OAI211_X1 U20045 ( .C1(n16834), .C2(n16833), .A(n16832), .B(n16831), .ZN(
        P3_U2667) );
  INV_X1 U20046 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18689) );
  AOI22_X1 U20047 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n16875), .B1(
        n16881), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n16847) );
  AOI21_X1 U20048 ( .B1(n18769), .B2(n18617), .A(n17156), .ZN(n18766) );
  AOI211_X1 U20049 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n16836), .A(n16835), .B(
        n16849), .ZN(n16845) );
  NAND2_X1 U20050 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16852) );
  INV_X1 U20051 ( .A(n16852), .ZN(n16854) );
  OAI21_X1 U20052 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n16854), .A(
        n16837), .ZN(n17799) );
  OAI21_X1 U20053 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16852), .A(
        n16838), .ZN(n16839) );
  XNOR2_X1 U20054 ( .A(n17799), .B(n16839), .ZN(n16842) );
  NAND2_X1 U20055 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16853) );
  NAND2_X1 U20056 ( .A1(n16872), .A2(n16840), .ZN(n16841) );
  OAI22_X1 U20057 ( .A1(n16843), .A2(n16842), .B1(n16853), .B2(n16841), .ZN(
        n16844) );
  AOI211_X1 U20058 ( .C1(n16882), .C2(n18766), .A(n16845), .B(n16844), .ZN(
        n16846) );
  OAI211_X1 U20059 ( .C1(n16848), .C2(n18689), .A(n16847), .B(n16846), .ZN(
        P3_U2668) );
  INV_X1 U20060 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17814) );
  NAND2_X1 U20061 ( .A1(n18777), .A2(n16868), .ZN(n18614) );
  AND2_X1 U20062 ( .A1(n18617), .A2(n18614), .ZN(n18773) );
  AOI22_X1 U20063 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n16869), .B1(n18773), 
        .B2(n16882), .ZN(n16865) );
  NOR2_X1 U20064 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16871) );
  INV_X1 U20065 ( .A(n16871), .ZN(n16851) );
  AOI211_X1 U20066 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16851), .A(n16850), .B(
        n16849), .ZN(n16862) );
  OAI21_X1 U20067 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16852), .ZN(n17810) );
  OAI211_X1 U20068 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16872), .B(n16853), .ZN(n16859) );
  NAND2_X1 U20069 ( .A1(n16854), .A2(n20887), .ZN(n16855) );
  OAI211_X1 U20070 ( .C1(n16857), .C2(n17810), .A(n16856), .B(n16855), .ZN(
        n16858) );
  OAI211_X1 U20071 ( .C1(n16860), .C2(n17810), .A(n16859), .B(n16858), .ZN(
        n16861) );
  AOI211_X1 U20072 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16863), .A(n16862), .B(
        n16861), .ZN(n16864) );
  OAI211_X1 U20073 ( .C1(n17814), .C2(n16866), .A(n16865), .B(n16864), .ZN(
        P3_U2669) );
  NAND2_X1 U20074 ( .A1(n16868), .A2(n16867), .ZN(n18632) );
  INV_X1 U20075 ( .A(n18632), .ZN(n18780) );
  AOI22_X1 U20076 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16869), .B1(n18780), 
        .B2(n16882), .ZN(n16879) );
  AOI22_X1 U20077 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(n16881), .B1(n16870), .B2(
        n17823), .ZN(n16878) );
  AOI21_X1 U20078 ( .B1(P3_EBX_REG_1__SCAN_IN), .B2(P3_EBX_REG_0__SCAN_IN), 
        .A(n16871), .ZN(n17183) );
  AOI22_X1 U20079 ( .A1(n16880), .A2(n17183), .B1(n16872), .B2(n20843), .ZN(
        n16877) );
  NOR2_X1 U20080 ( .A1(n9590), .A2(n20887), .ZN(n16874) );
  OAI221_X1 U20081 ( .B1(n16875), .B2(n16874), .C1(n16875), .C2(n18660), .A(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16876) );
  NAND4_X1 U20082 ( .A1(n16879), .A2(n16878), .A3(n16877), .A4(n16876), .ZN(
        P3_U2670) );
  NOR2_X1 U20083 ( .A1(n16881), .A2(n16880), .ZN(n16887) );
  INV_X1 U20084 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17190) );
  AOI22_X1 U20085 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16883), .B1(n16882), 
        .B2(n20806), .ZN(n16886) );
  INV_X1 U20086 ( .A(n18786), .ZN(n18763) );
  NAND3_X1 U20087 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18763), .A3(
        n16884), .ZN(n16885) );
  OAI211_X1 U20088 ( .C1(n16887), .C2(n17190), .A(n16886), .B(n16885), .ZN(
        P3_U2671) );
  NOR2_X1 U20089 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16888), .ZN(n16914) );
  AOI22_X1 U20090 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16898) );
  AOI22_X1 U20091 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n15648), .ZN(n16890) );
  AOI22_X1 U20092 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n9568), .ZN(n16889) );
  OAI211_X1 U20093 ( .C1(n17146), .C2(n18244), .A(n16890), .B(n16889), .ZN(
        n16896) );
  AOI22_X1 U20094 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17044), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16894) );
  AOI22_X1 U20095 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n17122), .ZN(n16893) );
  AOI22_X1 U20096 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n15684), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17143), .ZN(n16892) );
  NAND2_X1 U20097 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17149), .ZN(
        n16891) );
  NAND4_X1 U20098 ( .A1(n16894), .A2(n16893), .A3(n16892), .A4(n16891), .ZN(
        n16895) );
  AOI211_X1 U20099 ( .C1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .C2(n17156), .A(
        n16896), .B(n16895), .ZN(n16897) );
  OAI211_X1 U20100 ( .C1(n17041), .C2(n17108), .A(n16898), .B(n16897), .ZN(
        n16912) );
  AOI22_X1 U20101 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16910) );
  INV_X1 U20102 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16902) );
  AOI22_X1 U20103 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16901) );
  AOI22_X1 U20104 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16900) );
  OAI211_X1 U20105 ( .C1(n17090), .C2(n16902), .A(n16901), .B(n16900), .ZN(
        n16908) );
  AOI22_X1 U20106 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16906) );
  AOI22_X1 U20107 ( .A1(n15684), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16905) );
  AOI22_X1 U20108 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16904) );
  NAND2_X1 U20109 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n16903) );
  NAND4_X1 U20110 ( .A1(n16906), .A2(n16905), .A3(n16904), .A4(n16903), .ZN(
        n16907) );
  AOI211_X1 U20111 ( .C1(n17105), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n16908), .B(n16907), .ZN(n16909) );
  OAI211_X1 U20112 ( .C1(n12721), .C2(n18190), .A(n16910), .B(n16909), .ZN(
        n16917) );
  NAND3_X1 U20113 ( .A1(n16917), .A2(n16915), .A3(n16916), .ZN(n16911) );
  XOR2_X1 U20114 ( .A(n16912), .B(n16911), .Z(n17206) );
  OAI22_X1 U20115 ( .A1(n16914), .A2(n16913), .B1(n17206), .B2(n17186), .ZN(
        P3_U2673) );
  NAND2_X1 U20116 ( .A1(n16916), .A2(n16915), .ZN(n16918) );
  XNOR2_X1 U20117 ( .A(n16918), .B(n16917), .ZN(n17207) );
  NOR4_X1 U20118 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16947), .A3(n16920), .A4(
        n16919), .ZN(n16921) );
  AOI21_X1 U20119 ( .B1(n17188), .B2(n17207), .A(n16921), .ZN(n16922) );
  OAI21_X1 U20120 ( .B1(n16924), .B2(n16923), .A(n16922), .ZN(P3_U2674) );
  OAI221_X1 U20121 ( .B1(n16926), .B2(n16931), .C1(n16926), .C2(n16930), .A(
        n16925), .ZN(n17220) );
  AOI22_X1 U20122 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16932), .B1(n16928), 
        .B2(n16927), .ZN(n16929) );
  OAI21_X1 U20123 ( .B1(n17186), .B2(n17220), .A(n16929), .ZN(P3_U2676) );
  NAND2_X1 U20124 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16941), .ZN(n16937) );
  XOR2_X1 U20125 ( .A(n16931), .B(n16930), .Z(n17221) );
  AOI22_X1 U20126 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16932), .B1(n17188), 
        .B2(n17221), .ZN(n16933) );
  OAI21_X1 U20127 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n16937), .A(n16933), .ZN(
        P3_U2677) );
  OAI21_X1 U20128 ( .B1(n16936), .B2(n16935), .A(n16934), .ZN(n17229) );
  OAI211_X1 U20129 ( .C1(n16941), .C2(P3_EBX_REG_25__SCAN_IN), .A(n17186), .B(
        n16937), .ZN(n16938) );
  OAI21_X1 U20130 ( .B1(n17229), .B2(n17186), .A(n16938), .ZN(P3_U2678) );
  AOI21_X1 U20131 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17186), .A(n16946), .ZN(
        n16940) );
  XNOR2_X1 U20132 ( .A(n16939), .B(n16942), .ZN(n17234) );
  OAI22_X1 U20133 ( .A1(n16941), .A2(n16940), .B1(n17186), .B2(n17234), .ZN(
        P3_U2679) );
  AOI21_X1 U20134 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17186), .A(n16962), .ZN(
        n16945) );
  OAI21_X1 U20135 ( .B1(n16944), .B2(n16943), .A(n16942), .ZN(n17239) );
  OAI22_X1 U20136 ( .A1(n16946), .A2(n16945), .B1(n17186), .B2(n17239), .ZN(
        P3_U2680) );
  OAI21_X1 U20137 ( .B1(n16948), .B2(n17188), .A(n16947), .ZN(n16949) );
  INV_X1 U20138 ( .A(n16949), .ZN(n16961) );
  AOI22_X1 U20139 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16950) );
  OAI21_X1 U20140 ( .B1(n12721), .B2(n17060), .A(n16950), .ZN(n16960) );
  INV_X1 U20141 ( .A(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17058) );
  AOI22_X1 U20142 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16958) );
  OAI22_X1 U20143 ( .A1(n9564), .A2(n16951), .B1(n17113), .B2(n18190), .ZN(
        n16956) );
  AOI22_X1 U20144 ( .A1(n15684), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16954) );
  AOI22_X1 U20145 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16953) );
  AOI22_X1 U20146 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16952) );
  NAND3_X1 U20147 ( .A1(n16954), .A2(n16953), .A3(n16952), .ZN(n16955) );
  AOI211_X1 U20148 ( .C1(n16899), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n16956), .B(n16955), .ZN(n16957) );
  OAI211_X1 U20149 ( .C1(n17004), .C2(n17058), .A(n16958), .B(n16957), .ZN(
        n16959) );
  AOI211_X1 U20150 ( .C1(n17137), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n16960), .B(n16959), .ZN(n17243) );
  OAI22_X1 U20151 ( .A1(n16962), .A2(n16961), .B1(n17243), .B2(n17186), .ZN(
        P3_U2681) );
  NAND2_X1 U20152 ( .A1(n17186), .A2(n16963), .ZN(n16990) );
  AOI22_X1 U20153 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16974) );
  AOI22_X1 U20154 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17056), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16965) );
  AOI22_X1 U20155 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16964) );
  OAI211_X1 U20156 ( .C1(n17146), .C2(n16966), .A(n16965), .B(n16964), .ZN(
        n16972) );
  AOI22_X1 U20157 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16970) );
  AOI22_X1 U20158 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16969) );
  AOI22_X1 U20159 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16968) );
  NAND2_X1 U20160 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n16967) );
  NAND4_X1 U20161 ( .A1(n16970), .A2(n16969), .A3(n16968), .A4(n16967), .ZN(
        n16971) );
  AOI211_X1 U20162 ( .C1(n12701), .C2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n16972), .B(n16971), .ZN(n16973) );
  OAI211_X1 U20163 ( .C1(n17113), .C2(n18184), .A(n16974), .B(n16973), .ZN(
        n17248) );
  AOI22_X1 U20164 ( .A1(n17188), .A2(n17248), .B1(n16975), .B2(n16977), .ZN(
        n16976) );
  OAI21_X1 U20165 ( .B1(n16977), .B2(n16990), .A(n16976), .ZN(P3_U2682) );
  NOR2_X1 U20166 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n9657), .ZN(n16991) );
  INV_X1 U20167 ( .A(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16979) );
  AOI22_X1 U20168 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16978) );
  OAI21_X1 U20169 ( .B1(n16980), .B2(n16979), .A(n16978), .ZN(n16989) );
  AOI22_X1 U20170 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16987) );
  AOI22_X1 U20171 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16981) );
  OAI21_X1 U20172 ( .B1(n17090), .B2(n20874), .A(n16981), .ZN(n16985) );
  AOI22_X1 U20173 ( .A1(n9568), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15648), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16983) );
  AOI22_X1 U20174 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17056), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16982) );
  OAI211_X1 U20175 ( .C1(n17146), .C2(n17083), .A(n16983), .B(n16982), .ZN(
        n16984) );
  AOI211_X1 U20176 ( .C1(n17131), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n16985), .B(n16984), .ZN(n16986) );
  OAI211_X1 U20177 ( .C1(n17113), .C2(n18178), .A(n16987), .B(n16986), .ZN(
        n16988) );
  AOI211_X1 U20178 ( .C1(n17137), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n16989), .B(n16988), .ZN(n17256) );
  OAI22_X1 U20179 ( .A1(n16991), .A2(n16990), .B1(n17256), .B2(n17186), .ZN(
        P3_U2683) );
  AOI21_X1 U20180 ( .B1(n16993), .B2(n16992), .A(n17188), .ZN(n16994) );
  INV_X1 U20181 ( .A(n16994), .ZN(n17007) );
  AOI22_X1 U20182 ( .A1(n9568), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15648), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16995) );
  OAI21_X1 U20183 ( .B1(n10053), .B2(n17089), .A(n16995), .ZN(n17006) );
  INV_X1 U20184 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U20185 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17056), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17002) );
  OAI22_X1 U20186 ( .A1(n9565), .A2(n18232), .B1(n17113), .B2(n18172), .ZN(
        n17000) );
  AOI22_X1 U20187 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16998) );
  AOI22_X1 U20188 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16997) );
  AOI22_X1 U20189 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16996) );
  NAND3_X1 U20190 ( .A1(n16998), .A2(n16997), .A3(n16996), .ZN(n16999) );
  AOI211_X1 U20191 ( .C1(n17131), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n17000), .B(n16999), .ZN(n17001) );
  OAI211_X1 U20192 ( .C1(n17004), .C2(n17003), .A(n17002), .B(n17001), .ZN(
        n17005) );
  AOI211_X1 U20193 ( .C1(n17100), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n17006), .B(n17005), .ZN(n17261) );
  OAI22_X1 U20194 ( .A1(n9657), .A2(n17007), .B1(n17261), .B2(n17186), .ZN(
        P3_U2684) );
  NAND3_X1 U20195 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(P3_EBX_REG_16__SCAN_IN), 
        .A3(n17036), .ZN(n17021) );
  NOR2_X1 U20196 ( .A1(n17188), .A2(n17008), .ZN(n17019) );
  AOI22_X1 U20197 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17056), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17018) );
  AOI22_X1 U20198 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17009) );
  OAI21_X1 U20199 ( .B1(n17088), .B2(n20864), .A(n17009), .ZN(n17016) );
  OAI22_X1 U20200 ( .A1(n9565), .A2(n18228), .B1(n17090), .B2(n17118), .ZN(
        n17010) );
  AOI21_X1 U20201 ( .B1(n17149), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n17010), .ZN(n17014) );
  AOI22_X1 U20202 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17013) );
  AOI22_X1 U20203 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17012) );
  AOI22_X1 U20204 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17011) );
  NAND4_X1 U20205 ( .A1(n17014), .A2(n17013), .A3(n17012), .A4(n17011), .ZN(
        n17015) );
  AOI211_X1 U20206 ( .C1(n17137), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n17016), .B(n17015), .ZN(n17017) );
  OAI211_X1 U20207 ( .C1(n12721), .C2(n17112), .A(n17018), .B(n17017), .ZN(
        n17262) );
  AOI22_X1 U20208 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17019), .B1(n17188), 
        .B2(n17262), .ZN(n17020) );
  OAI21_X1 U20209 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17021), .A(n17020), .ZN(
        P3_U2685) );
  NAND2_X1 U20210 ( .A1(n17186), .A2(n17022), .ZN(n17053) );
  AOI22_X1 U20211 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15648), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17034) );
  AOI22_X1 U20212 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17023) );
  OAI21_X1 U20213 ( .B1(n9564), .B2(n17024), .A(n17023), .ZN(n17031) );
  OAI22_X1 U20214 ( .A1(n9565), .A2(n20773), .B1(n17113), .B2(n18154), .ZN(
        n17025) );
  AOI21_X1 U20215 ( .B1(n17105), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n17025), .ZN(n17029) );
  AOI22_X1 U20216 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15684), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20217 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17027) );
  AOI22_X1 U20218 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17026) );
  NAND4_X1 U20219 ( .A1(n17029), .A2(n17028), .A3(n17027), .A4(n17026), .ZN(
        n17030) );
  AOI211_X1 U20220 ( .C1(n17032), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n17031), .B(n17030), .ZN(n17033) );
  OAI211_X1 U20221 ( .C1(n12700), .C2(n17035), .A(n17034), .B(n17033), .ZN(
        n17273) );
  AOI22_X1 U20222 ( .A1(n17188), .A2(n17273), .B1(n17036), .B2(n17038), .ZN(
        n17037) );
  OAI21_X1 U20223 ( .B1(n17038), .B2(n17053), .A(n17037), .ZN(P3_U2687) );
  NOR2_X1 U20224 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17039), .ZN(n17054) );
  AOI22_X1 U20225 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n15648), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n12691), .ZN(n17040) );
  OAI21_X1 U20226 ( .B1(n17041), .B2(n9616), .A(n17040), .ZN(n17052) );
  AOI22_X1 U20227 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n9574), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17050) );
  AOI22_X1 U20228 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12701), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17156), .ZN(n17042) );
  OAI21_X1 U20229 ( .B1(n17113), .B2(n17043), .A(n17042), .ZN(n17048) );
  INV_X1 U20230 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18197) );
  AOI22_X1 U20231 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17046) );
  AOI22_X1 U20232 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n17044), .ZN(n17045) );
  OAI211_X1 U20233 ( .C1(n18197), .C2(n17146), .A(n17046), .B(n17045), .ZN(
        n17047) );
  AOI211_X1 U20234 ( .C1(n17131), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n17048), .B(n17047), .ZN(n17049) );
  OAI211_X1 U20235 ( .C1(n10053), .C2(n18244), .A(n17050), .B(n17049), .ZN(
        n17051) );
  AOI211_X1 U20236 ( .C1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .C2(n15684), .A(
        n17052), .B(n17051), .ZN(n17282) );
  OAI22_X1 U20237 ( .A1(n17054), .A2(n17053), .B1(n17282), .B2(n17186), .ZN(
        P3_U2688) );
  NAND3_X1 U20238 ( .A1(n18193), .A2(P3_EBX_REG_13__SCAN_IN), .A3(n17055), 
        .ZN(n17071) );
  AOI22_X1 U20239 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17056), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17057) );
  OAI21_X1 U20240 ( .B1(n9564), .B2(n17058), .A(n17057), .ZN(n17069) );
  AOI22_X1 U20241 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9574), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17066) );
  AOI22_X1 U20242 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17059) );
  OAI21_X1 U20243 ( .B1(n17113), .B2(n17060), .A(n17059), .ZN(n17064) );
  AOI22_X1 U20244 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17062) );
  AOI22_X1 U20245 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17061) );
  OAI211_X1 U20246 ( .C1(n17146), .C2(n18190), .A(n17062), .B(n17061), .ZN(
        n17063) );
  AOI211_X1 U20247 ( .C1(n17131), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n17064), .B(n17063), .ZN(n17065) );
  OAI211_X1 U20248 ( .C1(n17088), .C2(n17067), .A(n17066), .B(n17065), .ZN(
        n17068) );
  AOI211_X1 U20249 ( .C1(n16899), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n17069), .B(n17068), .ZN(n17287) );
  NAND3_X1 U20250 ( .A1(n17071), .A2(P3_EBX_REG_14__SCAN_IN), .A3(n17186), 
        .ZN(n17070) );
  OAI221_X1 U20251 ( .B1(n17071), .B2(P3_EBX_REG_14__SCAN_IN), .C1(n17186), 
        .C2(n17287), .A(n17070), .ZN(P3_U2689) );
  NAND2_X1 U20252 ( .A1(n17186), .A2(n17072), .ZN(n17101) );
  AOI22_X1 U20253 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17082) );
  AOI22_X1 U20254 ( .A1(n17122), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17074) );
  AOI22_X1 U20255 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17073) );
  OAI211_X1 U20256 ( .C1(n17146), .C2(n18178), .A(n17074), .B(n17073), .ZN(
        n17080) );
  AOI22_X1 U20257 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15684), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17078) );
  AOI22_X1 U20258 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15648), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17077) );
  AOI22_X1 U20259 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17076) );
  NAND2_X1 U20260 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n17075) );
  NAND4_X1 U20261 ( .A1(n17078), .A2(n17077), .A3(n17076), .A4(n17075), .ZN(
        n17079) );
  AOI211_X1 U20262 ( .C1(n17131), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n17080), .B(n17079), .ZN(n17081) );
  OAI211_X1 U20263 ( .C1(n9565), .C2(n17083), .A(n17082), .B(n17081), .ZN(
        n17292) );
  OAI22_X1 U20264 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17101), .B1(n17292), 
        .B2(n17186), .ZN(n17084) );
  NOR2_X1 U20265 ( .A1(n17085), .A2(n17084), .ZN(P3_U2691) );
  INV_X1 U20266 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17087) );
  AOI22_X1 U20267 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15684), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17086) );
  OAI21_X1 U20268 ( .B1(n17088), .B2(n17087), .A(n17086), .ZN(n17099) );
  AOI22_X1 U20269 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(n9568), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17097) );
  OAI22_X1 U20270 ( .A1(n17146), .A2(n18172), .B1(n17090), .B2(n17089), .ZN(
        n17095) );
  AOI22_X1 U20271 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17093) );
  AOI22_X1 U20272 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17092) );
  AOI22_X1 U20273 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17091) );
  NAND3_X1 U20274 ( .A1(n17093), .A2(n17092), .A3(n17091), .ZN(n17094) );
  AOI211_X1 U20275 ( .C1(n17149), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n17095), .B(n17094), .ZN(n17096) );
  OAI211_X1 U20276 ( .C1(n9618), .C2(n20809), .A(n17097), .B(n17096), .ZN(
        n17098) );
  AOI211_X1 U20277 ( .C1(n17100), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n17099), .B(n17098), .ZN(n17297) );
  NOR2_X1 U20278 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17121), .ZN(n17102) );
  OAI22_X1 U20279 ( .A1(n17297), .A2(n17186), .B1(n17102), .B2(n17101), .ZN(
        P3_U2692) );
  OAI21_X1 U20280 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17103), .A(n17186), .ZN(
        n17120) );
  AOI22_X1 U20281 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9574), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17117) );
  AOI22_X1 U20282 ( .A1(n15684), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17104) );
  OAI21_X1 U20283 ( .B1(n10053), .B2(n18228), .A(n17104), .ZN(n17115) );
  AOI22_X1 U20284 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17111) );
  AOI22_X1 U20285 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17107) );
  AOI22_X1 U20286 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15648), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17106) );
  OAI211_X1 U20287 ( .C1(n17108), .C2(n20864), .A(n17107), .B(n17106), .ZN(
        n17109) );
  AOI21_X1 U20288 ( .B1(n17156), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n17109), .ZN(n17110) );
  OAI211_X1 U20289 ( .C1(n17113), .C2(n17112), .A(n17111), .B(n17110), .ZN(
        n17114) );
  AOI211_X1 U20290 ( .C1(n17143), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n17115), .B(n17114), .ZN(n17116) );
  OAI211_X1 U20291 ( .C1(n12700), .C2(n17118), .A(n17117), .B(n17116), .ZN(
        n17300) );
  INV_X1 U20292 ( .A(n17300), .ZN(n17119) );
  OAI22_X1 U20293 ( .A1(n17121), .A2(n17120), .B1(n17119), .B2(n17186), .ZN(
        P3_U2693) );
  AOI22_X1 U20294 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17123) );
  OAI21_X1 U20295 ( .B1(n9618), .B2(n17124), .A(n17123), .ZN(n17136) );
  AOI22_X1 U20296 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n15684), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17133) );
  AOI22_X1 U20297 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12701), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17125) );
  OAI21_X1 U20298 ( .B1(n17146), .B2(n18160), .A(n17125), .ZN(n17130) );
  AOI22_X1 U20299 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15648), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20300 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17126) );
  OAI211_X1 U20301 ( .C1(n9565), .C2(n17128), .A(n17127), .B(n17126), .ZN(
        n17129) );
  AOI211_X1 U20302 ( .C1(n17131), .C2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n17130), .B(n17129), .ZN(n17132) );
  OAI211_X1 U20303 ( .C1(n9564), .C2(n17134), .A(n17133), .B(n17132), .ZN(
        n17135) );
  AOI211_X1 U20304 ( .C1(n17137), .C2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n17136), .B(n17135), .ZN(n17307) );
  OAI21_X1 U20305 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n9669), .A(n17138), .ZN(
        n17139) );
  AOI22_X1 U20306 ( .A1(n17188), .A2(n17307), .B1(n17139), .B2(n17186), .ZN(
        P3_U2694) );
  AOI22_X1 U20307 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17158) );
  AOI22_X1 U20308 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17145) );
  AOI22_X1 U20309 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17144) );
  OAI211_X1 U20310 ( .C1(n17146), .C2(n18154), .A(n17145), .B(n17144), .ZN(
        n17155) );
  AOI22_X1 U20311 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17153) );
  AOI22_X1 U20312 ( .A1(n15684), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17152) );
  AOI22_X1 U20313 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17151) );
  NAND2_X1 U20314 ( .A1(n12701), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n17150) );
  NAND4_X1 U20315 ( .A1(n17153), .A2(n17152), .A3(n17151), .A4(n17150), .ZN(
        n17154) );
  AOI211_X1 U20316 ( .C1(n17156), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n17155), .B(n17154), .ZN(n17157) );
  OAI211_X1 U20317 ( .C1(n10053), .C2(n20773), .A(n17158), .B(n17157), .ZN(
        n17310) );
  NAND3_X1 U20318 ( .A1(n17186), .A2(n17160), .A3(n17159), .ZN(n17161) );
  OAI21_X1 U20319 ( .B1(n17186), .B2(n17310), .A(n17161), .ZN(n17162) );
  AOI21_X1 U20320 ( .B1(n18193), .B2(n9669), .A(n17162), .ZN(P3_U2695) );
  NOR2_X1 U20321 ( .A1(n17188), .A2(n17164), .ZN(n17166) );
  OAI222_X1 U20322 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n18193), .B1(
        P3_EBX_REG_7__SCAN_IN), .B2(n17164), .C1(n17166), .C2(n17163), .ZN(
        n17165) );
  OAI21_X1 U20323 ( .B1(n18197), .B2(n17186), .A(n17165), .ZN(P3_U2696) );
  OAI21_X1 U20324 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17167), .A(n17166), .ZN(
        n17168) );
  OAI21_X1 U20325 ( .B1(n17186), .B2(n18190), .A(n17168), .ZN(P3_U2697) );
  OAI21_X1 U20326 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17170), .A(n17169), .ZN(
        n17171) );
  AOI22_X1 U20327 ( .A1(n17188), .A2(n18184), .B1(n17171), .B2(n17186), .ZN(
        P3_U2698) );
  AOI22_X1 U20328 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n17188), .B1(
        P3_EBX_REG_4__SCAN_IN), .B2(n17184), .ZN(n17175) );
  OAI211_X1 U20329 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17173), .A(n17187), .B(
        n17172), .ZN(n17174) );
  NAND2_X1 U20330 ( .A1(n17175), .A2(n17174), .ZN(P3_U2699) );
  NAND2_X1 U20331 ( .A1(n17176), .A2(n17187), .ZN(n17178) );
  NAND3_X1 U20332 ( .A1(n17178), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n17186), .ZN(
        n17177) );
  OAI221_X1 U20333 ( .B1(n17178), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n17186), 
        .C2(n18172), .A(n17177), .ZN(P3_U2700) );
  AND2_X1 U20334 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17179) );
  AOI21_X1 U20335 ( .B1(n17191), .B2(n17179), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n17182) );
  AOI21_X1 U20336 ( .B1(n18193), .B2(n17180), .A(n17184), .ZN(n17181) );
  INV_X1 U20337 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18166) );
  OAI22_X1 U20338 ( .A1(n17182), .A2(n17181), .B1(n18166), .B2(n17186), .ZN(
        P3_U2701) );
  AOI22_X1 U20339 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(n17184), .B1(n17187), .B2(
        n17183), .ZN(n17185) );
  OAI21_X1 U20340 ( .B1(n18160), .B2(n17186), .A(n17185), .ZN(P3_U2702) );
  AOI22_X1 U20341 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17188), .B1(
        n17187), .B2(n17190), .ZN(n17189) );
  OAI21_X1 U20342 ( .B1(n17191), .B2(n17190), .A(n17189), .ZN(P3_U2703) );
  INV_X1 U20343 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17353) );
  INV_X1 U20344 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17359) );
  NAND3_X1 U20345 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(n9585), .ZN(n17196) );
  NAND3_X1 U20346 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(P3_EAX_REG_2__SCAN_IN), .ZN(n17315) );
  NAND2_X1 U20347 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n17342) );
  INV_X1 U20348 ( .A(n17342), .ZN(n17193) );
  INV_X1 U20349 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17396) );
  NAND3_X1 U20350 ( .A1(n17194), .A2(n17193), .A3(P3_EAX_REG_5__SCAN_IN), .ZN(
        n17195) );
  NOR2_X2 U20351 ( .A1(n17196), .A2(n17195), .ZN(n17318) );
  NAND3_X1 U20352 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .ZN(n17283) );
  NOR2_X1 U20353 ( .A1(n17312), .A2(n17283), .ZN(n17197) );
  INV_X1 U20354 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17458) );
  NOR2_X2 U20355 ( .A1(n17284), .A2(n17458), .ZN(n17279) );
  NAND2_X1 U20356 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .ZN(n17241) );
  NAND4_X1 U20357 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_22__SCAN_IN), 
        .A3(P3_EAX_REG_20__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17198)
         );
  NAND2_X1 U20358 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17236), .ZN(n17235) );
  NOR2_X2 U20359 ( .A1(n17359), .A2(n17230), .ZN(n17225) );
  NAND2_X1 U20360 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17225), .ZN(n17222) );
  NAND2_X1 U20361 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17212), .ZN(n17208) );
  NAND2_X1 U20362 ( .A1(n17203), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17202) );
  NAND2_X1 U20363 ( .A1(n17199), .A2(n17305), .ZN(n17242) );
  OAI22_X1 U20364 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17326), .B1(n17305), 
        .B2(n17203), .ZN(n17200) );
  AOI22_X1 U20365 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17274), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17200), .ZN(n17201) );
  OAI21_X1 U20366 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17202), .A(n17201), .ZN(
        P3_U2704) );
  NAND2_X1 U20367 ( .A1(n18181), .A2(n17305), .ZN(n17278) );
  AOI22_X1 U20368 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17267), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17274), .ZN(n17205) );
  OAI211_X1 U20369 ( .C1(n17203), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17335), .B(
        n17202), .ZN(n17204) );
  OAI211_X1 U20370 ( .C1(n17206), .C2(n17346), .A(n17205), .B(n17204), .ZN(
        P3_U2705) );
  INV_X1 U20371 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18179) );
  AOI22_X1 U20372 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17267), .B1(n17207), .B2(
        n17311), .ZN(n17210) );
  OAI211_X1 U20373 ( .C1(n17212), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17335), .B(
        n17208), .ZN(n17209) );
  OAI211_X1 U20374 ( .C1(n17242), .C2(n18179), .A(n17210), .B(n17209), .ZN(
        P3_U2706) );
  INV_X1 U20375 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18174) );
  AOI22_X1 U20376 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17267), .B1(n17211), .B2(
        n17311), .ZN(n17215) );
  AOI211_X1 U20377 ( .C1(n17353), .C2(n17216), .A(n17212), .B(n17305), .ZN(
        n17213) );
  INV_X1 U20378 ( .A(n17213), .ZN(n17214) );
  OAI211_X1 U20379 ( .C1(n17242), .C2(n18174), .A(n17215), .B(n17214), .ZN(
        P3_U2707) );
  AOI22_X1 U20380 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17267), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17274), .ZN(n17219) );
  OAI211_X1 U20381 ( .C1(n17217), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17335), .B(
        n17216), .ZN(n17218) );
  OAI211_X1 U20382 ( .C1(n17346), .C2(n17220), .A(n17219), .B(n17218), .ZN(
        P3_U2708) );
  INV_X1 U20383 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18161) );
  AOI22_X1 U20384 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17267), .B1(n17221), .B2(
        n17311), .ZN(n17224) );
  OAI211_X1 U20385 ( .C1(n17225), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17335), .B(
        n17222), .ZN(n17223) );
  OAI211_X1 U20386 ( .C1(n17242), .C2(n18161), .A(n17224), .B(n17223), .ZN(
        P3_U2709) );
  AOI22_X1 U20387 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17267), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17274), .ZN(n17228) );
  AOI211_X1 U20388 ( .C1(n17359), .C2(n17230), .A(n17225), .B(n17305), .ZN(
        n17226) );
  INV_X1 U20389 ( .A(n17226), .ZN(n17227) );
  OAI211_X1 U20390 ( .C1(n17346), .C2(n17229), .A(n17228), .B(n17227), .ZN(
        P3_U2710) );
  AOI22_X1 U20391 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17267), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17274), .ZN(n17233) );
  OAI211_X1 U20392 ( .C1(n17231), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17335), .B(
        n17230), .ZN(n17232) );
  OAI211_X1 U20393 ( .C1(n17346), .C2(n17234), .A(n17233), .B(n17232), .ZN(
        P3_U2711) );
  AOI22_X1 U20394 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17267), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17274), .ZN(n17238) );
  OAI211_X1 U20395 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17236), .A(n17335), .B(
        n17235), .ZN(n17237) );
  OAI211_X1 U20396 ( .C1(n17346), .C2(n17239), .A(n17238), .B(n17237), .ZN(
        P3_U2712) );
  INV_X1 U20397 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n20824) );
  NAND2_X1 U20398 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17257), .ZN(n17253) );
  NOR2_X1 U20399 ( .A1(n20824), .A2(n17253), .ZN(n17252) );
  INV_X1 U20400 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17365) );
  INV_X1 U20401 ( .A(n17253), .ZN(n17247) );
  OAI22_X1 U20402 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17326), .B1(n17305), 
        .B2(n17247), .ZN(n17245) );
  INV_X1 U20403 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n20807) );
  OAI22_X1 U20404 ( .A1(n17243), .A2(n17346), .B1(n20807), .B2(n17242), .ZN(
        n17244) );
  AOI221_X1 U20405 ( .B1(n17252), .B2(n17365), .C1(n17245), .C2(
        P3_EAX_REG_22__SCAN_IN), .A(n17244), .ZN(n17246) );
  OAI21_X1 U20406 ( .B1(n18186), .B2(n17278), .A(n17246), .ZN(P3_U2713) );
  AOI21_X1 U20407 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17335), .A(n17247), .ZN(
        n17251) );
  AOI22_X1 U20408 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17267), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17274), .ZN(n17250) );
  NAND2_X1 U20409 ( .A1(n17311), .A2(n17248), .ZN(n17249) );
  OAI211_X1 U20410 ( .C1(n17252), .C2(n17251), .A(n17250), .B(n17249), .ZN(
        P3_U2714) );
  AOI22_X1 U20411 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17267), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17274), .ZN(n17255) );
  OAI211_X1 U20412 ( .C1(n17257), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17335), .B(
        n17253), .ZN(n17254) );
  OAI211_X1 U20413 ( .C1(n17256), .C2(n17346), .A(n17255), .B(n17254), .ZN(
        P3_U2715) );
  AOI22_X1 U20414 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17267), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17274), .ZN(n17260) );
  INV_X1 U20415 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17370) );
  INV_X1 U20416 ( .A(n17268), .ZN(n17264) );
  NAND2_X1 U20417 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17264), .ZN(n17263) );
  AOI211_X1 U20418 ( .C1(n17370), .C2(n17263), .A(n17257), .B(n17305), .ZN(
        n17258) );
  INV_X1 U20419 ( .A(n17258), .ZN(n17259) );
  OAI211_X1 U20420 ( .C1(n17261), .C2(n17346), .A(n17260), .B(n17259), .ZN(
        P3_U2716) );
  AOI22_X1 U20421 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17274), .B1(n17311), .B2(
        n17262), .ZN(n17266) );
  OAI211_X1 U20422 ( .C1(n17264), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17335), .B(
        n17263), .ZN(n17265) );
  OAI211_X1 U20423 ( .C1(n17278), .C2(n18162), .A(n17266), .B(n17265), .ZN(
        P3_U2717) );
  AOI22_X1 U20424 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17267), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17274), .ZN(n17271) );
  OAI211_X1 U20425 ( .C1(n17269), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17335), .B(
        n17268), .ZN(n17270) );
  OAI211_X1 U20426 ( .C1(n17272), .C2(n17346), .A(n17271), .B(n17270), .ZN(
        P3_U2718) );
  INV_X1 U20427 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18149) );
  AOI22_X1 U20428 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n17274), .B1(n17311), .B2(
        n17273), .ZN(n17277) );
  OAI211_X1 U20429 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17279), .A(n17335), .B(
        n17275), .ZN(n17276) );
  OAI211_X1 U20430 ( .C1(n17278), .C2(n18149), .A(n17277), .B(n17276), .ZN(
        P3_U2719) );
  AOI211_X1 U20431 ( .C1(n17458), .C2(n17284), .A(n17305), .B(n17279), .ZN(
        n17280) );
  AOI21_X1 U20432 ( .B1(n17341), .B2(BUF2_REG_15__SCAN_IN), .A(n17280), .ZN(
        n17281) );
  OAI21_X1 U20433 ( .B1(n17282), .B2(n17346), .A(n17281), .ZN(P3_U2720) );
  INV_X1 U20434 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17388) );
  NAND3_X1 U20435 ( .A1(n18193), .A2(P3_EAX_REG_8__SCAN_IN), .A3(n17318), .ZN(
        n17304) );
  NAND2_X1 U20436 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17309), .ZN(n17301) );
  NOR2_X1 U20437 ( .A1(n17283), .A2(n17301), .ZN(n17291) );
  INV_X1 U20438 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17453) );
  AOI22_X1 U20439 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17341), .B1(n17291), .B2(
        n17453), .ZN(n17286) );
  NAND3_X1 U20440 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17335), .A3(n17284), 
        .ZN(n17285) );
  OAI211_X1 U20441 ( .C1(n17287), .C2(n17346), .A(n17286), .B(n17285), .ZN(
        P3_U2721) );
  INV_X1 U20442 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17451) );
  NAND2_X1 U20443 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .ZN(n17288) );
  NOR2_X1 U20444 ( .A1(n17288), .A2(n17301), .ZN(n17295) );
  AOI21_X1 U20445 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17335), .A(n17295), .ZN(
        n17290) );
  OAI222_X1 U20446 ( .A1(n17339), .A2(n17451), .B1(n17291), .B2(n17290), .C1(
        n17346), .C2(n17289), .ZN(P3_U2722) );
  INV_X1 U20447 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17447) );
  INV_X1 U20448 ( .A(n17301), .ZN(n17296) );
  AOI22_X1 U20449 ( .A1(n17296), .A2(P3_EAX_REG_11__SCAN_IN), .B1(
        P3_EAX_REG_12__SCAN_IN), .B2(n17335), .ZN(n17294) );
  INV_X1 U20450 ( .A(n17292), .ZN(n17293) );
  OAI222_X1 U20451 ( .A1(n17339), .A2(n17447), .B1(n17295), .B2(n17294), .C1(
        n17346), .C2(n17293), .ZN(P3_U2723) );
  INV_X1 U20452 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17445) );
  INV_X1 U20453 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17384) );
  NOR2_X1 U20454 ( .A1(n17384), .A2(n17301), .ZN(n17299) );
  AOI21_X1 U20455 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17335), .A(n17296), .ZN(
        n17298) );
  OAI222_X1 U20456 ( .A1(n17339), .A2(n17445), .B1(n17299), .B2(n17298), .C1(
        n17346), .C2(n17297), .ZN(P3_U2724) );
  AOI22_X1 U20457 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17341), .B1(n17311), .B2(
        n17300), .ZN(n17303) );
  OAI211_X1 U20458 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17309), .A(n17335), .B(
        n17301), .ZN(n17302) );
  NAND2_X1 U20459 ( .A1(n17303), .A2(n17302), .ZN(P3_U2725) );
  OAI21_X1 U20460 ( .B1(n17388), .B2(n17305), .A(n17304), .ZN(n17306) );
  INV_X1 U20461 ( .A(n17306), .ZN(n17308) );
  OAI222_X1 U20462 ( .A1(n17339), .A2(n17441), .B1(n17309), .B2(n17308), .C1(
        n17346), .C2(n17307), .ZN(P3_U2726) );
  AOI22_X1 U20463 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17341), .B1(n17311), .B2(
        n17310), .ZN(n17314) );
  OAI211_X1 U20464 ( .C1(P3_EAX_REG_8__SCAN_IN), .C2(n17318), .A(n17335), .B(
        n17312), .ZN(n17313) );
  NAND2_X1 U20465 ( .A1(n17314), .A2(n17313), .ZN(P3_U2727) );
  INV_X1 U20466 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17394) );
  NOR3_X1 U20467 ( .A1(n17315), .A2(n17342), .A3(n17326), .ZN(n17328) );
  NAND2_X1 U20468 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17328), .ZN(n17319) );
  NOR2_X1 U20469 ( .A1(n17394), .A2(n17319), .ZN(n17321) );
  AOI21_X1 U20470 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17335), .A(n17321), .ZN(
        n17317) );
  OAI222_X1 U20471 ( .A1(n17339), .A2(n18191), .B1(n17318), .B2(n17317), .C1(
        n17346), .C2(n17316), .ZN(P3_U2728) );
  INV_X1 U20472 ( .A(n17319), .ZN(n17324) );
  AOI21_X1 U20473 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17335), .A(n17324), .ZN(
        n17322) );
  OAI222_X1 U20474 ( .A1(n17339), .A2(n18186), .B1(n17322), .B2(n17321), .C1(
        n17346), .C2(n17320), .ZN(P3_U2729) );
  INV_X1 U20475 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18180) );
  AOI21_X1 U20476 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17335), .A(n17328), .ZN(
        n17325) );
  OAI222_X1 U20477 ( .A1(n17339), .A2(n18180), .B1(n17325), .B2(n17324), .C1(
        n17346), .C2(n17323), .ZN(P3_U2730) );
  INV_X1 U20478 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17400) );
  NOR2_X1 U20479 ( .A1(n17342), .A2(n17326), .ZN(n17334) );
  NAND2_X1 U20480 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17334), .ZN(n17330) );
  NOR2_X1 U20481 ( .A1(n17400), .A2(n17330), .ZN(n17333) );
  AOI21_X1 U20482 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17335), .A(n17333), .ZN(
        n17329) );
  OAI222_X1 U20483 ( .A1(n17339), .A2(n18173), .B1(n17329), .B2(n17328), .C1(
        n17346), .C2(n17327), .ZN(P3_U2731) );
  INV_X1 U20484 ( .A(n17330), .ZN(n17338) );
  AOI21_X1 U20485 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17335), .A(n17338), .ZN(
        n17332) );
  OAI222_X1 U20486 ( .A1(n18167), .A2(n17339), .B1(n17333), .B2(n17332), .C1(
        n17346), .C2(n17331), .ZN(P3_U2732) );
  AOI21_X1 U20487 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17335), .A(n17334), .ZN(
        n17337) );
  OAI222_X1 U20488 ( .A1(n18162), .A2(n17339), .B1(n17338), .B2(n17337), .C1(
        n17346), .C2(n17336), .ZN(P3_U2733) );
  AOI22_X1 U20489 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17341), .B1(n17340), .B2(
        P3_EAX_REG_1__SCAN_IN), .ZN(n17345) );
  OAI211_X1 U20490 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(P3_EAX_REG_0__SCAN_IN), 
        .A(n17343), .B(n17342), .ZN(n17344) );
  OAI211_X1 U20491 ( .C1(n17347), .C2(n17346), .A(n17345), .B(n17344), .ZN(
        P3_U2734) );
  NAND2_X1 U20492 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17664), .ZN(n17362) );
  NOR2_X1 U20493 ( .A1(n17357), .A2(n17349), .ZN(P3_U2736) );
  INV_X1 U20494 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17428) );
  NOR2_X1 U20495 ( .A1(n17406), .A2(n18151), .ZN(n17360) );
  INV_X2 U20496 ( .A(n17362), .ZN(n17404) );
  AOI22_X1 U20497 ( .A1(n17404), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17350) );
  OAI21_X1 U20498 ( .B1(n17428), .B2(n17375), .A(n17350), .ZN(P3_U2737) );
  INV_X1 U20499 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n20793) );
  AOI22_X1 U20500 ( .A1(n17404), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17351) );
  OAI21_X1 U20501 ( .B1(n20793), .B2(n17375), .A(n17351), .ZN(P3_U2738) );
  AOI22_X1 U20502 ( .A1(n17404), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17352) );
  OAI21_X1 U20503 ( .B1(n17353), .B2(n17375), .A(n17352), .ZN(P3_U2739) );
  INV_X1 U20504 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17355) );
  AOI22_X1 U20505 ( .A1(n17404), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17354) );
  OAI21_X1 U20506 ( .B1(n17355), .B2(n17375), .A(n17354), .ZN(P3_U2740) );
  INV_X1 U20507 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n20820) );
  AOI22_X1 U20508 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17360), .B1(n17404), 
        .B2(P3_UWORD_REG_10__SCAN_IN), .ZN(n17356) );
  OAI21_X1 U20509 ( .B1(n20820), .B2(n17357), .A(n17356), .ZN(P3_U2741) );
  AOI22_X1 U20510 ( .A1(n17404), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17358) );
  OAI21_X1 U20511 ( .B1(n17359), .B2(n17375), .A(n17358), .ZN(P3_U2742) );
  INV_X1 U20512 ( .A(P3_UWORD_REG_8__SCAN_IN), .ZN(n20867) );
  AOI22_X1 U20513 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17360), .B1(n17392), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17361) );
  OAI21_X1 U20514 ( .B1(n17362), .B2(n20867), .A(n17361), .ZN(P3_U2743) );
  INV_X1 U20515 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20780) );
  AOI22_X1 U20516 ( .A1(n17404), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17363) );
  OAI21_X1 U20517 ( .B1(n20780), .B2(n17375), .A(n17363), .ZN(P3_U2744) );
  AOI22_X1 U20518 ( .A1(n17404), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17364) );
  OAI21_X1 U20519 ( .B1(n17365), .B2(n17375), .A(n17364), .ZN(P3_U2745) );
  AOI22_X1 U20520 ( .A1(n17404), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17366) );
  OAI21_X1 U20521 ( .B1(n20824), .B2(n17375), .A(n17366), .ZN(P3_U2746) );
  INV_X1 U20522 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17368) );
  AOI22_X1 U20523 ( .A1(n17404), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17367) );
  OAI21_X1 U20524 ( .B1(n17368), .B2(n17375), .A(n17367), .ZN(P3_U2747) );
  AOI22_X1 U20525 ( .A1(n17404), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17369) );
  OAI21_X1 U20526 ( .B1(n17370), .B2(n17375), .A(n17369), .ZN(P3_U2748) );
  INV_X1 U20527 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17372) );
  AOI22_X1 U20528 ( .A1(n17404), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17371) );
  OAI21_X1 U20529 ( .B1(n17372), .B2(n17375), .A(n17371), .ZN(P3_U2749) );
  INV_X1 U20530 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17413) );
  AOI22_X1 U20531 ( .A1(n17404), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17373) );
  OAI21_X1 U20532 ( .B1(n17413), .B2(n17375), .A(n17373), .ZN(P3_U2750) );
  INV_X1 U20533 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17376) );
  AOI22_X1 U20534 ( .A1(n17404), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17374) );
  OAI21_X1 U20535 ( .B1(n17376), .B2(n17375), .A(n17374), .ZN(P3_U2751) );
  AOI22_X1 U20536 ( .A1(n17404), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17377) );
  OAI21_X1 U20537 ( .B1(n17458), .B2(n17406), .A(n17377), .ZN(P3_U2752) );
  AOI22_X1 U20538 ( .A1(n17404), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17378) );
  OAI21_X1 U20539 ( .B1(n17453), .B2(n17406), .A(n17378), .ZN(P3_U2753) );
  INV_X1 U20540 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17380) );
  AOI22_X1 U20541 ( .A1(n17404), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17379) );
  OAI21_X1 U20542 ( .B1(n17380), .B2(n17406), .A(n17379), .ZN(P3_U2754) );
  INV_X1 U20543 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17382) );
  AOI22_X1 U20544 ( .A1(n17404), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17381) );
  OAI21_X1 U20545 ( .B1(n17382), .B2(n17406), .A(n17381), .ZN(P3_U2755) );
  AOI22_X1 U20546 ( .A1(n17404), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17383) );
  OAI21_X1 U20547 ( .B1(n17384), .B2(n17406), .A(n17383), .ZN(P3_U2756) );
  INV_X1 U20548 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17386) );
  AOI22_X1 U20549 ( .A1(n17404), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17385) );
  OAI21_X1 U20550 ( .B1(n17386), .B2(n17406), .A(n17385), .ZN(P3_U2757) );
  AOI22_X1 U20551 ( .A1(n17404), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17387) );
  OAI21_X1 U20552 ( .B1(n17388), .B2(n17406), .A(n17387), .ZN(P3_U2758) );
  INV_X1 U20553 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17439) );
  AOI22_X1 U20554 ( .A1(n17404), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17389) );
  OAI21_X1 U20555 ( .B1(n17439), .B2(n17406), .A(n17389), .ZN(P3_U2759) );
  INV_X1 U20556 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17391) );
  AOI22_X1 U20557 ( .A1(n17404), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17390) );
  OAI21_X1 U20558 ( .B1(n17391), .B2(n17406), .A(n17390), .ZN(P3_U2760) );
  AOI22_X1 U20559 ( .A1(n17404), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17393) );
  OAI21_X1 U20560 ( .B1(n17394), .B2(n17406), .A(n17393), .ZN(P3_U2761) );
  AOI22_X1 U20561 ( .A1(n17404), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17395) );
  OAI21_X1 U20562 ( .B1(n17396), .B2(n17406), .A(n17395), .ZN(P3_U2762) );
  INV_X1 U20563 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17398) );
  AOI22_X1 U20564 ( .A1(n17404), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17397) );
  OAI21_X1 U20565 ( .B1(n17398), .B2(n17406), .A(n17397), .ZN(P3_U2763) );
  AOI22_X1 U20566 ( .A1(n17404), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17399) );
  OAI21_X1 U20567 ( .B1(n17400), .B2(n17406), .A(n17399), .ZN(P3_U2764) );
  INV_X1 U20568 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17402) );
  AOI22_X1 U20569 ( .A1(n17404), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17401) );
  OAI21_X1 U20570 ( .B1(n17402), .B2(n17406), .A(n17401), .ZN(P3_U2765) );
  INV_X1 U20571 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17431) );
  AOI22_X1 U20572 ( .A1(n17404), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17403) );
  OAI21_X1 U20573 ( .B1(n17431), .B2(n17406), .A(n17403), .ZN(P3_U2766) );
  AOI22_X1 U20574 ( .A1(n17404), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17392), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17405) );
  OAI21_X1 U20575 ( .B1(n17407), .B2(n17406), .A(n17405), .ZN(P3_U2767) );
  INV_X1 U20576 ( .A(n17408), .ZN(n17410) );
  INV_X2 U20577 ( .A(n17421), .ZN(n17454) );
  INV_X2 U20578 ( .A(n17457), .ZN(n17448) );
  AOI22_X1 U20579 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17448), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17454), .ZN(n17411) );
  OAI21_X1 U20580 ( .B1(n18149), .B2(n17450), .A(n17411), .ZN(P3_U2768) );
  AOI22_X1 U20581 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17454), .ZN(n17412) );
  OAI21_X1 U20582 ( .B1(n17413), .B2(n17457), .A(n17412), .ZN(P3_U2769) );
  AOI22_X1 U20583 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17448), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17454), .ZN(n17414) );
  OAI21_X1 U20584 ( .B1(n18162), .B2(n17450), .A(n17414), .ZN(P3_U2770) );
  AOI22_X1 U20585 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17448), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17454), .ZN(n17415) );
  OAI21_X1 U20586 ( .B1(n18167), .B2(n17450), .A(n17415), .ZN(P3_U2771) );
  AOI22_X1 U20587 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17448), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17454), .ZN(n17416) );
  OAI21_X1 U20588 ( .B1(n18173), .B2(n17450), .A(n17416), .ZN(P3_U2772) );
  AOI22_X1 U20589 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17448), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17454), .ZN(n17417) );
  OAI21_X1 U20590 ( .B1(n18180), .B2(n17450), .A(n17417), .ZN(P3_U2773) );
  AOI22_X1 U20591 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17448), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17454), .ZN(n17418) );
  OAI21_X1 U20592 ( .B1(n18186), .B2(n17450), .A(n17418), .ZN(P3_U2774) );
  AOI22_X1 U20593 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17448), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17454), .ZN(n17419) );
  OAI21_X1 U20594 ( .B1(n18191), .B2(n17450), .A(n17419), .ZN(P3_U2775) );
  AOI22_X1 U20595 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17455), .B1(
        P3_EAX_REG_24__SCAN_IN), .B2(n17448), .ZN(n17420) );
  OAI21_X1 U20596 ( .B1(n17421), .B2(n20867), .A(n17420), .ZN(P3_U2776) );
  AOI22_X1 U20597 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17448), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17454), .ZN(n17422) );
  OAI21_X1 U20598 ( .B1(n17441), .B2(n17450), .A(n17422), .ZN(P3_U2777) );
  INV_X1 U20599 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17443) );
  AOI22_X1 U20600 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17448), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17454), .ZN(n17423) );
  OAI21_X1 U20601 ( .B1(n17443), .B2(n17450), .A(n17423), .ZN(P3_U2778) );
  AOI22_X1 U20602 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17448), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17454), .ZN(n17424) );
  OAI21_X1 U20603 ( .B1(n17445), .B2(n17450), .A(n17424), .ZN(P3_U2779) );
  AOI22_X1 U20604 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17448), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17454), .ZN(n17425) );
  OAI21_X1 U20605 ( .B1(n17447), .B2(n17450), .A(n17425), .ZN(P3_U2780) );
  AOI22_X1 U20606 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17448), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17454), .ZN(n17426) );
  OAI21_X1 U20607 ( .B1(n17451), .B2(n17450), .A(n17426), .ZN(P3_U2781) );
  AOI22_X1 U20608 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17454), .ZN(n17427) );
  OAI21_X1 U20609 ( .B1(n17428), .B2(n17457), .A(n17427), .ZN(P3_U2782) );
  AOI22_X1 U20610 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17448), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17454), .ZN(n17429) );
  OAI21_X1 U20611 ( .B1(n18149), .B2(n17450), .A(n17429), .ZN(P3_U2783) );
  AOI22_X1 U20612 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17454), .ZN(n17430) );
  OAI21_X1 U20613 ( .B1(n17431), .B2(n17457), .A(n17430), .ZN(P3_U2784) );
  AOI22_X1 U20614 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17448), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17454), .ZN(n17432) );
  OAI21_X1 U20615 ( .B1(n18162), .B2(n17450), .A(n17432), .ZN(P3_U2785) );
  AOI22_X1 U20616 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17448), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17454), .ZN(n17433) );
  OAI21_X1 U20617 ( .B1(n18167), .B2(n17450), .A(n17433), .ZN(P3_U2786) );
  AOI22_X1 U20618 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17448), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17454), .ZN(n17434) );
  OAI21_X1 U20619 ( .B1(n18173), .B2(n17450), .A(n17434), .ZN(P3_U2787) );
  AOI22_X1 U20620 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17448), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17454), .ZN(n17435) );
  OAI21_X1 U20621 ( .B1(n18180), .B2(n17450), .A(n17435), .ZN(P3_U2788) );
  AOI22_X1 U20622 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17448), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17454), .ZN(n17436) );
  OAI21_X1 U20623 ( .B1(n18186), .B2(n17450), .A(n17436), .ZN(P3_U2789) );
  AOI22_X1 U20624 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17448), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17454), .ZN(n17437) );
  OAI21_X1 U20625 ( .B1(n18191), .B2(n17450), .A(n17437), .ZN(P3_U2790) );
  AOI22_X1 U20626 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17454), .ZN(n17438) );
  OAI21_X1 U20627 ( .B1(n17439), .B2(n17457), .A(n17438), .ZN(P3_U2791) );
  AOI22_X1 U20628 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17448), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17454), .ZN(n17440) );
  OAI21_X1 U20629 ( .B1(n17441), .B2(n17450), .A(n17440), .ZN(P3_U2792) );
  AOI22_X1 U20630 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17448), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17454), .ZN(n17442) );
  OAI21_X1 U20631 ( .B1(n17443), .B2(n17450), .A(n17442), .ZN(P3_U2793) );
  AOI22_X1 U20632 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17448), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17454), .ZN(n17444) );
  OAI21_X1 U20633 ( .B1(n17445), .B2(n17450), .A(n17444), .ZN(P3_U2794) );
  AOI22_X1 U20634 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17448), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17454), .ZN(n17446) );
  OAI21_X1 U20635 ( .B1(n17447), .B2(n17450), .A(n17446), .ZN(P3_U2795) );
  AOI22_X1 U20636 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17448), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17454), .ZN(n17449) );
  OAI21_X1 U20637 ( .B1(n17451), .B2(n17450), .A(n17449), .ZN(P3_U2796) );
  AOI22_X1 U20638 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17454), .ZN(n17452) );
  OAI21_X1 U20639 ( .B1(n17453), .B2(n17457), .A(n17452), .ZN(P3_U2797) );
  AOI22_X1 U20640 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17454), .ZN(n17456) );
  OAI21_X1 U20641 ( .B1(n17458), .B2(n17457), .A(n17456), .ZN(P3_U2798) );
  AOI22_X1 U20642 ( .A1(n17462), .A2(n17788), .B1(n17459), .B2(n17664), .ZN(
        n17460) );
  AND2_X1 U20643 ( .A1(n17827), .A2(n17460), .ZN(n17488) );
  OAI21_X1 U20644 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17564), .A(
        n17488), .ZN(n17478) );
  NOR2_X1 U20645 ( .A1(n17739), .A2(n17816), .ZN(n17571) );
  OAI22_X1 U20646 ( .A1(n17834), .A2(n9615), .B1(n17461), .B2(n17832), .ZN(
        n17494) );
  NOR2_X1 U20647 ( .A1(n17484), .A2(n17494), .ZN(n17485) );
  NOR3_X1 U20648 ( .A1(n17571), .A2(n17485), .A3(n20916), .ZN(n17468) );
  NAND2_X1 U20649 ( .A1(n18044), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17465) );
  INV_X1 U20650 ( .A(n17617), .ZN(n17578) );
  NOR2_X1 U20651 ( .A1(n17578), .A2(n17462), .ZN(n17482) );
  OAI211_X1 U20652 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17482), .B(n17463), .ZN(n17464) );
  OAI211_X1 U20653 ( .C1(n17666), .C2(n17466), .A(n17465), .B(n17464), .ZN(
        n17467) );
  AOI211_X1 U20654 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17478), .A(
        n17468), .B(n17467), .ZN(n17473) );
  OAI211_X1 U20655 ( .C1(n17471), .C2(n17470), .A(n17722), .B(n17469), .ZN(
        n17472) );
  OAI211_X1 U20656 ( .C1(n9635), .C2(n17474), .A(n17473), .B(n17472), .ZN(
        P3_U2802) );
  NOR2_X1 U20657 ( .A1(n16400), .A2(n17475), .ZN(n17476) );
  XOR2_X1 U20658 ( .A(n17476), .B(n17632), .Z(n17842) );
  AOI22_X1 U20659 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17478), .B1(
        n17682), .B2(n17477), .ZN(n17479) );
  NAND2_X1 U20660 ( .A1(n18044), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17840) );
  OAI211_X1 U20661 ( .C1(n17842), .C2(n17737), .A(n17479), .B(n17840), .ZN(
        n17480) );
  AOI21_X1 U20662 ( .B1(n17482), .B2(n17481), .A(n17480), .ZN(n17483) );
  OAI221_X1 U20663 ( .B1(n17485), .B2(n17484), .C1(n17485), .C2(n9635), .A(
        n17483), .ZN(P3_U2803) );
  NAND3_X1 U20664 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n17843), .ZN(n17849) );
  NAND2_X1 U20665 ( .A1(n17497), .A2(n17599), .ZN(n17524) );
  INV_X1 U20666 ( .A(n17564), .ZN(n17490) );
  AOI21_X1 U20667 ( .B1(n17486), .B2(n18542), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17487) );
  OAI22_X1 U20668 ( .A1(n17488), .A2(n17487), .B1(n18137), .B2(n18735), .ZN(
        n17489) );
  AOI221_X1 U20669 ( .B1(n17682), .B2(n17491), .C1(n17490), .C2(n17491), .A(
        n17489), .ZN(n17496) );
  OAI21_X1 U20670 ( .B1(n17493), .B2(n17843), .A(n17492), .ZN(n17846) );
  AOI22_X1 U20671 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17494), .B1(
        n17722), .B2(n17846), .ZN(n17495) );
  OAI211_X1 U20672 ( .C1(n17849), .C2(n17524), .A(n17496), .B(n17495), .ZN(
        P3_U2804) );
  NAND2_X1 U20673 ( .A1(n17958), .A2(n17497), .ZN(n17865) );
  NOR2_X1 U20674 ( .A1(n17865), .A2(n17878), .ZN(n17498) );
  XOR2_X1 U20675 ( .A(n17498), .B(n17855), .Z(n17857) );
  OAI21_X1 U20676 ( .B1(n17499), .B2(n17828), .A(n17827), .ZN(n17500) );
  AOI21_X1 U20677 ( .B1(n18542), .B2(n17501), .A(n17500), .ZN(n17530) );
  OAI21_X1 U20678 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17828), .A(
        n17530), .ZN(n17516) );
  INV_X1 U20679 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17531) );
  NAND4_X1 U20680 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n9592), .A3(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A4(n17617), .ZN(n17532) );
  NOR2_X1 U20681 ( .A1(n17531), .A2(n17532), .ZN(n17518) );
  OAI211_X1 U20682 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17518), .B(n17502), .ZN(n17503) );
  NAND2_X1 U20683 ( .A1(n9577), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17862) );
  OAI211_X1 U20684 ( .C1(n17666), .C2(n17504), .A(n17503), .B(n17862), .ZN(
        n17505) );
  AOI21_X1 U20685 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n17516), .A(
        n17505), .ZN(n17512) );
  NOR2_X1 U20686 ( .A1(n17887), .A2(n17506), .ZN(n17868) );
  NAND2_X1 U20687 ( .A1(n17868), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17507) );
  XOR2_X1 U20688 ( .A(n17507), .B(n17855), .Z(n17860) );
  AOI21_X1 U20689 ( .B1(n17632), .B2(n17509), .A(n17508), .ZN(n17510) );
  XOR2_X1 U20690 ( .A(n17510), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17861) );
  AOI22_X1 U20691 ( .A1(n17816), .A2(n17860), .B1(n17722), .B2(n17861), .ZN(
        n17511) );
  OAI211_X1 U20692 ( .C1(n17857), .C2(n9615), .A(n17512), .B(n17511), .ZN(
        P3_U2805) );
  AOI22_X1 U20693 ( .A1(n9577), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n17682), 
        .B2(n17513), .ZN(n17514) );
  INV_X1 U20694 ( .A(n17514), .ZN(n17515) );
  AOI221_X1 U20695 ( .B1(n17518), .B2(n17517), .C1(n17516), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17515), .ZN(n17523) );
  INV_X1 U20696 ( .A(n17865), .ZN(n17519) );
  OAI22_X1 U20697 ( .A1(n17868), .A2(n17832), .B1(n17519), .B2(n9615), .ZN(
        n17534) );
  OAI21_X1 U20698 ( .B1(n17521), .B2(n17878), .A(n17520), .ZN(n17875) );
  AOI22_X1 U20699 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17534), .B1(
        n17722), .B2(n17875), .ZN(n17522) );
  OAI211_X1 U20700 ( .C1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n17524), .A(
        n17523), .B(n17522), .ZN(P3_U2806) );
  OAI21_X1 U20701 ( .B1(n17595), .B2(n17880), .A(n17539), .ZN(n17526) );
  OAI211_X1 U20702 ( .C1(n17632), .C2(n17896), .A(n17526), .B(n17525), .ZN(
        n17527) );
  XNOR2_X1 U20703 ( .A(n17870), .B(n17527), .ZN(n17886) );
  AOI22_X1 U20704 ( .A1(n18044), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n17682), 
        .B2(n17528), .ZN(n17529) );
  OAI221_X1 U20705 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17532), .C1(
        n17531), .C2(n17530), .A(n17529), .ZN(n17533) );
  AOI221_X1 U20706 ( .B1(n17535), .B2(n17870), .C1(n17534), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17533), .ZN(n17536) );
  OAI21_X1 U20707 ( .B1(n17737), .B2(n17886), .A(n17536), .ZN(P3_U2807) );
  INV_X1 U20708 ( .A(n17897), .ZN(n17537) );
  NAND2_X1 U20709 ( .A1(n17933), .A2(n17537), .ZN(n17541) );
  AOI221_X1 U20710 ( .B1(n17612), .B2(n17539), .C1(n17541), .C2(n17539), .A(
        n17538), .ZN(n17540) );
  XOR2_X1 U20711 ( .A(n17896), .B(n17540), .Z(n17902) );
  NOR2_X1 U20712 ( .A1(n17622), .A2(n17541), .ZN(n17550) );
  INV_X1 U20713 ( .A(n17541), .ZN(n17893) );
  NOR2_X1 U20714 ( .A1(n17958), .A2(n9615), .ZN(n17642) );
  AOI21_X1 U20715 ( .B1(n17816), .B2(n17887), .A(n17642), .ZN(n17623) );
  OAI21_X1 U20716 ( .B1(n17571), .B2(n17893), .A(n17623), .ZN(n17560) );
  NAND2_X1 U20717 ( .A1(n9592), .A2(n17617), .ZN(n17556) );
  NAND2_X1 U20718 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17542) );
  OAI21_X1 U20719 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17542), .ZN(n17548) );
  INV_X1 U20720 ( .A(n17788), .ZN(n17727) );
  OAI22_X1 U20721 ( .A1(n9592), .A2(n17727), .B1(n17543), .B2(n17828), .ZN(
        n17544) );
  NOR2_X1 U20722 ( .A1(n17786), .A2(n17544), .ZN(n17565) );
  OAI21_X1 U20723 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17564), .A(
        n17565), .ZN(n17558) );
  AOI22_X1 U20724 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17558), .B1(
        n17682), .B2(n17545), .ZN(n17547) );
  NAND2_X1 U20725 ( .A1(n18044), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17546) );
  OAI211_X1 U20726 ( .C1(n17556), .C2(n17548), .A(n17547), .B(n17546), .ZN(
        n17549) );
  AOI221_X1 U20727 ( .B1(n17550), .B2(n17896), .C1(n17560), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n17549), .ZN(n17551) );
  OAI21_X1 U20728 ( .B1(n17737), .B2(n17902), .A(n17551), .ZN(P3_U2808) );
  AND3_X1 U20729 ( .A1(n17632), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17552), .ZN(n17574) );
  AOI22_X1 U20730 ( .A1(n17894), .A2(n17574), .B1(n17553), .B2(n17595), .ZN(
        n17554) );
  XOR2_X1 U20731 ( .A(n17554), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .Z(
        n17912) );
  NOR2_X1 U20732 ( .A1(n18137), .A2(n18726), .ZN(n17909) );
  OAI22_X1 U20733 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17556), .B1(
        n17555), .B2(n17666), .ZN(n17557) );
  AOI211_X1 U20734 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n17558), .A(
        n17909), .B(n17557), .ZN(n17562) );
  NOR2_X1 U20735 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17559), .ZN(
        n17910) );
  NAND2_X1 U20736 ( .A1(n17933), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17891) );
  NOR2_X1 U20737 ( .A1(n17622), .A2(n17891), .ZN(n17585) );
  AOI22_X1 U20738 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17560), .B1(
        n17910), .B2(n17585), .ZN(n17561) );
  OAI211_X1 U20739 ( .C1(n17912), .C2(n17737), .A(n17562), .B(n17561), .ZN(
        P3_U2809) );
  OAI221_X1 U20740 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17593), 
        .C1(n17922), .C2(n17574), .A(n17525), .ZN(n17563) );
  XOR2_X1 U20741 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17563), .Z(
        n17921) );
  NAND2_X1 U20742 ( .A1(n17666), .A2(n17564), .ZN(n17819) );
  INV_X1 U20743 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18723) );
  NOR2_X1 U20744 ( .A1(n18137), .A2(n18723), .ZN(n17569) );
  AOI221_X1 U20745 ( .B1(n17567), .B2(n17566), .C1(n18313), .C2(n17566), .A(
        n17565), .ZN(n17568) );
  AOI211_X1 U20746 ( .C1(n17570), .C2(n17819), .A(n17569), .B(n17568), .ZN(
        n17573) );
  NOR2_X1 U20747 ( .A1(n17922), .A2(n17891), .ZN(n17914) );
  OAI21_X1 U20748 ( .B1(n17571), .B2(n17914), .A(n17623), .ZN(n17584) );
  NOR2_X1 U20749 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17922), .ZN(
        n17913) );
  AOI22_X1 U20750 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17584), .B1(
        n17585), .B2(n17913), .ZN(n17572) );
  OAI211_X1 U20751 ( .C1(n17737), .C2(n17921), .A(n17573), .B(n17572), .ZN(
        P3_U2810) );
  AOI21_X1 U20752 ( .B1(n17593), .B2(n17595), .A(n17574), .ZN(n17575) );
  XOR2_X1 U20753 ( .A(n17575), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n17927) );
  INV_X1 U20754 ( .A(n17824), .ZN(n17703) );
  OAI21_X1 U20755 ( .B1(n17786), .B2(n17577), .A(n17703), .ZN(n17600) );
  OAI21_X1 U20756 ( .B1(n17576), .B2(n17828), .A(n17600), .ZN(n17590) );
  AOI22_X1 U20757 ( .A1(n18044), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17590), .ZN(n17581) );
  NOR2_X1 U20758 ( .A1(n17578), .A2(n17577), .ZN(n17592) );
  NAND2_X1 U20759 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17579) );
  OAI211_X1 U20760 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17592), .B(n17579), .ZN(n17580) );
  OAI211_X1 U20761 ( .C1(n17666), .C2(n17582), .A(n17581), .B(n17580), .ZN(
        n17583) );
  AOI221_X1 U20762 ( .B1(n17585), .B2(n17922), .C1(n17584), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17583), .ZN(n17586) );
  OAI21_X1 U20763 ( .B1(n17927), .B2(n17737), .A(n17586), .ZN(P3_U2811) );
  OAI21_X1 U20764 ( .B1(n17622), .B2(n17933), .A(n17623), .ZN(n17587) );
  INV_X1 U20765 ( .A(n17587), .ZN(n17610) );
  INV_X1 U20766 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17904) );
  OAI22_X1 U20767 ( .A1(n18137), .A2(n18719), .B1(n17666), .B2(n17588), .ZN(
        n17589) );
  AOI221_X1 U20768 ( .B1(n17592), .B2(n17591), .C1(n17590), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17589), .ZN(n17598) );
  AOI21_X1 U20769 ( .B1(n17632), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17593), .ZN(n17594) );
  XOR2_X1 U20770 ( .A(n17595), .B(n17594), .Z(n17938) );
  NOR2_X1 U20771 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17596), .ZN(
        n17937) );
  AOI22_X1 U20772 ( .A1(n17722), .A2(n17938), .B1(n17599), .B2(n17937), .ZN(
        n17597) );
  OAI211_X1 U20773 ( .C1(n17610), .C2(n17904), .A(n17598), .B(n17597), .ZN(
        P3_U2812) );
  AOI21_X1 U20774 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17599), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17609) );
  AOI221_X1 U20775 ( .B1(n17602), .B2(n17601), .C1(n18313), .C2(n17601), .A(
        n17600), .ZN(n17603) );
  AOI21_X1 U20776 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n18044), .A(n17603), 
        .ZN(n17608) );
  OAI21_X1 U20777 ( .B1(n17605), .B2(n17943), .A(n17604), .ZN(n17941) );
  AOI22_X1 U20778 ( .A1(n17722), .A2(n17941), .B1(n17606), .B2(n17819), .ZN(
        n17607) );
  OAI211_X1 U20779 ( .C1(n17610), .C2(n17609), .A(n17608), .B(n17607), .ZN(
        P3_U2813) );
  NOR2_X1 U20780 ( .A1(n17734), .A2(n17611), .ZN(n17719) );
  AOI22_X1 U20781 ( .A1(n17719), .A2(n17888), .B1(n17612), .B2(n17734), .ZN(
        n17613) );
  XOR2_X1 U20782 ( .A(n17613), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .Z(
        n17957) );
  OAI21_X1 U20783 ( .B1(n17727), .B2(n17614), .A(n17827), .ZN(n17615) );
  INV_X1 U20784 ( .A(n17615), .ZN(n17651) );
  OAI21_X1 U20785 ( .B1(n17616), .B2(n17828), .A(n17651), .ZN(n17629) );
  NAND2_X1 U20786 ( .A1(n17661), .A2(n17617), .ZN(n17678) );
  NOR2_X1 U20787 ( .A1(n17618), .A2(n17678), .ZN(n17631) );
  NAND2_X1 U20788 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17619) );
  OAI211_X1 U20789 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17631), .B(n17619), .ZN(n17620) );
  NAND2_X1 U20790 ( .A1(n18044), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n17955) );
  OAI211_X1 U20791 ( .C1(n17666), .C2(n17621), .A(n17620), .B(n17955), .ZN(
        n17625) );
  AOI22_X1 U20792 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17623), .B1(
        n17622), .B2(n17952), .ZN(n17624) );
  AOI211_X1 U20793 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n17629), .A(
        n17625), .B(n17624), .ZN(n17626) );
  OAI21_X1 U20794 ( .B1(n17957), .B2(n17737), .A(n17626), .ZN(P3_U2814) );
  NAND2_X1 U20795 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17636) );
  INV_X1 U20796 ( .A(n17698), .ZN(n18009) );
  NOR2_X1 U20797 ( .A1(n17975), .A2(n18009), .ZN(n17670) );
  INV_X1 U20798 ( .A(n17670), .ZN(n17990) );
  NOR2_X1 U20799 ( .A1(n17636), .A2(n17990), .ZN(n17653) );
  NOR2_X1 U20800 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17653), .ZN(
        n17967) );
  NAND2_X1 U20801 ( .A1(n17816), .A2(n17887), .ZN(n17646) );
  NAND2_X1 U20802 ( .A1(n18044), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n17970) );
  OAI21_X1 U20803 ( .B1(n17666), .B2(n17627), .A(n17970), .ZN(n17628) );
  AOI221_X1 U20804 ( .B1(n17631), .B2(n17630), .C1(n17629), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17628), .ZN(n17645) );
  NAND2_X1 U20805 ( .A1(n17632), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17671) );
  INV_X1 U20806 ( .A(n17671), .ZN(n17638) );
  NOR2_X1 U20807 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17633), .ZN(
        n17720) );
  NAND2_X1 U20808 ( .A1(n17634), .A2(n17720), .ZN(n17683) );
  NOR2_X1 U20809 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17683), .ZN(
        n17655) );
  NAND2_X1 U20810 ( .A1(n18006), .A2(n17635), .ZN(n17672) );
  NOR2_X1 U20811 ( .A1(n17636), .A2(n17672), .ZN(n17637) );
  OAI22_X1 U20812 ( .A1(n17639), .A2(n17638), .B1(n17655), .B2(n17637), .ZN(
        n17640) );
  XOR2_X1 U20813 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17640), .Z(
        n17972) );
  INV_X1 U20814 ( .A(n17972), .ZN(n17643) );
  NAND2_X1 U20815 ( .A1(n17647), .A2(n17641), .ZN(n17959) );
  AOI22_X1 U20816 ( .A1(n17722), .A2(n17643), .B1(n17642), .B2(n17959), .ZN(
        n17644) );
  OAI211_X1 U20817 ( .C1(n17967), .C2(n17646), .A(n17645), .B(n17644), .ZN(
        P3_U2815) );
  OAI221_X1 U20818 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17993), .A(n17647), .ZN(
        n17978) );
  AND3_X1 U20819 ( .A1(n9684), .A2(n17648), .A3(n18542), .ZN(n17694) );
  AOI21_X1 U20820 ( .B1(n17660), .B2(n17694), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17650) );
  OAI22_X1 U20821 ( .A1(n17651), .A2(n17650), .B1(n17811), .B2(n17649), .ZN(
        n17652) );
  AOI21_X1 U20822 ( .B1(n18044), .B2(P3_REIP_REG_14__SCAN_IN), .A(n17652), 
        .ZN(n17659) );
  INV_X1 U20823 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17657) );
  AOI221_X1 U20824 ( .B1(n17654), .B2(n17657), .C1(n17990), .C2(n17657), .A(
        n17653), .ZN(n17982) );
  INV_X1 U20825 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17998) );
  AOI22_X1 U20826 ( .A1(n17719), .A2(n17977), .B1(n17655), .B2(n17998), .ZN(
        n17656) );
  XOR2_X1 U20827 ( .A(n17657), .B(n17656), .Z(n17983) );
  AOI22_X1 U20828 ( .A1(n17816), .A2(n17982), .B1(n17722), .B2(n17983), .ZN(
        n17658) );
  OAI211_X1 U20829 ( .C1(n9615), .C2(n17978), .A(n17659), .B(n17658), .ZN(
        P3_U2816) );
  OR2_X1 U20830 ( .A1(n17975), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17997) );
  AOI211_X1 U20831 ( .C1(n17677), .C2(n17667), .A(n17660), .B(n17678), .ZN(
        n17669) );
  OAI21_X1 U20832 ( .B1(n17661), .B2(n17727), .A(n17827), .ZN(n17662) );
  AOI21_X1 U20833 ( .B1(n17664), .B2(n17663), .A(n17662), .ZN(n17676) );
  OAI22_X1 U20834 ( .A1(n17676), .A2(n17667), .B1(n17666), .B2(n17665), .ZN(
        n17668) );
  AOI211_X1 U20835 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n9577), .A(n17669), .B(
        n17668), .ZN(n17675) );
  OAI22_X1 U20836 ( .A1(n17993), .A2(n9615), .B1(n17670), .B2(n17832), .ZN(
        n17686) );
  AOI22_X1 U20837 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17672), .B1(
        n17671), .B2(n17683), .ZN(n17673) );
  XOR2_X1 U20838 ( .A(n17673), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n17987) );
  AOI22_X1 U20839 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17686), .B1(
        n17722), .B2(n17987), .ZN(n17674) );
  OAI211_X1 U20840 ( .C1(n17726), .C2(n17997), .A(n17675), .B(n17674), .ZN(
        P3_U2817) );
  NOR3_X1 U20841 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17726), .A3(
        n17989), .ZN(n17680) );
  NAND2_X1 U20842 ( .A1(n9577), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18002) );
  OAI221_X1 U20843 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17678), .C1(
        n17677), .C2(n17676), .A(n18002), .ZN(n17679) );
  AOI211_X1 U20844 ( .C1(n17682), .C2(n17681), .A(n17680), .B(n17679), .ZN(
        n17688) );
  INV_X1 U20845 ( .A(n17719), .ZN(n17684) );
  OAI21_X1 U20846 ( .B1(n17684), .B2(n17989), .A(n17683), .ZN(n17685) );
  XOR2_X1 U20847 ( .A(n17685), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18001) );
  AOI22_X1 U20848 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17686), .B1(
        n17722), .B2(n18001), .ZN(n17687) );
  NAND2_X1 U20849 ( .A1(n17688), .A2(n17687), .ZN(P3_U2818) );
  INV_X1 U20850 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17690) );
  NAND2_X1 U20851 ( .A1(n17697), .A2(n17690), .ZN(n18019) );
  NOR2_X1 U20852 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17708) );
  AOI22_X1 U20853 ( .A1(n17697), .A2(n17719), .B1(n17708), .B2(n17720), .ZN(
        n17689) );
  XOR2_X1 U20854 ( .A(n17690), .B(n17689), .Z(n18005) );
  INV_X1 U20855 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18705) );
  NOR2_X1 U20856 ( .A1(n18137), .A2(n18705), .ZN(n17696) );
  NAND4_X1 U20857 ( .A1(n9684), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A4(n18542), .ZN(n17715) );
  NOR2_X1 U20858 ( .A1(n17691), .A2(n17715), .ZN(n17706) );
  AOI21_X1 U20859 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17703), .A(
        n17706), .ZN(n17693) );
  OAI22_X1 U20860 ( .A1(n17694), .A2(n17693), .B1(n17811), .B2(n17692), .ZN(
        n17695) );
  AOI211_X1 U20861 ( .C1(n17722), .C2(n18005), .A(n17696), .B(n17695), .ZN(
        n17701) );
  NOR2_X1 U20862 ( .A1(n17697), .A2(n17726), .ZN(n17710) );
  OAI22_X1 U20863 ( .A1(n17699), .A2(n9615), .B1(n17832), .B2(n17698), .ZN(
        n17723) );
  OAI21_X1 U20864 ( .B1(n17710), .B2(n17723), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17700) );
  OAI211_X1 U20865 ( .C1(n17726), .C2(n18019), .A(n17701), .B(n17700), .ZN(
        P3_U2819) );
  INV_X1 U20866 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18036) );
  AOI22_X1 U20867 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17719), .B1(
        n17720), .B2(n18036), .ZN(n17702) );
  XOR2_X1 U20868 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n17702), .Z(
        n18026) );
  NOR2_X1 U20869 ( .A1(n17714), .A2(n17715), .ZN(n17713) );
  AOI21_X1 U20870 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17703), .A(
        n17713), .ZN(n17705) );
  OAI22_X1 U20871 ( .A1(n17706), .A2(n17705), .B1(n17811), .B2(n17704), .ZN(
        n17707) );
  AOI21_X1 U20872 ( .B1(n18044), .B2(P3_REIP_REG_10__SCAN_IN), .A(n17707), 
        .ZN(n17712) );
  INV_X1 U20873 ( .A(n17708), .ZN(n17709) );
  AOI22_X1 U20874 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17723), .B1(
        n17710), .B2(n17709), .ZN(n17711) );
  OAI211_X1 U20875 ( .C1(n18026), .C2(n17737), .A(n17712), .B(n17711), .ZN(
        P3_U2820) );
  AOI211_X1 U20876 ( .C1(n17715), .C2(n17714), .A(n17824), .B(n17713), .ZN(
        n17717) );
  NOR2_X1 U20877 ( .A1(n18137), .A2(n18701), .ZN(n17716) );
  AOI211_X1 U20878 ( .C1(n17718), .C2(n17819), .A(n17717), .B(n17716), .ZN(
        n17725) );
  NOR2_X1 U20879 ( .A1(n17720), .A2(n17719), .ZN(n17721) );
  XOR2_X1 U20880 ( .A(n17721), .B(n18036), .Z(n18032) );
  AOI22_X1 U20881 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17723), .B1(
        n17722), .B2(n18032), .ZN(n17724) );
  OAI211_X1 U20882 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n17726), .A(
        n17725), .B(n17724), .ZN(P3_U2821) );
  OAI21_X1 U20883 ( .B1(n9684), .B2(n17727), .A(n17827), .ZN(n17747) );
  INV_X1 U20884 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17728) );
  AOI221_X1 U20885 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C1(n17729), .C2(n17728), .A(n18313), .ZN(n17731) );
  NOR2_X1 U20886 ( .A1(n18137), .A2(n18700), .ZN(n17730) );
  AOI211_X1 U20887 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17747), .A(
        n17731), .B(n17730), .ZN(n17741) );
  AOI21_X1 U20888 ( .B1(n17734), .B2(n18042), .A(n17733), .ZN(n18052) );
  OAI21_X1 U20889 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17736), .A(
        n17735), .ZN(n18039) );
  OAI22_X1 U20890 ( .A1(n18052), .A2(n17737), .B1(n17832), .B2(n18039), .ZN(
        n17738) );
  AOI21_X1 U20891 ( .B1(n17739), .B2(n9941), .A(n17738), .ZN(n17740) );
  OAI211_X1 U20892 ( .C1(n17811), .C2(n17742), .A(n17741), .B(n17740), .ZN(
        P3_U2822) );
  OAI21_X1 U20893 ( .B1(n17745), .B2(n17744), .A(n17743), .ZN(n17746) );
  XOR2_X1 U20894 ( .A(n17746), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18061) );
  AND2_X1 U20895 ( .A1(n9684), .A2(n18542), .ZN(n17749) );
  NOR2_X1 U20896 ( .A1(n18137), .A2(n18697), .ZN(n18053) );
  AOI221_X1 U20897 ( .B1(n17749), .B2(n17748), .C1(n17747), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18053), .ZN(n17754) );
  AOI21_X1 U20898 ( .B1(n18054), .B2(n17751), .A(n17750), .ZN(n18058) );
  AOI22_X1 U20899 ( .A1(n17820), .A2(n18058), .B1(n17752), .B2(n17819), .ZN(
        n17753) );
  OAI211_X1 U20900 ( .C1(n17832), .C2(n18061), .A(n17754), .B(n17753), .ZN(
        P3_U2823) );
  AOI21_X1 U20901 ( .B1(n17757), .B2(n17756), .A(n17755), .ZN(n18065) );
  NOR2_X1 U20902 ( .A1(n17758), .A2(n18313), .ZN(n17760) );
  AOI22_X1 U20903 ( .A1(n17820), .A2(n18065), .B1(n17760), .B2(n17759), .ZN(
        n17766) );
  NOR2_X1 U20904 ( .A1(n17824), .A2(n17760), .ZN(n17778) );
  OAI21_X1 U20905 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17762), .A(
        n17761), .ZN(n18068) );
  OAI22_X1 U20906 ( .A1(n17811), .A2(n17763), .B1(n17832), .B2(n18068), .ZN(
        n17764) );
  AOI21_X1 U20907 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17778), .A(
        n17764), .ZN(n17765) );
  OAI211_X1 U20908 ( .C1(n18137), .C2(n18695), .A(n17766), .B(n17765), .ZN(
        P3_U2824) );
  OAI21_X1 U20909 ( .B1(n17769), .B2(n17768), .A(n17767), .ZN(n18070) );
  OAI21_X1 U20910 ( .B1(n17786), .B2(n17770), .A(n9757), .ZN(n17777) );
  INV_X1 U20911 ( .A(n17820), .ZN(n17831) );
  OAI21_X1 U20912 ( .B1(n17773), .B2(n17772), .A(n17771), .ZN(n17774) );
  XOR2_X1 U20913 ( .A(n17774), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n18075) );
  OAI22_X1 U20914 ( .A1(n17811), .A2(n17775), .B1(n17831), .B2(n18075), .ZN(
        n17776) );
  AOI21_X1 U20915 ( .B1(n17778), .B2(n17777), .A(n17776), .ZN(n17779) );
  NAND2_X1 U20916 ( .A1(n18044), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18069) );
  OAI211_X1 U20917 ( .C1(n17832), .C2(n18070), .A(n17779), .B(n18069), .ZN(
        P3_U2825) );
  OAI21_X1 U20918 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n17781), .A(
        n17780), .ZN(n18088) );
  AOI22_X1 U20919 ( .A1(n9577), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18542), .B2(
        n17782), .ZN(n17793) );
  AOI21_X1 U20920 ( .B1(n17785), .B2(n17784), .A(n17783), .ZN(n18086) );
  AOI21_X1 U20921 ( .B1(n17788), .B2(n17787), .A(n17786), .ZN(n17801) );
  OAI22_X1 U20922 ( .A1(n17811), .A2(n17790), .B1(n17801), .B2(n17789), .ZN(
        n17791) );
  AOI21_X1 U20923 ( .B1(n17820), .B2(n18086), .A(n17791), .ZN(n17792) );
  OAI211_X1 U20924 ( .C1(n17832), .C2(n18088), .A(n17793), .B(n17792), .ZN(
        P3_U2826) );
  OAI21_X1 U20925 ( .B1(n17796), .B2(n17795), .A(n17794), .ZN(n18097) );
  AOI21_X1 U20926 ( .B1(n18093), .B2(n17798), .A(n17797), .ZN(n18095) );
  AOI21_X1 U20927 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17827), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17800) );
  OAI22_X1 U20928 ( .A1(n17801), .A2(n17800), .B1(n17811), .B2(n17799), .ZN(
        n17802) );
  AOI21_X1 U20929 ( .B1(n17820), .B2(n18095), .A(n17802), .ZN(n17803) );
  NAND2_X1 U20930 ( .A1(n9577), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18092) );
  OAI211_X1 U20931 ( .C1(n17832), .C2(n18097), .A(n17803), .B(n18092), .ZN(
        P3_U2827) );
  AOI21_X1 U20932 ( .B1(n17806), .B2(n17805), .A(n17804), .ZN(n18112) );
  INV_X1 U20933 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18687) );
  NOR2_X1 U20934 ( .A1(n18137), .A2(n18687), .ZN(n18113) );
  OAI21_X1 U20935 ( .B1(n17809), .B2(n17808), .A(n17807), .ZN(n18108) );
  OAI22_X1 U20936 ( .A1(n17811), .A2(n17810), .B1(n17832), .B2(n18108), .ZN(
        n17812) );
  AOI211_X1 U20937 ( .C1(n17820), .C2(n18112), .A(n18113), .B(n17812), .ZN(
        n17813) );
  OAI221_X1 U20938 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18313), .C1(
        n17814), .C2(n17827), .A(n17813), .ZN(P3_U2828) );
  NOR2_X1 U20939 ( .A1(n17826), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17815) );
  XNOR2_X1 U20940 ( .A(n17815), .B(n17818), .ZN(n18118) );
  AOI22_X1 U20941 ( .A1(n17816), .A2(n18118), .B1(n9577), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17822) );
  AOI21_X1 U20942 ( .B1(n17825), .B2(n17818), .A(n17817), .ZN(n18123) );
  AOI22_X1 U20943 ( .A1(n17820), .A2(n18123), .B1(n17823), .B2(n17819), .ZN(
        n17821) );
  OAI211_X1 U20944 ( .C1(n17824), .C2(n17823), .A(n17822), .B(n17821), .ZN(
        P3_U2829) );
  OAI21_X1 U20945 ( .B1(n17826), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17825), .ZN(n18133) );
  INV_X1 U20946 ( .A(n18133), .ZN(n18131) );
  NAND3_X1 U20947 ( .A1(n18770), .A2(n17828), .A3(n17827), .ZN(n17829) );
  AOI22_X1 U20948 ( .A1(n18044), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17829), .ZN(n17830) );
  OAI221_X1 U20949 ( .B1(n18131), .B2(n17832), .C1(n18133), .C2(n17831), .A(
        n17830), .ZN(P3_U2830) );
  NAND2_X1 U20950 ( .A1(n18137), .A2(n18116), .ZN(n18120) );
  OAI21_X1 U20951 ( .B1(n17834), .B2(n18041), .A(n17833), .ZN(n17835) );
  AOI21_X1 U20952 ( .B1(n18597), .B2(n17836), .A(n17835), .ZN(n17844) );
  AOI21_X1 U20953 ( .B1(n18129), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17837), .ZN(n17838) );
  AOI21_X1 U20954 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17844), .A(
        n17838), .ZN(n17839) );
  AOI21_X1 U20955 ( .B1(n18114), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17839), .ZN(n17841) );
  OAI211_X1 U20956 ( .C1(n17842), .C2(n18051), .A(n17841), .B(n17840), .ZN(
        P3_U2835) );
  OR2_X1 U20957 ( .A1(n17851), .A2(n17903), .ZN(n17879) );
  AOI211_X1 U20958 ( .C1(n18129), .C2(n17844), .A(n9577), .B(n17843), .ZN(
        n17845) );
  AOI21_X1 U20959 ( .B1(n18033), .B2(n17846), .A(n17845), .ZN(n17848) );
  NAND2_X1 U20960 ( .A1(n9577), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17847) );
  OAI211_X1 U20961 ( .C1(n17849), .C2(n17879), .A(n17848), .B(n17847), .ZN(
        P3_U2836) );
  NAND2_X1 U20962 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17855), .ZN(
        n17850) );
  NOR3_X1 U20963 ( .A1(n17852), .A2(n17851), .A3(n17850), .ZN(n17859) );
  NAND2_X1 U20964 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17854) );
  OAI21_X1 U20965 ( .B1(n17869), .B2(n18626), .A(n17866), .ZN(n17853) );
  AOI221_X1 U20966 ( .B1(n18609), .B2(n17854), .C1(n18078), .C2(n17854), .A(
        n17853), .ZN(n17856) );
  OAI22_X1 U20967 ( .A1(n17857), .A2(n18041), .B1(n17856), .B2(n17855), .ZN(
        n17858) );
  AOI211_X1 U20968 ( .C1(n18597), .C2(n17860), .A(n17859), .B(n17858), .ZN(
        n17864) );
  AOI22_X1 U20969 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18114), .B1(
        n18033), .B2(n17861), .ZN(n17863) );
  OAI211_X1 U20970 ( .C1(n17864), .C2(n18116), .A(n17863), .B(n17862), .ZN(
        P3_U2837) );
  AOI21_X1 U20971 ( .B1(n18008), .B2(n17865), .A(n18114), .ZN(n17867) );
  OAI211_X1 U20972 ( .C1(n17868), .C2(n18107), .A(n17867), .B(n17866), .ZN(
        n17873) );
  NOR2_X1 U20973 ( .A1(n17869), .A2(n18626), .ZN(n17871) );
  NOR3_X1 U20974 ( .A1(n17871), .A2(n17870), .A3(n17873), .ZN(n17872) );
  NOR2_X1 U20975 ( .A1(n17872), .A2(n18044), .ZN(n17881) );
  OAI21_X1 U20976 ( .B1(n17874), .B2(n17873), .A(n17881), .ZN(n17877) );
  AOI22_X1 U20977 ( .A1(n18044), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n18033), 
        .B2(n17875), .ZN(n17876) );
  OAI221_X1 U20978 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17879), 
        .C1(n17878), .C2(n17877), .A(n17876), .ZN(P3_U2838) );
  NAND2_X1 U20979 ( .A1(n9577), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17885) );
  NOR2_X1 U20980 ( .A1(n18114), .A2(n17880), .ZN(n17883) );
  OAI221_X1 U20981 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17883), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n17882), .A(n17881), .ZN(
        n17884) );
  OAI211_X1 U20982 ( .C1(n17886), .C2(n18051), .A(n17885), .B(n17884), .ZN(
        P3_U2839) );
  AOI22_X1 U20983 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18114), .B1(
        n9577), .B2(P3_REIP_REG_22__SCAN_IN), .ZN(n17901) );
  NAND2_X1 U20984 ( .A1(n18597), .A2(n17887), .ZN(n17968) );
  OAI21_X1 U20985 ( .B1(n17958), .B2(n18041), .A(n17968), .ZN(n17905) );
  NOR2_X1 U20986 ( .A1(n18787), .A2(n17949), .ZN(n18028) );
  NAND2_X1 U20987 ( .A1(n17888), .A2(n18028), .ZN(n17947) );
  AOI21_X1 U20988 ( .B1(n17889), .B2(n17914), .A(n18630), .ZN(n17890) );
  AOI221_X1 U20989 ( .B1(n17891), .B2(n18628), .C1(n17947), .C2(n18628), .A(
        n17890), .ZN(n17892) );
  OAI221_X1 U20990 ( .B1(n18626), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), 
        .C1(n18626), .C2(n17928), .A(n17892), .ZN(n17915) );
  NAND2_X1 U20991 ( .A1(n18107), .A2(n18041), .ZN(n18013) );
  INV_X1 U20992 ( .A(n18013), .ZN(n17932) );
  OAI22_X1 U20993 ( .A1(n9586), .A2(n17894), .B1(n17893), .B2(n17932), .ZN(
        n17895) );
  NOR2_X1 U20994 ( .A1(n17915), .A2(n17895), .ZN(n17907) );
  OAI211_X1 U20995 ( .C1(n9586), .C2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17907), .ZN(n17899) );
  OAI22_X1 U20996 ( .A1(n17897), .A2(n17903), .B1(n17896), .B2(n18116), .ZN(
        n17898) );
  OAI21_X1 U20997 ( .B1(n17905), .B2(n17899), .A(n17898), .ZN(n17900) );
  OAI211_X1 U20998 ( .C1(n18051), .C2(n17902), .A(n17901), .B(n17900), .ZN(
        P3_U2840) );
  NOR2_X1 U20999 ( .A1(n17904), .A2(n17903), .ZN(n17923) );
  AOI211_X1 U21000 ( .C1(n17951), .C2(n17907), .A(n9577), .B(n17906), .ZN(
        n17908) );
  AOI211_X1 U21001 ( .C1(n17910), .C2(n17923), .A(n17909), .B(n17908), .ZN(
        n17911) );
  OAI21_X1 U21002 ( .B1(n17912), .B2(n18051), .A(n17911), .ZN(P3_U2841) );
  AOI22_X1 U21003 ( .A1(n18044), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n17923), 
        .B2(n17913), .ZN(n17920) );
  INV_X1 U21004 ( .A(n17914), .ZN(n17916) );
  AOI21_X1 U21005 ( .B1(n17916), .B2(n18013), .A(n17915), .ZN(n17917) );
  AOI21_X1 U21006 ( .B1(n17951), .B2(n17917), .A(n9577), .ZN(n17924) );
  AND3_X1 U21007 ( .A1(n18119), .A2(n17922), .A3(P3_STATE2_REG_2__SCAN_IN), 
        .ZN(n17918) );
  OAI21_X1 U21008 ( .B1(n17924), .B2(n17918), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17919) );
  OAI211_X1 U21009 ( .C1(n18051), .C2(n17921), .A(n17920), .B(n17919), .ZN(
        P3_U2842) );
  AOI22_X1 U21010 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17924), .B1(
        n17923), .B2(n17922), .ZN(n17926) );
  NAND2_X1 U21011 ( .A1(n9577), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17925) );
  OAI211_X1 U21012 ( .C1(n17927), .C2(n18051), .A(n17926), .B(n17925), .ZN(
        P3_U2843) );
  NOR2_X1 U21013 ( .A1(n17928), .A2(n18626), .ZN(n17929) );
  AOI221_X1 U21014 ( .B1(n17952), .B2(n18078), .C1(n17930), .C2(n18078), .A(
        n17929), .ZN(n17931) );
  OAI211_X1 U21015 ( .C1(n17933), .C2(n17932), .A(n17951), .B(n17931), .ZN(
        n17942) );
  OAI221_X1 U21016 ( .B1(n17942), .B2(n17943), .C1(n17942), .C2(n18078), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17940) );
  OAI22_X1 U21017 ( .A1(n18079), .A2(n18626), .B1(n18077), .B2(n17934), .ZN(
        n18090) );
  NAND2_X1 U21018 ( .A1(n17935), .A2(n18090), .ZN(n18063) );
  NOR3_X1 U21019 ( .A1(n18055), .A2(n18054), .A3(n18063), .ZN(n18038) );
  NAND2_X1 U21020 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18038), .ZN(
        n17961) );
  NAND2_X1 U21021 ( .A1(n17936), .A2(n17961), .ZN(n18000) );
  NAND2_X1 U21022 ( .A1(n18129), .A2(n18000), .ZN(n18037) );
  NOR2_X1 U21023 ( .A1(n9944), .A2(n18037), .ZN(n17953) );
  AOI22_X1 U21024 ( .A1(n18033), .A2(n17938), .B1(n17953), .B2(n17937), .ZN(
        n17939) );
  OAI221_X1 U21025 ( .B1(n9577), .B2(n17940), .C1(n18137), .C2(n18719), .A(
        n17939), .ZN(P3_U2844) );
  AOI22_X1 U21026 ( .A1(n18044), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n18033), 
        .B2(n17941), .ZN(n17946) );
  NAND3_X1 U21027 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18137), .A3(
        n17942), .ZN(n17945) );
  NAND3_X1 U21028 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17953), .A3(
        n17943), .ZN(n17944) );
  NAND3_X1 U21029 ( .A1(n17946), .A2(n17945), .A3(n17944), .ZN(P3_U2845) );
  INV_X1 U21030 ( .A(n17947), .ZN(n17948) );
  AOI21_X1 U21031 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18029), .A(
        n17948), .ZN(n17950) );
  NAND2_X1 U21032 ( .A1(n18608), .A2(n17949), .ZN(n18027) );
  OAI21_X1 U21033 ( .B1(n18011), .B2(n18626), .A(n18027), .ZN(n17973) );
  AOI211_X1 U21034 ( .C1(n17960), .C2(n17988), .A(n17950), .B(n17973), .ZN(
        n17963) );
  AOI221_X1 U21035 ( .B1(n9586), .B2(n17951), .C1(n17963), .C2(n17951), .A(
        n9577), .ZN(n17954) );
  AOI22_X1 U21036 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17954), .B1(
        n17953), .B2(n17952), .ZN(n17956) );
  OAI211_X1 U21037 ( .C1(n17957), .C2(n18051), .A(n17956), .B(n17955), .ZN(
        P3_U2846) );
  OR2_X1 U21038 ( .A1(n18041), .A2(n17958), .ZN(n17966) );
  INV_X1 U21039 ( .A(n17959), .ZN(n17965) );
  INV_X1 U21040 ( .A(n17960), .ZN(n17962) );
  INV_X1 U21041 ( .A(n17961), .ZN(n17976) );
  AOI21_X1 U21042 ( .B1(n17962), .B2(n17976), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17964) );
  OAI222_X1 U21043 ( .A1(n17968), .A2(n17967), .B1(n17966), .B2(n17965), .C1(
        n17964), .C2(n17963), .ZN(n17969) );
  AOI22_X1 U21044 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18114), .B1(
        n18129), .B2(n17969), .ZN(n17971) );
  OAI211_X1 U21045 ( .C1(n17972), .C2(n18051), .A(n17971), .B(n17970), .ZN(
        P3_U2847) );
  INV_X1 U21046 ( .A(n18028), .ZN(n17974) );
  AOI221_X1 U21047 ( .B1(n17975), .B2(n18628), .C1(n17974), .C2(n18628), .A(
        n17973), .ZN(n17992) );
  OAI21_X1 U21048 ( .B1(n9586), .B2(n17977), .A(n17992), .ZN(n17981) );
  NAND2_X1 U21049 ( .A1(n17977), .A2(n17976), .ZN(n17979) );
  OAI22_X1 U21050 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17979), .B1(
        n17978), .B2(n18041), .ZN(n17980) );
  AOI21_X1 U21051 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17981), .A(
        n17980), .ZN(n17986) );
  AOI22_X1 U21052 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18114), .B1(
        n9577), .B2(P3_REIP_REG_14__SCAN_IN), .ZN(n17985) );
  AOI22_X1 U21053 ( .A1(n18033), .A2(n17983), .B1(n18134), .B2(n17982), .ZN(
        n17984) );
  OAI211_X1 U21054 ( .C1(n17986), .C2(n18116), .A(n17985), .B(n17984), .ZN(
        P3_U2848) );
  AOI22_X1 U21055 ( .A1(n9577), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18033), 
        .B2(n17987), .ZN(n17996) );
  AOI22_X1 U21056 ( .A1(n18597), .A2(n17990), .B1(n17989), .B2(n17988), .ZN(
        n17991) );
  OAI211_X1 U21057 ( .C1(n17993), .C2(n18041), .A(n17992), .B(n17991), .ZN(
        n17999) );
  OAI21_X1 U21058 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18022), .A(
        n18129), .ZN(n17994) );
  OAI211_X1 U21059 ( .C1(n17999), .C2(n17994), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18137), .ZN(n17995) );
  OAI211_X1 U21060 ( .C1(n17997), .C2(n18037), .A(n17996), .B(n17995), .ZN(
        P3_U2849) );
  OAI222_X1 U21061 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18006), 
        .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18000), .C1(n17999), 
        .C2(n17998), .ZN(n18004) );
  AOI22_X1 U21062 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18114), .B1(
        n18033), .B2(n18001), .ZN(n18003) );
  OAI211_X1 U21063 ( .C1(n18116), .C2(n18004), .A(n18003), .B(n18002), .ZN(
        P3_U2850) );
  AOI22_X1 U21064 ( .A1(n18044), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18033), 
        .B2(n18005), .ZN(n18018) );
  NOR2_X1 U21065 ( .A1(n18006), .A2(n18022), .ZN(n18016) );
  AOI21_X1 U21066 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18028), .A(
        n18029), .ZN(n18012) );
  AOI22_X1 U21067 ( .A1(n18597), .A2(n18009), .B1(n18008), .B2(n18007), .ZN(
        n18010) );
  OAI211_X1 U21068 ( .C1(n18011), .C2(n18626), .A(n18129), .B(n18010), .ZN(
        n18031) );
  AOI211_X1 U21069 ( .C1(n18014), .C2(n18013), .A(n18012), .B(n18031), .ZN(
        n18021) );
  OAI211_X1 U21070 ( .C1(n18029), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18021), .B(n18027), .ZN(n18015) );
  OAI211_X1 U21071 ( .C1(n18016), .C2(n18015), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18137), .ZN(n18017) );
  OAI211_X1 U21072 ( .C1(n18019), .C2(n18037), .A(n18018), .B(n18017), .ZN(
        P3_U2851) );
  NOR2_X1 U21073 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18037), .ZN(
        n18020) );
  AOI22_X1 U21074 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18020), .B1(
        n9577), .B2(P3_REIP_REG_10__SCAN_IN), .ZN(n18025) );
  OAI211_X1 U21075 ( .C1(n18022), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18027), .B(n18021), .ZN(n18023) );
  NAND3_X1 U21076 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18137), .A3(
        n18023), .ZN(n18024) );
  OAI211_X1 U21077 ( .C1(n18026), .C2(n18051), .A(n18025), .B(n18024), .ZN(
        P3_U2852) );
  OAI21_X1 U21078 ( .B1(n18029), .B2(n18028), .A(n18027), .ZN(n18030) );
  OAI21_X1 U21079 ( .B1(n18031), .B2(n18030), .A(n18137), .ZN(n18035) );
  AOI22_X1 U21080 ( .A1(n18044), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18033), 
        .B2(n18032), .ZN(n18034) );
  OAI221_X1 U21081 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18037), .C1(
        n18036), .C2(n18035), .A(n18034), .ZN(P3_U2853) );
  INV_X1 U21082 ( .A(n18038), .ZN(n18040) );
  OAI222_X1 U21083 ( .A1(n18042), .A2(n18041), .B1(n18040), .B2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C1(n18107), .C2(n18039), .ZN(
        n18043) );
  AOI22_X1 U21084 ( .A1(n18044), .A2(P3_REIP_REG_8__SCAN_IN), .B1(n18129), 
        .B2(n18043), .ZN(n18050) );
  OAI21_X1 U21085 ( .B1(n18099), .B2(n18045), .A(n18100), .ZN(n18046) );
  AOI21_X1 U21086 ( .B1(n18609), .B2(n18047), .A(n18046), .ZN(n18062) );
  OAI211_X1 U21087 ( .C1(n9586), .C2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n18062), .ZN(n18056) );
  OAI221_X1 U21088 ( .B1(n18114), .B2(n18124), .C1(n18114), .C2(n18056), .A(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18049) );
  OAI211_X1 U21089 ( .C1(n18052), .C2(n18051), .A(n18050), .B(n18049), .ZN(
        P3_U2854) );
  AOI21_X1 U21090 ( .B1(n18114), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18053), .ZN(n18060) );
  AOI221_X1 U21091 ( .B1(n18055), .B2(n18054), .C1(n18063), .C2(n18054), .A(
        n18116), .ZN(n18057) );
  AOI22_X1 U21092 ( .A1(n18132), .A2(n18058), .B1(n18057), .B2(n18056), .ZN(
        n18059) );
  OAI211_X1 U21093 ( .C1(n18127), .C2(n18061), .A(n18060), .B(n18059), .ZN(
        P3_U2855) );
  AOI21_X1 U21094 ( .B1(n18129), .B2(n18062), .A(n9577), .ZN(n18073) );
  AOI22_X1 U21095 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18073), .B1(
        n9577), .B2(P3_REIP_REG_6__SCAN_IN), .ZN(n18067) );
  NOR3_X1 U21096 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18116), .A3(
        n18063), .ZN(n18064) );
  AOI21_X1 U21097 ( .B1(n18065), .B2(n18132), .A(n18064), .ZN(n18066) );
  OAI211_X1 U21098 ( .C1(n18127), .C2(n18068), .A(n18067), .B(n18066), .ZN(
        P3_U2856) );
  NAND3_X1 U21099 ( .A1(n18129), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18090), .ZN(n18082) );
  NOR2_X1 U21100 ( .A1(n18081), .A2(n18082), .ZN(n18072) );
  OAI21_X1 U21101 ( .B1(n18127), .B2(n18070), .A(n18069), .ZN(n18071) );
  AOI221_X1 U21102 ( .B1(n18073), .B2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(
        n18072), .C2(n9820), .A(n18071), .ZN(n18074) );
  OAI21_X1 U21103 ( .B1(n18076), .B2(n18075), .A(n18074), .ZN(P3_U2857) );
  NOR2_X1 U21104 ( .A1(n18137), .A2(n18691), .ZN(n18085) );
  AOI22_X1 U21105 ( .A1(n18609), .A2(n18079), .B1(n18078), .B2(n18077), .ZN(
        n18080) );
  NAND3_X1 U21106 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18080), .A3(
        n18100), .ZN(n18089) );
  AOI21_X1 U21107 ( .B1(n18124), .B2(n18089), .A(n18114), .ZN(n18083) );
  AOI22_X1 U21108 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18083), .B1(
        n18082), .B2(n18081), .ZN(n18084) );
  AOI211_X1 U21109 ( .C1(n18086), .C2(n18132), .A(n18085), .B(n18084), .ZN(
        n18087) );
  OAI21_X1 U21110 ( .B1(n18127), .B2(n18088), .A(n18087), .ZN(P3_U2858) );
  OAI211_X1 U21111 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18090), .A(
        n18129), .B(n18089), .ZN(n18091) );
  OAI211_X1 U21112 ( .C1(n18120), .C2(n18093), .A(n18092), .B(n18091), .ZN(
        n18094) );
  AOI21_X1 U21113 ( .B1(n18132), .B2(n18095), .A(n18094), .ZN(n18096) );
  OAI21_X1 U21114 ( .B1(n18127), .B2(n18097), .A(n18096), .ZN(P3_U2859) );
  NOR2_X1 U21115 ( .A1(n18626), .A2(n18098), .ZN(n18110) );
  AOI21_X1 U21116 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18100), .A(
        n18099), .ZN(n18102) );
  NOR2_X1 U21117 ( .A1(n18771), .A2(n18787), .ZN(n18101) );
  OAI221_X1 U21118 ( .B1(n18102), .B2(n18609), .C1(n18102), .C2(n18101), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18106) );
  NAND3_X1 U21119 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18104), .A3(
        n18103), .ZN(n18105) );
  OAI211_X1 U21120 ( .C1(n18108), .C2(n18107), .A(n18106), .B(n18105), .ZN(
        n18109) );
  AOI211_X1 U21121 ( .C1(n18112), .C2(n18111), .A(n18110), .B(n18109), .ZN(
        n18117) );
  AOI21_X1 U21122 ( .B1(n18114), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n18113), .ZN(n18115) );
  OAI21_X1 U21123 ( .B1(n18117), .B2(n18116), .A(n18115), .ZN(P3_U2860) );
  INV_X1 U21124 ( .A(n18118), .ZN(n18128) );
  NOR2_X1 U21125 ( .A1(n18137), .A2(n20843), .ZN(n18122) );
  NAND3_X1 U21126 ( .A1(n18129), .A2(n18119), .A3(n18787), .ZN(n18135) );
  AOI21_X1 U21127 ( .B1(n18120), .B2(n18135), .A(n18771), .ZN(n18121) );
  AOI211_X1 U21128 ( .C1(n18123), .C2(n18132), .A(n18122), .B(n18121), .ZN(
        n18126) );
  OAI211_X1 U21129 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18608), .A(
        n18124), .B(n18771), .ZN(n18125) );
  OAI211_X1 U21130 ( .C1(n18128), .C2(n18127), .A(n18126), .B(n18125), .ZN(
        P3_U2861) );
  INV_X1 U21131 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18796) );
  AOI211_X1 U21132 ( .C1(n18630), .C2(n18129), .A(n9577), .B(n18787), .ZN(
        n18130) );
  AOI221_X1 U21133 ( .B1(n18134), .B2(n18133), .C1(n18132), .C2(n18131), .A(
        n18130), .ZN(n18136) );
  OAI211_X1 U21134 ( .C1(n18796), .C2(n18137), .A(n18136), .B(n18135), .ZN(
        P3_U2862) );
  AOI21_X1 U21135 ( .B1(n18140), .B2(n18139), .A(n18138), .ZN(n18654) );
  OAI21_X1 U21136 ( .B1(n18654), .B2(n18199), .A(n18145), .ZN(n18141) );
  OAI221_X1 U21137 ( .B1(n18407), .B2(n18811), .C1(n18407), .C2(n18145), .A(
        n18141), .ZN(P3_U2863) );
  NAND2_X1 U21138 ( .A1(n18640), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18433) );
  INV_X1 U21139 ( .A(n18433), .ZN(n18359) );
  NAND2_X1 U21140 ( .A1(n18643), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18291) );
  INV_X1 U21141 ( .A(n18291), .ZN(n18337) );
  NOR2_X1 U21142 ( .A1(n18359), .A2(n18337), .ZN(n18143) );
  OAI22_X1 U21143 ( .A1(n18144), .A2(n18643), .B1(n18143), .B2(n18142), .ZN(
        P3_U2866) );
  INV_X1 U21144 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18644) );
  NOR2_X1 U21145 ( .A1(n18644), .A2(n18145), .ZN(P3_U2867) );
  NOR2_X1 U21146 ( .A1(n18643), .A2(n18384), .ZN(n18540) );
  NAND2_X1 U21147 ( .A1(n18540), .A2(n18407), .ZN(n18535) );
  INV_X1 U21148 ( .A(n18535), .ZN(n18527) );
  NAND2_X1 U21149 ( .A1(n18635), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18386) );
  NAND2_X1 U21150 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18477) );
  NOR2_X1 U21151 ( .A1(n18527), .A2(n9560), .ZN(n18504) );
  NOR2_X1 U21152 ( .A1(n18407), .A2(n18759), .ZN(n18146) );
  NOR2_X1 U21153 ( .A1(n18635), .A2(n18407), .ZN(n18338) );
  INV_X1 U21154 ( .A(n18338), .ZN(n18634) );
  NOR2_X2 U21155 ( .A1(n18634), .A2(n18477), .ZN(n18581) );
  NOR2_X1 U21156 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18360) );
  INV_X1 U21157 ( .A(n18360), .ZN(n18636) );
  NAND2_X1 U21158 ( .A1(n18640), .A2(n18643), .ZN(n18219) );
  NOR2_X2 U21159 ( .A1(n18636), .A2(n18219), .ZN(n18265) );
  NOR2_X1 U21160 ( .A1(n18581), .A2(n18265), .ZN(n18220) );
  OAI22_X1 U21161 ( .A1(n18505), .A2(n18504), .B1(n18146), .B2(n18220), .ZN(
        n18147) );
  AND2_X1 U21162 ( .A1(n18147), .A2(n18508), .ZN(n18198) );
  INV_X1 U21163 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18148) );
  NOR2_X1 U21164 ( .A1(n18148), .A2(n18313), .ZN(n18503) );
  NOR2_X2 U21165 ( .A1(n18312), .A2(n18149), .ZN(n18537) );
  NAND2_X1 U21166 ( .A1(n18805), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18536) );
  INV_X1 U21167 ( .A(n18536), .ZN(n18502) );
  NOR2_X1 U21168 ( .A1(n18502), .A2(n18220), .ZN(n18192) );
  AOI22_X1 U21169 ( .A1(n18503), .A2(n9560), .B1(n18537), .B2(n18192), .ZN(
        n18153) );
  OR3_X1 U21170 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18150), .A3(n18759), 
        .ZN(n18194) );
  NOR2_X2 U21171 ( .A1(n18151), .A2(n18194), .ZN(n18543) );
  NAND2_X1 U21172 ( .A1(n18542), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18511) );
  INV_X1 U21173 ( .A(n18511), .ZN(n18538) );
  AOI22_X1 U21174 ( .A1(n18543), .A2(n18265), .B1(n18538), .B2(n18527), .ZN(
        n18152) );
  OAI211_X1 U21175 ( .C1(n18198), .C2(n18154), .A(n18153), .B(n18152), .ZN(
        P3_U2868) );
  INV_X1 U21176 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18155) );
  NOR2_X1 U21177 ( .A1(n18155), .A2(n18313), .ZN(n18548) );
  NOR2_X2 U21178 ( .A1(n18312), .A2(n18156), .ZN(n18547) );
  AOI22_X1 U21179 ( .A1(n18548), .A2(n9560), .B1(n18547), .B2(n18192), .ZN(
        n18159) );
  NOR2_X2 U21180 ( .A1(n18157), .A2(n18194), .ZN(n18549) );
  NAND2_X1 U21181 ( .A1(n18542), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18553) );
  INV_X1 U21182 ( .A(n18553), .ZN(n18483) );
  AOI22_X1 U21183 ( .A1(n18549), .A2(n18265), .B1(n18483), .B2(n18527), .ZN(
        n18158) );
  OAI211_X1 U21184 ( .C1(n18198), .C2(n18160), .A(n18159), .B(n18158), .ZN(
        P3_U2869) );
  NOR2_X1 U21185 ( .A1(n18161), .A2(n18313), .ZN(n18414) );
  NOR2_X2 U21186 ( .A1(n18312), .A2(n18162), .ZN(n18555) );
  AOI22_X1 U21187 ( .A1(n18414), .A2(n9560), .B1(n18555), .B2(n18192), .ZN(
        n18165) );
  NOR2_X2 U21188 ( .A1(n18163), .A2(n18194), .ZN(n18556) );
  NAND2_X1 U21189 ( .A1(n18542), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18417) );
  INV_X1 U21190 ( .A(n18417), .ZN(n18554) );
  AOI22_X1 U21191 ( .A1(n18556), .A2(n18265), .B1(n18554), .B2(n18527), .ZN(
        n18164) );
  OAI211_X1 U21192 ( .C1(n18198), .C2(n18166), .A(n18165), .B(n18164), .ZN(
        P3_U2870) );
  NOR2_X2 U21193 ( .A1(n18312), .A2(n18167), .ZN(n18560) );
  INV_X1 U21194 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n18168) );
  NOR2_X2 U21195 ( .A1(n18168), .A2(n18313), .ZN(n18562) );
  AOI22_X1 U21196 ( .A1(n18560), .A2(n18192), .B1(n18562), .B2(n9560), .ZN(
        n18171) );
  AND2_X1 U21197 ( .A1(n18542), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18561) );
  NOR2_X1 U21198 ( .A1(n18194), .A2(n18169), .ZN(n18229) );
  AOI22_X1 U21199 ( .A1(n18561), .A2(n18527), .B1(n18229), .B2(n18265), .ZN(
        n18170) );
  OAI211_X1 U21200 ( .C1(n18198), .C2(n18172), .A(n18171), .B(n18170), .ZN(
        P3_U2871) );
  NOR2_X2 U21201 ( .A1(n18173), .A2(n18312), .ZN(n18566) );
  NOR2_X2 U21202 ( .A1(n18174), .A2(n18313), .ZN(n18568) );
  AOI22_X1 U21203 ( .A1(n18566), .A2(n18192), .B1(n18568), .B2(n9560), .ZN(
        n18177) );
  INV_X1 U21204 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n20844) );
  NOR2_X2 U21205 ( .A1(n20844), .A2(n18313), .ZN(n18567) );
  NOR2_X1 U21206 ( .A1(n18194), .A2(n18175), .ZN(n18208) );
  AOI22_X1 U21207 ( .A1(n18567), .A2(n18527), .B1(n18208), .B2(n18265), .ZN(
        n18176) );
  OAI211_X1 U21208 ( .C1(n18198), .C2(n18178), .A(n18177), .B(n18176), .ZN(
        P3_U2872) );
  NOR2_X1 U21209 ( .A1(n18179), .A2(n18313), .ZN(n18521) );
  NOR2_X2 U21210 ( .A1(n18180), .A2(n18312), .ZN(n18573) );
  AOI22_X1 U21211 ( .A1(n18521), .A2(n9560), .B1(n18573), .B2(n18192), .ZN(
        n18183) );
  NOR2_X2 U21212 ( .A1(n18181), .A2(n18194), .ZN(n18574) );
  NAND2_X1 U21213 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18542), .ZN(n18524) );
  INV_X1 U21214 ( .A(n18524), .ZN(n18572) );
  AOI22_X1 U21215 ( .A1(n18574), .A2(n18265), .B1(n18572), .B2(n18527), .ZN(
        n18182) );
  OAI211_X1 U21216 ( .C1(n18198), .C2(n18184), .A(n18183), .B(n18182), .ZN(
        P3_U2873) );
  INV_X1 U21217 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18185) );
  NOR2_X1 U21218 ( .A1(n18185), .A2(n18313), .ZN(n18525) );
  NOR2_X2 U21219 ( .A1(n18186), .A2(n18312), .ZN(n18578) );
  AOI22_X1 U21220 ( .A1(n18525), .A2(n9560), .B1(n18578), .B2(n18192), .ZN(
        n18189) );
  NOR2_X2 U21221 ( .A1(n18187), .A2(n18194), .ZN(n18582) );
  NAND2_X1 U21222 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18542), .ZN(n18530) );
  INV_X1 U21223 ( .A(n18530), .ZN(n18580) );
  AOI22_X1 U21224 ( .A1(n18582), .A2(n18265), .B1(n18580), .B2(n18527), .ZN(
        n18188) );
  OAI211_X1 U21225 ( .C1(n18198), .C2(n18190), .A(n18189), .B(n18188), .ZN(
        P3_U2874) );
  NOR2_X2 U21226 ( .A1(n20856), .A2(n18313), .ZN(n18589) );
  NOR2_X2 U21227 ( .A1(n18191), .A2(n18312), .ZN(n18588) );
  AOI22_X1 U21228 ( .A1(n18589), .A2(n9560), .B1(n18588), .B2(n18192), .ZN(
        n18196) );
  NOR2_X2 U21229 ( .A1(n19218), .A2(n18313), .ZN(n18591) );
  NOR2_X1 U21230 ( .A1(n18194), .A2(n18193), .ZN(n18241) );
  AOI22_X1 U21231 ( .A1(n18591), .A2(n18527), .B1(n18241), .B2(n18265), .ZN(
        n18195) );
  OAI211_X1 U21232 ( .C1(n18198), .C2(n18197), .A(n18196), .B(n18195), .ZN(
        P3_U2875) );
  INV_X1 U21233 ( .A(n18503), .ZN(n18546) );
  NAND2_X1 U21234 ( .A1(n18635), .A2(n18536), .ZN(n18476) );
  NOR2_X1 U21235 ( .A1(n18219), .A2(n18476), .ZN(n18215) );
  AOI22_X1 U21236 ( .A1(n18538), .A2(n18581), .B1(n18537), .B2(n18215), .ZN(
        n18201) );
  INV_X1 U21237 ( .A(n18219), .ZN(n18247) );
  NOR2_X1 U21238 ( .A1(n18312), .A2(n18199), .ZN(n18539) );
  AND2_X1 U21239 ( .A1(n18635), .A2(n18539), .ZN(n18478) );
  AOI22_X1 U21240 ( .A1(n18542), .A2(n18540), .B1(n18247), .B2(n18478), .ZN(
        n18216) );
  NOR2_X2 U21241 ( .A1(n18386), .A2(n18219), .ZN(n18286) );
  AOI22_X1 U21242 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18216), .B1(
        n18543), .B2(n18286), .ZN(n18200) );
  OAI211_X1 U21243 ( .C1(n18546), .C2(n18535), .A(n18201), .B(n18200), .ZN(
        P3_U2876) );
  INV_X1 U21244 ( .A(n18581), .ZN(n18595) );
  AOI22_X1 U21245 ( .A1(n18548), .A2(n18527), .B1(n18547), .B2(n18215), .ZN(
        n18203) );
  AOI22_X1 U21246 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18216), .B1(
        n18549), .B2(n18286), .ZN(n18202) );
  OAI211_X1 U21247 ( .C1(n18553), .C2(n18595), .A(n18203), .B(n18202), .ZN(
        P3_U2877) );
  AOI22_X1 U21248 ( .A1(n18414), .A2(n18527), .B1(n18555), .B2(n18215), .ZN(
        n18205) );
  AOI22_X1 U21249 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18216), .B1(
        n18556), .B2(n18286), .ZN(n18204) );
  OAI211_X1 U21250 ( .C1(n18417), .C2(n18595), .A(n18205), .B(n18204), .ZN(
        P3_U2878) );
  INV_X1 U21251 ( .A(n18286), .ZN(n18274) );
  AOI22_X1 U21252 ( .A1(n18561), .A2(n18581), .B1(n18560), .B2(n18215), .ZN(
        n18207) );
  AOI22_X1 U21253 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18216), .B1(
        n18562), .B2(n18527), .ZN(n18206) );
  OAI211_X1 U21254 ( .C1(n18565), .C2(n18274), .A(n18207), .B(n18206), .ZN(
        P3_U2879) );
  AOI22_X1 U21255 ( .A1(n18566), .A2(n18215), .B1(n18568), .B2(n18527), .ZN(
        n18210) );
  AOI22_X1 U21256 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18216), .B1(
        n18567), .B2(n18581), .ZN(n18209) );
  OAI211_X1 U21257 ( .C1(n18571), .C2(n18274), .A(n18210), .B(n18209), .ZN(
        P3_U2880) );
  INV_X1 U21258 ( .A(n18521), .ZN(n18577) );
  AOI22_X1 U21259 ( .A1(n18573), .A2(n18215), .B1(n18572), .B2(n18581), .ZN(
        n18212) );
  AOI22_X1 U21260 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18216), .B1(
        n18574), .B2(n18286), .ZN(n18211) );
  OAI211_X1 U21261 ( .C1(n18577), .C2(n18535), .A(n18212), .B(n18211), .ZN(
        P3_U2881) );
  INV_X1 U21262 ( .A(n18525), .ZN(n18585) );
  AOI22_X1 U21263 ( .A1(n18580), .A2(n18581), .B1(n18578), .B2(n18215), .ZN(
        n18214) );
  AOI22_X1 U21264 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18216), .B1(
        n18582), .B2(n18286), .ZN(n18213) );
  OAI211_X1 U21265 ( .C1(n18585), .C2(n18535), .A(n18214), .B(n18213), .ZN(
        P3_U2882) );
  INV_X1 U21266 ( .A(n18241), .ZN(n18596) );
  AOI22_X1 U21267 ( .A1(n18589), .A2(n18527), .B1(n18588), .B2(n18215), .ZN(
        n18218) );
  AOI22_X1 U21268 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18216), .B1(
        n18591), .B2(n18581), .ZN(n18217) );
  OAI211_X1 U21269 ( .C1(n18596), .C2(n18274), .A(n18218), .B(n18217), .ZN(
        P3_U2883) );
  NOR2_X1 U21270 ( .A1(n18635), .A2(n18219), .ZN(n18290) );
  NAND2_X1 U21271 ( .A1(n18290), .A2(n18407), .ZN(n18306) );
  INV_X1 U21272 ( .A(n18306), .ZN(n18308) );
  NOR2_X1 U21273 ( .A1(n18286), .A2(n18308), .ZN(n18268) );
  OAI21_X1 U21274 ( .B1(n18505), .B2(n18220), .A(n18268), .ZN(n18221) );
  OAI211_X1 U21275 ( .C1(n18759), .C2(n18308), .A(n18221), .B(n18508), .ZN(
        n18237) );
  INV_X1 U21276 ( .A(n18237), .ZN(n18245) );
  NOR2_X1 U21277 ( .A1(n18502), .A2(n18268), .ZN(n18240) );
  AOI22_X1 U21278 ( .A1(n18503), .A2(n18581), .B1(n18537), .B2(n18240), .ZN(
        n18223) );
  AOI22_X1 U21279 ( .A1(n18543), .A2(n18308), .B1(n18538), .B2(n18265), .ZN(
        n18222) );
  OAI211_X1 U21280 ( .C1(n18245), .C2(n20773), .A(n18223), .B(n18222), .ZN(
        P3_U2884) );
  INV_X1 U21281 ( .A(n18265), .ZN(n18262) );
  AOI22_X1 U21282 ( .A1(n18548), .A2(n18581), .B1(n18547), .B2(n18240), .ZN(
        n18225) );
  AOI22_X1 U21283 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18237), .B1(
        n18549), .B2(n18308), .ZN(n18224) );
  OAI211_X1 U21284 ( .C1(n18553), .C2(n18262), .A(n18225), .B(n18224), .ZN(
        P3_U2885) );
  AOI22_X1 U21285 ( .A1(n18414), .A2(n18581), .B1(n18555), .B2(n18240), .ZN(
        n18227) );
  AOI22_X1 U21286 ( .A1(n18556), .A2(n18308), .B1(n18554), .B2(n18265), .ZN(
        n18226) );
  OAI211_X1 U21287 ( .C1(n18245), .C2(n18228), .A(n18227), .B(n18226), .ZN(
        P3_U2886) );
  AOI22_X1 U21288 ( .A1(n18561), .A2(n18265), .B1(n18560), .B2(n18240), .ZN(
        n18231) );
  AOI22_X1 U21289 ( .A1(n18229), .A2(n18308), .B1(n18562), .B2(n18581), .ZN(
        n18230) );
  OAI211_X1 U21290 ( .C1(n18245), .C2(n18232), .A(n18231), .B(n18230), .ZN(
        P3_U2887) );
  AOI22_X1 U21291 ( .A1(n18566), .A2(n18240), .B1(n18568), .B2(n18581), .ZN(
        n18234) );
  AOI22_X1 U21292 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18237), .B1(
        n18567), .B2(n18265), .ZN(n18233) );
  OAI211_X1 U21293 ( .C1(n18571), .C2(n18306), .A(n18234), .B(n18233), .ZN(
        P3_U2888) );
  AOI22_X1 U21294 ( .A1(n18521), .A2(n18581), .B1(n18573), .B2(n18240), .ZN(
        n18236) );
  AOI22_X1 U21295 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18237), .B1(
        n18574), .B2(n18308), .ZN(n18235) );
  OAI211_X1 U21296 ( .C1(n18524), .C2(n18262), .A(n18236), .B(n18235), .ZN(
        P3_U2889) );
  AOI22_X1 U21297 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18237), .B1(
        n18578), .B2(n18240), .ZN(n18239) );
  AOI22_X1 U21298 ( .A1(n18582), .A2(n18308), .B1(n18580), .B2(n18265), .ZN(
        n18238) );
  OAI211_X1 U21299 ( .C1(n18585), .C2(n18595), .A(n18239), .B(n18238), .ZN(
        P3_U2890) );
  AOI22_X1 U21300 ( .A1(n18591), .A2(n18265), .B1(n18588), .B2(n18240), .ZN(
        n18243) );
  AOI22_X1 U21301 ( .A1(n18241), .A2(n18308), .B1(n18589), .B2(n18581), .ZN(
        n18242) );
  OAI211_X1 U21302 ( .C1(n18245), .C2(n18244), .A(n18243), .B(n18242), .ZN(
        P3_U2891) );
  AND2_X1 U21303 ( .A1(n18536), .A2(n18290), .ZN(n18263) );
  AOI22_X1 U21304 ( .A1(n18503), .A2(n18265), .B1(n18537), .B2(n18263), .ZN(
        n18249) );
  OAI211_X1 U21305 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18246), .A(
        n18247), .B(n18539), .ZN(n18264) );
  NAND2_X1 U21306 ( .A1(n18338), .A2(n18247), .ZN(n18328) );
  INV_X1 U21307 ( .A(n18328), .ZN(n18332) );
  AOI22_X1 U21308 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18264), .B1(
        n18543), .B2(n18332), .ZN(n18248) );
  OAI211_X1 U21309 ( .C1(n18511), .C2(n18274), .A(n18249), .B(n18248), .ZN(
        P3_U2892) );
  INV_X1 U21310 ( .A(n18548), .ZN(n18486) );
  AOI22_X1 U21311 ( .A1(n18483), .A2(n18286), .B1(n18547), .B2(n18263), .ZN(
        n18251) );
  AOI22_X1 U21312 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18264), .B1(
        n18549), .B2(n18332), .ZN(n18250) );
  OAI211_X1 U21313 ( .C1(n18486), .C2(n18262), .A(n18251), .B(n18250), .ZN(
        P3_U2893) );
  INV_X1 U21314 ( .A(n18414), .ZN(n18559) );
  AOI22_X1 U21315 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18264), .B1(
        n18555), .B2(n18263), .ZN(n18253) );
  AOI22_X1 U21316 ( .A1(n18556), .A2(n18332), .B1(n18554), .B2(n18286), .ZN(
        n18252) );
  OAI211_X1 U21317 ( .C1(n18559), .C2(n18262), .A(n18253), .B(n18252), .ZN(
        P3_U2894) );
  AOI22_X1 U21318 ( .A1(n18560), .A2(n18263), .B1(n18562), .B2(n18265), .ZN(
        n18255) );
  AOI22_X1 U21319 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18264), .B1(
        n18561), .B2(n18286), .ZN(n18254) );
  OAI211_X1 U21320 ( .C1(n18565), .C2(n18328), .A(n18255), .B(n18254), .ZN(
        P3_U2895) );
  AOI22_X1 U21321 ( .A1(n18566), .A2(n18263), .B1(n18568), .B2(n18265), .ZN(
        n18257) );
  AOI22_X1 U21322 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18264), .B1(
        n18567), .B2(n18286), .ZN(n18256) );
  OAI211_X1 U21323 ( .C1(n18571), .C2(n18328), .A(n18257), .B(n18256), .ZN(
        P3_U2896) );
  AOI22_X1 U21324 ( .A1(n18521), .A2(n18265), .B1(n18573), .B2(n18263), .ZN(
        n18259) );
  AOI22_X1 U21325 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18264), .B1(
        n18574), .B2(n18332), .ZN(n18258) );
  OAI211_X1 U21326 ( .C1(n18524), .C2(n18274), .A(n18259), .B(n18258), .ZN(
        P3_U2897) );
  AOI22_X1 U21327 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18264), .B1(
        n18578), .B2(n18263), .ZN(n18261) );
  AOI22_X1 U21328 ( .A1(n18582), .A2(n18332), .B1(n18580), .B2(n18286), .ZN(
        n18260) );
  OAI211_X1 U21329 ( .C1(n18585), .C2(n18262), .A(n18261), .B(n18260), .ZN(
        P3_U2898) );
  AOI22_X1 U21330 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18264), .B1(
        n18588), .B2(n18263), .ZN(n18267) );
  AOI22_X1 U21331 ( .A1(n18591), .A2(n18286), .B1(n18589), .B2(n18265), .ZN(
        n18266) );
  OAI211_X1 U21332 ( .C1(n18596), .C2(n18328), .A(n18267), .B(n18266), .ZN(
        P3_U2899) );
  NAND2_X1 U21333 ( .A1(n18360), .A2(n18337), .ZN(n18353) );
  INV_X1 U21334 ( .A(n18353), .ZN(n18356) );
  NOR2_X1 U21335 ( .A1(n18332), .A2(n18356), .ZN(n18314) );
  NOR2_X1 U21336 ( .A1(n18502), .A2(n18314), .ZN(n18285) );
  AOI22_X1 U21337 ( .A1(n18538), .A2(n18308), .B1(n18537), .B2(n18285), .ZN(
        n18271) );
  OAI22_X1 U21338 ( .A1(n18268), .A2(n18313), .B1(n18314), .B2(n18312), .ZN(
        n18269) );
  OAI21_X1 U21339 ( .B1(n18356), .B2(n18759), .A(n18269), .ZN(n18287) );
  AOI22_X1 U21340 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18287), .B1(
        n18543), .B2(n18356), .ZN(n18270) );
  OAI211_X1 U21341 ( .C1(n18546), .C2(n18274), .A(n18271), .B(n18270), .ZN(
        P3_U2900) );
  AOI22_X1 U21342 ( .A1(n18483), .A2(n18308), .B1(n18547), .B2(n18285), .ZN(
        n18273) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18287), .B1(
        n18549), .B2(n18356), .ZN(n18272) );
  OAI211_X1 U21344 ( .C1(n18486), .C2(n18274), .A(n18273), .B(n18272), .ZN(
        P3_U2901) );
  AOI22_X1 U21345 ( .A1(n18414), .A2(n18286), .B1(n18555), .B2(n18285), .ZN(
        n18276) );
  AOI22_X1 U21346 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18287), .B1(
        n18556), .B2(n18356), .ZN(n18275) );
  OAI211_X1 U21347 ( .C1(n18417), .C2(n18306), .A(n18276), .B(n18275), .ZN(
        P3_U2902) );
  AOI22_X1 U21348 ( .A1(n18561), .A2(n18308), .B1(n18560), .B2(n18285), .ZN(
        n18278) );
  AOI22_X1 U21349 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18287), .B1(
        n18562), .B2(n18286), .ZN(n18277) );
  OAI211_X1 U21350 ( .C1(n18565), .C2(n18353), .A(n18278), .B(n18277), .ZN(
        P3_U2903) );
  AOI22_X1 U21351 ( .A1(n18567), .A2(n18308), .B1(n18566), .B2(n18285), .ZN(
        n18280) );
  AOI22_X1 U21352 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18287), .B1(
        n18568), .B2(n18286), .ZN(n18279) );
  OAI211_X1 U21353 ( .C1(n18571), .C2(n18353), .A(n18280), .B(n18279), .ZN(
        P3_U2904) );
  AOI22_X1 U21354 ( .A1(n18521), .A2(n18286), .B1(n18573), .B2(n18285), .ZN(
        n18282) );
  AOI22_X1 U21355 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18287), .B1(
        n18574), .B2(n18356), .ZN(n18281) );
  OAI211_X1 U21356 ( .C1(n18524), .C2(n18306), .A(n18282), .B(n18281), .ZN(
        P3_U2905) );
  AOI22_X1 U21357 ( .A1(n18525), .A2(n18286), .B1(n18578), .B2(n18285), .ZN(
        n18284) );
  AOI22_X1 U21358 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18287), .B1(
        n18582), .B2(n18356), .ZN(n18283) );
  OAI211_X1 U21359 ( .C1(n18530), .C2(n18306), .A(n18284), .B(n18283), .ZN(
        P3_U2906) );
  AOI22_X1 U21360 ( .A1(n18589), .A2(n18286), .B1(n18588), .B2(n18285), .ZN(
        n18289) );
  AOI22_X1 U21361 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18287), .B1(
        n18591), .B2(n18308), .ZN(n18288) );
  OAI211_X1 U21362 ( .C1(n18596), .C2(n18353), .A(n18289), .B(n18288), .ZN(
        P3_U2907) );
  NOR2_X1 U21363 ( .A1(n18291), .A2(n18476), .ZN(n18307) );
  AOI22_X1 U21364 ( .A1(n18538), .A2(n18332), .B1(n18537), .B2(n18307), .ZN(
        n18293) );
  AOI22_X1 U21365 ( .A1(n18542), .A2(n18290), .B1(n18337), .B2(n18478), .ZN(
        n18309) );
  NOR2_X2 U21366 ( .A1(n18291), .A2(n18386), .ZN(n18380) );
  AOI22_X1 U21367 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18309), .B1(
        n18543), .B2(n18380), .ZN(n18292) );
  OAI211_X1 U21368 ( .C1(n18546), .C2(n18306), .A(n18293), .B(n18292), .ZN(
        P3_U2908) );
  AOI22_X1 U21369 ( .A1(n18483), .A2(n18332), .B1(n18547), .B2(n18307), .ZN(
        n18295) );
  AOI22_X1 U21370 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18309), .B1(
        n18549), .B2(n18380), .ZN(n18294) );
  OAI211_X1 U21371 ( .C1(n18486), .C2(n18306), .A(n18295), .B(n18294), .ZN(
        P3_U2909) );
  AOI22_X1 U21372 ( .A1(n18414), .A2(n18308), .B1(n18555), .B2(n18307), .ZN(
        n18297) );
  AOI22_X1 U21373 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18309), .B1(
        n18556), .B2(n18380), .ZN(n18296) );
  OAI211_X1 U21374 ( .C1(n18417), .C2(n18328), .A(n18297), .B(n18296), .ZN(
        P3_U2910) );
  INV_X1 U21375 ( .A(n18380), .ZN(n18378) );
  AOI22_X1 U21376 ( .A1(n18561), .A2(n18332), .B1(n18560), .B2(n18307), .ZN(
        n18299) );
  AOI22_X1 U21377 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18309), .B1(
        n18562), .B2(n18308), .ZN(n18298) );
  OAI211_X1 U21378 ( .C1(n18565), .C2(n18378), .A(n18299), .B(n18298), .ZN(
        P3_U2911) );
  AOI22_X1 U21379 ( .A1(n18567), .A2(n18332), .B1(n18566), .B2(n18307), .ZN(
        n18301) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18309), .B1(
        n18568), .B2(n18308), .ZN(n18300) );
  OAI211_X1 U21381 ( .C1(n18571), .C2(n18378), .A(n18301), .B(n18300), .ZN(
        P3_U2912) );
  AOI22_X1 U21382 ( .A1(n18573), .A2(n18307), .B1(n18572), .B2(n18332), .ZN(
        n18303) );
  AOI22_X1 U21383 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18309), .B1(
        n18574), .B2(n18380), .ZN(n18302) );
  OAI211_X1 U21384 ( .C1(n18577), .C2(n18306), .A(n18303), .B(n18302), .ZN(
        P3_U2913) );
  AOI22_X1 U21385 ( .A1(n18580), .A2(n18332), .B1(n18578), .B2(n18307), .ZN(
        n18305) );
  AOI22_X1 U21386 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18309), .B1(
        n18582), .B2(n18380), .ZN(n18304) );
  OAI211_X1 U21387 ( .C1(n18585), .C2(n18306), .A(n18305), .B(n18304), .ZN(
        P3_U2914) );
  AOI22_X1 U21388 ( .A1(n18591), .A2(n18332), .B1(n18588), .B2(n18307), .ZN(
        n18311) );
  AOI22_X1 U21389 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18309), .B1(
        n18589), .B2(n18308), .ZN(n18310) );
  OAI211_X1 U21390 ( .C1(n18596), .C2(n18378), .A(n18311), .B(n18310), .ZN(
        P3_U2915) );
  NOR3_X1 U21391 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n18384), .ZN(n18391) );
  INV_X1 U21392 ( .A(n18391), .ZN(n18375) );
  INV_X1 U21393 ( .A(n18375), .ZN(n18398) );
  NOR2_X1 U21394 ( .A1(n18380), .A2(n18398), .ZN(n18361) );
  NOR2_X1 U21395 ( .A1(n18502), .A2(n18361), .ZN(n18331) );
  AOI22_X1 U21396 ( .A1(n18503), .A2(n18332), .B1(n18537), .B2(n18331), .ZN(
        n18317) );
  OAI22_X1 U21397 ( .A1(n18314), .A2(n18313), .B1(n18361), .B2(n18312), .ZN(
        n18315) );
  OAI21_X1 U21398 ( .B1(n18398), .B2(n18759), .A(n18315), .ZN(n18333) );
  AOI22_X1 U21399 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18333), .B1(
        n18543), .B2(n18391), .ZN(n18316) );
  OAI211_X1 U21400 ( .C1(n18511), .C2(n18353), .A(n18317), .B(n18316), .ZN(
        P3_U2916) );
  AOI22_X1 U21401 ( .A1(n18548), .A2(n18332), .B1(n18547), .B2(n18331), .ZN(
        n18319) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18333), .B1(
        n18549), .B2(n18391), .ZN(n18318) );
  OAI211_X1 U21403 ( .C1(n18553), .C2(n18353), .A(n18319), .B(n18318), .ZN(
        P3_U2917) );
  AOI22_X1 U21404 ( .A1(n18555), .A2(n18331), .B1(n18554), .B2(n18356), .ZN(
        n18321) );
  AOI22_X1 U21405 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18333), .B1(
        n18556), .B2(n18398), .ZN(n18320) );
  OAI211_X1 U21406 ( .C1(n18559), .C2(n18328), .A(n18321), .B(n18320), .ZN(
        P3_U2918) );
  AOI22_X1 U21407 ( .A1(n18560), .A2(n18331), .B1(n18562), .B2(n18332), .ZN(
        n18323) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18333), .B1(
        n18561), .B2(n18356), .ZN(n18322) );
  OAI211_X1 U21409 ( .C1(n18565), .C2(n18375), .A(n18323), .B(n18322), .ZN(
        P3_U2919) );
  AOI22_X1 U21410 ( .A1(n18566), .A2(n18331), .B1(n18568), .B2(n18332), .ZN(
        n18325) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18333), .B1(
        n18567), .B2(n18356), .ZN(n18324) );
  OAI211_X1 U21412 ( .C1(n18571), .C2(n18375), .A(n18325), .B(n18324), .ZN(
        P3_U2920) );
  AOI22_X1 U21413 ( .A1(n18573), .A2(n18331), .B1(n18572), .B2(n18356), .ZN(
        n18327) );
  AOI22_X1 U21414 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18333), .B1(
        n18574), .B2(n18391), .ZN(n18326) );
  OAI211_X1 U21415 ( .C1(n18577), .C2(n18328), .A(n18327), .B(n18326), .ZN(
        P3_U2921) );
  AOI22_X1 U21416 ( .A1(n18525), .A2(n18332), .B1(n18578), .B2(n18331), .ZN(
        n18330) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18333), .B1(
        n18582), .B2(n18398), .ZN(n18329) );
  OAI211_X1 U21418 ( .C1(n18530), .C2(n18353), .A(n18330), .B(n18329), .ZN(
        P3_U2922) );
  AOI22_X1 U21419 ( .A1(n18591), .A2(n18356), .B1(n18588), .B2(n18331), .ZN(
        n18335) );
  AOI22_X1 U21420 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18333), .B1(
        n18589), .B2(n18332), .ZN(n18334) );
  OAI211_X1 U21421 ( .C1(n18596), .C2(n18375), .A(n18335), .B(n18334), .ZN(
        P3_U2923) );
  AOI22_X1 U21422 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18634), .B1(n18635), 
        .B2(n18505), .ZN(n18336) );
  NAND3_X1 U21423 ( .A1(n18508), .A2(n18337), .A3(n18336), .ZN(n18355) );
  AOI22_X1 U21424 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18355), .B1(
        n18537), .B2(n18354), .ZN(n18340) );
  NAND2_X1 U21425 ( .A1(n18338), .A2(n18337), .ZN(n18424) );
  INV_X1 U21426 ( .A(n18424), .ZN(n18428) );
  AOI22_X1 U21427 ( .A1(n18503), .A2(n18356), .B1(n18543), .B2(n18428), .ZN(
        n18339) );
  OAI211_X1 U21428 ( .C1(n18511), .C2(n18378), .A(n18340), .B(n18339), .ZN(
        P3_U2924) );
  AOI22_X1 U21429 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18355), .B1(
        n18547), .B2(n18354), .ZN(n18342) );
  AOI22_X1 U21430 ( .A1(n18548), .A2(n18356), .B1(n18549), .B2(n18428), .ZN(
        n18341) );
  OAI211_X1 U21431 ( .C1(n18553), .C2(n18378), .A(n18342), .B(n18341), .ZN(
        P3_U2925) );
  AOI22_X1 U21432 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18355), .B1(
        n18555), .B2(n18354), .ZN(n18344) );
  AOI22_X1 U21433 ( .A1(n18556), .A2(n18428), .B1(n18554), .B2(n18380), .ZN(
        n18343) );
  OAI211_X1 U21434 ( .C1(n18559), .C2(n18353), .A(n18344), .B(n18343), .ZN(
        P3_U2926) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18355), .B1(
        n18560), .B2(n18354), .ZN(n18346) );
  AOI22_X1 U21436 ( .A1(n18561), .A2(n18380), .B1(n18562), .B2(n18356), .ZN(
        n18345) );
  OAI211_X1 U21437 ( .C1(n18565), .C2(n18424), .A(n18346), .B(n18345), .ZN(
        P3_U2927) );
  AOI22_X1 U21438 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18355), .B1(
        n18566), .B2(n18354), .ZN(n18348) );
  AOI22_X1 U21439 ( .A1(n18567), .A2(n18380), .B1(n18568), .B2(n18356), .ZN(
        n18347) );
  OAI211_X1 U21440 ( .C1(n18571), .C2(n18424), .A(n18348), .B(n18347), .ZN(
        P3_U2928) );
  AOI22_X1 U21441 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18355), .B1(
        n18573), .B2(n18354), .ZN(n18350) );
  AOI22_X1 U21442 ( .A1(n18521), .A2(n18356), .B1(n18574), .B2(n18428), .ZN(
        n18349) );
  OAI211_X1 U21443 ( .C1(n18524), .C2(n18378), .A(n18350), .B(n18349), .ZN(
        P3_U2929) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18355), .B1(
        n18578), .B2(n18354), .ZN(n18352) );
  AOI22_X1 U21445 ( .A1(n18582), .A2(n18428), .B1(n18580), .B2(n18380), .ZN(
        n18351) );
  OAI211_X1 U21446 ( .C1(n18585), .C2(n18353), .A(n18352), .B(n18351), .ZN(
        P3_U2930) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18355), .B1(
        n18588), .B2(n18354), .ZN(n18358) );
  AOI22_X1 U21448 ( .A1(n18591), .A2(n18380), .B1(n18589), .B2(n18356), .ZN(
        n18357) );
  OAI211_X1 U21449 ( .C1(n18596), .C2(n18424), .A(n18358), .B(n18357), .ZN(
        P3_U2931) );
  NAND2_X1 U21450 ( .A1(n18360), .A2(n18359), .ZN(n18448) );
  INV_X1 U21451 ( .A(n18448), .ZN(n18450) );
  NOR2_X1 U21452 ( .A1(n18428), .A2(n18450), .ZN(n18408) );
  NOR2_X1 U21453 ( .A1(n18502), .A2(n18408), .ZN(n18379) );
  AOI22_X1 U21454 ( .A1(n18503), .A2(n18380), .B1(n18537), .B2(n18379), .ZN(
        n18364) );
  OAI21_X1 U21455 ( .B1(n18361), .B2(n18505), .A(n18408), .ZN(n18362) );
  OAI211_X1 U21456 ( .C1(n18450), .C2(n18759), .A(n18508), .B(n18362), .ZN(
        n18381) );
  AOI22_X1 U21457 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18381), .B1(
        n18543), .B2(n18450), .ZN(n18363) );
  OAI211_X1 U21458 ( .C1(n18511), .C2(n18375), .A(n18364), .B(n18363), .ZN(
        P3_U2932) );
  AOI22_X1 U21459 ( .A1(n18548), .A2(n18380), .B1(n18547), .B2(n18379), .ZN(
        n18366) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18381), .B1(
        n18549), .B2(n18450), .ZN(n18365) );
  OAI211_X1 U21461 ( .C1(n18553), .C2(n18375), .A(n18366), .B(n18365), .ZN(
        P3_U2933) );
  AOI22_X1 U21462 ( .A1(n18555), .A2(n18379), .B1(n18554), .B2(n18398), .ZN(
        n18368) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18381), .B1(
        n18556), .B2(n18450), .ZN(n18367) );
  OAI211_X1 U21464 ( .C1(n18559), .C2(n18378), .A(n18368), .B(n18367), .ZN(
        P3_U2934) );
  AOI22_X1 U21465 ( .A1(n18560), .A2(n18379), .B1(n18562), .B2(n18380), .ZN(
        n18370) );
  AOI22_X1 U21466 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18381), .B1(
        n18561), .B2(n18398), .ZN(n18369) );
  OAI211_X1 U21467 ( .C1(n18565), .C2(n18448), .A(n18370), .B(n18369), .ZN(
        P3_U2935) );
  AOI22_X1 U21468 ( .A1(n18567), .A2(n18391), .B1(n18566), .B2(n18379), .ZN(
        n18372) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18381), .B1(
        n18568), .B2(n18380), .ZN(n18371) );
  OAI211_X1 U21470 ( .C1(n18571), .C2(n18448), .A(n18372), .B(n18371), .ZN(
        P3_U2936) );
  AOI22_X1 U21471 ( .A1(n18521), .A2(n18380), .B1(n18573), .B2(n18379), .ZN(
        n18374) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18381), .B1(
        n18574), .B2(n18450), .ZN(n18373) );
  OAI211_X1 U21473 ( .C1(n18524), .C2(n18375), .A(n18374), .B(n18373), .ZN(
        P3_U2937) );
  AOI22_X1 U21474 ( .A1(n18580), .A2(n18398), .B1(n18578), .B2(n18379), .ZN(
        n18377) );
  AOI22_X1 U21475 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18381), .B1(
        n18582), .B2(n18450), .ZN(n18376) );
  OAI211_X1 U21476 ( .C1(n18585), .C2(n18378), .A(n18377), .B(n18376), .ZN(
        P3_U2938) );
  AOI22_X1 U21477 ( .A1(n18591), .A2(n18398), .B1(n18588), .B2(n18379), .ZN(
        n18383) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18381), .B1(
        n18589), .B2(n18380), .ZN(n18382) );
  OAI211_X1 U21479 ( .C1(n18596), .C2(n18448), .A(n18383), .B(n18382), .ZN(
        P3_U2939) );
  NOR2_X1 U21480 ( .A1(n18433), .A2(n18476), .ZN(n18403) );
  AOI22_X1 U21481 ( .A1(n18503), .A2(n18398), .B1(n18537), .B2(n18403), .ZN(
        n18388) );
  NOR2_X1 U21482 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18384), .ZN(
        n18385) );
  NOR2_X1 U21483 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18433), .ZN(
        n18432) );
  AOI22_X1 U21484 ( .A1(n18542), .A2(n18385), .B1(n18539), .B2(n18432), .ZN(
        n18404) );
  NOR2_X2 U21485 ( .A1(n18433), .A2(n18386), .ZN(n18472) );
  AOI22_X1 U21486 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18404), .B1(
        n18472), .B2(n18543), .ZN(n18387) );
  OAI211_X1 U21487 ( .C1(n18511), .C2(n18424), .A(n18388), .B(n18387), .ZN(
        P3_U2940) );
  AOI22_X1 U21488 ( .A1(n18548), .A2(n18391), .B1(n18547), .B2(n18403), .ZN(
        n18390) );
  AOI22_X1 U21489 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18404), .B1(
        n18472), .B2(n18549), .ZN(n18389) );
  OAI211_X1 U21490 ( .C1(n18553), .C2(n18424), .A(n18390), .B(n18389), .ZN(
        P3_U2941) );
  AOI22_X1 U21491 ( .A1(n18414), .A2(n18391), .B1(n18555), .B2(n18403), .ZN(
        n18393) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18404), .B1(
        n18472), .B2(n18556), .ZN(n18392) );
  OAI211_X1 U21493 ( .C1(n18417), .C2(n18424), .A(n18393), .B(n18392), .ZN(
        P3_U2942) );
  INV_X1 U21494 ( .A(n18472), .ZN(n18470) );
  AOI22_X1 U21495 ( .A1(n18561), .A2(n18428), .B1(n18560), .B2(n18403), .ZN(
        n18395) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18404), .B1(
        n18562), .B2(n18398), .ZN(n18394) );
  OAI211_X1 U21497 ( .C1(n18470), .C2(n18565), .A(n18395), .B(n18394), .ZN(
        P3_U2943) );
  AOI22_X1 U21498 ( .A1(n18566), .A2(n18403), .B1(n18568), .B2(n18398), .ZN(
        n18397) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18404), .B1(
        n18567), .B2(n18428), .ZN(n18396) );
  OAI211_X1 U21500 ( .C1(n18470), .C2(n18571), .A(n18397), .B(n18396), .ZN(
        P3_U2944) );
  AOI22_X1 U21501 ( .A1(n18521), .A2(n18398), .B1(n18573), .B2(n18403), .ZN(
        n18400) );
  AOI22_X1 U21502 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18404), .B1(
        n18472), .B2(n18574), .ZN(n18399) );
  OAI211_X1 U21503 ( .C1(n18524), .C2(n18424), .A(n18400), .B(n18399), .ZN(
        P3_U2945) );
  AOI22_X1 U21504 ( .A1(n18525), .A2(n18398), .B1(n18578), .B2(n18403), .ZN(
        n18402) );
  AOI22_X1 U21505 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18404), .B1(
        n18472), .B2(n18582), .ZN(n18401) );
  OAI211_X1 U21506 ( .C1(n18530), .C2(n18424), .A(n18402), .B(n18401), .ZN(
        P3_U2946) );
  AOI22_X1 U21507 ( .A1(n18589), .A2(n18398), .B1(n18588), .B2(n18403), .ZN(
        n18406) );
  AOI22_X1 U21508 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18404), .B1(
        n18591), .B2(n18428), .ZN(n18405) );
  OAI211_X1 U21509 ( .C1(n18470), .C2(n18596), .A(n18406), .B(n18405), .ZN(
        P3_U2947) );
  NOR2_X1 U21510 ( .A1(n18635), .A2(n18433), .ZN(n18480) );
  NAND2_X1 U21511 ( .A1(n18407), .A2(n18480), .ZN(n18495) );
  NOR2_X1 U21512 ( .A1(n18472), .A2(n18498), .ZN(n18454) );
  NOR2_X1 U21513 ( .A1(n18454), .A2(n18502), .ZN(n18427) );
  AOI22_X1 U21514 ( .A1(n18503), .A2(n18428), .B1(n18537), .B2(n18427), .ZN(
        n18411) );
  OAI21_X1 U21515 ( .B1(n18408), .B2(n18505), .A(n18454), .ZN(n18409) );
  OAI211_X1 U21516 ( .C1(n18498), .C2(n18759), .A(n18508), .B(n18409), .ZN(
        n18429) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18429), .B1(
        n18498), .B2(n18543), .ZN(n18410) );
  OAI211_X1 U21518 ( .C1(n18511), .C2(n18448), .A(n18411), .B(n18410), .ZN(
        P3_U2948) );
  AOI22_X1 U21519 ( .A1(n18548), .A2(n18428), .B1(n18547), .B2(n18427), .ZN(
        n18413) );
  AOI22_X1 U21520 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18429), .B1(
        n18498), .B2(n18549), .ZN(n18412) );
  OAI211_X1 U21521 ( .C1(n18553), .C2(n18448), .A(n18413), .B(n18412), .ZN(
        P3_U2949) );
  AOI22_X1 U21522 ( .A1(n18414), .A2(n18428), .B1(n18555), .B2(n18427), .ZN(
        n18416) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18429), .B1(
        n18498), .B2(n18556), .ZN(n18415) );
  OAI211_X1 U21524 ( .C1(n18417), .C2(n18448), .A(n18416), .B(n18415), .ZN(
        P3_U2950) );
  AOI22_X1 U21525 ( .A1(n18561), .A2(n18450), .B1(n18560), .B2(n18427), .ZN(
        n18419) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18429), .B1(
        n18562), .B2(n18428), .ZN(n18418) );
  OAI211_X1 U21527 ( .C1(n18495), .C2(n18565), .A(n18419), .B(n18418), .ZN(
        P3_U2951) );
  AOI22_X1 U21528 ( .A1(n18567), .A2(n18450), .B1(n18566), .B2(n18427), .ZN(
        n18421) );
  AOI22_X1 U21529 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18429), .B1(
        n18568), .B2(n18428), .ZN(n18420) );
  OAI211_X1 U21530 ( .C1(n18495), .C2(n18571), .A(n18421), .B(n18420), .ZN(
        P3_U2952) );
  AOI22_X1 U21531 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18429), .B1(
        n18573), .B2(n18427), .ZN(n18423) );
  AOI22_X1 U21532 ( .A1(n18498), .A2(n18574), .B1(n18572), .B2(n18450), .ZN(
        n18422) );
  OAI211_X1 U21533 ( .C1(n18577), .C2(n18424), .A(n18423), .B(n18422), .ZN(
        P3_U2953) );
  AOI22_X1 U21534 ( .A1(n18525), .A2(n18428), .B1(n18578), .B2(n18427), .ZN(
        n18426) );
  AOI22_X1 U21535 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18429), .B1(
        n18498), .B2(n18582), .ZN(n18425) );
  OAI211_X1 U21536 ( .C1(n18530), .C2(n18448), .A(n18426), .B(n18425), .ZN(
        P3_U2954) );
  AOI22_X1 U21537 ( .A1(n18589), .A2(n18428), .B1(n18588), .B2(n18427), .ZN(
        n18431) );
  AOI22_X1 U21538 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18429), .B1(
        n18591), .B2(n18450), .ZN(n18430) );
  OAI211_X1 U21539 ( .C1(n18495), .C2(n18596), .A(n18431), .B(n18430), .ZN(
        P3_U2955) );
  AND2_X1 U21540 ( .A1(n18536), .A2(n18480), .ZN(n18449) );
  AOI22_X1 U21541 ( .A1(n18503), .A2(n18450), .B1(n18537), .B2(n18449), .ZN(
        n18435) );
  AOI22_X1 U21542 ( .A1(n18542), .A2(n18432), .B1(n18480), .B2(n18539), .ZN(
        n18451) );
  AOI22_X1 U21543 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18451), .B1(
        n18526), .B2(n18543), .ZN(n18434) );
  OAI211_X1 U21544 ( .C1(n18470), .C2(n18511), .A(n18435), .B(n18434), .ZN(
        P3_U2956) );
  AOI22_X1 U21545 ( .A1(n18472), .A2(n18483), .B1(n18547), .B2(n18449), .ZN(
        n18437) );
  AOI22_X1 U21546 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18451), .B1(
        n18526), .B2(n18549), .ZN(n18436) );
  OAI211_X1 U21547 ( .C1(n18486), .C2(n18448), .A(n18437), .B(n18436), .ZN(
        P3_U2957) );
  AOI22_X1 U21548 ( .A1(n18472), .A2(n18554), .B1(n18555), .B2(n18449), .ZN(
        n18439) );
  AOI22_X1 U21549 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18451), .B1(
        n18526), .B2(n18556), .ZN(n18438) );
  OAI211_X1 U21550 ( .C1(n18559), .C2(n18448), .A(n18439), .B(n18438), .ZN(
        P3_U2958) );
  INV_X1 U21551 ( .A(n18526), .ZN(n18516) );
  AOI22_X1 U21552 ( .A1(n18472), .A2(n18561), .B1(n18560), .B2(n18449), .ZN(
        n18441) );
  AOI22_X1 U21553 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18451), .B1(
        n18562), .B2(n18450), .ZN(n18440) );
  OAI211_X1 U21554 ( .C1(n18516), .C2(n18565), .A(n18441), .B(n18440), .ZN(
        P3_U2959) );
  AOI22_X1 U21555 ( .A1(n18566), .A2(n18449), .B1(n18568), .B2(n18450), .ZN(
        n18443) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18451), .B1(
        n18472), .B2(n18567), .ZN(n18442) );
  OAI211_X1 U21557 ( .C1(n18516), .C2(n18571), .A(n18443), .B(n18442), .ZN(
        P3_U2960) );
  AOI22_X1 U21558 ( .A1(n18472), .A2(n18572), .B1(n18573), .B2(n18449), .ZN(
        n18445) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18451), .B1(
        n18526), .B2(n18574), .ZN(n18444) );
  OAI211_X1 U21560 ( .C1(n18577), .C2(n18448), .A(n18445), .B(n18444), .ZN(
        P3_U2961) );
  AOI22_X1 U21561 ( .A1(n18472), .A2(n18580), .B1(n18578), .B2(n18449), .ZN(
        n18447) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18451), .B1(
        n18526), .B2(n18582), .ZN(n18446) );
  OAI211_X1 U21563 ( .C1(n18585), .C2(n18448), .A(n18447), .B(n18446), .ZN(
        P3_U2962) );
  AOI22_X1 U21564 ( .A1(n18472), .A2(n18591), .B1(n18588), .B2(n18449), .ZN(
        n18453) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18451), .B1(
        n18589), .B2(n18450), .ZN(n18452) );
  OAI211_X1 U21566 ( .C1(n18516), .C2(n18596), .A(n18453), .B(n18452), .ZN(
        P3_U2963) );
  NOR2_X2 U21567 ( .A1(n18636), .A2(n18477), .ZN(n18590) );
  INV_X1 U21568 ( .A(n18590), .ZN(n18586) );
  AOI21_X1 U21569 ( .B1(n18586), .B2(n18516), .A(n18502), .ZN(n18471) );
  AOI22_X1 U21570 ( .A1(n18498), .A2(n18538), .B1(n18537), .B2(n18471), .ZN(
        n18457) );
  AOI221_X1 U21571 ( .B1(n18454), .B2(n18516), .C1(n18505), .C2(n18516), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18455) );
  OAI21_X1 U21572 ( .B1(n18590), .B2(n18455), .A(n18508), .ZN(n18473) );
  AOI22_X1 U21573 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18473), .B1(
        n18590), .B2(n18543), .ZN(n18456) );
  OAI211_X1 U21574 ( .C1(n18546), .C2(n18470), .A(n18457), .B(n18456), .ZN(
        P3_U2964) );
  AOI22_X1 U21575 ( .A1(n18498), .A2(n18483), .B1(n18471), .B2(n18547), .ZN(
        n18459) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18473), .B1(
        n18590), .B2(n18549), .ZN(n18458) );
  OAI211_X1 U21577 ( .C1(n18470), .C2(n18486), .A(n18459), .B(n18458), .ZN(
        P3_U2965) );
  AOI22_X1 U21578 ( .A1(n18498), .A2(n18554), .B1(n18471), .B2(n18555), .ZN(
        n18461) );
  AOI22_X1 U21579 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18473), .B1(
        n18590), .B2(n18556), .ZN(n18460) );
  OAI211_X1 U21580 ( .C1(n18470), .C2(n18559), .A(n18461), .B(n18460), .ZN(
        P3_U2966) );
  AOI22_X1 U21581 ( .A1(n18472), .A2(n18562), .B1(n18471), .B2(n18560), .ZN(
        n18463) );
  AOI22_X1 U21582 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18473), .B1(
        n18498), .B2(n18561), .ZN(n18462) );
  OAI211_X1 U21583 ( .C1(n18586), .C2(n18565), .A(n18463), .B(n18462), .ZN(
        P3_U2967) );
  AOI22_X1 U21584 ( .A1(n18472), .A2(n18568), .B1(n18471), .B2(n18566), .ZN(
        n18465) );
  AOI22_X1 U21585 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18473), .B1(
        n18498), .B2(n18567), .ZN(n18464) );
  OAI211_X1 U21586 ( .C1(n18586), .C2(n18571), .A(n18465), .B(n18464), .ZN(
        P3_U2968) );
  AOI22_X1 U21587 ( .A1(n18498), .A2(n18572), .B1(n18471), .B2(n18573), .ZN(
        n18467) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18473), .B1(
        n18590), .B2(n18574), .ZN(n18466) );
  OAI211_X1 U21589 ( .C1(n18470), .C2(n18577), .A(n18467), .B(n18466), .ZN(
        P3_U2969) );
  AOI22_X1 U21590 ( .A1(n18498), .A2(n18580), .B1(n18471), .B2(n18578), .ZN(
        n18469) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18473), .B1(
        n18590), .B2(n18582), .ZN(n18468) );
  OAI211_X1 U21592 ( .C1(n18470), .C2(n18585), .A(n18469), .B(n18468), .ZN(
        P3_U2970) );
  AOI22_X1 U21593 ( .A1(n18472), .A2(n18589), .B1(n18471), .B2(n18588), .ZN(
        n18475) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18473), .B1(
        n18498), .B2(n18591), .ZN(n18474) );
  OAI211_X1 U21595 ( .C1(n18586), .C2(n18596), .A(n18475), .B(n18474), .ZN(
        P3_U2971) );
  NOR2_X1 U21596 ( .A1(n18477), .A2(n18476), .ZN(n18541) );
  AOI22_X1 U21597 ( .A1(n18526), .A2(n18538), .B1(n18537), .B2(n18541), .ZN(
        n18482) );
  INV_X1 U21598 ( .A(n18477), .ZN(n18479) );
  AOI22_X1 U21599 ( .A1(n18542), .A2(n18480), .B1(n18479), .B2(n18478), .ZN(
        n18499) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18499), .B1(
        n18543), .B2(n9560), .ZN(n18481) );
  OAI211_X1 U21601 ( .C1(n18546), .C2(n18495), .A(n18482), .B(n18481), .ZN(
        P3_U2972) );
  AOI22_X1 U21602 ( .A1(n18526), .A2(n18483), .B1(n18547), .B2(n18541), .ZN(
        n18485) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18499), .B1(
        n18549), .B2(n9560), .ZN(n18484) );
  OAI211_X1 U21604 ( .C1(n18495), .C2(n18486), .A(n18485), .B(n18484), .ZN(
        P3_U2973) );
  AOI22_X1 U21605 ( .A1(n18526), .A2(n18554), .B1(n18555), .B2(n18541), .ZN(
        n18488) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18499), .B1(
        n18556), .B2(n9560), .ZN(n18487) );
  OAI211_X1 U21607 ( .C1(n18495), .C2(n18559), .A(n18488), .B(n18487), .ZN(
        P3_U2974) );
  INV_X1 U21608 ( .A(n9560), .ZN(n18552) );
  AOI22_X1 U21609 ( .A1(n18526), .A2(n18561), .B1(n18560), .B2(n18541), .ZN(
        n18490) );
  AOI22_X1 U21610 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18499), .B1(
        n18498), .B2(n18562), .ZN(n18489) );
  OAI211_X1 U21611 ( .C1(n18565), .C2(n18552), .A(n18490), .B(n18489), .ZN(
        P3_U2975) );
  AOI22_X1 U21612 ( .A1(n18498), .A2(n18568), .B1(n18566), .B2(n18541), .ZN(
        n18492) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18499), .B1(
        n18526), .B2(n18567), .ZN(n18491) );
  OAI211_X1 U21614 ( .C1(n18571), .C2(n18552), .A(n18492), .B(n18491), .ZN(
        P3_U2976) );
  AOI22_X1 U21615 ( .A1(n18526), .A2(n18572), .B1(n18573), .B2(n18541), .ZN(
        n18494) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18499), .B1(
        n18574), .B2(n9560), .ZN(n18493) );
  OAI211_X1 U21617 ( .C1(n18495), .C2(n18577), .A(n18494), .B(n18493), .ZN(
        P3_U2977) );
  AOI22_X1 U21618 ( .A1(n18498), .A2(n18525), .B1(n18578), .B2(n18541), .ZN(
        n18497) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18499), .B1(
        n18582), .B2(n9560), .ZN(n18496) );
  OAI211_X1 U21620 ( .C1(n18516), .C2(n18530), .A(n18497), .B(n18496), .ZN(
        P3_U2978) );
  AOI22_X1 U21621 ( .A1(n18498), .A2(n18589), .B1(n18588), .B2(n18541), .ZN(
        n18501) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18499), .B1(
        n18526), .B2(n18591), .ZN(n18500) );
  OAI211_X1 U21623 ( .C1(n18596), .C2(n18552), .A(n18501), .B(n18500), .ZN(
        P3_U2979) );
  NOR2_X1 U21624 ( .A1(n18502), .A2(n18504), .ZN(n18531) );
  AOI22_X1 U21625 ( .A1(n18503), .A2(n18526), .B1(n18537), .B2(n18531), .ZN(
        n18510) );
  NOR2_X1 U21626 ( .A1(n18590), .A2(n18526), .ZN(n18506) );
  OAI21_X1 U21627 ( .B1(n18506), .B2(n18505), .A(n18504), .ZN(n18507) );
  OAI211_X1 U21628 ( .C1(n18527), .C2(n18759), .A(n18508), .B(n18507), .ZN(
        n18532) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18532), .B1(
        n18543), .B2(n18527), .ZN(n18509) );
  OAI211_X1 U21630 ( .C1(n18586), .C2(n18511), .A(n18510), .B(n18509), .ZN(
        P3_U2980) );
  AOI22_X1 U21631 ( .A1(n18526), .A2(n18548), .B1(n18547), .B2(n18531), .ZN(
        n18513) );
  AOI22_X1 U21632 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18532), .B1(
        n18549), .B2(n18527), .ZN(n18512) );
  OAI211_X1 U21633 ( .C1(n18586), .C2(n18553), .A(n18513), .B(n18512), .ZN(
        P3_U2981) );
  AOI22_X1 U21634 ( .A1(n18590), .A2(n18554), .B1(n18555), .B2(n18531), .ZN(
        n18515) );
  AOI22_X1 U21635 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18532), .B1(
        n18556), .B2(n18527), .ZN(n18514) );
  OAI211_X1 U21636 ( .C1(n18516), .C2(n18559), .A(n18515), .B(n18514), .ZN(
        P3_U2982) );
  AOI22_X1 U21637 ( .A1(n18526), .A2(n18562), .B1(n18560), .B2(n18531), .ZN(
        n18518) );
  AOI22_X1 U21638 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18532), .B1(
        n18590), .B2(n18561), .ZN(n18517) );
  OAI211_X1 U21639 ( .C1(n18565), .C2(n18535), .A(n18518), .B(n18517), .ZN(
        P3_U2983) );
  AOI22_X1 U21640 ( .A1(n18526), .A2(n18568), .B1(n18566), .B2(n18531), .ZN(
        n18520) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18532), .B1(
        n18590), .B2(n18567), .ZN(n18519) );
  OAI211_X1 U21642 ( .C1(n18571), .C2(n18535), .A(n18520), .B(n18519), .ZN(
        P3_U2984) );
  AOI22_X1 U21643 ( .A1(n18526), .A2(n18521), .B1(n18573), .B2(n18531), .ZN(
        n18523) );
  AOI22_X1 U21644 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18532), .B1(
        n18574), .B2(n18527), .ZN(n18522) );
  OAI211_X1 U21645 ( .C1(n18586), .C2(n18524), .A(n18523), .B(n18522), .ZN(
        P3_U2985) );
  AOI22_X1 U21646 ( .A1(n18526), .A2(n18525), .B1(n18578), .B2(n18531), .ZN(
        n18529) );
  AOI22_X1 U21647 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18532), .B1(
        n18582), .B2(n18527), .ZN(n18528) );
  OAI211_X1 U21648 ( .C1(n18586), .C2(n18530), .A(n18529), .B(n18528), .ZN(
        P3_U2986) );
  AOI22_X1 U21649 ( .A1(n18590), .A2(n18591), .B1(n18588), .B2(n18531), .ZN(
        n18534) );
  AOI22_X1 U21650 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18532), .B1(
        n18526), .B2(n18589), .ZN(n18533) );
  OAI211_X1 U21651 ( .C1(n18596), .C2(n18535), .A(n18534), .B(n18533), .ZN(
        P3_U2987) );
  AND2_X1 U21652 ( .A1(n18536), .A2(n18540), .ZN(n18587) );
  AOI22_X1 U21653 ( .A1(n18538), .A2(n9560), .B1(n18537), .B2(n18587), .ZN(
        n18545) );
  AOI22_X1 U21654 ( .A1(n18542), .A2(n18541), .B1(n18540), .B2(n18539), .ZN(
        n18592) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18592), .B1(
        n18543), .B2(n18581), .ZN(n18544) );
  OAI211_X1 U21656 ( .C1(n18546), .C2(n18586), .A(n18545), .B(n18544), .ZN(
        P3_U2988) );
  AOI22_X1 U21657 ( .A1(n18590), .A2(n18548), .B1(n18547), .B2(n18587), .ZN(
        n18551) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18592), .B1(
        n18549), .B2(n18581), .ZN(n18550) );
  OAI211_X1 U21659 ( .C1(n18553), .C2(n18552), .A(n18551), .B(n18550), .ZN(
        P3_U2989) );
  AOI22_X1 U21660 ( .A1(n18555), .A2(n18587), .B1(n18554), .B2(n9560), .ZN(
        n18558) );
  AOI22_X1 U21661 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18592), .B1(
        n18556), .B2(n18581), .ZN(n18557) );
  OAI211_X1 U21662 ( .C1(n18586), .C2(n18559), .A(n18558), .B(n18557), .ZN(
        P3_U2990) );
  AOI22_X1 U21663 ( .A1(n18561), .A2(n9560), .B1(n18560), .B2(n18587), .ZN(
        n18564) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18592), .B1(
        n18590), .B2(n18562), .ZN(n18563) );
  OAI211_X1 U21665 ( .C1(n18565), .C2(n18595), .A(n18564), .B(n18563), .ZN(
        P3_U2991) );
  AOI22_X1 U21666 ( .A1(n18567), .A2(n9560), .B1(n18566), .B2(n18587), .ZN(
        n18570) );
  AOI22_X1 U21667 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18592), .B1(
        n18590), .B2(n18568), .ZN(n18569) );
  OAI211_X1 U21668 ( .C1(n18571), .C2(n18595), .A(n18570), .B(n18569), .ZN(
        P3_U2992) );
  AOI22_X1 U21669 ( .A1(n18573), .A2(n18587), .B1(n18572), .B2(n9560), .ZN(
        n18576) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18592), .B1(
        n18574), .B2(n18581), .ZN(n18575) );
  OAI211_X1 U21671 ( .C1(n18586), .C2(n18577), .A(n18576), .B(n18575), .ZN(
        P3_U2993) );
  AOI22_X1 U21672 ( .A1(n18580), .A2(n9560), .B1(n18578), .B2(n18587), .ZN(
        n18584) );
  AOI22_X1 U21673 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18592), .B1(
        n18582), .B2(n18581), .ZN(n18583) );
  OAI211_X1 U21674 ( .C1(n18586), .C2(n18585), .A(n18584), .B(n18583), .ZN(
        P3_U2994) );
  AOI22_X1 U21675 ( .A1(n18590), .A2(n18589), .B1(n18588), .B2(n18587), .ZN(
        n18594) );
  AOI22_X1 U21676 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18592), .B1(
        n18591), .B2(n9560), .ZN(n18593) );
  OAI211_X1 U21677 ( .C1(n18596), .C2(n18595), .A(n18594), .B(n18593), .ZN(
        P3_U2995) );
  NOR2_X1 U21678 ( .A1(n18609), .A2(n18597), .ZN(n18600) );
  OAI222_X1 U21679 ( .A1(n18603), .A2(n18602), .B1(n18601), .B2(n18600), .C1(
        n18599), .C2(n18598), .ZN(n18802) );
  OAI21_X1 U21680 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18604), .ZN(n18605) );
  OAI211_X1 U21681 ( .C1(n18607), .C2(n18627), .A(n18606), .B(n18605), .ZN(
        n18649) );
  AOI21_X1 U21682 ( .B1(n18628), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n18608), .ZN(n18631) );
  INV_X1 U21683 ( .A(n18631), .ZN(n18621) );
  AOI22_X1 U21684 ( .A1(n18613), .A2(n18621), .B1(n18609), .B2(n18614), .ZN(
        n18764) );
  NOR2_X1 U21685 ( .A1(n18638), .A2(n18764), .ZN(n18619) );
  AOI21_X1 U21686 ( .B1(n18612), .B2(n18611), .A(n18610), .ZN(n18622) );
  OAI21_X1 U21687 ( .B1(n18613), .B2(n18630), .A(n18622), .ZN(n18616) );
  INV_X1 U21688 ( .A(n18614), .ZN(n18615) );
  AOI21_X1 U21689 ( .B1(n18617), .B2(n18616), .A(n18615), .ZN(n18761) );
  NAND2_X1 U21690 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18761), .ZN(
        n18618) );
  OAI22_X1 U21691 ( .A1(n18619), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n18638), .B2(n18618), .ZN(n18647) );
  OAI211_X1 U21692 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18621), .B(n18620), .ZN(
        n18625) );
  OR3_X1 U21693 ( .A1(n18777), .A2(n18623), .A3(n18622), .ZN(n18624) );
  OAI211_X1 U21694 ( .C1(n18773), .C2(n18626), .A(n18625), .B(n18624), .ZN(
        n18775) );
  MUX2_X1 U21695 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n18775), .S(
        n18627), .Z(n18642) );
  NOR2_X1 U21696 ( .A1(n18629), .A2(n18628), .ZN(n18633) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18630), .B1(
        n18633), .B2(n20806), .ZN(n18785) );
  OAI22_X1 U21698 ( .A1(n18633), .A2(n18632), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18631), .ZN(n18781) );
  AOI222_X1 U21699 ( .A1(n18785), .A2(n18781), .B1(n18785), .B2(n18635), .C1(
        n18781), .C2(n18634), .ZN(n18637) );
  OAI21_X1 U21700 ( .B1(n18638), .B2(n18637), .A(n18636), .ZN(n18641) );
  AND2_X1 U21701 ( .A1(n18642), .A2(n18641), .ZN(n18639) );
  OAI221_X1 U21702 ( .B1(n18642), .B2(n18641), .C1(n18640), .C2(n18639), .A(
        n18644), .ZN(n18646) );
  AOI21_X1 U21703 ( .B1(n18644), .B2(n18643), .A(n18642), .ZN(n18645) );
  AOI222_X1 U21704 ( .A1(n18647), .A2(n18646), .B1(n18647), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18646), .C2(n18645), .ZN(
        n18648) );
  NOR4_X1 U21705 ( .A1(n18650), .A2(n18802), .A3(n18649), .A4(n18648), .ZN(
        n18658) );
  AOI22_X1 U21706 ( .A1(n18784), .A2(n18666), .B1(n18806), .B2(n17404), .ZN(
        n18655) );
  AOI21_X1 U21707 ( .B1(n18652), .B2(n18651), .A(n18657), .ZN(n18653) );
  AOI21_X1 U21708 ( .B1(n18658), .B2(n18653), .A(n18809), .ZN(n18760) );
  NAND2_X1 U21709 ( .A1(n18806), .A2(n18805), .ZN(n18659) );
  OAI211_X1 U21710 ( .C1(n18808), .C2(n18759), .A(n18760), .B(n18659), .ZN(
        n18662) );
  OAI22_X1 U21711 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18655), .B1(n18654), 
        .B2(n18662), .ZN(n18656) );
  OAI21_X1 U21712 ( .B1(n18658), .B2(n18657), .A(n18656), .ZN(P3_U2996) );
  NOR3_X1 U21713 ( .A1(n18809), .A2(n18770), .A3(n18659), .ZN(n18664) );
  AOI211_X1 U21714 ( .C1(n18806), .C2(n17404), .A(n18660), .B(n18664), .ZN(
        n18661) );
  OAI21_X1 U21715 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n18662), .A(n18661), 
        .ZN(P3_U2997) );
  NOR4_X1 U21716 ( .A1(n18666), .A2(n18665), .A3(n18664), .A4(n18663), .ZN(
        P3_U2998) );
  INV_X1 U21717 ( .A(n18757), .ZN(n18754) );
  AND2_X1 U21718 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18754), .ZN(
        P3_U2999) );
  AND2_X1 U21719 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18754), .ZN(
        P3_U3000) );
  AND2_X1 U21720 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18754), .ZN(
        P3_U3001) );
  AND2_X1 U21721 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18754), .ZN(
        P3_U3002) );
  AND2_X1 U21722 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18754), .ZN(
        P3_U3003) );
  AND2_X1 U21723 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18754), .ZN(
        P3_U3004) );
  AND2_X1 U21724 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18754), .ZN(
        P3_U3005) );
  AND2_X1 U21725 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18754), .ZN(
        P3_U3006) );
  AND2_X1 U21726 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18754), .ZN(
        P3_U3007) );
  AND2_X1 U21727 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18754), .ZN(
        P3_U3008) );
  AND2_X1 U21728 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18754), .ZN(
        P3_U3009) );
  AND2_X1 U21729 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18754), .ZN(
        P3_U3010) );
  AND2_X1 U21730 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18754), .ZN(
        P3_U3011) );
  AND2_X1 U21731 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18754), .ZN(
        P3_U3012) );
  AND2_X1 U21732 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18754), .ZN(
        P3_U3013) );
  AND2_X1 U21733 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18754), .ZN(
        P3_U3014) );
  AND2_X1 U21734 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18754), .ZN(
        P3_U3015) );
  AND2_X1 U21735 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18754), .ZN(
        P3_U3016) );
  AND2_X1 U21736 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18754), .ZN(
        P3_U3017) );
  AND2_X1 U21737 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18754), .ZN(
        P3_U3018) );
  AND2_X1 U21738 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18754), .ZN(
        P3_U3019) );
  AND2_X1 U21739 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18754), .ZN(
        P3_U3020) );
  AND2_X1 U21740 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18754), .ZN(P3_U3021) );
  AND2_X1 U21741 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18754), .ZN(P3_U3022) );
  AND2_X1 U21742 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18754), .ZN(P3_U3023) );
  AND2_X1 U21743 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18754), .ZN(P3_U3024) );
  AND2_X1 U21744 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18754), .ZN(P3_U3025) );
  AND2_X1 U21745 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18754), .ZN(P3_U3026) );
  AND2_X1 U21746 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18754), .ZN(P3_U3027) );
  AND2_X1 U21747 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18754), .ZN(P3_U3028) );
  OAI21_X1 U21748 ( .B1(n20684), .B2(n18667), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18668) );
  INV_X1 U21749 ( .A(n18668), .ZN(n18671) );
  NAND2_X1 U21750 ( .A1(n18806), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18678) );
  INV_X1 U21751 ( .A(n18678), .ZN(n18673) );
  NOR2_X1 U21752 ( .A1(n18673), .A2(n18682), .ZN(n18684) );
  INV_X1 U21753 ( .A(NA), .ZN(n20694) );
  OAI21_X1 U21754 ( .B1(n20694), .B2(n18669), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18683) );
  INV_X1 U21755 ( .A(n18683), .ZN(n18670) );
  OAI22_X1 U21756 ( .A1(n18800), .A2(n18671), .B1(n18684), .B2(n18670), .ZN(
        P3_U3029) );
  NOR2_X1 U21757 ( .A1(n18685), .A2(n20684), .ZN(n18680) );
  INV_X1 U21758 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18672) );
  NOR3_X1 U21759 ( .A1(n18680), .A2(n18672), .A3(n18682), .ZN(n18674) );
  NOR2_X1 U21760 ( .A1(n18674), .A2(n18673), .ZN(n18676) );
  OAI211_X1 U21761 ( .C1(n20684), .C2(n18677), .A(n18676), .B(n18675), .ZN(
        P3_U3030) );
  OAI22_X1 U21762 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18678), .ZN(n18679) );
  OAI22_X1 U21763 ( .A1(n18680), .A2(n18679), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18681) );
  OAI22_X1 U21764 ( .A1(n18684), .A2(n18683), .B1(n18682), .B2(n18681), .ZN(
        P3_U3031) );
  OAI222_X1 U21765 ( .A1(n20843), .A2(n18739), .B1(n18686), .B2(n18800), .C1(
        n18687), .C2(n18743), .ZN(P3_U3032) );
  OAI222_X1 U21766 ( .A1(n18743), .A2(n18689), .B1(n18688), .B2(n18800), .C1(
        n18687), .C2(n18747), .ZN(P3_U3033) );
  OAI222_X1 U21767 ( .A1(n18743), .A2(n18691), .B1(n18690), .B2(n18800), .C1(
        n18689), .C2(n18739), .ZN(P3_U3034) );
  INV_X1 U21768 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18694) );
  OAI222_X1 U21769 ( .A1(n18743), .A2(n18694), .B1(n18692), .B2(n18800), .C1(
        n18691), .C2(n18739), .ZN(P3_U3035) );
  OAI222_X1 U21770 ( .A1(n18694), .A2(n18739), .B1(n18693), .B2(n18800), .C1(
        n18695), .C2(n18743), .ZN(P3_U3036) );
  OAI222_X1 U21771 ( .A1(n18743), .A2(n18697), .B1(n18696), .B2(n18800), .C1(
        n18695), .C2(n18739), .ZN(P3_U3037) );
  OAI222_X1 U21772 ( .A1(n18743), .A2(n18700), .B1(n18698), .B2(n18800), .C1(
        n18697), .C2(n18739), .ZN(P3_U3038) );
  OAI222_X1 U21773 ( .A1(n18700), .A2(n18739), .B1(n18699), .B2(n18800), .C1(
        n18701), .C2(n18743), .ZN(P3_U3039) );
  OAI222_X1 U21774 ( .A1(n18743), .A2(n18703), .B1(n18702), .B2(n18800), .C1(
        n18701), .C2(n18739), .ZN(P3_U3040) );
  OAI222_X1 U21775 ( .A1(n18743), .A2(n18705), .B1(n18704), .B2(n18800), .C1(
        n18703), .C2(n18739), .ZN(P3_U3041) );
  OAI222_X1 U21776 ( .A1(n18743), .A2(n18707), .B1(n18706), .B2(n18800), .C1(
        n18705), .C2(n18739), .ZN(P3_U3042) );
  OAI222_X1 U21777 ( .A1(n18743), .A2(n18709), .B1(n18708), .B2(n18800), .C1(
        n18707), .C2(n18739), .ZN(P3_U3043) );
  INV_X1 U21778 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18712) );
  OAI222_X1 U21779 ( .A1(n18743), .A2(n18712), .B1(n18710), .B2(n18800), .C1(
        n18709), .C2(n18739), .ZN(P3_U3044) );
  OAI222_X1 U21780 ( .A1(n18712), .A2(n18739), .B1(n18711), .B2(n18800), .C1(
        n18713), .C2(n18743), .ZN(P3_U3045) );
  INV_X1 U21781 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18715) );
  OAI222_X1 U21782 ( .A1(n18743), .A2(n18715), .B1(n18714), .B2(n18800), .C1(
        n18713), .C2(n18747), .ZN(P3_U3046) );
  OAI222_X1 U21783 ( .A1(n18743), .A2(n18718), .B1(n18716), .B2(n18800), .C1(
        n18715), .C2(n18747), .ZN(P3_U3047) );
  OAI222_X1 U21784 ( .A1(n18718), .A2(n18739), .B1(n18717), .B2(n18800), .C1(
        n18719), .C2(n18743), .ZN(P3_U3048) );
  OAI222_X1 U21785 ( .A1(n18743), .A2(n18722), .B1(n18720), .B2(n18800), .C1(
        n18719), .C2(n18747), .ZN(P3_U3049) );
  OAI222_X1 U21786 ( .A1(n18722), .A2(n18739), .B1(n18721), .B2(n18800), .C1(
        n18723), .C2(n18743), .ZN(P3_U3050) );
  OAI222_X1 U21787 ( .A1(n18743), .A2(n18726), .B1(n18724), .B2(n18800), .C1(
        n18723), .C2(n18747), .ZN(P3_U3051) );
  INV_X1 U21788 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18727) );
  OAI222_X1 U21789 ( .A1(n18726), .A2(n18739), .B1(n18725), .B2(n18800), .C1(
        n18727), .C2(n18743), .ZN(P3_U3052) );
  OAI222_X1 U21790 ( .A1(n18743), .A2(n18730), .B1(n18728), .B2(n18800), .C1(
        n18727), .C2(n18747), .ZN(P3_U3053) );
  OAI222_X1 U21791 ( .A1(n18730), .A2(n18739), .B1(n18729), .B2(n18800), .C1(
        n18731), .C2(n18743), .ZN(P3_U3054) );
  OAI222_X1 U21792 ( .A1(n18743), .A2(n18733), .B1(n18732), .B2(n18800), .C1(
        n18731), .C2(n18747), .ZN(P3_U3055) );
  OAI222_X1 U21793 ( .A1(n18743), .A2(n18735), .B1(n18734), .B2(n18800), .C1(
        n18733), .C2(n18747), .ZN(P3_U3056) );
  OAI222_X1 U21794 ( .A1(n18743), .A2(n18736), .B1(n20868), .B2(n18800), .C1(
        n18735), .C2(n18739), .ZN(P3_U3057) );
  INV_X1 U21795 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18740) );
  OAI222_X1 U21796 ( .A1(n18743), .A2(n18740), .B1(n18737), .B2(n18800), .C1(
        n18736), .C2(n18739), .ZN(P3_U3058) );
  OAI222_X1 U21797 ( .A1(n18740), .A2(n18739), .B1(n18738), .B2(n18800), .C1(
        n18741), .C2(n18743), .ZN(P3_U3059) );
  OAI222_X1 U21798 ( .A1(n18743), .A2(n18746), .B1(n18742), .B2(n18800), .C1(
        n18741), .C2(n18747), .ZN(P3_U3060) );
  OAI222_X1 U21799 ( .A1(n18747), .A2(n18746), .B1(n18745), .B2(n18800), .C1(
        n18744), .C2(n18743), .ZN(P3_U3061) );
  OAI22_X1 U21800 ( .A1(n18817), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18800), .ZN(n18748) );
  INV_X1 U21801 ( .A(n18748), .ZN(P3_U3274) );
  OAI22_X1 U21802 ( .A1(n18817), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18800), .ZN(n18749) );
  INV_X1 U21803 ( .A(n18749), .ZN(P3_U3275) );
  OAI22_X1 U21804 ( .A1(n18817), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18800), .ZN(n18750) );
  INV_X1 U21805 ( .A(n18750), .ZN(P3_U3276) );
  OAI22_X1 U21806 ( .A1(n18817), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18800), .ZN(n18751) );
  INV_X1 U21807 ( .A(n18751), .ZN(P3_U3277) );
  INV_X1 U21808 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18753) );
  INV_X1 U21809 ( .A(n18755), .ZN(n18752) );
  AOI21_X1 U21810 ( .B1(n18754), .B2(n18753), .A(n18752), .ZN(P3_U3280) );
  OAI21_X1 U21811 ( .B1(n18757), .B2(n18756), .A(n18755), .ZN(P3_U3281) );
  OAI21_X1 U21812 ( .B1(n18760), .B2(n18759), .A(n18758), .ZN(P3_U3282) );
  NOR2_X1 U21813 ( .A1(n18761), .A2(n18763), .ZN(n18762) );
  NOR2_X1 U21814 ( .A1(n18762), .A2(n18790), .ZN(n18768) );
  NOR3_X1 U21815 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18764), .A3(
        n18763), .ZN(n18765) );
  AOI21_X1 U21816 ( .B1(n18766), .B2(n18784), .A(n18765), .ZN(n18767) );
  OAI22_X1 U21817 ( .A1(n18769), .A2(n18768), .B1(n18790), .B2(n18767), .ZN(
        P3_U3285) );
  NOR2_X1 U21818 ( .A1(n18770), .A2(n18787), .ZN(n18778) );
  OAI22_X1 U21819 ( .A1(n18772), .A2(n18771), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18779) );
  INV_X1 U21820 ( .A(n18779), .ZN(n18774) );
  AOI222_X1 U21821 ( .A1(n18775), .A2(n18786), .B1(n18778), .B2(n18774), .C1(
        n18784), .C2(n18773), .ZN(n18776) );
  AOI22_X1 U21822 ( .A1(n18790), .A2(n18777), .B1(n18776), .B2(n18788), .ZN(
        P3_U3288) );
  AOI222_X1 U21823 ( .A1(n18781), .A2(n18786), .B1(n18784), .B2(n18780), .C1(
        n18779), .C2(n18778), .ZN(n18782) );
  AOI22_X1 U21824 ( .A1(n18790), .A2(n18783), .B1(n18782), .B2(n18788), .ZN(
        P3_U3289) );
  AOI222_X1 U21825 ( .A1(n18787), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18786), 
        .B2(n18785), .C1(n20806), .C2(n18784), .ZN(n18789) );
  AOI22_X1 U21826 ( .A1(n18790), .A2(n20806), .B1(n18789), .B2(n18788), .ZN(
        P3_U3290) );
  AOI21_X1 U21827 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18791) );
  AOI22_X1 U21828 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18791), .B2(n20843), .ZN(n18793) );
  INV_X1 U21829 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18792) );
  AOI22_X1 U21830 ( .A1(n18794), .A2(n18793), .B1(n18792), .B2(n18797), .ZN(
        P3_U3292) );
  INV_X1 U21831 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18798) );
  NOR2_X1 U21832 ( .A1(n18797), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18795) );
  AOI22_X1 U21833 ( .A1(n18798), .A2(n18797), .B1(n18796), .B2(n18795), .ZN(
        P3_U3293) );
  INV_X1 U21834 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18799) );
  AOI22_X1 U21835 ( .A1(n18800), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18799), 
        .B2(n18817), .ZN(P3_U3294) );
  MUX2_X1 U21836 ( .A(P3_MORE_REG_SCAN_IN), .B(n18802), .S(n18801), .Z(
        P3_U3295) );
  OAI21_X1 U21837 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18804), .A(n18803), 
        .ZN(n18807) );
  AOI211_X1 U21838 ( .C1(n18820), .C2(n18807), .A(n18806), .B(n18805), .ZN(
        n18810) );
  OAI21_X1 U21839 ( .B1(n18810), .B2(n18809), .A(n18808), .ZN(n18816) );
  OAI21_X1 U21840 ( .B1(n18812), .B2(n18811), .A(n18821), .ZN(n18813) );
  AOI21_X1 U21841 ( .B1(n17404), .B2(n18814), .A(n18813), .ZN(n18815) );
  MUX2_X1 U21842 ( .A(n18816), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n18815), 
        .Z(P3_U3296) );
  MUX2_X1 U21843 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .B(P3_M_IO_N_REG_SCAN_IN), 
        .S(n18817), .Z(P3_U3297) );
  INV_X1 U21844 ( .A(n18818), .ZN(n18822) );
  OAI21_X1 U21845 ( .B1(n18822), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n18821), 
        .ZN(n18819) );
  OAI21_X1 U21846 ( .B1(n18821), .B2(n18820), .A(n18819), .ZN(P3_U3298) );
  NOR2_X1 U21847 ( .A1(n18822), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18824)
         );
  OAI21_X1 U21848 ( .B1(n18825), .B2(n18824), .A(n18823), .ZN(P3_U3299) );
  INV_X1 U21849 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19739) );
  NAND2_X1 U21850 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19739), .ZN(n19732) );
  OR2_X1 U21851 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19729) );
  OAI21_X1 U21852 ( .B1(n19728), .B2(n19732), .A(n19729), .ZN(n19798) );
  AOI21_X1 U21853 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19798), .ZN(n18826) );
  INV_X1 U21854 ( .A(n18826), .ZN(P2_U2815) );
  INV_X1 U21855 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n20812) );
  OAI22_X1 U21856 ( .A1(n18829), .A2(n20812), .B1(n18828), .B2(n18827), .ZN(
        P2_U2816) );
  AOI22_X1 U21857 ( .A1(n19868), .A2(n20812), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n19869), .ZN(n18830) );
  OAI21_X1 U21858 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19733), .A(n18830), 
        .ZN(P2_U2817) );
  OAI21_X1 U21859 ( .B1(n19723), .B2(BS16), .A(n19798), .ZN(n19796) );
  OAI21_X1 U21860 ( .B1(n19798), .B2(n19446), .A(n19796), .ZN(P2_U2818) );
  NOR2_X1 U21861 ( .A1(n18831), .A2(n19714), .ZN(n19840) );
  OAI21_X1 U21862 ( .B1(n19840), .B2(n18833), .A(n18832), .ZN(P2_U2819) );
  NOR4_X1 U21863 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18837) );
  NOR4_X1 U21864 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18836) );
  NOR4_X1 U21865 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18835) );
  NOR4_X1 U21866 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18834) );
  NAND4_X1 U21867 ( .A1(n18837), .A2(n18836), .A3(n18835), .A4(n18834), .ZN(
        n18843) );
  NOR4_X1 U21868 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18841) );
  AOI211_X1 U21869 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_21__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18840) );
  NOR4_X1 U21870 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18839) );
  NOR4_X1 U21871 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18838) );
  NAND4_X1 U21872 ( .A1(n18841), .A2(n18840), .A3(n18839), .A4(n18838), .ZN(
        n18842) );
  NOR2_X1 U21873 ( .A1(n18843), .A2(n18842), .ZN(n18854) );
  INV_X1 U21874 ( .A(n18854), .ZN(n18845) );
  NOR2_X1 U21875 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18845), .ZN(n18847) );
  INV_X1 U21876 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18844) );
  AOI22_X1 U21877 ( .A1(n18847), .A2(n18848), .B1(n18845), .B2(n18844), .ZN(
        P2_U2820) );
  NOR2_X1 U21878 ( .A1(n18854), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18846)
         );
  OR4_X1 U21879 ( .A1(n18845), .A2(P2_REIP_REG_0__SCAN_IN), .A3(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A4(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n18852) );
  OAI21_X1 U21880 ( .B1(n18847), .B2(n18846), .A(n18852), .ZN(P2_U2821) );
  INV_X1 U21881 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19797) );
  NAND2_X1 U21882 ( .A1(n18847), .A2(n19797), .ZN(n18851) );
  OAI21_X1 U21883 ( .B1(n19740), .B2(n18848), .A(n18854), .ZN(n18849) );
  OAI21_X1 U21884 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18854), .A(n18849), 
        .ZN(n18850) );
  OAI221_X1 U21885 ( .B1(n18851), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18851), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18850), .ZN(P2_U2822) );
  INV_X1 U21886 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18853) );
  OAI211_X1 U21887 ( .C1(n18854), .C2(n18853), .A(n18852), .B(n18851), .ZN(
        P2_U2823) );
  OAI22_X1 U21888 ( .A1(n18858), .A2(n18857), .B1(n18856), .B2(n18855), .ZN(
        n18867) );
  INV_X1 U21889 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19774) );
  OAI222_X1 U21890 ( .A1(n19008), .A2(n18860), .B1(n19009), .B2(n18859), .C1(
        n18993), .C2(n19774), .ZN(n18861) );
  AOI21_X1 U21891 ( .B1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n19041), .A(
        n18861), .ZN(n18866) );
  OAI22_X1 U21892 ( .A1(n18863), .A2(n19006), .B1(n18862), .B2(n19011), .ZN(
        n18864) );
  INV_X1 U21893 ( .A(n18864), .ZN(n18865) );
  OAI211_X1 U21894 ( .C1(n19720), .C2(n18867), .A(n18866), .B(n18865), .ZN(
        P2_U2834) );
  NAND2_X1 U21895 ( .A1(n13017), .A2(n18868), .ZN(n18869) );
  XOR2_X1 U21896 ( .A(n18870), .B(n18869), .Z(n18879) );
  AOI22_X1 U21897 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n19041), .B1(
        P2_REIP_REG_19__SCAN_IN), .B2(n19031), .ZN(n18871) );
  OAI21_X1 U21898 ( .B1(n18872), .B2(n19008), .A(n18871), .ZN(n18873) );
  AOI211_X1 U21899 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19025), .A(n19155), .B(
        n18873), .ZN(n18878) );
  OAI22_X1 U21900 ( .A1(n18875), .A2(n19006), .B1(n18874), .B2(n19011), .ZN(
        n18876) );
  INV_X1 U21901 ( .A(n18876), .ZN(n18877) );
  OAI211_X1 U21902 ( .C1(n19720), .C2(n18879), .A(n18878), .B(n18877), .ZN(
        P2_U2836) );
  AOI22_X1 U21903 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19041), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19031), .ZN(n18892) );
  INV_X1 U21904 ( .A(n18880), .ZN(n18882) );
  OAI22_X1 U21905 ( .A1(n18882), .A2(n19008), .B1(n18881), .B2(n18887), .ZN(
        n18883) );
  AOI211_X1 U21906 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19025), .A(n19155), .B(
        n18883), .ZN(n18891) );
  AOI22_X1 U21907 ( .A1(n18885), .A2(n19027), .B1(n18884), .B2(n19022), .ZN(
        n18890) );
  OAI21_X1 U21908 ( .B1(n18888), .B2(n18887), .A(n18886), .ZN(n18889) );
  NAND4_X1 U21909 ( .A1(n18892), .A2(n18891), .A3(n18890), .A4(n18889), .ZN(
        P2_U2838) );
  NOR2_X1 U21910 ( .A1(n13016), .A2(n18893), .ZN(n18895) );
  XOR2_X1 U21911 ( .A(n18895), .B(n18894), .Z(n18906) );
  INV_X1 U21912 ( .A(n18896), .ZN(n18897) );
  AOI22_X1 U21913 ( .A1(n18897), .A2(n19030), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19041), .ZN(n18898) );
  OAI211_X1 U21914 ( .C1(n18899), .C2(n19009), .A(n18898), .B(n18992), .ZN(
        n18900) );
  AOI21_X1 U21915 ( .B1(P2_REIP_REG_16__SCAN_IN), .B2(n19031), .A(n18900), 
        .ZN(n18905) );
  INV_X1 U21916 ( .A(n18901), .ZN(n18902) );
  OAI22_X1 U21917 ( .A1(n19055), .A2(n19006), .B1(n18902), .B2(n19011), .ZN(
        n18903) );
  INV_X1 U21918 ( .A(n18903), .ZN(n18904) );
  OAI211_X1 U21919 ( .C1(n19720), .C2(n18906), .A(n18905), .B(n18904), .ZN(
        P2_U2839) );
  NAND2_X1 U21920 ( .A1(n13017), .A2(n18907), .ZN(n18909) );
  XNOR2_X1 U21921 ( .A(n18909), .B(n18908), .ZN(n18916) );
  AOI22_X1 U21922 ( .A1(n18910), .A2(n19030), .B1(P2_REIP_REG_15__SCAN_IN), 
        .B2(n19031), .ZN(n18911) );
  OAI211_X1 U21923 ( .C1(n10814), .C2(n19009), .A(n18911), .B(n18992), .ZN(
        n18914) );
  OAI22_X1 U21924 ( .A1(n19061), .A2(n19006), .B1(n18912), .B2(n19011), .ZN(
        n18913) );
  AOI211_X1 U21925 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n19041), .A(
        n18914), .B(n18913), .ZN(n18915) );
  OAI21_X1 U21926 ( .B1(n18916), .B2(n19720), .A(n18915), .ZN(P2_U2840) );
  OAI21_X1 U21927 ( .B1(n10805), .B2(n19009), .A(n18992), .ZN(n18920) );
  OAI22_X1 U21928 ( .A1(n18918), .A2(n19008), .B1(n18991), .B2(n18917), .ZN(
        n18919) );
  AOI211_X1 U21929 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n19031), .A(n18920), 
        .B(n18919), .ZN(n18927) );
  NAND2_X1 U21930 ( .A1(n13017), .A2(n18921), .ZN(n18922) );
  XNOR2_X1 U21931 ( .A(n18923), .B(n18922), .ZN(n18925) );
  AOI22_X1 U21932 ( .A1(n18925), .A2(n19002), .B1(n19022), .B2(n18924), .ZN(
        n18926) );
  OAI211_X1 U21933 ( .C1(n19067), .C2(n19006), .A(n18927), .B(n18926), .ZN(
        P2_U2842) );
  NOR2_X1 U21934 ( .A1(n13016), .A2(n18928), .ZN(n18930) );
  XOR2_X1 U21935 ( .A(n18930), .B(n18929), .Z(n18937) );
  AOI22_X1 U21936 ( .A1(n19025), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19041), .ZN(n18931) );
  OAI21_X1 U21937 ( .B1(n18932), .B2(n19008), .A(n18931), .ZN(n18933) );
  AOI211_X1 U21938 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19031), .A(n19155), 
        .B(n18933), .ZN(n18936) );
  AOI22_X1 U21939 ( .A1(n19068), .A2(n19027), .B1(n19022), .B2(n18934), .ZN(
        n18935) );
  OAI211_X1 U21940 ( .C1(n19720), .C2(n18937), .A(n18936), .B(n18935), .ZN(
        P2_U2843) );
  NAND2_X1 U21941 ( .A1(n13017), .A2(n18938), .ZN(n18940) );
  XOR2_X1 U21942 ( .A(n18940), .B(n18939), .Z(n18949) );
  INV_X1 U21943 ( .A(n18941), .ZN(n18942) );
  AOI22_X1 U21944 ( .A1(n18942), .A2(n19030), .B1(n19031), .B2(
        P2_REIP_REG_11__SCAN_IN), .ZN(n18943) );
  OAI211_X1 U21945 ( .C1(n18944), .C2(n19009), .A(n18943), .B(n18992), .ZN(
        n18947) );
  OAI22_X1 U21946 ( .A1(n19073), .A2(n19006), .B1(n19011), .B2(n18945), .ZN(
        n18946) );
  AOI211_X1 U21947 ( .C1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n19041), .A(
        n18947), .B(n18946), .ZN(n18948) );
  OAI21_X1 U21948 ( .B1(n18949), .B2(n19720), .A(n18948), .ZN(P2_U2844) );
  INV_X1 U21949 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18960) );
  OAI22_X1 U21950 ( .A1(n18950), .A2(n19008), .B1(n19757), .B2(n18993), .ZN(
        n18951) );
  AOI211_X1 U21951 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n19025), .A(n19155), .B(
        n18951), .ZN(n18959) );
  NOR2_X1 U21952 ( .A1(n13016), .A2(n18952), .ZN(n18953) );
  XNOR2_X1 U21953 ( .A(n18954), .B(n18953), .ZN(n18957) );
  OAI22_X1 U21954 ( .A1(n19076), .A2(n19006), .B1(n19011), .B2(n18955), .ZN(
        n18956) );
  AOI21_X1 U21955 ( .B1(n18957), .B2(n19002), .A(n18956), .ZN(n18958) );
  OAI211_X1 U21956 ( .C1(n18960), .C2(n18991), .A(n18959), .B(n18958), .ZN(
        P2_U2845) );
  NAND2_X1 U21957 ( .A1(n13017), .A2(n18961), .ZN(n18963) );
  XOR2_X1 U21958 ( .A(n18963), .B(n18962), .Z(n18970) );
  AOI22_X1 U21959 ( .A1(n18964), .A2(n19030), .B1(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19041), .ZN(n18965) );
  OAI211_X1 U21960 ( .C1(n19755), .C2(n18993), .A(n18965), .B(n18992), .ZN(
        n18968) );
  OAI22_X1 U21961 ( .A1(n19078), .A2(n19006), .B1(n19011), .B2(n18966), .ZN(
        n18967) );
  AOI211_X1 U21962 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n19025), .A(n18968), .B(
        n18967), .ZN(n18969) );
  OAI21_X1 U21963 ( .B1(n18970), .B2(n19720), .A(n18969), .ZN(P2_U2846) );
  NAND2_X1 U21964 ( .A1(n13017), .A2(n18971), .ZN(n18973) );
  XOR2_X1 U21965 ( .A(n18973), .B(n18972), .Z(n18980) );
  AOI22_X1 U21966 ( .A1(n18974), .A2(n19030), .B1(P2_REIP_REG_7__SCAN_IN), 
        .B2(n19031), .ZN(n18975) );
  OAI211_X1 U21967 ( .C1(n10786), .C2(n19009), .A(n18975), .B(n18992), .ZN(
        n18978) );
  OAI22_X1 U21968 ( .A1(n19082), .A2(n19006), .B1(n19011), .B2(n18976), .ZN(
        n18977) );
  AOI211_X1 U21969 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19041), .A(
        n18978), .B(n18977), .ZN(n18979) );
  OAI21_X1 U21970 ( .B1(n18980), .B2(n19720), .A(n18979), .ZN(P2_U2848) );
  OAI22_X1 U21971 ( .A1(n18981), .A2(n19008), .B1(n18993), .B2(n19749), .ZN(
        n18982) );
  AOI211_X1 U21972 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n19025), .A(n19155), .B(
        n18982), .ZN(n18990) );
  NOR2_X1 U21973 ( .A1(n13016), .A2(n18983), .ZN(n18984) );
  XNOR2_X1 U21974 ( .A(n18985), .B(n18984), .ZN(n18988) );
  OAI22_X1 U21975 ( .A1(n19084), .A2(n19006), .B1(n19011), .B2(n18986), .ZN(
        n18987) );
  AOI21_X1 U21976 ( .B1(n18988), .B2(n19002), .A(n18987), .ZN(n18989) );
  OAI211_X1 U21977 ( .C1(n9963), .C2(n18991), .A(n18990), .B(n18989), .ZN(
        P2_U2849) );
  OAI21_X1 U21978 ( .B1(n19748), .B2(n18993), .A(n18992), .ZN(n18997) );
  OAI22_X1 U21979 ( .A1(n18995), .A2(n19008), .B1(n19009), .B2(n18994), .ZN(
        n18996) );
  AOI211_X1 U21980 ( .C1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n19041), .A(
        n18997), .B(n18996), .ZN(n19005) );
  NAND2_X1 U21981 ( .A1(n13017), .A2(n18998), .ZN(n18999) );
  XNOR2_X1 U21982 ( .A(n19000), .B(n18999), .ZN(n19003) );
  AOI22_X1 U21983 ( .A1(n19003), .A2(n19002), .B1(n19022), .B2(n19001), .ZN(
        n19004) );
  OAI211_X1 U21984 ( .C1(n19006), .C2(n19094), .A(n19005), .B(n19004), .ZN(
        P2_U2850) );
  OAI22_X1 U21985 ( .A1(n10774), .A2(n19009), .B1(n19008), .B2(n19007), .ZN(
        n19010) );
  AOI211_X1 U21986 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19031), .A(n19155), .B(
        n19010), .ZN(n19021) );
  AOI22_X1 U21987 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19041), .B1(
        n19027), .B2(n19097), .ZN(n19020) );
  OAI22_X1 U21988 ( .A1(n19098), .A2(n19012), .B1(n19011), .B2(n19160), .ZN(
        n19013) );
  INV_X1 U21989 ( .A(n19013), .ZN(n19019) );
  INV_X1 U21990 ( .A(n19164), .ZN(n19017) );
  NOR2_X1 U21991 ( .A1(n13016), .A2(n19014), .ZN(n19016) );
  AOI21_X1 U21992 ( .B1(n19017), .B2(n19016), .A(n19720), .ZN(n19015) );
  OAI21_X1 U21993 ( .B1(n19017), .B2(n19016), .A(n19015), .ZN(n19018) );
  NAND4_X1 U21994 ( .A1(n19021), .A2(n19020), .A3(n19019), .A4(n19018), .ZN(
        P2_U2851) );
  NAND2_X1 U21995 ( .A1(n19023), .A2(n19022), .ZN(n19035) );
  INV_X1 U21996 ( .A(n19024), .ZN(n19026) );
  AOI22_X1 U21997 ( .A1(n19027), .A2(n19026), .B1(P2_EBX_REG_0__SCAN_IN), .B2(
        n19025), .ZN(n19034) );
  INV_X1 U21998 ( .A(n19028), .ZN(n19029) );
  NAND2_X1 U21999 ( .A1(n19030), .A2(n19029), .ZN(n19033) );
  NAND2_X1 U22000 ( .A1(n19031), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n19032) );
  AND4_X1 U22001 ( .A1(n19035), .A2(n19034), .A3(n19033), .A4(n19032), .ZN(
        n19044) );
  INV_X1 U22002 ( .A(n19036), .ZN(n19037) );
  AOI22_X1 U22003 ( .A1(n19231), .A2(n19039), .B1(n19038), .B2(n19037), .ZN(
        n19043) );
  OAI21_X1 U22004 ( .B1(n19041), .B2(n19040), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19042) );
  NAND3_X1 U22005 ( .A1(n19044), .A2(n19043), .A3(n19042), .ZN(P2_U2855) );
  INV_X1 U22006 ( .A(n19045), .ZN(n19046) );
  AOI22_X1 U22007 ( .A1(n19046), .A2(n19111), .B1(n19051), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n19048) );
  AOI22_X1 U22008 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19110), .B1(n19052), 
        .B2(BUF2_REG_31__SCAN_IN), .ZN(n19047) );
  NAND2_X1 U22009 ( .A1(n19048), .A2(n19047), .ZN(P2_U2888) );
  AOI22_X1 U22010 ( .A1(n19050), .A2(n19049), .B1(n19110), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19059) );
  AOI22_X1 U22011 ( .A1(n19052), .A2(BUF2_REG_16__SCAN_IN), .B1(n19051), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19058) );
  OAI22_X1 U22012 ( .A1(n19055), .A2(n19054), .B1(n19115), .B2(n19053), .ZN(
        n19056) );
  INV_X1 U22013 ( .A(n19056), .ZN(n19057) );
  NAND3_X1 U22014 ( .A1(n19059), .A2(n19058), .A3(n19057), .ZN(P2_U2903) );
  INV_X1 U22015 ( .A(n19085), .ZN(n19119) );
  OAI222_X1 U22016 ( .A1(n19061), .A2(n19095), .B1(n13151), .B2(n19083), .C1(
        n19060), .C2(n19119), .ZN(P2_U2904) );
  INV_X1 U22017 ( .A(n19062), .ZN(n19065) );
  AOI22_X1 U22018 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19110), .B1(n19063), 
        .B2(n19085), .ZN(n19064) );
  OAI21_X1 U22019 ( .B1(n19095), .B2(n19065), .A(n19064), .ZN(P2_U2905) );
  INV_X1 U22020 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19125) );
  OAI222_X1 U22021 ( .A1(n19067), .A2(n19095), .B1(n19125), .B2(n19083), .C1(
        n19119), .C2(n19066), .ZN(P2_U2906) );
  INV_X1 U22022 ( .A(n19068), .ZN(n19071) );
  AOI22_X1 U22023 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19110), .B1(n19069), 
        .B2(n19085), .ZN(n19070) );
  OAI21_X1 U22024 ( .B1(n19095), .B2(n19071), .A(n19070), .ZN(P2_U2907) );
  INV_X1 U22025 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19129) );
  OAI222_X1 U22026 ( .A1(n19073), .A2(n19095), .B1(n19129), .B2(n19083), .C1(
        n19119), .C2(n19072), .ZN(P2_U2908) );
  AOI22_X1 U22027 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19110), .B1(n19074), 
        .B2(n19085), .ZN(n19075) );
  OAI21_X1 U22028 ( .B1(n19095), .B2(n19076), .A(n19075), .ZN(P2_U2909) );
  INV_X1 U22029 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19133) );
  OAI222_X1 U22030 ( .A1(n19078), .A2(n19095), .B1(n19133), .B2(n19083), .C1(
        n19119), .C2(n19077), .ZN(P2_U2910) );
  INV_X1 U22031 ( .A(n19079), .ZN(n19081) );
  INV_X1 U22032 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19135) );
  OAI222_X1 U22033 ( .A1(n19081), .A2(n19095), .B1(n19135), .B2(n19083), .C1(
        n19119), .C2(n19080), .ZN(P2_U2911) );
  INV_X1 U22034 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19137) );
  OAI222_X1 U22035 ( .A1(n19082), .A2(n19095), .B1(n19137), .B2(n19083), .C1(
        n19119), .C2(n19225), .ZN(P2_U2912) );
  INV_X1 U22036 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19139) );
  OAI222_X1 U22037 ( .A1(n19084), .A2(n19095), .B1(n19139), .B2(n19083), .C1(
        n19119), .C2(n19214), .ZN(P2_U2913) );
  AOI22_X1 U22038 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19110), .B1(n19086), .B2(
        n19085), .ZN(n19093) );
  AOI21_X1 U22039 ( .B1(n19812), .B2(n19810), .A(n19087), .ZN(n19106) );
  XNOR2_X1 U22040 ( .A(n19235), .B(n19088), .ZN(n19105) );
  NOR2_X1 U22041 ( .A1(n19106), .A2(n19105), .ZN(n19104) );
  NOR2_X1 U22042 ( .A1(n19805), .A2(n19804), .ZN(n19090) );
  OAI21_X1 U22043 ( .B1(n19104), .B2(n19090), .A(n19089), .ZN(n19099) );
  INV_X1 U22044 ( .A(n19098), .ZN(n19091) );
  NAND3_X1 U22045 ( .A1(n19099), .A2(n19091), .A3(n19100), .ZN(n19092) );
  OAI211_X1 U22046 ( .C1(n19095), .C2(n19094), .A(n19093), .B(n19092), .ZN(
        P2_U2914) );
  INV_X1 U22047 ( .A(n19096), .ZN(n19207) );
  AOI22_X1 U22048 ( .A1(n19111), .A2(n19097), .B1(n19110), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19103) );
  XNOR2_X1 U22049 ( .A(n19099), .B(n19098), .ZN(n19101) );
  NAND2_X1 U22050 ( .A1(n19101), .A2(n19100), .ZN(n19102) );
  OAI211_X1 U22051 ( .C1(n19207), .C2(n19119), .A(n19103), .B(n19102), .ZN(
        P2_U2915) );
  AOI22_X1 U22052 ( .A1(n19804), .A2(n19111), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19110), .ZN(n19109) );
  AOI21_X1 U22053 ( .B1(n19106), .B2(n19105), .A(n19104), .ZN(n19107) );
  OR2_X1 U22054 ( .A1(n19107), .A2(n19115), .ZN(n19108) );
  OAI211_X1 U22055 ( .C1(n19202), .C2(n19119), .A(n19109), .B(n19108), .ZN(
        P2_U2916) );
  AOI22_X1 U22056 ( .A1(n19111), .A2(n19826), .B1(n19110), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19118) );
  AOI21_X1 U22057 ( .B1(n19114), .B2(n19113), .A(n19112), .ZN(n19116) );
  OR2_X1 U22058 ( .A1(n19116), .A2(n19115), .ZN(n19117) );
  OAI211_X1 U22059 ( .C1(n19197), .C2(n19119), .A(n19118), .B(n19117), .ZN(
        P2_U2918) );
  NOR2_X1 U22060 ( .A1(n19147), .A2(n19120), .ZN(P2_U2920) );
  AOI22_X1 U22061 ( .A1(n19152), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19121) );
  OAI21_X1 U22062 ( .B1(n13151), .B2(n19154), .A(n19121), .ZN(P2_U2936) );
  AOI22_X1 U22063 ( .A1(n19152), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19122) );
  OAI21_X1 U22064 ( .B1(n19123), .B2(n19154), .A(n19122), .ZN(P2_U2937) );
  AOI22_X1 U22065 ( .A1(n19152), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19124) );
  OAI21_X1 U22066 ( .B1(n19125), .B2(n19154), .A(n19124), .ZN(P2_U2938) );
  AOI22_X1 U22067 ( .A1(n19152), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19126) );
  OAI21_X1 U22068 ( .B1(n19127), .B2(n19154), .A(n19126), .ZN(P2_U2939) );
  AOI22_X1 U22069 ( .A1(n19152), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19128) );
  OAI21_X1 U22070 ( .B1(n19129), .B2(n19154), .A(n19128), .ZN(P2_U2940) );
  AOI22_X1 U22071 ( .A1(n19152), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19130) );
  OAI21_X1 U22072 ( .B1(n19131), .B2(n19154), .A(n19130), .ZN(P2_U2941) );
  AOI22_X1 U22073 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n19151), .B1(n19152), 
        .B2(P2_LWORD_REG_9__SCAN_IN), .ZN(n19132) );
  OAI21_X1 U22074 ( .B1(n19133), .B2(n19154), .A(n19132), .ZN(P2_U2942) );
  AOI22_X1 U22075 ( .A1(n19152), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19134) );
  OAI21_X1 U22076 ( .B1(n19135), .B2(n19154), .A(n19134), .ZN(P2_U2943) );
  AOI22_X1 U22077 ( .A1(n19152), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19136) );
  OAI21_X1 U22078 ( .B1(n19137), .B2(n19154), .A(n19136), .ZN(P2_U2944) );
  AOI22_X1 U22079 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n19151), .B1(n19152), 
        .B2(P2_LWORD_REG_6__SCAN_IN), .ZN(n19138) );
  OAI21_X1 U22080 ( .B1(n19139), .B2(n19154), .A(n19138), .ZN(P2_U2945) );
  INV_X1 U22081 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19141) );
  AOI22_X1 U22082 ( .A1(n19152), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19140) );
  OAI21_X1 U22083 ( .B1(n19141), .B2(n19154), .A(n19140), .ZN(P2_U2946) );
  INV_X1 U22084 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19143) );
  AOI22_X1 U22085 ( .A1(n19152), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19142) );
  OAI21_X1 U22086 ( .B1(n19143), .B2(n19154), .A(n19142), .ZN(P2_U2947) );
  AOI22_X1 U22087 ( .A1(P2_EAX_REG_3__SCAN_IN), .A2(n19144), .B1(n19152), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n19145) );
  OAI21_X1 U22088 ( .B1(n20838), .B2(n19147), .A(n19145), .ZN(P2_U2948) );
  INV_X1 U22089 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n20850) );
  INV_X1 U22090 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19148) );
  OAI222_X1 U22091 ( .A1(n19864), .A2(n20850), .B1(n19154), .B2(n19148), .C1(
        n19147), .C2(n19146), .ZN(P2_U2949) );
  INV_X1 U22092 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19150) );
  AOI22_X1 U22093 ( .A1(n19152), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19149) );
  OAI21_X1 U22094 ( .B1(n19150), .B2(n19154), .A(n19149), .ZN(P2_U2950) );
  AOI22_X1 U22095 ( .A1(n19152), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19151), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19153) );
  OAI21_X1 U22096 ( .B1(n13263), .B2(n19154), .A(n19153), .ZN(P2_U2951) );
  AOI22_X1 U22097 ( .A1(n19166), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19155), .ZN(n19163) );
  NAND2_X1 U22098 ( .A1(n19156), .A2(n19169), .ZN(n19159) );
  NAND2_X1 U22099 ( .A1(n19157), .A2(n19167), .ZN(n19158) );
  OAI211_X1 U22100 ( .C1(n19179), .C2(n19160), .A(n19159), .B(n19158), .ZN(
        n19161) );
  INV_X1 U22101 ( .A(n19161), .ZN(n19162) );
  OAI211_X1 U22102 ( .C1(n19165), .C2(n19164), .A(n19163), .B(n19162), .ZN(
        P2_U3010) );
  AOI22_X1 U22103 ( .A1(n19168), .A2(n19167), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19166), .ZN(n19182) );
  NAND2_X1 U22104 ( .A1(n19170), .A2(n19169), .ZN(n19177) );
  INV_X1 U22105 ( .A(n19171), .ZN(n19174) );
  INV_X1 U22106 ( .A(n19172), .ZN(n19173) );
  AOI21_X1 U22107 ( .B1(n19175), .B2(n19174), .A(n19173), .ZN(n19176) );
  OAI211_X1 U22108 ( .C1(n19179), .C2(n19178), .A(n19177), .B(n19176), .ZN(
        n19180) );
  INV_X1 U22109 ( .A(n19180), .ZN(n19181) );
  NAND2_X1 U22110 ( .A1(n19182), .A2(n19181), .ZN(P2_U3012) );
  NAND2_X1 U22111 ( .A1(n19184), .A2(n19652), .ZN(n19680) );
  NAND2_X1 U22112 ( .A1(n16335), .A2(n19819), .ZN(n19288) );
  NOR2_X1 U22113 ( .A1(n19445), .A2(n19288), .ZN(n19224) );
  AOI22_X1 U22114 ( .A1(n19658), .A2(n19705), .B1(n19649), .B2(n19224), .ZN(
        n19195) );
  OAI21_X1 U22115 ( .B1(n19705), .B2(n19256), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19185) );
  NAND2_X1 U22116 ( .A1(n19185), .A2(n19802), .ZN(n19193) );
  NOR2_X1 U22117 ( .A1(n19186), .A2(n16335), .ZN(n19701) );
  NOR2_X1 U22118 ( .A1(n19701), .A2(n19224), .ZN(n19192) );
  INV_X1 U22119 ( .A(n19192), .ZN(n19190) );
  INV_X1 U22120 ( .A(n19224), .ZN(n19187) );
  OAI211_X1 U22121 ( .C1(n19188), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19187), 
        .B(n19609), .ZN(n19189) );
  OAI211_X1 U22122 ( .C1(n19193), .C2(n19190), .A(n19656), .B(n19189), .ZN(
        n19227) );
  OAI21_X1 U22123 ( .B1(n10403), .B2(n19224), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19191) );
  AOI22_X1 U22124 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19227), .B1(
        n19650), .B2(n19226), .ZN(n19194) );
  OAI211_X1 U22125 ( .C1(n19661), .C2(n19230), .A(n19195), .B(n19194), .ZN(
        P2_U3048) );
  AOI22_X1 U22126 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19222), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19221), .ZN(n19667) );
  AOI22_X1 U22127 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19221), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19222), .ZN(n19624) );
  INV_X1 U22128 ( .A(n19624), .ZN(n19664) );
  AOI22_X1 U22129 ( .A1(n19664), .A2(n19705), .B1(n19662), .B2(n19224), .ZN(
        n19199) );
  NOR2_X2 U22130 ( .A1(n19197), .A2(n19421), .ZN(n19663) );
  AOI22_X1 U22131 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19227), .B1(
        n19663), .B2(n19226), .ZN(n19198) );
  OAI211_X1 U22132 ( .C1(n19667), .C2(n19230), .A(n19199), .B(n19198), .ZN(
        P2_U3049) );
  AOI22_X1 U22133 ( .A1(n19670), .A2(n19705), .B1(n19668), .B2(n19224), .ZN(
        n19201) );
  AOI22_X1 U22134 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19227), .B1(
        n19669), .B2(n19226), .ZN(n19200) );
  OAI211_X1 U22135 ( .C1(n19673), .C2(n19230), .A(n19201), .B(n19200), .ZN(
        P2_U3050) );
  AOI22_X1 U22136 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19222), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19221), .ZN(n19681) );
  AOI22_X1 U22137 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19221), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19222), .ZN(n19630) );
  INV_X1 U22138 ( .A(n19630), .ZN(n19676) );
  AOI22_X1 U22139 ( .A1(n19676), .A2(n19705), .B1(n9562), .B2(n19224), .ZN(
        n19204) );
  NOR2_X2 U22140 ( .A1(n19202), .A2(n19421), .ZN(n19675) );
  AOI22_X1 U22141 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19227), .B1(
        n19675), .B2(n19226), .ZN(n19203) );
  OAI211_X1 U22142 ( .C1(n19681), .C2(n19230), .A(n19204), .B(n19203), .ZN(
        P2_U3051) );
  AOI22_X1 U22143 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19222), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19221), .ZN(n19687) );
  INV_X1 U22144 ( .A(n19687), .ZN(n19587) );
  NOR2_X2 U22145 ( .A1(n19206), .A2(n19205), .ZN(n19682) );
  AOI22_X1 U22146 ( .A1(n19587), .A2(n19705), .B1(n19682), .B2(n19224), .ZN(
        n19209) );
  NOR2_X2 U22147 ( .A1(n19207), .A2(n19421), .ZN(n19683) );
  AOI22_X1 U22148 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19227), .B1(
        n19683), .B2(n19226), .ZN(n19208) );
  OAI211_X1 U22149 ( .C1(n19590), .C2(n19230), .A(n19209), .B(n19208), .ZN(
        P2_U3052) );
  AOI22_X1 U22150 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19222), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19221), .ZN(n19693) );
  AOI22_X1 U22151 ( .A1(n19634), .A2(n19705), .B1(n19688), .B2(n19224), .ZN(
        n19212) );
  NOR2_X2 U22152 ( .A1(n19210), .A2(n19421), .ZN(n19689) );
  AOI22_X1 U22153 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19227), .B1(
        n19689), .B2(n19226), .ZN(n19211) );
  OAI211_X1 U22154 ( .C1(n19637), .C2(n19230), .A(n19212), .B(n19211), .ZN(
        P2_U3053) );
  AOI22_X1 U22155 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19221), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19222), .ZN(n19699) );
  INV_X1 U22156 ( .A(n19699), .ZN(n19594) );
  AND2_X1 U22157 ( .A1(n19213), .A2(n19223), .ZN(n19694) );
  AOI22_X1 U22158 ( .A1(n19594), .A2(n19705), .B1(n19694), .B2(n19224), .ZN(
        n19216) );
  NOR2_X2 U22159 ( .A1(n19214), .A2(n19421), .ZN(n19695) );
  AOI22_X1 U22160 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19227), .B1(
        n19695), .B2(n19226), .ZN(n19215) );
  OAI211_X1 U22161 ( .C1(n19538), .C2(n19230), .A(n19216), .B(n19215), .ZN(
        P2_U3054) );
  AOI22_X1 U22162 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19222), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19221), .ZN(n19710) );
  INV_X1 U22163 ( .A(n19710), .ZN(n19598) );
  AND2_X1 U22164 ( .A1(n9583), .A2(n19223), .ZN(n19700) );
  AOI22_X1 U22165 ( .A1(n19598), .A2(n19705), .B1(n19700), .B2(n19224), .ZN(
        n19229) );
  NOR2_X2 U22166 ( .A1(n19225), .A2(n19421), .ZN(n19702) );
  AOI22_X1 U22167 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19227), .B1(
        n19702), .B2(n19226), .ZN(n19228) );
  OAI211_X1 U22168 ( .C1(n19545), .C2(n19230), .A(n19229), .B(n19228), .ZN(
        P2_U3055) );
  OR2_X1 U22169 ( .A1(n19288), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19236) );
  INV_X1 U22170 ( .A(n10399), .ZN(n19233) );
  NOR2_X1 U22171 ( .A1(n19837), .A2(n19236), .ZN(n19254) );
  OAI21_X1 U22172 ( .B1(n19233), .B2(n19254), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19234) );
  OAI21_X1 U22173 ( .B1(n19236), .B2(n19609), .A(n19234), .ZN(n19255) );
  AOI22_X1 U22174 ( .A1(n19255), .A2(n19650), .B1(n19649), .B2(n19254), .ZN(
        n19241) );
  AOI21_X1 U22175 ( .B1(n10399), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19239) );
  NAND2_X1 U22176 ( .A1(n19235), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19420) );
  OAI21_X1 U22177 ( .B1(n19420), .B2(n19237), .A(n19236), .ZN(n19238) );
  OAI211_X1 U22178 ( .C1(n19254), .C2(n19239), .A(n19238), .B(n19656), .ZN(
        n19257) );
  AOI22_X1 U22179 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19257), .B1(
        n19256), .B2(n19658), .ZN(n19240) );
  OAI211_X1 U22180 ( .C1(n19661), .C2(n19287), .A(n19241), .B(n19240), .ZN(
        P2_U3056) );
  AOI22_X1 U22181 ( .A1(n19255), .A2(n19663), .B1(n19662), .B2(n19254), .ZN(
        n19243) );
  AOI22_X1 U22182 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19257), .B1(
        n19256), .B2(n19664), .ZN(n19242) );
  OAI211_X1 U22183 ( .C1(n19667), .C2(n19287), .A(n19243), .B(n19242), .ZN(
        P2_U3057) );
  AOI22_X1 U22184 ( .A1(n19255), .A2(n19669), .B1(n19668), .B2(n19254), .ZN(
        n19245) );
  AOI22_X1 U22185 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19257), .B1(
        n19256), .B2(n19670), .ZN(n19244) );
  OAI211_X1 U22186 ( .C1(n19673), .C2(n19287), .A(n19245), .B(n19244), .ZN(
        P2_U3058) );
  AOI22_X1 U22187 ( .A1(n19255), .A2(n19675), .B1(n9562), .B2(n19254), .ZN(
        n19247) );
  AOI22_X1 U22188 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19257), .B1(
        n19256), .B2(n19676), .ZN(n19246) );
  OAI211_X1 U22189 ( .C1(n19681), .C2(n19287), .A(n19247), .B(n19246), .ZN(
        P2_U3059) );
  AOI22_X1 U22190 ( .A1(n19255), .A2(n19683), .B1(n19682), .B2(n19254), .ZN(
        n19249) );
  AOI22_X1 U22191 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19257), .B1(
        n19256), .B2(n19587), .ZN(n19248) );
  OAI211_X1 U22192 ( .C1(n19590), .C2(n19287), .A(n19249), .B(n19248), .ZN(
        P2_U3060) );
  AOI22_X1 U22193 ( .A1(n19255), .A2(n19689), .B1(n19688), .B2(n19254), .ZN(
        n19251) );
  AOI22_X1 U22194 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19257), .B1(
        n19256), .B2(n19634), .ZN(n19250) );
  OAI211_X1 U22195 ( .C1(n19637), .C2(n19287), .A(n19251), .B(n19250), .ZN(
        P2_U3061) );
  AOI22_X1 U22196 ( .A1(n19255), .A2(n19695), .B1(n19694), .B2(n19254), .ZN(
        n19253) );
  AOI22_X1 U22197 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19257), .B1(
        n19256), .B2(n19594), .ZN(n19252) );
  OAI211_X1 U22198 ( .C1(n19538), .C2(n19287), .A(n19253), .B(n19252), .ZN(
        P2_U3062) );
  AOI22_X1 U22199 ( .A1(n19255), .A2(n19702), .B1(n19700), .B2(n19254), .ZN(
        n19259) );
  AOI22_X1 U22200 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19257), .B1(
        n19256), .B2(n19598), .ZN(n19258) );
  OAI211_X1 U22201 ( .C1(n19545), .C2(n19287), .A(n19259), .B(n19258), .ZN(
        P2_U3063) );
  NOR2_X1 U22202 ( .A1(n19828), .A2(n19288), .ZN(n19291) );
  INV_X1 U22203 ( .A(n19291), .ZN(n19296) );
  NOR2_X1 U22204 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19296), .ZN(
        n19282) );
  OAI21_X1 U22205 ( .B1(n19262), .B2(n19282), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19261) );
  NOR2_X1 U22206 ( .A1(n19496), .A2(n19288), .ZN(n19263) );
  INV_X1 U22207 ( .A(n19263), .ZN(n19260) );
  NAND2_X1 U22208 ( .A1(n19261), .A2(n19260), .ZN(n19283) );
  AOI22_X1 U22209 ( .A1(n19283), .A2(n19650), .B1(n19649), .B2(n19282), .ZN(
        n19269) );
  AOI21_X1 U22210 ( .B1(n19262), .B2(n10900), .A(n19282), .ZN(n19266) );
  AOI21_X1 U22211 ( .B1(n19318), .B2(n19287), .A(n19446), .ZN(n19264) );
  NOR2_X1 U22212 ( .A1(n19264), .A2(n19263), .ZN(n19265) );
  MUX2_X1 U22213 ( .A(n19266), .B(n19265), .S(n19802), .Z(n19267) );
  AOI22_X1 U22214 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19284), .B1(
        n19308), .B2(n19606), .ZN(n19268) );
  OAI211_X1 U22215 ( .C1(n19620), .C2(n19287), .A(n19269), .B(n19268), .ZN(
        P2_U3064) );
  AOI22_X1 U22216 ( .A1(n19283), .A2(n19663), .B1(n19662), .B2(n19282), .ZN(
        n19271) );
  INV_X1 U22217 ( .A(n19667), .ZN(n19621) );
  AOI22_X1 U22218 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19284), .B1(
        n19308), .B2(n19621), .ZN(n19270) );
  OAI211_X1 U22219 ( .C1(n19624), .C2(n19287), .A(n19271), .B(n19270), .ZN(
        P2_U3065) );
  AOI22_X1 U22220 ( .A1(n19283), .A2(n19669), .B1(n19668), .B2(n19282), .ZN(
        n19273) );
  AOI22_X1 U22221 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19284), .B1(
        n19308), .B2(n19562), .ZN(n19272) );
  OAI211_X1 U22222 ( .C1(n19565), .C2(n19287), .A(n19273), .B(n19272), .ZN(
        P2_U3066) );
  AOI22_X1 U22223 ( .A1(n19283), .A2(n19675), .B1(n9562), .B2(n19282), .ZN(
        n19275) );
  INV_X1 U22224 ( .A(n19681), .ZN(n19627) );
  AOI22_X1 U22225 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19284), .B1(
        n19308), .B2(n19627), .ZN(n19274) );
  OAI211_X1 U22226 ( .C1(n19630), .C2(n19287), .A(n19275), .B(n19274), .ZN(
        P2_U3067) );
  AOI22_X1 U22227 ( .A1(n19283), .A2(n19683), .B1(n19682), .B2(n19282), .ZN(
        n19277) );
  AOI22_X1 U22228 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19284), .B1(
        n19308), .B2(n19684), .ZN(n19276) );
  OAI211_X1 U22229 ( .C1(n19687), .C2(n19287), .A(n19277), .B(n19276), .ZN(
        P2_U3068) );
  AOI22_X1 U22230 ( .A1(n19283), .A2(n19689), .B1(n19688), .B2(n19282), .ZN(
        n19279) );
  INV_X1 U22231 ( .A(n19637), .ZN(n19690) );
  AOI22_X1 U22232 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19284), .B1(
        n19308), .B2(n19690), .ZN(n19278) );
  OAI211_X1 U22233 ( .C1(n19693), .C2(n19287), .A(n19279), .B(n19278), .ZN(
        P2_U3069) );
  AOI22_X1 U22234 ( .A1(n19283), .A2(n19695), .B1(n19694), .B2(n19282), .ZN(
        n19281) );
  AOI22_X1 U22235 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19284), .B1(
        n19308), .B2(n19696), .ZN(n19280) );
  OAI211_X1 U22236 ( .C1(n19699), .C2(n19287), .A(n19281), .B(n19280), .ZN(
        P2_U3070) );
  AOI22_X1 U22237 ( .A1(n19283), .A2(n19702), .B1(n19700), .B2(n19282), .ZN(
        n19286) );
  AOI22_X1 U22238 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19284), .B1(
        n19308), .B2(n19704), .ZN(n19285) );
  OAI211_X1 U22239 ( .C1(n19710), .C2(n19287), .A(n19286), .B(n19285), .ZN(
        P2_U3071) );
  INV_X1 U22240 ( .A(n19288), .ZN(n19289) );
  AND2_X1 U22241 ( .A1(n19388), .A2(n19289), .ZN(n19313) );
  AOI22_X1 U22242 ( .A1(n19658), .A2(n19308), .B1(n19649), .B2(n19313), .ZN(
        n19299) );
  OAI21_X1 U22243 ( .B1(n19420), .B2(n19290), .A(n19802), .ZN(n19297) );
  NOR2_X1 U22244 ( .A1(n19297), .A2(n19291), .ZN(n19292) );
  OAI21_X1 U22245 ( .B1(n19293), .B2(n19313), .A(n19656), .ZN(n19315) );
  OAI21_X1 U22246 ( .B1(n19294), .B2(n19313), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19295) );
  OAI21_X1 U22247 ( .B1(n19297), .B2(n19296), .A(n19295), .ZN(n19314) );
  AOI22_X1 U22248 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19315), .B1(
        n19650), .B2(n19314), .ZN(n19298) );
  OAI211_X1 U22249 ( .C1(n19661), .C2(n19326), .A(n19299), .B(n19298), .ZN(
        P2_U3072) );
  AOI22_X1 U22250 ( .A1(n19621), .A2(n19348), .B1(n19313), .B2(n19662), .ZN(
        n19301) );
  AOI22_X1 U22251 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19315), .B1(
        n19663), .B2(n19314), .ZN(n19300) );
  OAI211_X1 U22252 ( .C1(n19624), .C2(n19318), .A(n19301), .B(n19300), .ZN(
        P2_U3073) );
  AOI22_X1 U22253 ( .A1(n19562), .A2(n19348), .B1(n19668), .B2(n19313), .ZN(
        n19303) );
  AOI22_X1 U22254 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19315), .B1(
        n19669), .B2(n19314), .ZN(n19302) );
  OAI211_X1 U22255 ( .C1(n19565), .C2(n19318), .A(n19303), .B(n19302), .ZN(
        P2_U3074) );
  AOI22_X1 U22256 ( .A1(n19627), .A2(n19348), .B1(n19313), .B2(n9562), .ZN(
        n19305) );
  AOI22_X1 U22257 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19315), .B1(
        n19675), .B2(n19314), .ZN(n19304) );
  OAI211_X1 U22258 ( .C1(n19630), .C2(n19318), .A(n19305), .B(n19304), .ZN(
        P2_U3075) );
  AOI22_X1 U22259 ( .A1(n19587), .A2(n19308), .B1(n19313), .B2(n19682), .ZN(
        n19307) );
  AOI22_X1 U22260 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19315), .B1(
        n19683), .B2(n19314), .ZN(n19306) );
  OAI211_X1 U22261 ( .C1(n19590), .C2(n19326), .A(n19307), .B(n19306), .ZN(
        P2_U3076) );
  AOI22_X1 U22262 ( .A1(n19634), .A2(n19308), .B1(n19313), .B2(n19688), .ZN(
        n19310) );
  AOI22_X1 U22263 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19315), .B1(
        n19689), .B2(n19314), .ZN(n19309) );
  OAI211_X1 U22264 ( .C1(n19637), .C2(n19326), .A(n19310), .B(n19309), .ZN(
        P2_U3077) );
  AOI22_X1 U22265 ( .A1(n19696), .A2(n19348), .B1(n19313), .B2(n19694), .ZN(
        n19312) );
  AOI22_X1 U22266 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19315), .B1(
        n19695), .B2(n19314), .ZN(n19311) );
  OAI211_X1 U22267 ( .C1(n19699), .C2(n19318), .A(n19312), .B(n19311), .ZN(
        P2_U3078) );
  AOI22_X1 U22268 ( .A1(n19704), .A2(n19348), .B1(n19313), .B2(n19700), .ZN(
        n19317) );
  AOI22_X1 U22269 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19315), .B1(
        n19702), .B2(n19314), .ZN(n19316) );
  OAI211_X1 U22270 ( .C1(n19710), .C2(n19318), .A(n19317), .B(n19316), .ZN(
        P2_U3079) );
  OR2_X1 U22271 ( .A1(n19321), .A2(n19320), .ZN(n19553) );
  NOR2_X1 U22272 ( .A1(n19553), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19331) );
  INV_X1 U22273 ( .A(n19331), .ZN(n19325) );
  AND2_X1 U22274 ( .A1(n19390), .A2(n19322), .ZN(n19346) );
  OAI21_X1 U22275 ( .B1(n19323), .B2(n19346), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19324) );
  OAI21_X1 U22276 ( .B1(n19609), .B2(n19325), .A(n19324), .ZN(n19347) );
  AOI22_X1 U22277 ( .A1(n19347), .A2(n19650), .B1(n19649), .B2(n19346), .ZN(
        n19333) );
  AOI21_X1 U22278 ( .B1(n19326), .B2(n19372), .A(n19446), .ZN(n19330) );
  INV_X1 U22279 ( .A(n19346), .ZN(n19327) );
  OAI211_X1 U22280 ( .C1(n19328), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19327), 
        .B(n19609), .ZN(n19329) );
  OAI211_X1 U22281 ( .C1(n19331), .C2(n19330), .A(n19329), .B(n19656), .ZN(
        n19349) );
  AOI22_X1 U22282 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19349), .B1(
        n19348), .B2(n19658), .ZN(n19332) );
  OAI211_X1 U22283 ( .C1(n19661), .C2(n19372), .A(n19333), .B(n19332), .ZN(
        P2_U3080) );
  AOI22_X1 U22284 ( .A1(n19347), .A2(n19663), .B1(n19662), .B2(n19346), .ZN(
        n19335) );
  AOI22_X1 U22285 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19349), .B1(
        n19348), .B2(n19664), .ZN(n19334) );
  OAI211_X1 U22286 ( .C1(n19667), .C2(n19372), .A(n19335), .B(n19334), .ZN(
        P2_U3081) );
  AOI22_X1 U22287 ( .A1(n19347), .A2(n19669), .B1(n19668), .B2(n19346), .ZN(
        n19337) );
  AOI22_X1 U22288 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19349), .B1(
        n19348), .B2(n19670), .ZN(n19336) );
  OAI211_X1 U22289 ( .C1(n19673), .C2(n19372), .A(n19337), .B(n19336), .ZN(
        P2_U3082) );
  AOI22_X1 U22290 ( .A1(n19347), .A2(n19675), .B1(n9562), .B2(n19346), .ZN(
        n19339) );
  AOI22_X1 U22291 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19349), .B1(
        n19348), .B2(n19676), .ZN(n19338) );
  OAI211_X1 U22292 ( .C1(n19681), .C2(n19372), .A(n19339), .B(n19338), .ZN(
        P2_U3083) );
  AOI22_X1 U22293 ( .A1(n19347), .A2(n19683), .B1(n19682), .B2(n19346), .ZN(
        n19341) );
  AOI22_X1 U22294 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19349), .B1(
        n19348), .B2(n19587), .ZN(n19340) );
  OAI211_X1 U22295 ( .C1(n19590), .C2(n19372), .A(n19341), .B(n19340), .ZN(
        P2_U3084) );
  AOI22_X1 U22296 ( .A1(n19347), .A2(n19689), .B1(n19688), .B2(n19346), .ZN(
        n19343) );
  AOI22_X1 U22297 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19349), .B1(
        n19348), .B2(n19634), .ZN(n19342) );
  OAI211_X1 U22298 ( .C1(n19637), .C2(n19372), .A(n19343), .B(n19342), .ZN(
        P2_U3085) );
  AOI22_X1 U22299 ( .A1(n19347), .A2(n19695), .B1(n19694), .B2(n19346), .ZN(
        n19345) );
  AOI22_X1 U22300 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19349), .B1(
        n19348), .B2(n19594), .ZN(n19344) );
  OAI211_X1 U22301 ( .C1(n19538), .C2(n19372), .A(n19345), .B(n19344), .ZN(
        P2_U3086) );
  AOI22_X1 U22302 ( .A1(n19347), .A2(n19702), .B1(n19700), .B2(n19346), .ZN(
        n19351) );
  AOI22_X1 U22303 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19349), .B1(
        n19348), .B2(n19598), .ZN(n19350) );
  OAI211_X1 U22304 ( .C1(n19545), .C2(n19372), .A(n19351), .B(n19350), .ZN(
        P2_U3087) );
  AND3_X1 U22305 ( .A1(n19828), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(
        n19390), .ZN(n19377) );
  AOI22_X1 U22306 ( .A1(n19606), .A2(n19411), .B1(n19649), .B2(n19377), .ZN(
        n19363) );
  OAI21_X1 U22307 ( .B1(n19420), .B2(n19353), .A(n19802), .ZN(n19361) );
  NAND2_X1 U22308 ( .A1(n19828), .A2(n19390), .ZN(n19360) );
  INV_X1 U22309 ( .A(n19360), .ZN(n19356) );
  INV_X1 U22310 ( .A(n19377), .ZN(n19354) );
  OAI211_X1 U22311 ( .C1(n19357), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19354), 
        .B(n19609), .ZN(n19355) );
  OAI211_X1 U22312 ( .C1(n19361), .C2(n19356), .A(n19656), .B(n19355), .ZN(
        n19380) );
  INV_X1 U22313 ( .A(n19357), .ZN(n19358) );
  OAI21_X1 U22314 ( .B1(n19358), .B2(n19377), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19359) );
  OAI21_X1 U22315 ( .B1(n19361), .B2(n19360), .A(n19359), .ZN(n19379) );
  AOI22_X1 U22316 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19380), .B1(
        n19650), .B2(n19379), .ZN(n19362) );
  OAI211_X1 U22317 ( .C1(n19620), .C2(n19372), .A(n19363), .B(n19362), .ZN(
        P2_U3088) );
  AOI22_X1 U22318 ( .A1(n19621), .A2(n19411), .B1(n19377), .B2(n19662), .ZN(
        n19365) );
  AOI22_X1 U22319 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19380), .B1(
        n19663), .B2(n19379), .ZN(n19364) );
  OAI211_X1 U22320 ( .C1(n19624), .C2(n19372), .A(n19365), .B(n19364), .ZN(
        P2_U3089) );
  INV_X1 U22321 ( .A(n19372), .ZN(n19378) );
  AOI22_X1 U22322 ( .A1(n19670), .A2(n19378), .B1(n19668), .B2(n19377), .ZN(
        n19367) );
  AOI22_X1 U22323 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19380), .B1(
        n19669), .B2(n19379), .ZN(n19366) );
  OAI211_X1 U22324 ( .C1(n19673), .C2(n19392), .A(n19367), .B(n19366), .ZN(
        P2_U3090) );
  AOI22_X1 U22325 ( .A1(n19676), .A2(n19378), .B1(n19377), .B2(n9562), .ZN(
        n19369) );
  AOI22_X1 U22326 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19380), .B1(
        n19675), .B2(n19379), .ZN(n19368) );
  OAI211_X1 U22327 ( .C1(n19681), .C2(n19392), .A(n19369), .B(n19368), .ZN(
        P2_U3091) );
  AOI22_X1 U22328 ( .A1(n19684), .A2(n19411), .B1(n19377), .B2(n19682), .ZN(
        n19371) );
  AOI22_X1 U22329 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19380), .B1(
        n19683), .B2(n19379), .ZN(n19370) );
  OAI211_X1 U22330 ( .C1(n19687), .C2(n19372), .A(n19371), .B(n19370), .ZN(
        P2_U3092) );
  AOI22_X1 U22331 ( .A1(n19634), .A2(n19378), .B1(n19377), .B2(n19688), .ZN(
        n19374) );
  AOI22_X1 U22332 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19380), .B1(
        n19689), .B2(n19379), .ZN(n19373) );
  OAI211_X1 U22333 ( .C1(n19637), .C2(n19392), .A(n19374), .B(n19373), .ZN(
        P2_U3093) );
  AOI22_X1 U22334 ( .A1(n19594), .A2(n19378), .B1(n19377), .B2(n19694), .ZN(
        n19376) );
  AOI22_X1 U22335 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19380), .B1(
        n19695), .B2(n19379), .ZN(n19375) );
  OAI211_X1 U22336 ( .C1(n19538), .C2(n19392), .A(n19376), .B(n19375), .ZN(
        P2_U3094) );
  AOI22_X1 U22337 ( .A1(n19598), .A2(n19378), .B1(n19377), .B2(n19700), .ZN(
        n19382) );
  AOI22_X1 U22338 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19380), .B1(
        n19702), .B2(n19379), .ZN(n19381) );
  OAI211_X1 U22339 ( .C1(n19545), .C2(n19392), .A(n19382), .B(n19381), .ZN(
        P2_U3095) );
  INV_X1 U22340 ( .A(n19390), .ZN(n19385) );
  NAND2_X1 U22341 ( .A1(n19605), .A2(n16335), .ZN(n19423) );
  NOR2_X1 U22342 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19423), .ZN(
        n19409) );
  OAI21_X1 U22343 ( .B1(n19386), .B2(n19409), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19384) );
  OAI21_X1 U22344 ( .B1(n19496), .B2(n19385), .A(n19384), .ZN(n19410) );
  AOI22_X1 U22345 ( .A1(n19410), .A2(n19650), .B1(n19649), .B2(n19409), .ZN(
        n19396) );
  INV_X1 U22346 ( .A(n19386), .ZN(n19387) );
  AOI21_X1 U22347 ( .B1(n19387), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19394) );
  INV_X1 U22348 ( .A(n19388), .ZN(n19389) );
  NAND3_X1 U22349 ( .A1(n19390), .A2(n19445), .A3(n19389), .ZN(n19391) );
  OAI221_X1 U22350 ( .B1(n19446), .B2(n19392), .C1(n19446), .C2(n19415), .A(
        n19391), .ZN(n19393) );
  OAI211_X1 U22351 ( .C1(n19394), .C2(n19409), .A(n19656), .B(n19393), .ZN(
        n19412) );
  AOI22_X1 U22352 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19658), .ZN(n19395) );
  OAI211_X1 U22353 ( .C1(n19661), .C2(n19415), .A(n19396), .B(n19395), .ZN(
        P2_U3096) );
  AOI22_X1 U22354 ( .A1(n19410), .A2(n19663), .B1(n19662), .B2(n19409), .ZN(
        n19398) );
  AOI22_X1 U22355 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19664), .ZN(n19397) );
  OAI211_X1 U22356 ( .C1(n19667), .C2(n19415), .A(n19398), .B(n19397), .ZN(
        P2_U3097) );
  AOI22_X1 U22357 ( .A1(n19410), .A2(n19669), .B1(n19668), .B2(n19409), .ZN(
        n19400) );
  AOI22_X1 U22358 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19670), .ZN(n19399) );
  OAI211_X1 U22359 ( .C1(n19673), .C2(n19415), .A(n19400), .B(n19399), .ZN(
        P2_U3098) );
  AOI22_X1 U22360 ( .A1(n19410), .A2(n19675), .B1(n9562), .B2(n19409), .ZN(
        n19402) );
  AOI22_X1 U22361 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19676), .ZN(n19401) );
  OAI211_X1 U22362 ( .C1(n19681), .C2(n19415), .A(n19402), .B(n19401), .ZN(
        P2_U3099) );
  AOI22_X1 U22363 ( .A1(n19410), .A2(n19683), .B1(n19682), .B2(n19409), .ZN(
        n19404) );
  AOI22_X1 U22364 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19587), .ZN(n19403) );
  OAI211_X1 U22365 ( .C1(n19590), .C2(n19415), .A(n19404), .B(n19403), .ZN(
        P2_U3100) );
  AOI22_X1 U22366 ( .A1(n19410), .A2(n19689), .B1(n19688), .B2(n19409), .ZN(
        n19406) );
  AOI22_X1 U22367 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19634), .ZN(n19405) );
  OAI211_X1 U22368 ( .C1(n19637), .C2(n19415), .A(n19406), .B(n19405), .ZN(
        P2_U3101) );
  AOI22_X1 U22369 ( .A1(n19410), .A2(n19695), .B1(n19694), .B2(n19409), .ZN(
        n19408) );
  AOI22_X1 U22370 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19594), .ZN(n19407) );
  OAI211_X1 U22371 ( .C1(n19538), .C2(n19415), .A(n19408), .B(n19407), .ZN(
        P2_U3102) );
  AOI22_X1 U22372 ( .A1(n19410), .A2(n19702), .B1(n19700), .B2(n19409), .ZN(
        n19414) );
  AOI22_X1 U22373 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19598), .ZN(n19413) );
  OAI211_X1 U22374 ( .C1(n19545), .C2(n19415), .A(n19414), .B(n19413), .ZN(
        P2_U3103) );
  INV_X1 U22375 ( .A(n10398), .ZN(n19417) );
  NOR3_X1 U22376 ( .A1(n19417), .A2(n19452), .A3(n19860), .ZN(n19422) );
  INV_X1 U22377 ( .A(n19423), .ZN(n19418) );
  AOI21_X1 U22378 ( .B1(n10900), .B2(n19418), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19419) );
  NOR2_X1 U22379 ( .A1(n19422), .A2(n19419), .ZN(n19440) );
  AOI22_X1 U22380 ( .A1(n19440), .A2(n19650), .B1(n19452), .B2(n19649), .ZN(
        n19427) );
  NOR2_X1 U22381 ( .A1(n19420), .A2(n19603), .ZN(n19799) );
  INV_X1 U22382 ( .A(n19799), .ZN(n19424) );
  AOI211_X1 U22383 ( .C1(n19424), .C2(n19423), .A(n19422), .B(n19421), .ZN(
        n19425) );
  OAI21_X1 U22384 ( .B1(n19452), .B2(n10900), .A(n19425), .ZN(n19442) );
  AOI22_X1 U22385 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19658), .ZN(n19426) );
  OAI211_X1 U22386 ( .C1(n19661), .C2(n19475), .A(n19427), .B(n19426), .ZN(
        P2_U3104) );
  AOI22_X1 U22387 ( .A1(n19440), .A2(n19663), .B1(n19452), .B2(n19662), .ZN(
        n19429) );
  AOI22_X1 U22388 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19664), .ZN(n19428) );
  OAI211_X1 U22389 ( .C1(n19667), .C2(n19475), .A(n19429), .B(n19428), .ZN(
        P2_U3105) );
  AOI22_X1 U22390 ( .A1(n19440), .A2(n19669), .B1(n19452), .B2(n19668), .ZN(
        n19431) );
  AOI22_X1 U22391 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19670), .ZN(n19430) );
  OAI211_X1 U22392 ( .C1(n19673), .C2(n19475), .A(n19431), .B(n19430), .ZN(
        P2_U3106) );
  AOI22_X1 U22393 ( .A1(n19440), .A2(n19675), .B1(n19452), .B2(n9562), .ZN(
        n19433) );
  AOI22_X1 U22394 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19676), .ZN(n19432) );
  OAI211_X1 U22395 ( .C1(n19681), .C2(n19475), .A(n19433), .B(n19432), .ZN(
        P2_U3107) );
  AOI22_X1 U22396 ( .A1(n19440), .A2(n19683), .B1(n19452), .B2(n19682), .ZN(
        n19435) );
  AOI22_X1 U22397 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19587), .ZN(n19434) );
  OAI211_X1 U22398 ( .C1(n19590), .C2(n19475), .A(n19435), .B(n19434), .ZN(
        P2_U3108) );
  AOI22_X1 U22399 ( .A1(n19440), .A2(n19689), .B1(n19452), .B2(n19688), .ZN(
        n19437) );
  AOI22_X1 U22400 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19634), .ZN(n19436) );
  OAI211_X1 U22401 ( .C1(n19637), .C2(n19475), .A(n19437), .B(n19436), .ZN(
        P2_U3109) );
  AOI22_X1 U22402 ( .A1(n19440), .A2(n19695), .B1(n19452), .B2(n19694), .ZN(
        n19439) );
  AOI22_X1 U22403 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19594), .ZN(n19438) );
  OAI211_X1 U22404 ( .C1(n19538), .C2(n19475), .A(n19439), .B(n19438), .ZN(
        P2_U3110) );
  AOI22_X1 U22405 ( .A1(n19440), .A2(n19702), .B1(n19452), .B2(n19700), .ZN(
        n19444) );
  AOI22_X1 U22406 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19598), .ZN(n19443) );
  OAI211_X1 U22407 ( .C1(n19545), .C2(n19475), .A(n19444), .B(n19443), .ZN(
        P2_U3111) );
  NOR2_X1 U22408 ( .A1(n19445), .A2(n19497), .ZN(n19470) );
  AOI22_X1 U22409 ( .A1(n19606), .A2(n19489), .B1(n19649), .B2(n19470), .ZN(
        n19457) );
  AOI21_X1 U22410 ( .B1(n19482), .B2(n19475), .A(n19446), .ZN(n19447) );
  NOR2_X1 U22411 ( .A1(n19447), .A2(n19609), .ZN(n19451) );
  AOI21_X1 U22412 ( .B1(n10417), .B2(n10900), .A(n19802), .ZN(n19448) );
  AOI21_X1 U22413 ( .B1(n19451), .B2(n19449), .A(n19448), .ZN(n19450) );
  OAI21_X1 U22414 ( .B1(n19450), .B2(n19470), .A(n19656), .ZN(n19472) );
  INV_X1 U22415 ( .A(n19451), .ZN(n19455) );
  OAI21_X1 U22416 ( .B1(n10417), .B2(n19470), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19454) );
  NOR3_X1 U22417 ( .A1(n19452), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19470), 
        .ZN(n19453) );
  AOI22_X1 U22418 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19472), .B1(
        n19650), .B2(n19471), .ZN(n19456) );
  OAI211_X1 U22419 ( .C1(n19620), .C2(n19475), .A(n19457), .B(n19456), .ZN(
        P2_U3112) );
  AOI22_X1 U22420 ( .A1(n19621), .A2(n19489), .B1(n19662), .B2(n19470), .ZN(
        n19459) );
  AOI22_X1 U22421 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19472), .B1(
        n19663), .B2(n19471), .ZN(n19458) );
  OAI211_X1 U22422 ( .C1(n19624), .C2(n19475), .A(n19459), .B(n19458), .ZN(
        P2_U3113) );
  AOI22_X1 U22423 ( .A1(n19562), .A2(n19489), .B1(n19668), .B2(n19470), .ZN(
        n19461) );
  AOI22_X1 U22424 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19472), .B1(
        n19669), .B2(n19471), .ZN(n19460) );
  OAI211_X1 U22425 ( .C1(n19565), .C2(n19475), .A(n19461), .B(n19460), .ZN(
        P2_U3114) );
  AOI22_X1 U22426 ( .A1(n19627), .A2(n19489), .B1(n9562), .B2(n19470), .ZN(
        n19463) );
  AOI22_X1 U22427 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19472), .B1(
        n19675), .B2(n19471), .ZN(n19462) );
  OAI211_X1 U22428 ( .C1(n19630), .C2(n19475), .A(n19463), .B(n19462), .ZN(
        P2_U3115) );
  AOI22_X1 U22429 ( .A1(n19684), .A2(n19489), .B1(n19682), .B2(n19470), .ZN(
        n19465) );
  AOI22_X1 U22430 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19472), .B1(
        n19683), .B2(n19471), .ZN(n19464) );
  OAI211_X1 U22431 ( .C1(n19687), .C2(n19475), .A(n19465), .B(n19464), .ZN(
        P2_U3116) );
  AOI22_X1 U22432 ( .A1(n19690), .A2(n19489), .B1(n19688), .B2(n19470), .ZN(
        n19467) );
  AOI22_X1 U22433 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19472), .B1(
        n19689), .B2(n19471), .ZN(n19466) );
  OAI211_X1 U22434 ( .C1(n19693), .C2(n19475), .A(n19467), .B(n19466), .ZN(
        P2_U3117) );
  AOI22_X1 U22435 ( .A1(n19696), .A2(n19489), .B1(n19694), .B2(n19470), .ZN(
        n19469) );
  AOI22_X1 U22436 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19472), .B1(
        n19695), .B2(n19471), .ZN(n19468) );
  OAI211_X1 U22437 ( .C1(n19699), .C2(n19475), .A(n19469), .B(n19468), .ZN(
        P2_U3118) );
  AOI22_X1 U22438 ( .A1(n19704), .A2(n19489), .B1(n19700), .B2(n19470), .ZN(
        n19474) );
  AOI22_X1 U22439 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19472), .B1(
        n19702), .B2(n19471), .ZN(n19473) );
  OAI211_X1 U22440 ( .C1(n19710), .C2(n19475), .A(n19474), .B(n19473), .ZN(
        P2_U3119) );
  AOI22_X1 U22441 ( .A1(n19621), .A2(n19499), .B1(n19498), .B2(n19662), .ZN(
        n19477) );
  AOI22_X1 U22442 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19491), .B1(
        n19663), .B2(n19490), .ZN(n19476) );
  OAI211_X1 U22443 ( .C1(n19624), .C2(n19482), .A(n19477), .B(n19476), .ZN(
        P2_U3121) );
  AOI22_X1 U22444 ( .A1(n19562), .A2(n19499), .B1(n19668), .B2(n19498), .ZN(
        n19479) );
  AOI22_X1 U22445 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19491), .B1(
        n19669), .B2(n19490), .ZN(n19478) );
  OAI211_X1 U22446 ( .C1(n19565), .C2(n19482), .A(n19479), .B(n19478), .ZN(
        P2_U3122) );
  AOI22_X1 U22447 ( .A1(n19627), .A2(n19499), .B1(n19498), .B2(n9562), .ZN(
        n19481) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19491), .B1(
        n19675), .B2(n19490), .ZN(n19480) );
  OAI211_X1 U22449 ( .C1(n19630), .C2(n19482), .A(n19481), .B(n19480), .ZN(
        P2_U3123) );
  AOI22_X1 U22450 ( .A1(n19587), .A2(n19489), .B1(n19498), .B2(n19682), .ZN(
        n19484) );
  AOI22_X1 U22451 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19491), .B1(
        n19683), .B2(n19490), .ZN(n19483) );
  OAI211_X1 U22452 ( .C1(n19590), .C2(n19523), .A(n19484), .B(n19483), .ZN(
        P2_U3124) );
  AOI22_X1 U22453 ( .A1(n19634), .A2(n19489), .B1(n19498), .B2(n19688), .ZN(
        n19486) );
  AOI22_X1 U22454 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19491), .B1(
        n19689), .B2(n19490), .ZN(n19485) );
  OAI211_X1 U22455 ( .C1(n19637), .C2(n19523), .A(n19486), .B(n19485), .ZN(
        P2_U3125) );
  AOI22_X1 U22456 ( .A1(n19594), .A2(n19489), .B1(n19498), .B2(n19694), .ZN(
        n19488) );
  AOI22_X1 U22457 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19491), .B1(
        n19695), .B2(n19490), .ZN(n19487) );
  OAI211_X1 U22458 ( .C1(n19538), .C2(n19523), .A(n19488), .B(n19487), .ZN(
        P2_U3126) );
  AOI22_X1 U22459 ( .A1(n19598), .A2(n19489), .B1(n19498), .B2(n19700), .ZN(
        n19493) );
  AOI22_X1 U22460 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19491), .B1(
        n19702), .B2(n19490), .ZN(n19492) );
  OAI211_X1 U22461 ( .C1(n19545), .C2(n19523), .A(n19493), .B(n19492), .ZN(
        P2_U3127) );
  NOR3_X2 U22462 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19828), .A3(
        n19497), .ZN(n19518) );
  OAI21_X1 U22463 ( .B1(n19494), .B2(n19518), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19495) );
  OAI21_X1 U22464 ( .B1(n19497), .B2(n19496), .A(n19495), .ZN(n19519) );
  AOI22_X1 U22465 ( .A1(n19519), .A2(n19650), .B1(n19649), .B2(n19518), .ZN(
        n19505) );
  AOI221_X1 U22466 ( .B1(n19499), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19541), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19498), .ZN(n19501) );
  MUX2_X1 U22467 ( .A(n19501), .B(n19500), .S(P2_STATE2_REG_2__SCAN_IN), .Z(
        n19502) );
  NOR2_X1 U22468 ( .A1(n19502), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19503) );
  AOI22_X1 U22469 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19520), .B1(
        n19541), .B2(n19606), .ZN(n19504) );
  OAI211_X1 U22470 ( .C1(n19620), .C2(n19523), .A(n19505), .B(n19504), .ZN(
        P2_U3128) );
  AOI22_X1 U22471 ( .A1(n19519), .A2(n19663), .B1(n19662), .B2(n19518), .ZN(
        n19507) );
  AOI22_X1 U22472 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19520), .B1(
        n19541), .B2(n19621), .ZN(n19506) );
  OAI211_X1 U22473 ( .C1(n19624), .C2(n19523), .A(n19507), .B(n19506), .ZN(
        P2_U3129) );
  AOI22_X1 U22474 ( .A1(n19519), .A2(n19669), .B1(n19668), .B2(n19518), .ZN(
        n19509) );
  AOI22_X1 U22475 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19520), .B1(
        n19541), .B2(n19562), .ZN(n19508) );
  OAI211_X1 U22476 ( .C1(n19565), .C2(n19523), .A(n19509), .B(n19508), .ZN(
        P2_U3130) );
  AOI22_X1 U22477 ( .A1(n19519), .A2(n19675), .B1(n9562), .B2(n19518), .ZN(
        n19511) );
  AOI22_X1 U22478 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19520), .B1(
        n19541), .B2(n19627), .ZN(n19510) );
  OAI211_X1 U22479 ( .C1(n19630), .C2(n19523), .A(n19511), .B(n19510), .ZN(
        P2_U3131) );
  AOI22_X1 U22480 ( .A1(n19519), .A2(n19683), .B1(n19682), .B2(n19518), .ZN(
        n19513) );
  AOI22_X1 U22481 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19520), .B1(
        n19541), .B2(n19684), .ZN(n19512) );
  OAI211_X1 U22482 ( .C1(n19687), .C2(n19523), .A(n19513), .B(n19512), .ZN(
        P2_U3132) );
  AOI22_X1 U22483 ( .A1(n19519), .A2(n19689), .B1(n19688), .B2(n19518), .ZN(
        n19515) );
  AOI22_X1 U22484 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19520), .B1(
        n19541), .B2(n19690), .ZN(n19514) );
  OAI211_X1 U22485 ( .C1(n19693), .C2(n19523), .A(n19515), .B(n19514), .ZN(
        P2_U3133) );
  AOI22_X1 U22486 ( .A1(n19519), .A2(n19695), .B1(n19694), .B2(n19518), .ZN(
        n19517) );
  AOI22_X1 U22487 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19520), .B1(
        n19541), .B2(n19696), .ZN(n19516) );
  OAI211_X1 U22488 ( .C1(n19699), .C2(n19523), .A(n19517), .B(n19516), .ZN(
        P2_U3134) );
  AOI22_X1 U22489 ( .A1(n19519), .A2(n19702), .B1(n19700), .B2(n19518), .ZN(
        n19522) );
  AOI22_X1 U22490 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19520), .B1(
        n19541), .B2(n19704), .ZN(n19521) );
  OAI211_X1 U22491 ( .C1(n19710), .C2(n19523), .A(n19522), .B(n19521), .ZN(
        P2_U3135) );
  AOI22_X1 U22492 ( .A1(n19540), .A2(n19650), .B1(n19649), .B2(n19539), .ZN(
        n19525) );
  AOI22_X1 U22493 ( .A1(n19541), .A2(n19658), .B1(n19551), .B2(n19606), .ZN(
        n19524) );
  OAI211_X1 U22494 ( .C1(n19527), .C2(n19526), .A(n19525), .B(n19524), .ZN(
        P2_U3136) );
  AOI22_X1 U22495 ( .A1(n19540), .A2(n19663), .B1(n19539), .B2(n19662), .ZN(
        n19529) );
  AOI22_X1 U22496 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19542), .B1(
        n19541), .B2(n19664), .ZN(n19528) );
  OAI211_X1 U22497 ( .C1(n19667), .C2(n19579), .A(n19529), .B(n19528), .ZN(
        P2_U3137) );
  AOI22_X1 U22498 ( .A1(n19540), .A2(n19675), .B1(n19539), .B2(n9562), .ZN(
        n19531) );
  AOI22_X1 U22499 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19542), .B1(
        n19541), .B2(n19676), .ZN(n19530) );
  OAI211_X1 U22500 ( .C1(n19681), .C2(n19579), .A(n19531), .B(n19530), .ZN(
        P2_U3139) );
  AOI22_X1 U22501 ( .A1(n19540), .A2(n19683), .B1(n19539), .B2(n19682), .ZN(
        n19533) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19542), .B1(
        n19541), .B2(n19587), .ZN(n19532) );
  OAI211_X1 U22503 ( .C1(n19590), .C2(n19579), .A(n19533), .B(n19532), .ZN(
        P2_U3140) );
  AOI22_X1 U22504 ( .A1(n19540), .A2(n19689), .B1(n19539), .B2(n19688), .ZN(
        n19535) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19542), .B1(
        n19541), .B2(n19634), .ZN(n19534) );
  OAI211_X1 U22506 ( .C1(n19637), .C2(n19579), .A(n19535), .B(n19534), .ZN(
        P2_U3141) );
  AOI22_X1 U22507 ( .A1(n19540), .A2(n19695), .B1(n19539), .B2(n19694), .ZN(
        n19537) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19542), .B1(
        n19541), .B2(n19594), .ZN(n19536) );
  OAI211_X1 U22509 ( .C1(n19538), .C2(n19579), .A(n19537), .B(n19536), .ZN(
        P2_U3142) );
  AOI22_X1 U22510 ( .A1(n19540), .A2(n19702), .B1(n19539), .B2(n19700), .ZN(
        n19544) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19542), .B1(
        n19541), .B2(n19598), .ZN(n19543) );
  OAI211_X1 U22512 ( .C1(n19545), .C2(n19579), .A(n19544), .B(n19543), .ZN(
        P2_U3143) );
  INV_X1 U22513 ( .A(n19546), .ZN(n19550) );
  NOR2_X1 U22514 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19547), .ZN(
        n19574) );
  OAI21_X1 U22515 ( .B1(n19548), .B2(n19574), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19549) );
  OAI21_X1 U22516 ( .B1(n19550), .B2(n19553), .A(n19549), .ZN(n19575) );
  AOI22_X1 U22517 ( .A1(n19575), .A2(n19650), .B1(n19649), .B2(n19574), .ZN(
        n19559) );
  OAI21_X1 U22518 ( .B1(n19599), .B2(n19551), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19552) );
  OAI21_X1 U22519 ( .B1(n19553), .B2(n16335), .A(n19552), .ZN(n19557) );
  INV_X1 U22520 ( .A(n19574), .ZN(n19554) );
  OAI211_X1 U22521 ( .C1(n19555), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19554), 
        .B(n19609), .ZN(n19556) );
  NAND3_X1 U22522 ( .A1(n19557), .A2(n19656), .A3(n19556), .ZN(n19576) );
  AOI22_X1 U22523 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19576), .B1(
        n19599), .B2(n19606), .ZN(n19558) );
  OAI211_X1 U22524 ( .C1(n19620), .C2(n19579), .A(n19559), .B(n19558), .ZN(
        P2_U3144) );
  AOI22_X1 U22525 ( .A1(n19575), .A2(n19663), .B1(n19662), .B2(n19574), .ZN(
        n19561) );
  AOI22_X1 U22526 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19576), .B1(
        n19599), .B2(n19621), .ZN(n19560) );
  OAI211_X1 U22527 ( .C1(n19624), .C2(n19579), .A(n19561), .B(n19560), .ZN(
        P2_U3145) );
  AOI22_X1 U22528 ( .A1(n19575), .A2(n19669), .B1(n19668), .B2(n19574), .ZN(
        n19564) );
  AOI22_X1 U22529 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19576), .B1(
        n19599), .B2(n19562), .ZN(n19563) );
  OAI211_X1 U22530 ( .C1(n19565), .C2(n19579), .A(n19564), .B(n19563), .ZN(
        P2_U3146) );
  AOI22_X1 U22531 ( .A1(n19575), .A2(n19675), .B1(n9562), .B2(n19574), .ZN(
        n19567) );
  AOI22_X1 U22532 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19576), .B1(
        n19599), .B2(n19627), .ZN(n19566) );
  OAI211_X1 U22533 ( .C1(n19630), .C2(n19579), .A(n19567), .B(n19566), .ZN(
        P2_U3147) );
  AOI22_X1 U22534 ( .A1(n19575), .A2(n19683), .B1(n19682), .B2(n19574), .ZN(
        n19569) );
  AOI22_X1 U22535 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19576), .B1(
        n19599), .B2(n19684), .ZN(n19568) );
  OAI211_X1 U22536 ( .C1(n19687), .C2(n19579), .A(n19569), .B(n19568), .ZN(
        P2_U3148) );
  AOI22_X1 U22537 ( .A1(n19575), .A2(n19689), .B1(n19688), .B2(n19574), .ZN(
        n19571) );
  AOI22_X1 U22538 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19576), .B1(
        n19599), .B2(n19690), .ZN(n19570) );
  OAI211_X1 U22539 ( .C1(n19693), .C2(n19579), .A(n19571), .B(n19570), .ZN(
        P2_U3149) );
  AOI22_X1 U22540 ( .A1(n19575), .A2(n19695), .B1(n19694), .B2(n19574), .ZN(
        n19573) );
  AOI22_X1 U22541 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19576), .B1(
        n19599), .B2(n19696), .ZN(n19572) );
  OAI211_X1 U22542 ( .C1(n19699), .C2(n19579), .A(n19573), .B(n19572), .ZN(
        P2_U3150) );
  AOI22_X1 U22543 ( .A1(n19575), .A2(n19702), .B1(n19700), .B2(n19574), .ZN(
        n19578) );
  AOI22_X1 U22544 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19576), .B1(
        n19599), .B2(n19704), .ZN(n19577) );
  OAI211_X1 U22545 ( .C1(n19710), .C2(n19579), .A(n19578), .B(n19577), .ZN(
        P2_U3151) );
  AOI22_X1 U22546 ( .A1(n19597), .A2(n19663), .B1(n19608), .B2(n19662), .ZN(
        n19581) );
  AOI22_X1 U22547 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19591), .B1(
        n19599), .B2(n19664), .ZN(n19580) );
  OAI211_X1 U22548 ( .C1(n19667), .C2(n19645), .A(n19581), .B(n19580), .ZN(
        P2_U3153) );
  AOI22_X1 U22549 ( .A1(n19597), .A2(n19669), .B1(n19608), .B2(n19668), .ZN(
        n19583) );
  AOI22_X1 U22550 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19591), .B1(
        n19599), .B2(n19670), .ZN(n19582) );
  OAI211_X1 U22551 ( .C1(n19673), .C2(n19645), .A(n19583), .B(n19582), .ZN(
        P2_U3154) );
  INV_X1 U22552 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n19586) );
  AOI22_X1 U22553 ( .A1(n19597), .A2(n19675), .B1(n19608), .B2(n9562), .ZN(
        n19585) );
  AOI22_X1 U22554 ( .A1(n19599), .A2(n19676), .B1(n19633), .B2(n19627), .ZN(
        n19584) );
  OAI211_X1 U22555 ( .C1(n19602), .C2(n19586), .A(n19585), .B(n19584), .ZN(
        P2_U3155) );
  AOI22_X1 U22556 ( .A1(n19597), .A2(n19683), .B1(n19608), .B2(n19682), .ZN(
        n19589) );
  AOI22_X1 U22557 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19591), .B1(
        n19599), .B2(n19587), .ZN(n19588) );
  OAI211_X1 U22558 ( .C1(n19590), .C2(n19645), .A(n19589), .B(n19588), .ZN(
        P2_U3156) );
  AOI22_X1 U22559 ( .A1(n19597), .A2(n19689), .B1(n19608), .B2(n19688), .ZN(
        n19593) );
  AOI22_X1 U22560 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19591), .B1(
        n19599), .B2(n19634), .ZN(n19592) );
  OAI211_X1 U22561 ( .C1(n19637), .C2(n19645), .A(n19593), .B(n19592), .ZN(
        P2_U3157) );
  AOI22_X1 U22562 ( .A1(n19597), .A2(n19695), .B1(n19608), .B2(n19694), .ZN(
        n19596) );
  AOI22_X1 U22563 ( .A1(n19599), .A2(n19594), .B1(n19633), .B2(n19696), .ZN(
        n19595) );
  OAI211_X1 U22564 ( .C1(n19602), .C2(n10512), .A(n19596), .B(n19595), .ZN(
        P2_U3158) );
  AOI22_X1 U22565 ( .A1(n19597), .A2(n19702), .B1(n19608), .B2(n19700), .ZN(
        n19601) );
  AOI22_X1 U22566 ( .A1(n19599), .A2(n19598), .B1(n19633), .B2(n19704), .ZN(
        n19600) );
  OAI211_X1 U22567 ( .C1(n19602), .C2(n12386), .A(n19601), .B(n19600), .ZN(
        P2_U3159) );
  NAND2_X1 U22568 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19605), .ZN(
        n19654) );
  NOR2_X1 U22569 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19654), .ZN(
        n19640) );
  AOI22_X1 U22570 ( .A1(n19606), .A2(n19677), .B1(n19649), .B2(n19640), .ZN(
        n19619) );
  OAI21_X1 U22571 ( .B1(n19633), .B2(n19677), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19607) );
  NAND2_X1 U22572 ( .A1(n19607), .A2(n19802), .ZN(n19617) );
  NOR2_X1 U22573 ( .A1(n19640), .A2(n19608), .ZN(n19616) );
  INV_X1 U22574 ( .A(n19616), .ZN(n19613) );
  INV_X1 U22575 ( .A(n19640), .ZN(n19610) );
  OAI211_X1 U22576 ( .C1(n19611), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19610), 
        .B(n19609), .ZN(n19612) );
  OAI211_X1 U22577 ( .C1(n19617), .C2(n19613), .A(n19656), .B(n19612), .ZN(
        n19642) );
  OAI21_X1 U22578 ( .B1(n19614), .B2(n19640), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19615) );
  AOI22_X1 U22579 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19642), .B1(
        n19650), .B2(n19641), .ZN(n19618) );
  OAI211_X1 U22580 ( .C1(n19620), .C2(n19645), .A(n19619), .B(n19618), .ZN(
        P2_U3160) );
  AOI22_X1 U22581 ( .A1(n19621), .A2(n19677), .B1(n19662), .B2(n19640), .ZN(
        n19623) );
  AOI22_X1 U22582 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19642), .B1(
        n19663), .B2(n19641), .ZN(n19622) );
  OAI211_X1 U22583 ( .C1(n19624), .C2(n19645), .A(n19623), .B(n19622), .ZN(
        P2_U3161) );
  AOI22_X1 U22584 ( .A1(n19670), .A2(n19633), .B1(n19668), .B2(n19640), .ZN(
        n19626) );
  AOI22_X1 U22585 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19642), .B1(
        n19669), .B2(n19641), .ZN(n19625) );
  OAI211_X1 U22586 ( .C1(n19673), .C2(n19709), .A(n19626), .B(n19625), .ZN(
        P2_U3162) );
  AOI22_X1 U22587 ( .A1(n19627), .A2(n19677), .B1(n9562), .B2(n19640), .ZN(
        n19629) );
  AOI22_X1 U22588 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19642), .B1(
        n19675), .B2(n19641), .ZN(n19628) );
  OAI211_X1 U22589 ( .C1(n19630), .C2(n19645), .A(n19629), .B(n19628), .ZN(
        P2_U3163) );
  AOI22_X1 U22590 ( .A1(n19684), .A2(n19677), .B1(n19682), .B2(n19640), .ZN(
        n19632) );
  AOI22_X1 U22591 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19642), .B1(
        n19683), .B2(n19641), .ZN(n19631) );
  OAI211_X1 U22592 ( .C1(n19687), .C2(n19645), .A(n19632), .B(n19631), .ZN(
        P2_U3164) );
  AOI22_X1 U22593 ( .A1(n19634), .A2(n19633), .B1(n19688), .B2(n19640), .ZN(
        n19636) );
  AOI22_X1 U22594 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19642), .B1(
        n19689), .B2(n19641), .ZN(n19635) );
  OAI211_X1 U22595 ( .C1(n19637), .C2(n19709), .A(n19636), .B(n19635), .ZN(
        P2_U3165) );
  AOI22_X1 U22596 ( .A1(n19696), .A2(n19677), .B1(n19694), .B2(n19640), .ZN(
        n19639) );
  AOI22_X1 U22597 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19642), .B1(
        n19695), .B2(n19641), .ZN(n19638) );
  OAI211_X1 U22598 ( .C1(n19699), .C2(n19645), .A(n19639), .B(n19638), .ZN(
        P2_U3166) );
  AOI22_X1 U22599 ( .A1(n19704), .A2(n19677), .B1(n19700), .B2(n19640), .ZN(
        n19644) );
  AOI22_X1 U22600 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19642), .B1(
        n19702), .B2(n19641), .ZN(n19643) );
  OAI211_X1 U22601 ( .C1(n19710), .C2(n19645), .A(n19644), .B(n19643), .ZN(
        P2_U3167) );
  INV_X1 U22602 ( .A(n19701), .ZN(n19646) );
  NAND3_X1 U22603 ( .A1(n19647), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19646), 
        .ZN(n19655) );
  OAI21_X1 U22604 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19654), .A(n19860), 
        .ZN(n19648) );
  AND2_X1 U22605 ( .A1(n19655), .A2(n19648), .ZN(n19703) );
  AOI22_X1 U22606 ( .A1(n19703), .A2(n19650), .B1(n19649), .B2(n19701), .ZN(
        n19660) );
  NOR2_X1 U22607 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10900), .ZN(
        n19831) );
  NAND3_X1 U22608 ( .A1(n19652), .A2(n19651), .A3(n10900), .ZN(n19653) );
  OAI21_X1 U22609 ( .B1(n19831), .B2(n19654), .A(n19653), .ZN(n19657) );
  NAND3_X1 U22610 ( .A1(n19657), .A2(n19656), .A3(n19655), .ZN(n19706) );
  AOI22_X1 U22611 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19706), .B1(
        n19677), .B2(n19658), .ZN(n19659) );
  OAI211_X1 U22612 ( .C1(n19661), .C2(n19680), .A(n19660), .B(n19659), .ZN(
        P2_U3168) );
  AOI22_X1 U22613 ( .A1(n19703), .A2(n19663), .B1(n19701), .B2(n19662), .ZN(
        n19666) );
  AOI22_X1 U22614 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19706), .B1(
        n19677), .B2(n19664), .ZN(n19665) );
  OAI211_X1 U22615 ( .C1(n19667), .C2(n19680), .A(n19666), .B(n19665), .ZN(
        P2_U3169) );
  AOI22_X1 U22616 ( .A1(n19703), .A2(n19669), .B1(n19668), .B2(n19701), .ZN(
        n19672) );
  AOI22_X1 U22617 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19706), .B1(
        n19677), .B2(n19670), .ZN(n19671) );
  OAI211_X1 U22618 ( .C1(n19673), .C2(n19680), .A(n19672), .B(n19671), .ZN(
        P2_U3170) );
  AOI22_X1 U22619 ( .A1(n19703), .A2(n19675), .B1(n19701), .B2(n9562), .ZN(
        n19679) );
  AOI22_X1 U22620 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19706), .B1(
        n19677), .B2(n19676), .ZN(n19678) );
  OAI211_X1 U22621 ( .C1(n19681), .C2(n19680), .A(n19679), .B(n19678), .ZN(
        P2_U3171) );
  AOI22_X1 U22622 ( .A1(n19703), .A2(n19683), .B1(n19701), .B2(n19682), .ZN(
        n19686) );
  AOI22_X1 U22623 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19706), .B1(
        n19705), .B2(n19684), .ZN(n19685) );
  OAI211_X1 U22624 ( .C1(n19687), .C2(n19709), .A(n19686), .B(n19685), .ZN(
        P2_U3172) );
  AOI22_X1 U22625 ( .A1(n19703), .A2(n19689), .B1(n19701), .B2(n19688), .ZN(
        n19692) );
  AOI22_X1 U22626 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19706), .B1(
        n19705), .B2(n19690), .ZN(n19691) );
  OAI211_X1 U22627 ( .C1(n19693), .C2(n19709), .A(n19692), .B(n19691), .ZN(
        P2_U3173) );
  AOI22_X1 U22628 ( .A1(n19703), .A2(n19695), .B1(n19701), .B2(n19694), .ZN(
        n19698) );
  AOI22_X1 U22629 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19706), .B1(
        n19705), .B2(n19696), .ZN(n19697) );
  OAI211_X1 U22630 ( .C1(n19699), .C2(n19709), .A(n19698), .B(n19697), .ZN(
        P2_U3174) );
  AOI22_X1 U22631 ( .A1(n19703), .A2(n19702), .B1(n19701), .B2(n19700), .ZN(
        n19708) );
  AOI22_X1 U22632 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19706), .B1(
        n19705), .B2(n19704), .ZN(n19707) );
  OAI211_X1 U22633 ( .C1(n19710), .C2(n19709), .A(n19708), .B(n19707), .ZN(
        P2_U3175) );
  NAND4_X1 U22634 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19712), .A3(n10900), 
        .A4(n19711), .ZN(n19713) );
  NAND2_X1 U22635 ( .A1(n19714), .A2(n19713), .ZN(n19718) );
  NAND2_X1 U22636 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19865), .ZN(n19715) );
  AOI21_X1 U22637 ( .B1(n19716), .B2(n19719), .A(n19715), .ZN(n19717) );
  AOI21_X1 U22638 ( .B1(n19719), .B2(n19718), .A(n19717), .ZN(n19721) );
  NAND2_X1 U22639 ( .A1(n19721), .A2(n19720), .ZN(P2_U3177) );
  AND2_X1 U22640 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19722), .ZN(
        P2_U3179) );
  AND2_X1 U22641 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19722), .ZN(
        P2_U3180) );
  AND2_X1 U22642 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19722), .ZN(
        P2_U3181) );
  AND2_X1 U22643 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19722), .ZN(
        P2_U3182) );
  AND2_X1 U22644 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19722), .ZN(
        P2_U3183) );
  AND2_X1 U22645 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19722), .ZN(
        P2_U3184) );
  AND2_X1 U22646 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19722), .ZN(
        P2_U3185) );
  AND2_X1 U22647 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19722), .ZN(
        P2_U3186) );
  AND2_X1 U22648 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19722), .ZN(
        P2_U3187) );
  AND2_X1 U22649 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19722), .ZN(
        P2_U3188) );
  INV_X1 U22650 ( .A(P2_DATAWIDTH_REG_21__SCAN_IN), .ZN(n20851) );
  NOR2_X1 U22651 ( .A1(n20851), .A2(n19798), .ZN(P2_U3189) );
  AND2_X1 U22652 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19722), .ZN(
        P2_U3190) );
  AND2_X1 U22653 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19722), .ZN(
        P2_U3191) );
  AND2_X1 U22654 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19722), .ZN(
        P2_U3192) );
  AND2_X1 U22655 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19722), .ZN(
        P2_U3193) );
  AND2_X1 U22656 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19722), .ZN(
        P2_U3194) );
  AND2_X1 U22657 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19722), .ZN(
        P2_U3195) );
  AND2_X1 U22658 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19722), .ZN(
        P2_U3196) );
  AND2_X1 U22659 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19722), .ZN(
        P2_U3197) );
  AND2_X1 U22660 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19722), .ZN(
        P2_U3198) );
  AND2_X1 U22661 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19722), .ZN(
        P2_U3199) );
  AND2_X1 U22662 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19722), .ZN(
        P2_U3200) );
  AND2_X1 U22663 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19722), .ZN(P2_U3201) );
  AND2_X1 U22664 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19722), .ZN(P2_U3202) );
  AND2_X1 U22665 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19722), .ZN(P2_U3203) );
  AND2_X1 U22666 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19722), .ZN(P2_U3204) );
  AND2_X1 U22667 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19722), .ZN(P2_U3205) );
  AND2_X1 U22668 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19722), .ZN(P2_U3206) );
  AND2_X1 U22669 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19722), .ZN(P2_U3207) );
  AND2_X1 U22670 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19722), .ZN(P2_U3208) );
  OAI21_X1 U22671 ( .B1(n20694), .B2(n19729), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19738) );
  NAND2_X1 U22672 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19865), .ZN(n19736) );
  NAND3_X1 U22673 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19736), .ZN(n19725) );
  AOI211_X1 U22674 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20684), .A(
        n19868), .B(n19723), .ZN(n19724) );
  AOI21_X1 U22675 ( .B1(n19738), .B2(n19725), .A(n19724), .ZN(n19726) );
  INV_X1 U22676 ( .A(n19726), .ZN(P2_U3209) );
  AND2_X1 U22677 ( .A1(n19727), .A2(n19736), .ZN(n19731) );
  NOR2_X1 U22678 ( .A1(HOLD), .A2(n19728), .ZN(n19737) );
  OAI211_X1 U22679 ( .C1(n19737), .C2(n19739), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .B(n19729), .ZN(n19730) );
  OAI211_X1 U22680 ( .C1(n19732), .C2(n20684), .A(n19731), .B(n19730), .ZN(
        P2_U3210) );
  OAI22_X1 U22681 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19733), .B1(NA), 
        .B2(n19736), .ZN(n19734) );
  OAI211_X1 U22682 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19734), .ZN(n19735) );
  OAI221_X1 U22683 ( .B1(n19738), .B2(n19737), .C1(n19738), .C2(n19736), .A(
        n19735), .ZN(P2_U3211) );
  OAI222_X1 U22684 ( .A1(n19792), .A2(n19742), .B1(n19741), .B2(n19868), .C1(
        n19740), .C2(n19790), .ZN(P2_U3212) );
  OAI222_X1 U22685 ( .A1(n19792), .A2(n19744), .B1(n19743), .B2(n19868), .C1(
        n19742), .C2(n19790), .ZN(P2_U3213) );
  INV_X1 U22686 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19746) );
  OAI222_X1 U22687 ( .A1(n19792), .A2(n19746), .B1(n19745), .B2(n19868), .C1(
        n19744), .C2(n19790), .ZN(P2_U3214) );
  OAI222_X1 U22688 ( .A1(n19792), .A2(n19748), .B1(n19747), .B2(n19868), .C1(
        n19746), .C2(n19790), .ZN(P2_U3215) );
  OAI222_X1 U22689 ( .A1(n19792), .A2(n19749), .B1(n20810), .B2(n19868), .C1(
        n19748), .C2(n19790), .ZN(P2_U3216) );
  OAI222_X1 U22690 ( .A1(n19792), .A2(n19751), .B1(n19750), .B2(n19868), .C1(
        n19749), .C2(n19790), .ZN(P2_U3217) );
  OAI222_X1 U22691 ( .A1(n19792), .A2(n19753), .B1(n19752), .B2(n19868), .C1(
        n19751), .C2(n19790), .ZN(P2_U3218) );
  OAI222_X1 U22692 ( .A1(n19792), .A2(n19755), .B1(n19754), .B2(n19868), .C1(
        n19753), .C2(n19790), .ZN(P2_U3219) );
  OAI222_X1 U22693 ( .A1(n19792), .A2(n19757), .B1(n19756), .B2(n19868), .C1(
        n19755), .C2(n19790), .ZN(P2_U3220) );
  OAI222_X1 U22694 ( .A1(n19792), .A2(n15452), .B1(n19758), .B2(n19868), .C1(
        n19757), .C2(n19790), .ZN(P2_U3221) );
  INV_X1 U22695 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19760) );
  OAI222_X1 U22696 ( .A1(n19792), .A2(n19760), .B1(n19759), .B2(n19868), .C1(
        n15452), .C2(n19790), .ZN(P2_U3222) );
  OAI222_X1 U22697 ( .A1(n19792), .A2(n20796), .B1(n19761), .B2(n19868), .C1(
        n19760), .C2(n19790), .ZN(P2_U3223) );
  OAI222_X1 U22698 ( .A1(n19792), .A2(n19763), .B1(n19762), .B2(n19868), .C1(
        n20796), .C2(n19790), .ZN(P2_U3224) );
  OAI222_X1 U22699 ( .A1(n19792), .A2(n15211), .B1(n19764), .B2(n19868), .C1(
        n19763), .C2(n19790), .ZN(P2_U3225) );
  OAI222_X1 U22700 ( .A1(n19792), .A2(n19765), .B1(n20873), .B2(n19868), .C1(
        n15211), .C2(n19790), .ZN(P2_U3226) );
  OAI222_X1 U22701 ( .A1(n19792), .A2(n19767), .B1(n19766), .B2(n19868), .C1(
        n19765), .C2(n19790), .ZN(P2_U3227) );
  OAI222_X1 U22702 ( .A1(n19792), .A2(n19769), .B1(n19768), .B2(n19868), .C1(
        n19767), .C2(n19790), .ZN(P2_U3228) );
  INV_X1 U22703 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19771) );
  OAI222_X1 U22704 ( .A1(n19792), .A2(n19771), .B1(n19770), .B2(n19868), .C1(
        n19769), .C2(n19790), .ZN(P2_U3229) );
  OAI222_X1 U22705 ( .A1(n19792), .A2(n19772), .B1(n20783), .B2(n19868), .C1(
        n19771), .C2(n19790), .ZN(P2_U3230) );
  OAI222_X1 U22706 ( .A1(n19792), .A2(n19774), .B1(n19773), .B2(n19868), .C1(
        n19772), .C2(n19790), .ZN(P2_U3231) );
  OAI222_X1 U22707 ( .A1(n19792), .A2(n15751), .B1(n19775), .B2(n19868), .C1(
        n19774), .C2(n19790), .ZN(P2_U3232) );
  OAI222_X1 U22708 ( .A1(n19792), .A2(n19777), .B1(n19776), .B2(n19868), .C1(
        n15751), .C2(n19790), .ZN(P2_U3233) );
  OAI222_X1 U22709 ( .A1(n19792), .A2(n19779), .B1(n19778), .B2(n19868), .C1(
        n19777), .C2(n19790), .ZN(P2_U3234) );
  OAI222_X1 U22710 ( .A1(n19792), .A2(n19781), .B1(n19780), .B2(n19868), .C1(
        n19779), .C2(n19790), .ZN(P2_U3235) );
  OAI222_X1 U22711 ( .A1(n19792), .A2(n19783), .B1(n19782), .B2(n19868), .C1(
        n19781), .C2(n19790), .ZN(P2_U3236) );
  OAI222_X1 U22712 ( .A1(n19792), .A2(n19786), .B1(n19784), .B2(n19868), .C1(
        n19783), .C2(n19790), .ZN(P2_U3237) );
  INV_X1 U22713 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19787) );
  OAI222_X1 U22714 ( .A1(n19790), .A2(n19786), .B1(n19785), .B2(n19868), .C1(
        n19787), .C2(n19792), .ZN(P2_U3238) );
  INV_X1 U22715 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19789) );
  OAI222_X1 U22716 ( .A1(n19792), .A2(n19789), .B1(n19788), .B2(n19868), .C1(
        n19787), .C2(n19790), .ZN(P2_U3239) );
  OAI222_X1 U22717 ( .A1(n19792), .A2(n10899), .B1(n20865), .B2(n19868), .C1(
        n19789), .C2(n19790), .ZN(P2_U3240) );
  OAI222_X1 U22718 ( .A1(n19792), .A2(n14255), .B1(n19791), .B2(n19868), .C1(
        n10899), .C2(n19790), .ZN(P2_U3241) );
  OAI22_X1 U22719 ( .A1(n19869), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19868), .ZN(n19793) );
  INV_X1 U22720 ( .A(n19793), .ZN(P2_U3585) );
  MUX2_X1 U22721 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19869), .Z(P2_U3586) );
  MUX2_X1 U22722 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .B(P2_BE_N_REG_1__SCAN_IN), .S(n19869), .Z(P2_U3587) );
  OAI22_X1 U22723 ( .A1(n19869), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19868), .ZN(n19794) );
  INV_X1 U22724 ( .A(n19794), .ZN(P2_U3588) );
  OAI21_X1 U22725 ( .B1(n19798), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19796), 
        .ZN(n19795) );
  INV_X1 U22726 ( .A(n19795), .ZN(P2_U3591) );
  OAI21_X1 U22727 ( .B1(n19798), .B2(n19797), .A(n19796), .ZN(P2_U3592) );
  NAND2_X1 U22728 ( .A1(n19799), .A2(n19802), .ZN(n19808) );
  AND2_X1 U22729 ( .A1(n19802), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19824) );
  NAND2_X1 U22730 ( .A1(n19800), .A2(n19824), .ZN(n19813) );
  NAND2_X1 U22731 ( .A1(n19822), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19803) );
  AOI21_X1 U22732 ( .B1(n19803), .B2(n19802), .A(n19801), .ZN(n19811) );
  NAND2_X1 U22733 ( .A1(n19813), .A2(n19811), .ZN(n19806) );
  AOI22_X1 U22734 ( .A1(n19806), .A2(n19805), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19804), .ZN(n19807) );
  AND2_X1 U22735 ( .A1(n19808), .A2(n19807), .ZN(n19809) );
  AOI22_X1 U22736 ( .A1(n19838), .A2(n16335), .B1(n19809), .B2(n19835), .ZN(
        P2_U3602) );
  INV_X1 U22737 ( .A(n19810), .ZN(n19817) );
  INV_X1 U22738 ( .A(n19811), .ZN(n19816) );
  NOR2_X1 U22739 ( .A1(n19812), .A2(n10900), .ZN(n19815) );
  INV_X1 U22740 ( .A(n19813), .ZN(n19814) );
  AOI211_X1 U22741 ( .C1(n19817), .C2(n19816), .A(n19815), .B(n19814), .ZN(
        n19818) );
  AOI22_X1 U22742 ( .A1(n19838), .A2(n19819), .B1(n19818), .B2(n19835), .ZN(
        P2_U3603) );
  INV_X1 U22743 ( .A(n19820), .ZN(n19829) );
  AND2_X1 U22744 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19821) );
  NOR2_X1 U22745 ( .A1(n19829), .A2(n19821), .ZN(n19823) );
  MUX2_X1 U22746 ( .A(n19824), .B(n19823), .S(n19822), .Z(n19825) );
  AOI21_X1 U22747 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19826), .A(n19825), 
        .ZN(n19827) );
  AOI22_X1 U22748 ( .A1(n19838), .A2(n19828), .B1(n19827), .B2(n19835), .ZN(
        P2_U3604) );
  NOR2_X1 U22749 ( .A1(n19830), .A2(n19829), .ZN(n19832) );
  AOI211_X1 U22750 ( .C1(n19834), .C2(n19833), .A(n19832), .B(n19831), .ZN(
        n19836) );
  AOI22_X1 U22751 ( .A1(n19838), .A2(n19837), .B1(n19836), .B2(n19835), .ZN(
        P2_U3605) );
  INV_X1 U22752 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19839) );
  AOI22_X1 U22753 ( .A1(n19868), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19839), 
        .B2(n19869), .ZN(P2_U3608) );
  INV_X1 U22754 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n19850) );
  INV_X1 U22755 ( .A(n19840), .ZN(n19849) );
  INV_X1 U22756 ( .A(n19841), .ZN(n19845) );
  AOI22_X1 U22757 ( .A1(n19845), .A2(n19844), .B1(n19843), .B2(n19842), .ZN(
        n19848) );
  NOR2_X1 U22758 ( .A1(n19849), .A2(n19846), .ZN(n19847) );
  AOI22_X1 U22759 ( .A1(n19850), .A2(n19849), .B1(n19848), .B2(n19847), .ZN(
        P2_U3609) );
  AOI21_X1 U22760 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19854), .A(n19851), 
        .ZN(n19856) );
  NOR3_X1 U22761 ( .A1(n19854), .A2(n19853), .A3(n19852), .ZN(n19855) );
  OAI21_X1 U22762 ( .B1(n19856), .B2(n19855), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19859) );
  OAI22_X1 U22763 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19857), .B1(n19865), 
        .B2(n19860), .ZN(n19858) );
  NAND2_X1 U22764 ( .A1(n19859), .A2(n19858), .ZN(n19867) );
  OAI21_X1 U22765 ( .B1(n19861), .B2(n19860), .A(n10900), .ZN(n19863) );
  OAI211_X1 U22766 ( .C1(n19865), .C2(n19864), .A(n19863), .B(n19862), .ZN(
        n19866) );
  MUX2_X1 U22767 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n19867), .S(n19866), 
        .Z(P2_U3610) );
  OAI22_X1 U22768 ( .A1(n19869), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19868), .ZN(n19870) );
  INV_X1 U22769 ( .A(n19870), .ZN(P2_U3611) );
  NOR2_X1 U22770 ( .A1(n19878), .A2(n20695), .ZN(n19872) );
  INV_X1 U22771 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19871) );
  AOI21_X1 U22772 ( .B1(n19872), .B2(n19871), .A(n20757), .ZN(P1_U2802) );
  OAI21_X1 U22773 ( .B1(n19874), .B2(n19873), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19875) );
  OAI21_X1 U22774 ( .B1(n19876), .B2(n20676), .A(n19875), .ZN(P1_U2803) );
  INV_X2 U22775 ( .A(n20757), .ZN(n20771) );
  NOR2_X1 U22776 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20683) );
  OAI21_X1 U22777 ( .B1(n20683), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20771), .ZN(
        n19877) );
  OAI21_X1 U22778 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20771), .A(n19877), 
        .ZN(P1_U2804) );
  OAI21_X1 U22779 ( .B1(n20695), .B2(n19878), .A(n20771), .ZN(n20681) );
  INV_X1 U22780 ( .A(n20681), .ZN(n20748) );
  OAI21_X1 U22781 ( .B1(BS16), .B2(n20683), .A(n20748), .ZN(n20746) );
  OAI21_X1 U22782 ( .B1(n20748), .B2(n20777), .A(n20746), .ZN(P1_U2805) );
  OAI21_X1 U22783 ( .B1(n19881), .B2(n19880), .A(n19879), .ZN(P1_U2806) );
  NOR4_X1 U22784 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19885) );
  NOR4_X1 U22785 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19884) );
  NOR4_X1 U22786 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19883) );
  NOR4_X1 U22787 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19882) );
  NAND4_X1 U22788 ( .A1(n19885), .A2(n19884), .A3(n19883), .A4(n19882), .ZN(
        n19891) );
  NOR4_X1 U22789 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19889) );
  AOI211_X1 U22790 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_7__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19888) );
  NOR4_X1 U22791 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19887) );
  NOR4_X1 U22792 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19886) );
  NAND4_X1 U22793 ( .A1(n19889), .A2(n19888), .A3(n19887), .A4(n19886), .ZN(
        n19890) );
  NOR2_X1 U22794 ( .A1(n19891), .A2(n19890), .ZN(n20756) );
  INV_X1 U22795 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19893) );
  NOR3_X1 U22796 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19894) );
  OAI21_X1 U22797 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19894), .A(n20756), .ZN(
        n19892) );
  OAI21_X1 U22798 ( .B1(n20756), .B2(n19893), .A(n19892), .ZN(P1_U2807) );
  INV_X1 U22799 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20747) );
  AOI21_X1 U22800 ( .B1(n20749), .B2(n20747), .A(n19894), .ZN(n19896) );
  INV_X1 U22801 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19895) );
  INV_X1 U22802 ( .A(n20756), .ZN(n20751) );
  AOI22_X1 U22803 ( .A1(n20756), .A2(n19896), .B1(n19895), .B2(n20751), .ZN(
        P1_U2808) );
  INV_X1 U22804 ( .A(n19897), .ZN(n19899) );
  NAND2_X1 U22805 ( .A1(n19913), .A2(n19898), .ZN(n19954) );
  OAI21_X1 U22806 ( .B1(n19899), .B2(n19954), .A(n19955), .ZN(n19926) );
  NOR3_X1 U22807 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19901), .A3(n19900), .ZN(
        n19902) );
  AOI211_X1 U22808 ( .C1(n19969), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n19968), .B(n19902), .ZN(n19906) );
  INV_X1 U22809 ( .A(n19903), .ZN(n19904) );
  AOI22_X1 U22810 ( .A1(n19974), .A2(P1_EBX_REG_9__SCAN_IN), .B1(n19942), .B2(
        n19904), .ZN(n19905) );
  AND2_X1 U22811 ( .A1(n19906), .A2(n19905), .ZN(n19912) );
  INV_X1 U22812 ( .A(n19907), .ZN(n19910) );
  AOI22_X1 U22813 ( .A1(n19910), .A2(n19936), .B1(n19909), .B2(n19908), .ZN(
        n19911) );
  OAI211_X1 U22814 ( .C1(n14028), .C2(n19926), .A(n19912), .B(n19911), .ZN(
        P1_U2831) );
  NAND2_X1 U22815 ( .A1(n19914), .A2(n19913), .ZN(n19962) );
  NOR3_X1 U22816 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n19915), .A3(n19962), .ZN(
        n19922) );
  NAND2_X1 U22817 ( .A1(n19969), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n19916) );
  OAI211_X1 U22818 ( .C1(n19986), .C2(n19917), .A(n19944), .B(n19916), .ZN(
        n19918) );
  AOI21_X1 U22819 ( .B1(n19974), .B2(P1_EBX_REG_8__SCAN_IN), .A(n19918), .ZN(
        n19919) );
  OAI21_X1 U22820 ( .B1(n19920), .B2(n19946), .A(n19919), .ZN(n19921) );
  AOI211_X1 U22821 ( .C1(n19924), .C2(n19923), .A(n19922), .B(n19921), .ZN(
        n19925) );
  OAI21_X1 U22822 ( .B1(n13990), .B2(n19926), .A(n19925), .ZN(P1_U2832) );
  INV_X1 U22823 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n19940) );
  NAND2_X1 U22824 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19927) );
  OAI21_X1 U22825 ( .B1(n19927), .B2(n19954), .A(n19955), .ZN(n19952) );
  NOR3_X1 U22826 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19927), .A3(n19962), .ZN(
        n19930) );
  INV_X1 U22827 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n19928) );
  NOR2_X1 U22828 ( .A1(n19960), .A2(n19928), .ZN(n19929) );
  NOR2_X1 U22829 ( .A1(n19930), .A2(n19929), .ZN(n19939) );
  NAND2_X1 U22830 ( .A1(n19942), .A2(n19931), .ZN(n19933) );
  AOI21_X1 U22831 ( .B1(n19969), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n19968), .ZN(n19932) );
  OAI211_X1 U22832 ( .C1(n19986), .C2(n19934), .A(n19933), .B(n19932), .ZN(
        n19935) );
  AOI21_X1 U22833 ( .B1(n19937), .B2(n19936), .A(n19935), .ZN(n19938) );
  OAI211_X1 U22834 ( .C1(n19940), .C2(n19952), .A(n19939), .B(n19938), .ZN(
        P1_U2833) );
  INV_X1 U22835 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n19953) );
  NOR2_X1 U22836 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n19962), .ZN(n19941) );
  AOI22_X1 U22837 ( .A1(n19942), .A2(n19988), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n19941), .ZN(n19951) );
  NAND2_X1 U22838 ( .A1(n19969), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19943) );
  OAI211_X1 U22839 ( .C1(n19986), .C2(n19945), .A(n19944), .B(n19943), .ZN(
        n19949) );
  NOR2_X1 U22840 ( .A1(n19947), .A2(n19946), .ZN(n19948) );
  AOI211_X1 U22841 ( .C1(n19974), .C2(P1_EBX_REG_6__SCAN_IN), .A(n19949), .B(
        n19948), .ZN(n19950) );
  OAI211_X1 U22842 ( .C1(n19953), .C2(n19952), .A(n19951), .B(n19950), .ZN(
        P1_U2834) );
  NAND2_X1 U22843 ( .A1(n19955), .A2(n19954), .ZN(n19978) );
  OAI22_X1 U22844 ( .A1(n19957), .A2(n19986), .B1(n19977), .B2(n19956), .ZN(
        n19958) );
  AOI211_X1 U22845 ( .C1(n19969), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n19968), .B(n19958), .ZN(n19966) );
  INV_X1 U22846 ( .A(n19959), .ZN(n19964) );
  OAI22_X1 U22847 ( .A1(n19962), .A2(P1_REIP_REG_5__SCAN_IN), .B1(n19961), 
        .B2(n19960), .ZN(n19963) );
  AOI21_X1 U22848 ( .B1(n19964), .B2(n19983), .A(n19963), .ZN(n19965) );
  OAI211_X1 U22849 ( .C1(n13781), .C2(n19978), .A(n19966), .B(n19965), .ZN(
        P1_U2835) );
  INV_X1 U22850 ( .A(n19967), .ZN(n19971) );
  AOI21_X1 U22851 ( .B1(n19969), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n19968), .ZN(n19970) );
  OAI21_X1 U22852 ( .B1(n19972), .B2(n19971), .A(n19970), .ZN(n19973) );
  AOI21_X1 U22853 ( .B1(n19974), .B2(P1_EBX_REG_4__SCAN_IN), .A(n19973), .ZN(
        n19975) );
  OAI21_X1 U22854 ( .B1(n19977), .B2(n19976), .A(n19975), .ZN(n19982) );
  AOI221_X1 U22855 ( .B1(n19980), .B2(n20840), .C1(n19979), .C2(n20840), .A(
        n19978), .ZN(n19981) );
  AOI211_X1 U22856 ( .C1(n19984), .C2(n19983), .A(n19982), .B(n19981), .ZN(
        n19985) );
  OAI21_X1 U22857 ( .B1(n19987), .B2(n19986), .A(n19985), .ZN(P1_U2836) );
  AOI22_X1 U22858 ( .A1(n19991), .A2(n19990), .B1(n19989), .B2(n19988), .ZN(
        n19992) );
  OAI21_X1 U22859 ( .B1(n19994), .B2(n19993), .A(n19992), .ZN(P1_U2866) );
  AOI22_X1 U22860 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19995) );
  OAI21_X1 U22861 ( .B1(n19996), .B2(n20023), .A(n19995), .ZN(P1_U2921) );
  INV_X1 U22862 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n19998) );
  AOI22_X1 U22863 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19997) );
  OAI21_X1 U22864 ( .B1(n19998), .B2(n20023), .A(n19997), .ZN(P1_U2922) );
  INV_X1 U22865 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20000) );
  AOI22_X1 U22866 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20021), .B1(n20007), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19999) );
  OAI21_X1 U22867 ( .B1(n20000), .B2(n20023), .A(n19999), .ZN(P1_U2923) );
  INV_X1 U22868 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20002) );
  AOI22_X1 U22869 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20021), .B1(n20007), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20001) );
  OAI21_X1 U22870 ( .B1(n20002), .B2(n20023), .A(n20001), .ZN(P1_U2924) );
  INV_X1 U22871 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20004) );
  AOI22_X1 U22872 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20021), .B1(n20007), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20003) );
  OAI21_X1 U22873 ( .B1(n20004), .B2(n20023), .A(n20003), .ZN(P1_U2925) );
  INV_X1 U22874 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20006) );
  AOI22_X1 U22875 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20021), .B1(n20007), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20005) );
  OAI21_X1 U22876 ( .B1(n20006), .B2(n20023), .A(n20005), .ZN(P1_U2926) );
  INV_X1 U22877 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20009) );
  AOI22_X1 U22878 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20021), .B1(n20007), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20008) );
  OAI21_X1 U22879 ( .B1(n20009), .B2(n20023), .A(n20008), .ZN(P1_U2927) );
  AOI22_X1 U22880 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20010) );
  OAI21_X1 U22881 ( .B1(n13748), .B2(n20023), .A(n20010), .ZN(P1_U2929) );
  AOI22_X1 U22882 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20011) );
  OAI21_X1 U22883 ( .B1(n11757), .B2(n20023), .A(n20011), .ZN(P1_U2930) );
  AOI22_X1 U22884 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20012) );
  OAI21_X1 U22885 ( .B1(n20013), .B2(n20023), .A(n20012), .ZN(P1_U2931) );
  AOI22_X1 U22886 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20014) );
  OAI21_X1 U22887 ( .B1(n20015), .B2(n20023), .A(n20014), .ZN(P1_U2932) );
  AOI22_X1 U22888 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20016) );
  OAI21_X1 U22889 ( .B1(n20017), .B2(n20023), .A(n20016), .ZN(P1_U2933) );
  AOI22_X1 U22890 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20018) );
  OAI21_X1 U22891 ( .B1(n13515), .B2(n20023), .A(n20018), .ZN(P1_U2934) );
  AOI22_X1 U22892 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20019) );
  OAI21_X1 U22893 ( .B1(n20020), .B2(n20023), .A(n20019), .ZN(P1_U2935) );
  AOI22_X1 U22894 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20021), .B1(n20924), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20022) );
  OAI21_X1 U22895 ( .B1(n20024), .B2(n20023), .A(n20022), .ZN(P1_U2936) );
  AOI22_X1 U22896 ( .A1(n20053), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20052), .ZN(n20026) );
  NAND2_X1 U22897 ( .A1(n20038), .A2(n20025), .ZN(n20040) );
  NAND2_X1 U22898 ( .A1(n20026), .A2(n20040), .ZN(P1_U2945) );
  AOI22_X1 U22899 ( .A1(n20053), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20052), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n20028) );
  NAND2_X1 U22900 ( .A1(n20038), .A2(n20027), .ZN(n20042) );
  NAND2_X1 U22901 ( .A1(n20028), .A2(n20042), .ZN(P1_U2946) );
  AOI22_X1 U22902 ( .A1(n20053), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20052), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20030) );
  NAND2_X1 U22903 ( .A1(n20038), .A2(n20029), .ZN(n20044) );
  NAND2_X1 U22904 ( .A1(n20030), .A2(n20044), .ZN(P1_U2947) );
  AOI22_X1 U22905 ( .A1(n20053), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20052), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n20032) );
  NAND2_X1 U22906 ( .A1(n20038), .A2(n20031), .ZN(n20046) );
  NAND2_X1 U22907 ( .A1(n20032), .A2(n20046), .ZN(P1_U2948) );
  AOI22_X1 U22908 ( .A1(n20053), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20052), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20034) );
  NAND2_X1 U22909 ( .A1(n20038), .A2(n20033), .ZN(n20048) );
  NAND2_X1 U22910 ( .A1(n20034), .A2(n20048), .ZN(P1_U2949) );
  AOI22_X1 U22911 ( .A1(n20053), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20052), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20036) );
  NAND2_X1 U22912 ( .A1(n20038), .A2(n20035), .ZN(n20050) );
  NAND2_X1 U22913 ( .A1(n20036), .A2(n20050), .ZN(P1_U2950) );
  AOI22_X1 U22914 ( .A1(n20053), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20052), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20039) );
  NAND2_X1 U22915 ( .A1(n20038), .A2(n20037), .ZN(n20054) );
  NAND2_X1 U22916 ( .A1(n20039), .A2(n20054), .ZN(P1_U2951) );
  AOI22_X1 U22917 ( .A1(n20053), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20052), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n20041) );
  NAND2_X1 U22918 ( .A1(n20041), .A2(n20040), .ZN(P1_U2960) );
  AOI22_X1 U22919 ( .A1(n20053), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20052), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20043) );
  NAND2_X1 U22920 ( .A1(n20043), .A2(n20042), .ZN(P1_U2961) );
  AOI22_X1 U22921 ( .A1(n20053), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20052), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20045) );
  NAND2_X1 U22922 ( .A1(n20045), .A2(n20044), .ZN(P1_U2962) );
  AOI22_X1 U22923 ( .A1(n20053), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20052), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20047) );
  NAND2_X1 U22924 ( .A1(n20047), .A2(n20046), .ZN(P1_U2963) );
  AOI22_X1 U22925 ( .A1(n20053), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20052), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20049) );
  NAND2_X1 U22926 ( .A1(n20049), .A2(n20048), .ZN(P1_U2964) );
  AOI22_X1 U22927 ( .A1(n20053), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20052), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20051) );
  NAND2_X1 U22928 ( .A1(n20051), .A2(n20050), .ZN(P1_U2965) );
  AOI22_X1 U22929 ( .A1(n20053), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20052), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20055) );
  NAND2_X1 U22930 ( .A1(n20055), .A2(n20054), .ZN(P1_U2966) );
  INV_X1 U22931 ( .A(n20056), .ZN(n20061) );
  OR2_X1 U22932 ( .A1(n20058), .A2(n20057), .ZN(n20059) );
  AOI22_X1 U22933 ( .A1(n20061), .A2(n20060), .B1(n20059), .B2(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20063) );
  OAI211_X1 U22934 ( .C1(n20064), .C2(n20081), .A(n20063), .B(n20062), .ZN(
        P1_U2999) );
  AOI21_X1 U22935 ( .B1(n20067), .B2(n20066), .A(n20065), .ZN(n20068) );
  OAI21_X1 U22936 ( .B1(n20069), .B2(n11573), .A(n20068), .ZN(n20070) );
  AOI21_X1 U22937 ( .B1(n20072), .B2(n20071), .A(n20070), .ZN(n20076) );
  OAI211_X1 U22938 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20074), .B(n20073), .ZN(n20075) );
  NAND2_X1 U22939 ( .A1(n20076), .A2(n20075), .ZN(P1_U3027) );
  NOR2_X1 U22940 ( .A1(n20078), .A2(n20077), .ZN(P1_U3032) );
  NOR2_X2 U22941 ( .A1(n20079), .A2(n20081), .ZN(n20132) );
  NOR2_X2 U22942 ( .A1(n20081), .A2(n20080), .ZN(n20131) );
  AOI22_X1 U22943 ( .A1(DATAI_16_), .A2(n20132), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20131), .ZN(n20578) );
  AOI22_X1 U22944 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20131), .B1(DATAI_24_), 
        .B2(n20132), .ZN(n20628) );
  INV_X1 U22945 ( .A(n20628), .ZN(n20575) );
  NAND2_X1 U22946 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20088), .ZN(n20117) );
  OR2_X1 U22947 ( .A1(n20084), .A2(n20117), .ZN(n20425) );
  NOR2_X1 U22948 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20209) );
  INV_X1 U22949 ( .A(n20507), .ZN(n20085) );
  NAND2_X1 U22950 ( .A1(n20209), .A2(n20085), .ZN(n20135) );
  NOR2_X1 U22951 ( .A1(n20425), .A2(n20135), .ZN(n20086) );
  AOI21_X1 U22952 ( .B1(n20670), .B2(n20575), .A(n20086), .ZN(n20101) );
  INV_X1 U22953 ( .A(n20430), .ZN(n20087) );
  NOR2_X1 U22954 ( .A1(n20087), .A2(n20373), .ZN(n20097) );
  OR2_X1 U22955 ( .A1(n20095), .A2(n20679), .ZN(n20566) );
  AND2_X1 U22956 ( .A1(n20088), .A2(n20566), .ZN(n20433) );
  INV_X1 U22957 ( .A(n20670), .ZN(n20089) );
  NAND2_X1 U22958 ( .A1(n20089), .A2(n20164), .ZN(n20090) );
  AOI21_X1 U22959 ( .B1(n20090), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20620), 
        .ZN(n20094) );
  OR2_X1 U22960 ( .A1(n13328), .A2(n20091), .ZN(n20212) );
  INV_X1 U22961 ( .A(n20212), .ZN(n20175) );
  NAND2_X1 U22962 ( .A1(n20175), .A2(n20372), .ZN(n20098) );
  AOI22_X1 U22963 ( .A1(n20094), .A2(n20098), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20135), .ZN(n20092) );
  OAI211_X1 U22964 ( .C1(n20097), .C2(n20679), .A(n20433), .B(n20092), .ZN(
        n20139) );
  NOR2_X2 U22965 ( .A1(n20093), .A2(n20257), .ZN(n20619) );
  INV_X1 U22966 ( .A(n20094), .ZN(n20099) );
  INV_X1 U22967 ( .A(n20095), .ZN(n20096) );
  NOR2_X1 U22968 ( .A1(n20096), .A2(n20679), .ZN(n20256) );
  INV_X1 U22969 ( .A(n20256), .ZN(n20436) );
  INV_X1 U22970 ( .A(n20097), .ZN(n20251) );
  OAI22_X1 U22971 ( .A1(n20099), .A2(n20098), .B1(n20436), .B2(n20251), .ZN(
        n20138) );
  AOI22_X1 U22972 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20139), .B1(
        n20619), .B2(n20138), .ZN(n20100) );
  OAI211_X1 U22973 ( .C1(n20578), .C2(n20164), .A(n20101), .B(n20100), .ZN(
        P1_U3033) );
  AOI22_X1 U22974 ( .A1(DATAI_17_), .A2(n20132), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20131), .ZN(n20582) );
  AOI22_X1 U22975 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20131), .B1(DATAI_25_), 
        .B2(n20132), .ZN(n20634) );
  INV_X1 U22976 ( .A(n20634), .ZN(n20579) );
  NAND2_X1 U22977 ( .A1(n20102), .A2(n20133), .ZN(n20441) );
  NOR2_X1 U22978 ( .A1(n20441), .A2(n20135), .ZN(n20103) );
  AOI21_X1 U22979 ( .B1(n20670), .B2(n20579), .A(n20103), .ZN(n20106) );
  NOR2_X2 U22980 ( .A1(n20104), .A2(n20257), .ZN(n20630) );
  AOI22_X1 U22981 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20139), .B1(
        n20630), .B2(n20138), .ZN(n20105) );
  OAI211_X1 U22982 ( .C1(n20582), .C2(n20164), .A(n20106), .B(n20105), .ZN(
        P1_U3034) );
  AOI22_X1 U22983 ( .A1(DATAI_18_), .A2(n20132), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20131), .ZN(n20586) );
  AOI22_X1 U22984 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20131), .B1(DATAI_26_), 
        .B2(n20132), .ZN(n20640) );
  INV_X1 U22985 ( .A(n20640), .ZN(n20583) );
  NAND2_X1 U22986 ( .A1(n20107), .A2(n20133), .ZN(n20445) );
  NOR2_X1 U22987 ( .A1(n20445), .A2(n20135), .ZN(n20108) );
  AOI21_X1 U22988 ( .B1(n20670), .B2(n20583), .A(n20108), .ZN(n20111) );
  NOR2_X2 U22989 ( .A1(n20109), .A2(n20257), .ZN(n20636) );
  AOI22_X1 U22990 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20139), .B1(
        n20636), .B2(n20138), .ZN(n20110) );
  OAI211_X1 U22991 ( .C1(n20586), .C2(n20164), .A(n20111), .B(n20110), .ZN(
        P1_U3035) );
  AOI22_X1 U22992 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20131), .B1(DATAI_27_), 
        .B2(n20132), .ZN(n20646) );
  INV_X1 U22993 ( .A(n20646), .ZN(n20587) );
  NAND2_X1 U22994 ( .A1(n20112), .A2(n20133), .ZN(n20449) );
  NOR2_X1 U22995 ( .A1(n20449), .A2(n20135), .ZN(n20113) );
  AOI21_X1 U22996 ( .B1(n20670), .B2(n20587), .A(n20113), .ZN(n20116) );
  NOR2_X2 U22997 ( .A1(n20114), .A2(n20257), .ZN(n20642) );
  AOI22_X1 U22998 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20139), .B1(
        n20642), .B2(n20138), .ZN(n20115) );
  OAI211_X1 U22999 ( .C1(n20590), .C2(n20164), .A(n20116), .B(n20115), .ZN(
        P1_U3036) );
  AOI22_X1 U23000 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20131), .B1(DATAI_28_), 
        .B2(n20132), .ZN(n20652) );
  INV_X1 U23001 ( .A(n20652), .ZN(n20591) );
  OR2_X1 U23002 ( .A1(n11326), .A2(n20117), .ZN(n20453) );
  NOR2_X1 U23003 ( .A1(n20453), .A2(n20135), .ZN(n20118) );
  AOI21_X1 U23004 ( .B1(n20670), .B2(n20591), .A(n20118), .ZN(n20121) );
  NOR2_X2 U23005 ( .A1(n20119), .A2(n20257), .ZN(n20648) );
  AOI22_X1 U23006 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20139), .B1(
        n20648), .B2(n20138), .ZN(n20120) );
  OAI211_X1 U23007 ( .C1(n20594), .C2(n20164), .A(n20121), .B(n20120), .ZN(
        P1_U3037) );
  AOI22_X1 U23008 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20131), .B1(DATAI_29_), 
        .B2(n20132), .ZN(n20658) );
  INV_X1 U23009 ( .A(n20658), .ZN(n20595) );
  NAND2_X1 U23010 ( .A1(n20122), .A2(n20133), .ZN(n20457) );
  NOR2_X1 U23011 ( .A1(n20457), .A2(n20135), .ZN(n20123) );
  AOI21_X1 U23012 ( .B1(n20670), .B2(n20595), .A(n20123), .ZN(n20126) );
  NOR2_X2 U23013 ( .A1(n20124), .A2(n20257), .ZN(n20654) );
  AOI22_X1 U23014 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20139), .B1(
        n20654), .B2(n20138), .ZN(n20125) );
  OAI211_X1 U23015 ( .C1(n20598), .C2(n20164), .A(n20126), .B(n20125), .ZN(
        P1_U3038) );
  AOI22_X1 U23016 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20131), .B1(DATAI_22_), 
        .B2(n20132), .ZN(n20602) );
  AOI22_X1 U23017 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20131), .B1(DATAI_30_), 
        .B2(n20132), .ZN(n20664) );
  INV_X1 U23018 ( .A(n20664), .ZN(n20599) );
  NAND2_X1 U23019 ( .A1(n11695), .A2(n20133), .ZN(n20461) );
  NOR2_X1 U23020 ( .A1(n20461), .A2(n20135), .ZN(n20127) );
  AOI21_X1 U23021 ( .B1(n20670), .B2(n20599), .A(n20127), .ZN(n20130) );
  NOR2_X2 U23022 ( .A1(n20128), .A2(n20257), .ZN(n20660) );
  AOI22_X1 U23023 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20139), .B1(
        n20660), .B2(n20138), .ZN(n20129) );
  OAI211_X1 U23024 ( .C1(n20602), .C2(n20164), .A(n20130), .B(n20129), .ZN(
        P1_U3039) );
  AOI22_X1 U23025 ( .A1(DATAI_31_), .A2(n20132), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20131), .ZN(n20675) );
  INV_X1 U23026 ( .A(n20675), .ZN(n20605) );
  NAND2_X1 U23027 ( .A1(n20134), .A2(n20133), .ZN(n20466) );
  NOR2_X1 U23028 ( .A1(n20466), .A2(n20135), .ZN(n20136) );
  AOI21_X1 U23029 ( .B1(n20670), .B2(n20605), .A(n20136), .ZN(n20141) );
  NOR2_X2 U23030 ( .A1(n20137), .A2(n20257), .ZN(n20668) );
  AOI22_X1 U23031 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20139), .B1(
        n20668), .B2(n20138), .ZN(n20140) );
  OAI211_X1 U23032 ( .C1(n20610), .C2(n20164), .A(n20141), .B(n20140), .ZN(
        P1_U3040) );
  OR2_X1 U23033 ( .A1(n20142), .A2(n20620), .ZN(n20539) );
  INV_X1 U23034 ( .A(n20209), .ZN(n20143) );
  NOR3_X2 U23035 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20536), .A3(
        n20143), .ZN(n20165) );
  INV_X1 U23036 ( .A(n20165), .ZN(n20145) );
  NOR2_X1 U23037 ( .A1(n20143), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20147) );
  INV_X1 U23038 ( .A(n20147), .ZN(n20144) );
  OAI222_X1 U23039 ( .A1(n20212), .A2(n20539), .B1(n20145), .B2(n20620), .C1(
        n20679), .C2(n20144), .ZN(n20166) );
  AOI22_X1 U23040 ( .A1(n20619), .A2(n20166), .B1(n20618), .B2(n20165), .ZN(
        n20150) );
  INV_X1 U23041 ( .A(n20146), .ZN(n20400) );
  NOR2_X1 U23042 ( .A1(n20214), .A2(n20400), .ZN(n20148) );
  OAI21_X1 U23043 ( .B1(n20148), .B2(n20147), .A(n20622), .ZN(n20168) );
  INV_X1 U23044 ( .A(n20164), .ZN(n20167) );
  AOI22_X1 U23045 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20168), .B1(
        n20167), .B2(n20575), .ZN(n20149) );
  OAI211_X1 U23046 ( .C1(n20578), .C2(n20206), .A(n20150), .B(n20149), .ZN(
        P1_U3041) );
  AOI22_X1 U23047 ( .A1(n20630), .A2(n20166), .B1(n20629), .B2(n20165), .ZN(
        n20152) );
  AOI22_X1 U23048 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20168), .B1(
        n20167), .B2(n20579), .ZN(n20151) );
  OAI211_X1 U23049 ( .C1(n20582), .C2(n20206), .A(n20152), .B(n20151), .ZN(
        P1_U3042) );
  AOI22_X1 U23050 ( .A1(n20636), .A2(n20166), .B1(n20635), .B2(n20165), .ZN(
        n20154) );
  INV_X1 U23051 ( .A(n20206), .ZN(n20161) );
  INV_X1 U23052 ( .A(n20586), .ZN(n20637) );
  AOI22_X1 U23053 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20168), .B1(
        n20161), .B2(n20637), .ZN(n20153) );
  OAI211_X1 U23054 ( .C1(n20640), .C2(n20164), .A(n20154), .B(n20153), .ZN(
        P1_U3043) );
  AOI22_X1 U23055 ( .A1(n20642), .A2(n20166), .B1(n20641), .B2(n20165), .ZN(
        n20156) );
  AOI22_X1 U23056 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20168), .B1(
        n20167), .B2(n20587), .ZN(n20155) );
  OAI211_X1 U23057 ( .C1(n20590), .C2(n20206), .A(n20156), .B(n20155), .ZN(
        P1_U3044) );
  AOI22_X1 U23058 ( .A1(n20648), .A2(n20166), .B1(n20647), .B2(n20165), .ZN(
        n20158) );
  AOI22_X1 U23059 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20168), .B1(
        n20167), .B2(n20591), .ZN(n20157) );
  OAI211_X1 U23060 ( .C1(n20594), .C2(n20206), .A(n20158), .B(n20157), .ZN(
        P1_U3045) );
  AOI22_X1 U23061 ( .A1(n20654), .A2(n20166), .B1(n20653), .B2(n20165), .ZN(
        n20160) );
  AOI22_X1 U23062 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20168), .B1(
        n20167), .B2(n20595), .ZN(n20159) );
  OAI211_X1 U23063 ( .C1(n20598), .C2(n20206), .A(n20160), .B(n20159), .ZN(
        P1_U3046) );
  AOI22_X1 U23064 ( .A1(n20660), .A2(n20166), .B1(n20659), .B2(n20165), .ZN(
        n20163) );
  INV_X1 U23065 ( .A(n20602), .ZN(n20661) );
  AOI22_X1 U23066 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20168), .B1(
        n20161), .B2(n20661), .ZN(n20162) );
  OAI211_X1 U23067 ( .C1(n20664), .C2(n20164), .A(n20163), .B(n20162), .ZN(
        P1_U3047) );
  AOI22_X1 U23068 ( .A1(n20668), .A2(n20166), .B1(n20666), .B2(n20165), .ZN(
        n20170) );
  AOI22_X1 U23069 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20168), .B1(
        n20167), .B2(n20605), .ZN(n20169) );
  OAI211_X1 U23070 ( .C1(n20610), .C2(n20206), .A(n20170), .B(n20169), .ZN(
        P1_U3048) );
  NAND2_X1 U23071 ( .A1(n20172), .A2(n20171), .ZN(n20424) );
  NAND3_X1 U23072 ( .A1(n20536), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        n20209), .ZN(n20200) );
  OAI22_X1 U23073 ( .A1(n20206), .A2(n20628), .B1(n20425), .B2(n20200), .ZN(
        n20173) );
  INV_X1 U23074 ( .A(n20173), .ZN(n20181) );
  NAND2_X1 U23075 ( .A1(n20242), .A2(n20206), .ZN(n20174) );
  AOI21_X1 U23076 ( .B1(n20174), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20620), 
        .ZN(n20177) );
  NAND2_X1 U23077 ( .A1(n20175), .A2(n11447), .ZN(n20178) );
  AOI22_X1 U23078 ( .A1(n20177), .A2(n20178), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20200), .ZN(n20176) );
  OR2_X1 U23079 ( .A1(n20430), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20310) );
  NAND2_X1 U23080 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20310), .ZN(n20307) );
  NAND3_X1 U23081 ( .A1(n20433), .A2(n20176), .A3(n20307), .ZN(n20203) );
  INV_X1 U23082 ( .A(n20177), .ZN(n20179) );
  OAI22_X1 U23083 ( .A1(n20179), .A2(n20178), .B1(n20310), .B2(n20436), .ZN(
        n20202) );
  AOI22_X1 U23084 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20203), .B1(
        n20619), .B2(n20202), .ZN(n20180) );
  OAI211_X1 U23085 ( .C1(n20578), .C2(n20242), .A(n20181), .B(n20180), .ZN(
        P1_U3049) );
  OAI22_X1 U23086 ( .A1(n20206), .A2(n20634), .B1(n20441), .B2(n20200), .ZN(
        n20182) );
  INV_X1 U23087 ( .A(n20182), .ZN(n20184) );
  AOI22_X1 U23088 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20203), .B1(
        n20630), .B2(n20202), .ZN(n20183) );
  OAI211_X1 U23089 ( .C1(n20582), .C2(n20242), .A(n20184), .B(n20183), .ZN(
        P1_U3050) );
  OAI22_X1 U23090 ( .A1(n20206), .A2(n20640), .B1(n20445), .B2(n20200), .ZN(
        n20185) );
  INV_X1 U23091 ( .A(n20185), .ZN(n20187) );
  AOI22_X1 U23092 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20203), .B1(
        n20636), .B2(n20202), .ZN(n20186) );
  OAI211_X1 U23093 ( .C1(n20586), .C2(n20242), .A(n20187), .B(n20186), .ZN(
        P1_U3051) );
  OAI22_X1 U23094 ( .A1(n20242), .A2(n20590), .B1(n20449), .B2(n20200), .ZN(
        n20188) );
  INV_X1 U23095 ( .A(n20188), .ZN(n20190) );
  AOI22_X1 U23096 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20203), .B1(
        n20642), .B2(n20202), .ZN(n20189) );
  OAI211_X1 U23097 ( .C1(n20646), .C2(n20206), .A(n20190), .B(n20189), .ZN(
        P1_U3052) );
  OAI22_X1 U23098 ( .A1(n20242), .A2(n20594), .B1(n20453), .B2(n20200), .ZN(
        n20191) );
  INV_X1 U23099 ( .A(n20191), .ZN(n20193) );
  AOI22_X1 U23100 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20203), .B1(
        n20648), .B2(n20202), .ZN(n20192) );
  OAI211_X1 U23101 ( .C1(n20652), .C2(n20206), .A(n20193), .B(n20192), .ZN(
        P1_U3053) );
  OAI22_X1 U23102 ( .A1(n20242), .A2(n20598), .B1(n20457), .B2(n20200), .ZN(
        n20194) );
  INV_X1 U23103 ( .A(n20194), .ZN(n20196) );
  AOI22_X1 U23104 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20203), .B1(
        n20654), .B2(n20202), .ZN(n20195) );
  OAI211_X1 U23105 ( .C1(n20658), .C2(n20206), .A(n20196), .B(n20195), .ZN(
        P1_U3054) );
  OAI22_X1 U23106 ( .A1(n20242), .A2(n20602), .B1(n20461), .B2(n20200), .ZN(
        n20197) );
  INV_X1 U23107 ( .A(n20197), .ZN(n20199) );
  AOI22_X1 U23108 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20203), .B1(
        n20660), .B2(n20202), .ZN(n20198) );
  OAI211_X1 U23109 ( .C1(n20664), .C2(n20206), .A(n20199), .B(n20198), .ZN(
        P1_U3055) );
  OAI22_X1 U23110 ( .A1(n20242), .A2(n20610), .B1(n20466), .B2(n20200), .ZN(
        n20201) );
  INV_X1 U23111 ( .A(n20201), .ZN(n20205) );
  AOI22_X1 U23112 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20203), .B1(
        n20668), .B2(n20202), .ZN(n20204) );
  OAI211_X1 U23113 ( .C1(n20675), .C2(n20206), .A(n20205), .B(n20204), .ZN(
        P1_U3056) );
  INV_X1 U23114 ( .A(n20482), .ZN(n20347) );
  NAND2_X1 U23115 ( .A1(n20209), .A2(n20207), .ZN(n20241) );
  OAI22_X1 U23116 ( .A1(n20252), .A2(n20578), .B1(n20425), .B2(n20241), .ZN(
        n20208) );
  INV_X1 U23117 ( .A(n20208), .ZN(n20222) );
  NAND2_X1 U23118 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20209), .ZN(
        n20218) );
  AND2_X1 U23119 ( .A1(n11712), .A2(n20210), .ZN(n20612) );
  INV_X1 U23120 ( .A(n20612), .ZN(n20211) );
  OR2_X1 U23121 ( .A1(n20212), .A2(n20211), .ZN(n20213) );
  AND2_X1 U23122 ( .A1(n20213), .A2(n20241), .ZN(n20220) );
  INV_X1 U23123 ( .A(n20220), .ZN(n20215) );
  OAI21_X1 U23124 ( .B1(n20214), .B2(n20477), .A(n20481), .ZN(n20219) );
  OAI21_X1 U23125 ( .B1(n20215), .B2(n20219), .A(n20622), .ZN(n20216) );
  AOI21_X1 U23126 ( .B1(n20620), .B2(n20218), .A(n20216), .ZN(n20217) );
  OAI22_X1 U23127 ( .A1(n20220), .A2(n20219), .B1(n20679), .B2(n20218), .ZN(
        n20244) );
  AOI22_X1 U23128 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20245), .B1(
        n20619), .B2(n20244), .ZN(n20221) );
  OAI211_X1 U23129 ( .C1(n20628), .C2(n20242), .A(n20222), .B(n20221), .ZN(
        P1_U3057) );
  OAI22_X1 U23130 ( .A1(n20242), .A2(n20634), .B1(n20441), .B2(n20241), .ZN(
        n20223) );
  INV_X1 U23131 ( .A(n20223), .ZN(n20225) );
  AOI22_X1 U23132 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20245), .B1(
        n20630), .B2(n20244), .ZN(n20224) );
  OAI211_X1 U23133 ( .C1(n20582), .C2(n20252), .A(n20225), .B(n20224), .ZN(
        P1_U3058) );
  OAI22_X1 U23134 ( .A1(n20242), .A2(n20640), .B1(n20445), .B2(n20241), .ZN(
        n20226) );
  INV_X1 U23135 ( .A(n20226), .ZN(n20228) );
  AOI22_X1 U23136 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20245), .B1(
        n20636), .B2(n20244), .ZN(n20227) );
  OAI211_X1 U23137 ( .C1(n20586), .C2(n20252), .A(n20228), .B(n20227), .ZN(
        P1_U3059) );
  OAI22_X1 U23138 ( .A1(n20252), .A2(n20590), .B1(n20449), .B2(n20241), .ZN(
        n20229) );
  INV_X1 U23139 ( .A(n20229), .ZN(n20231) );
  AOI22_X1 U23140 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20245), .B1(
        n20642), .B2(n20244), .ZN(n20230) );
  OAI211_X1 U23141 ( .C1(n20646), .C2(n20242), .A(n20231), .B(n20230), .ZN(
        P1_U3060) );
  OAI22_X1 U23142 ( .A1(n20242), .A2(n20652), .B1(n20453), .B2(n20241), .ZN(
        n20232) );
  INV_X1 U23143 ( .A(n20232), .ZN(n20234) );
  AOI22_X1 U23144 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20245), .B1(
        n20648), .B2(n20244), .ZN(n20233) );
  OAI211_X1 U23145 ( .C1(n20594), .C2(n20252), .A(n20234), .B(n20233), .ZN(
        P1_U3061) );
  OAI22_X1 U23146 ( .A1(n20252), .A2(n20598), .B1(n20457), .B2(n20241), .ZN(
        n20235) );
  INV_X1 U23147 ( .A(n20235), .ZN(n20237) );
  AOI22_X1 U23148 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20245), .B1(
        n20654), .B2(n20244), .ZN(n20236) );
  OAI211_X1 U23149 ( .C1(n20658), .C2(n20242), .A(n20237), .B(n20236), .ZN(
        P1_U3062) );
  OAI22_X1 U23150 ( .A1(n20242), .A2(n20664), .B1(n20461), .B2(n20241), .ZN(
        n20238) );
  INV_X1 U23151 ( .A(n20238), .ZN(n20240) );
  AOI22_X1 U23152 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20245), .B1(
        n20660), .B2(n20244), .ZN(n20239) );
  OAI211_X1 U23153 ( .C1(n20602), .C2(n20252), .A(n20240), .B(n20239), .ZN(
        P1_U3063) );
  OAI22_X1 U23154 ( .A1(n20242), .A2(n20675), .B1(n20466), .B2(n20241), .ZN(
        n20243) );
  INV_X1 U23155 ( .A(n20243), .ZN(n20247) );
  AOI22_X1 U23156 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20245), .B1(
        n20668), .B2(n20244), .ZN(n20246) );
  OAI211_X1 U23157 ( .C1(n20610), .C2(n20252), .A(n20247), .B(n20246), .ZN(
        P1_U3064) );
  INV_X1 U23158 ( .A(n20348), .ZN(n20249) );
  NOR2_X1 U23159 ( .A1(n13572), .A2(n20250), .ZN(n20341) );
  NAND2_X1 U23160 ( .A1(n20341), .A2(n20372), .ZN(n20254) );
  OAI22_X1 U23161 ( .A1(n20254), .A2(n20620), .B1(n20251), .B2(n20566), .ZN(
        n20273) );
  AOI22_X1 U23162 ( .A1(n20619), .A2(n20273), .B1(n20618), .B2(n9682), .ZN(
        n20260) );
  INV_X1 U23163 ( .A(n20303), .ZN(n20253) );
  OAI21_X1 U23164 ( .B1(n20274), .B2(n20253), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20255) );
  NAND2_X1 U23165 ( .A1(n20255), .A2(n20254), .ZN(n20258) );
  NOR2_X1 U23166 ( .A1(n20257), .A2(n20256), .ZN(n20573) );
  OAI221_X1 U23167 ( .B1(n9682), .B2(n20841), .C1(n9682), .C2(n20258), .A(
        n20573), .ZN(n20275) );
  AOI22_X1 U23168 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20275), .B1(
        n20274), .B2(n20575), .ZN(n20259) );
  OAI211_X1 U23169 ( .C1(n20578), .C2(n20303), .A(n20260), .B(n20259), .ZN(
        P1_U3065) );
  AOI22_X1 U23170 ( .A1(n20630), .A2(n20273), .B1(n20629), .B2(n9682), .ZN(
        n20262) );
  AOI22_X1 U23171 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20275), .B1(
        n20274), .B2(n20579), .ZN(n20261) );
  OAI211_X1 U23172 ( .C1(n20582), .C2(n20303), .A(n20262), .B(n20261), .ZN(
        P1_U3066) );
  AOI22_X1 U23173 ( .A1(n20636), .A2(n20273), .B1(n20635), .B2(n9682), .ZN(
        n20264) );
  AOI22_X1 U23174 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20275), .B1(
        n20274), .B2(n20583), .ZN(n20263) );
  OAI211_X1 U23175 ( .C1(n20586), .C2(n20303), .A(n20264), .B(n20263), .ZN(
        P1_U3067) );
  AOI22_X1 U23176 ( .A1(n20642), .A2(n20273), .B1(n20641), .B2(n9682), .ZN(
        n20266) );
  AOI22_X1 U23177 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20275), .B1(
        n20274), .B2(n20587), .ZN(n20265) );
  OAI211_X1 U23178 ( .C1(n20590), .C2(n20303), .A(n20266), .B(n20265), .ZN(
        P1_U3068) );
  AOI22_X1 U23179 ( .A1(n20648), .A2(n20273), .B1(n20647), .B2(n9682), .ZN(
        n20268) );
  AOI22_X1 U23180 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20275), .B1(
        n20274), .B2(n20591), .ZN(n20267) );
  OAI211_X1 U23181 ( .C1(n20594), .C2(n20303), .A(n20268), .B(n20267), .ZN(
        P1_U3069) );
  AOI22_X1 U23182 ( .A1(n20654), .A2(n20273), .B1(n20653), .B2(n9682), .ZN(
        n20270) );
  AOI22_X1 U23183 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20275), .B1(
        n20274), .B2(n20595), .ZN(n20269) );
  OAI211_X1 U23184 ( .C1(n20598), .C2(n20303), .A(n20270), .B(n20269), .ZN(
        P1_U3070) );
  AOI22_X1 U23185 ( .A1(n20660), .A2(n20273), .B1(n20659), .B2(n9682), .ZN(
        n20272) );
  AOI22_X1 U23186 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20275), .B1(
        n20274), .B2(n20599), .ZN(n20271) );
  OAI211_X1 U23187 ( .C1(n20602), .C2(n20303), .A(n20272), .B(n20271), .ZN(
        P1_U3071) );
  AOI22_X1 U23188 ( .A1(n20668), .A2(n20273), .B1(n20666), .B2(n9682), .ZN(
        n20277) );
  AOI22_X1 U23189 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20275), .B1(
        n20274), .B2(n20605), .ZN(n20276) );
  OAI211_X1 U23190 ( .C1(n20610), .C2(n20303), .A(n20277), .B(n20276), .ZN(
        P1_U3072) );
  INV_X1 U23191 ( .A(n20142), .ZN(n20278) );
  NOR2_X1 U23192 ( .A1(n20304), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20282) );
  INV_X1 U23193 ( .A(n20282), .ZN(n20279) );
  NOR2_X1 U23194 ( .A1(n20536), .A2(n20279), .ZN(n20297) );
  AOI21_X1 U23195 ( .B1(n20341), .B2(n20278), .A(n20297), .ZN(n20280) );
  OAI22_X1 U23196 ( .A1(n20280), .A2(n20620), .B1(n20279), .B2(n20679), .ZN(
        n20298) );
  AOI22_X1 U23197 ( .A1(n20619), .A2(n20298), .B1(n20618), .B2(n20297), .ZN(
        n20284) );
  OAI21_X1 U23198 ( .B1(n20348), .B2(n20777), .A(n20280), .ZN(n20281) );
  OAI221_X1 U23199 ( .B1(n20481), .B2(n20282), .C1(n20620), .C2(n20281), .A(
        n20622), .ZN(n20300) );
  INV_X1 U23200 ( .A(n20578), .ZN(n20625) );
  AOI22_X1 U23201 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20300), .B1(
        n20299), .B2(n20625), .ZN(n20283) );
  OAI211_X1 U23202 ( .C1(n20628), .C2(n20303), .A(n20284), .B(n20283), .ZN(
        P1_U3073) );
  AOI22_X1 U23203 ( .A1(n20630), .A2(n20298), .B1(n20629), .B2(n20297), .ZN(
        n20286) );
  INV_X1 U23204 ( .A(n20582), .ZN(n20631) );
  AOI22_X1 U23205 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20300), .B1(
        n20299), .B2(n20631), .ZN(n20285) );
  OAI211_X1 U23206 ( .C1(n20634), .C2(n20303), .A(n20286), .B(n20285), .ZN(
        P1_U3074) );
  AOI22_X1 U23207 ( .A1(n20636), .A2(n20298), .B1(n20635), .B2(n20297), .ZN(
        n20288) );
  AOI22_X1 U23208 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20300), .B1(
        n20299), .B2(n20637), .ZN(n20287) );
  OAI211_X1 U23209 ( .C1(n20640), .C2(n20303), .A(n20288), .B(n20287), .ZN(
        P1_U3075) );
  AOI22_X1 U23210 ( .A1(n20642), .A2(n20298), .B1(n20641), .B2(n20297), .ZN(
        n20290) );
  INV_X1 U23211 ( .A(n20590), .ZN(n20643) );
  AOI22_X1 U23212 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20300), .B1(
        n20299), .B2(n20643), .ZN(n20289) );
  OAI211_X1 U23213 ( .C1(n20646), .C2(n20303), .A(n20290), .B(n20289), .ZN(
        P1_U3076) );
  AOI22_X1 U23214 ( .A1(n20648), .A2(n20298), .B1(n20647), .B2(n20297), .ZN(
        n20292) );
  INV_X1 U23215 ( .A(n20594), .ZN(n20649) );
  AOI22_X1 U23216 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20300), .B1(
        n20299), .B2(n20649), .ZN(n20291) );
  OAI211_X1 U23217 ( .C1(n20652), .C2(n20303), .A(n20292), .B(n20291), .ZN(
        P1_U3077) );
  AOI22_X1 U23218 ( .A1(n20654), .A2(n20298), .B1(n20653), .B2(n20297), .ZN(
        n20294) );
  INV_X1 U23219 ( .A(n20598), .ZN(n20655) );
  AOI22_X1 U23220 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20300), .B1(
        n20299), .B2(n20655), .ZN(n20293) );
  OAI211_X1 U23221 ( .C1(n20658), .C2(n20303), .A(n20294), .B(n20293), .ZN(
        P1_U3078) );
  AOI22_X1 U23222 ( .A1(n20660), .A2(n20298), .B1(n20659), .B2(n20297), .ZN(
        n20296) );
  AOI22_X1 U23223 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20300), .B1(
        n20299), .B2(n20661), .ZN(n20295) );
  OAI211_X1 U23224 ( .C1(n20664), .C2(n20303), .A(n20296), .B(n20295), .ZN(
        P1_U3079) );
  AOI22_X1 U23225 ( .A1(n20668), .A2(n20298), .B1(n20666), .B2(n20297), .ZN(
        n20302) );
  INV_X1 U23226 ( .A(n20610), .ZN(n20669) );
  AOI22_X1 U23227 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20300), .B1(
        n20299), .B2(n20669), .ZN(n20301) );
  OAI211_X1 U23228 ( .C1(n20675), .C2(n20303), .A(n20302), .B(n20301), .ZN(
        P1_U3080) );
  NOR2_X1 U23229 ( .A1(n20615), .A2(n20304), .ZN(n20346) );
  NAND2_X1 U23230 ( .A1(n20536), .A2(n20346), .ZN(n20333) );
  OAI22_X1 U23231 ( .A1(n20334), .A2(n20628), .B1(n20425), .B2(n20333), .ZN(
        n20305) );
  INV_X1 U23232 ( .A(n20305), .ZN(n20314) );
  NAND2_X1 U23233 ( .A1(n20370), .A2(n20334), .ZN(n20306) );
  AOI21_X1 U23234 ( .B1(n20306), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20620), 
        .ZN(n20309) );
  NAND2_X1 U23235 ( .A1(n20341), .A2(n11447), .ZN(n20311) );
  AOI22_X1 U23236 ( .A1(n20309), .A2(n20311), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20333), .ZN(n20308) );
  NAND3_X1 U23237 ( .A1(n20573), .A2(n20308), .A3(n20307), .ZN(n20337) );
  INV_X1 U23238 ( .A(n20309), .ZN(n20312) );
  OAI22_X1 U23239 ( .A1(n20312), .A2(n20311), .B1(n20566), .B2(n20310), .ZN(
        n20336) );
  AOI22_X1 U23240 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20337), .B1(
        n20619), .B2(n20336), .ZN(n20313) );
  OAI211_X1 U23241 ( .C1(n20578), .C2(n20370), .A(n20314), .B(n20313), .ZN(
        P1_U3081) );
  OAI22_X1 U23242 ( .A1(n20334), .A2(n20634), .B1(n20333), .B2(n20441), .ZN(
        n20315) );
  INV_X1 U23243 ( .A(n20315), .ZN(n20317) );
  AOI22_X1 U23244 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20337), .B1(
        n20630), .B2(n20336), .ZN(n20316) );
  OAI211_X1 U23245 ( .C1(n20582), .C2(n20370), .A(n20317), .B(n20316), .ZN(
        P1_U3082) );
  OAI22_X1 U23246 ( .A1(n20334), .A2(n20640), .B1(n20333), .B2(n20445), .ZN(
        n20318) );
  INV_X1 U23247 ( .A(n20318), .ZN(n20320) );
  AOI22_X1 U23248 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20337), .B1(
        n20636), .B2(n20336), .ZN(n20319) );
  OAI211_X1 U23249 ( .C1(n20586), .C2(n20370), .A(n20320), .B(n20319), .ZN(
        P1_U3083) );
  OAI22_X1 U23250 ( .A1(n20370), .A2(n20590), .B1(n20333), .B2(n20449), .ZN(
        n20321) );
  INV_X1 U23251 ( .A(n20321), .ZN(n20323) );
  AOI22_X1 U23252 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20337), .B1(
        n20642), .B2(n20336), .ZN(n20322) );
  OAI211_X1 U23253 ( .C1(n20646), .C2(n20334), .A(n20323), .B(n20322), .ZN(
        P1_U3084) );
  OAI22_X1 U23254 ( .A1(n20334), .A2(n20652), .B1(n20333), .B2(n20453), .ZN(
        n20324) );
  INV_X1 U23255 ( .A(n20324), .ZN(n20326) );
  AOI22_X1 U23256 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20337), .B1(
        n20648), .B2(n20336), .ZN(n20325) );
  OAI211_X1 U23257 ( .C1(n20594), .C2(n20370), .A(n20326), .B(n20325), .ZN(
        P1_U3085) );
  OAI22_X1 U23258 ( .A1(n20334), .A2(n20658), .B1(n20333), .B2(n20457), .ZN(
        n20327) );
  INV_X1 U23259 ( .A(n20327), .ZN(n20329) );
  AOI22_X1 U23260 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20337), .B1(
        n20654), .B2(n20336), .ZN(n20328) );
  OAI211_X1 U23261 ( .C1(n20598), .C2(n20370), .A(n20329), .B(n20328), .ZN(
        P1_U3086) );
  OAI22_X1 U23262 ( .A1(n20370), .A2(n20602), .B1(n20333), .B2(n20461), .ZN(
        n20330) );
  INV_X1 U23263 ( .A(n20330), .ZN(n20332) );
  AOI22_X1 U23264 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20337), .B1(
        n20660), .B2(n20336), .ZN(n20331) );
  OAI211_X1 U23265 ( .C1(n20664), .C2(n20334), .A(n20332), .B(n20331), .ZN(
        P1_U3087) );
  OAI22_X1 U23266 ( .A1(n20334), .A2(n20675), .B1(n20333), .B2(n20466), .ZN(
        n20335) );
  INV_X1 U23267 ( .A(n20335), .ZN(n20339) );
  AOI22_X1 U23268 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20337), .B1(
        n20668), .B2(n20336), .ZN(n20338) );
  OAI211_X1 U23269 ( .C1(n20610), .C2(n20370), .A(n20339), .B(n20338), .ZN(
        P1_U3088) );
  INV_X1 U23270 ( .A(n20340), .ZN(n20365) );
  AOI21_X1 U23271 ( .B1(n20341), .B2(n20612), .A(n20365), .ZN(n20344) );
  INV_X1 U23272 ( .A(n20346), .ZN(n20342) );
  OAI22_X1 U23273 ( .A1(n20344), .A2(n20620), .B1(n20342), .B2(n20679), .ZN(
        n20366) );
  AOI22_X1 U23274 ( .A1(n20619), .A2(n20366), .B1(n20365), .B2(n20618), .ZN(
        n20350) );
  INV_X1 U23275 ( .A(n20477), .ZN(n20343) );
  NAND2_X1 U23276 ( .A1(n9587), .A2(n20343), .ZN(n20621) );
  OAI211_X1 U23277 ( .C1(n11721), .C2(n20621), .A(n20481), .B(n20344), .ZN(
        n20345) );
  OAI211_X1 U23278 ( .C1(n20481), .C2(n20346), .A(n20622), .B(n20345), .ZN(
        n20367) );
  AOI22_X1 U23279 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20367), .B1(
        n20393), .B2(n20625), .ZN(n20349) );
  OAI211_X1 U23280 ( .C1(n20628), .C2(n20370), .A(n20350), .B(n20349), .ZN(
        P1_U3089) );
  AOI22_X1 U23281 ( .A1(n20630), .A2(n20366), .B1(n20365), .B2(n20629), .ZN(
        n20352) );
  AOI22_X1 U23282 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20367), .B1(
        n20393), .B2(n20631), .ZN(n20351) );
  OAI211_X1 U23283 ( .C1(n20634), .C2(n20370), .A(n20352), .B(n20351), .ZN(
        P1_U3090) );
  AOI22_X1 U23284 ( .A1(n20636), .A2(n20366), .B1(n20365), .B2(n20635), .ZN(
        n20354) );
  AOI22_X1 U23285 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20367), .B1(
        n20393), .B2(n20637), .ZN(n20353) );
  OAI211_X1 U23286 ( .C1(n20640), .C2(n20370), .A(n20354), .B(n20353), .ZN(
        P1_U3091) );
  AOI22_X1 U23287 ( .A1(n20642), .A2(n20366), .B1(n20365), .B2(n20641), .ZN(
        n20356) );
  INV_X1 U23288 ( .A(n20370), .ZN(n20361) );
  AOI22_X1 U23289 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20367), .B1(
        n20361), .B2(n20587), .ZN(n20355) );
  OAI211_X1 U23290 ( .C1(n20590), .C2(n20364), .A(n20356), .B(n20355), .ZN(
        P1_U3092) );
  AOI22_X1 U23291 ( .A1(n20648), .A2(n20366), .B1(n20365), .B2(n20647), .ZN(
        n20358) );
  AOI22_X1 U23292 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20367), .B1(
        n20361), .B2(n20591), .ZN(n20357) );
  OAI211_X1 U23293 ( .C1(n20594), .C2(n20364), .A(n20358), .B(n20357), .ZN(
        P1_U3093) );
  AOI22_X1 U23294 ( .A1(n20654), .A2(n20366), .B1(n20365), .B2(n20653), .ZN(
        n20360) );
  AOI22_X1 U23295 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20367), .B1(
        n20361), .B2(n20595), .ZN(n20359) );
  OAI211_X1 U23296 ( .C1(n20598), .C2(n20364), .A(n20360), .B(n20359), .ZN(
        P1_U3094) );
  AOI22_X1 U23297 ( .A1(n20660), .A2(n20366), .B1(n20365), .B2(n20659), .ZN(
        n20363) );
  AOI22_X1 U23298 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20367), .B1(
        n20361), .B2(n20599), .ZN(n20362) );
  OAI211_X1 U23299 ( .C1(n20602), .C2(n20364), .A(n20363), .B(n20362), .ZN(
        P1_U3095) );
  AOI22_X1 U23300 ( .A1(n20668), .A2(n20366), .B1(n20365), .B2(n20666), .ZN(
        n20369) );
  AOI22_X1 U23301 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20367), .B1(
        n20393), .B2(n20669), .ZN(n20368) );
  OAI211_X1 U23302 ( .C1(n20675), .C2(n20370), .A(n20369), .B(n20368), .ZN(
        P1_U3096) );
  AND2_X1 U23303 ( .A1(n13328), .A2(n13572), .ZN(n20474) );
  NAND2_X1 U23304 ( .A1(n20371), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20473) );
  AOI21_X1 U23305 ( .B1(n20474), .B2(n20372), .A(n10064), .ZN(n20375) );
  NAND2_X1 U23306 ( .A1(n20373), .A2(n20430), .ZN(n20513) );
  OAI22_X1 U23307 ( .A1(n20375), .A2(n20620), .B1(n20513), .B2(n20436), .ZN(
        n20392) );
  AOI22_X1 U23308 ( .A1(n20619), .A2(n20392), .B1(n10064), .B2(n20618), .ZN(
        n20379) );
  INV_X1 U23309 ( .A(n20423), .ZN(n20374) );
  OAI21_X1 U23310 ( .B1(n20374), .B2(n20393), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20376) );
  NAND2_X1 U23311 ( .A1(n20376), .A2(n20375), .ZN(n20377) );
  OAI211_X1 U23312 ( .C1(n10064), .C2(n20841), .A(n20433), .B(n20377), .ZN(
        n20394) );
  AOI22_X1 U23313 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20394), .B1(
        n20393), .B2(n20575), .ZN(n20378) );
  OAI211_X1 U23314 ( .C1(n20578), .C2(n20423), .A(n20379), .B(n20378), .ZN(
        P1_U3097) );
  AOI22_X1 U23315 ( .A1(n20630), .A2(n20392), .B1(n10064), .B2(n20629), .ZN(
        n20381) );
  AOI22_X1 U23316 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20394), .B1(
        n20393), .B2(n20579), .ZN(n20380) );
  OAI211_X1 U23317 ( .C1(n20582), .C2(n20423), .A(n20381), .B(n20380), .ZN(
        P1_U3098) );
  AOI22_X1 U23318 ( .A1(n20636), .A2(n20392), .B1(n10064), .B2(n20635), .ZN(
        n20383) );
  AOI22_X1 U23319 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20394), .B1(
        n20393), .B2(n20583), .ZN(n20382) );
  OAI211_X1 U23320 ( .C1(n20586), .C2(n20423), .A(n20383), .B(n20382), .ZN(
        P1_U3099) );
  AOI22_X1 U23321 ( .A1(n20642), .A2(n20392), .B1(n10064), .B2(n20641), .ZN(
        n20385) );
  AOI22_X1 U23322 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20394), .B1(
        n20393), .B2(n20587), .ZN(n20384) );
  OAI211_X1 U23323 ( .C1(n20590), .C2(n20423), .A(n20385), .B(n20384), .ZN(
        P1_U3100) );
  AOI22_X1 U23324 ( .A1(n20648), .A2(n20392), .B1(n10064), .B2(n20647), .ZN(
        n20387) );
  AOI22_X1 U23325 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20394), .B1(
        n20393), .B2(n20591), .ZN(n20386) );
  OAI211_X1 U23326 ( .C1(n20594), .C2(n20423), .A(n20387), .B(n20386), .ZN(
        P1_U3101) );
  AOI22_X1 U23327 ( .A1(n20654), .A2(n20392), .B1(n10064), .B2(n20653), .ZN(
        n20389) );
  AOI22_X1 U23328 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20394), .B1(
        n20393), .B2(n20595), .ZN(n20388) );
  OAI211_X1 U23329 ( .C1(n20598), .C2(n20423), .A(n20389), .B(n20388), .ZN(
        P1_U3102) );
  AOI22_X1 U23330 ( .A1(n20660), .A2(n20392), .B1(n10064), .B2(n20659), .ZN(
        n20391) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20394), .B1(
        n20393), .B2(n20599), .ZN(n20390) );
  OAI211_X1 U23332 ( .C1(n20602), .C2(n20423), .A(n20391), .B(n20390), .ZN(
        P1_U3103) );
  AOI22_X1 U23333 ( .A1(n20668), .A2(n20392), .B1(n10064), .B2(n20666), .ZN(
        n20396) );
  AOI22_X1 U23334 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20394), .B1(
        n20393), .B2(n20605), .ZN(n20395) );
  OAI211_X1 U23335 ( .C1(n20610), .C2(n20423), .A(n20396), .B(n20395), .ZN(
        P1_U3104) );
  INV_X1 U23336 ( .A(n20474), .ZN(n20399) );
  NOR2_X1 U23337 ( .A1(n20473), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20401) );
  INV_X1 U23338 ( .A(n20401), .ZN(n20397) );
  NOR2_X1 U23339 ( .A1(n20536), .A2(n20397), .ZN(n20418) );
  INV_X1 U23340 ( .A(n20418), .ZN(n20398) );
  OAI222_X1 U23341 ( .A1(n20399), .A2(n20539), .B1(n20398), .B2(n20620), .C1(
        n20679), .C2(n20397), .ZN(n20419) );
  AOI22_X1 U23342 ( .A1(n20619), .A2(n20419), .B1(n20618), .B2(n20418), .ZN(
        n20405) );
  INV_X1 U23343 ( .A(n20483), .ZN(n20478) );
  NOR2_X1 U23344 ( .A1(n20478), .A2(n20400), .ZN(n20402) );
  OAI21_X1 U23345 ( .B1(n20402), .B2(n20401), .A(n20622), .ZN(n20420) );
  AOI22_X1 U23346 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20420), .B1(
        n20427), .B2(n20625), .ZN(n20404) );
  OAI211_X1 U23347 ( .C1(n20628), .C2(n20423), .A(n20405), .B(n20404), .ZN(
        P1_U3105) );
  AOI22_X1 U23348 ( .A1(n20630), .A2(n20419), .B1(n20629), .B2(n20418), .ZN(
        n20407) );
  AOI22_X1 U23349 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20420), .B1(
        n20427), .B2(n20631), .ZN(n20406) );
  OAI211_X1 U23350 ( .C1(n20634), .C2(n20423), .A(n20407), .B(n20406), .ZN(
        P1_U3106) );
  AOI22_X1 U23351 ( .A1(n20636), .A2(n20419), .B1(n20635), .B2(n20418), .ZN(
        n20409) );
  AOI22_X1 U23352 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20420), .B1(
        n20427), .B2(n20637), .ZN(n20408) );
  OAI211_X1 U23353 ( .C1(n20640), .C2(n20423), .A(n20409), .B(n20408), .ZN(
        P1_U3107) );
  AOI22_X1 U23354 ( .A1(n20642), .A2(n20419), .B1(n20641), .B2(n20418), .ZN(
        n20411) );
  AOI22_X1 U23355 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20420), .B1(
        n20427), .B2(n20643), .ZN(n20410) );
  OAI211_X1 U23356 ( .C1(n20646), .C2(n20423), .A(n20411), .B(n20410), .ZN(
        P1_U3108) );
  AOI22_X1 U23357 ( .A1(n20648), .A2(n20419), .B1(n20647), .B2(n20418), .ZN(
        n20413) );
  AOI22_X1 U23358 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20420), .B1(
        n20427), .B2(n20649), .ZN(n20412) );
  OAI211_X1 U23359 ( .C1(n20652), .C2(n20423), .A(n20413), .B(n20412), .ZN(
        P1_U3109) );
  AOI22_X1 U23360 ( .A1(n20654), .A2(n20419), .B1(n20653), .B2(n20418), .ZN(
        n20415) );
  AOI22_X1 U23361 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20420), .B1(
        n20427), .B2(n20655), .ZN(n20414) );
  OAI211_X1 U23362 ( .C1(n20658), .C2(n20423), .A(n20415), .B(n20414), .ZN(
        P1_U3110) );
  AOI22_X1 U23363 ( .A1(n20660), .A2(n20419), .B1(n20659), .B2(n20418), .ZN(
        n20417) );
  AOI22_X1 U23364 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20420), .B1(
        n20427), .B2(n20661), .ZN(n20416) );
  OAI211_X1 U23365 ( .C1(n20664), .C2(n20423), .A(n20417), .B(n20416), .ZN(
        P1_U3111) );
  AOI22_X1 U23366 ( .A1(n20668), .A2(n20419), .B1(n20666), .B2(n20418), .ZN(
        n20422) );
  AOI22_X1 U23367 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20420), .B1(
        n20427), .B2(n20669), .ZN(n20421) );
  OAI211_X1 U23368 ( .C1(n20675), .C2(n20423), .A(n20422), .B(n20421), .ZN(
        P1_U3112) );
  INV_X1 U23369 ( .A(n20424), .ZN(n20563) );
  NOR2_X1 U23370 ( .A1(n20615), .A2(n20473), .ZN(n20480) );
  INV_X1 U23371 ( .A(n20480), .ZN(n20475) );
  NOR2_X1 U23372 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20475), .ZN(
        n20431) );
  INV_X1 U23373 ( .A(n20431), .ZN(n20465) );
  OAI22_X1 U23374 ( .A1(n20472), .A2(n20628), .B1(n20425), .B2(n20465), .ZN(
        n20426) );
  INV_X1 U23375 ( .A(n20426), .ZN(n20440) );
  OAI21_X1 U23376 ( .B1(n20502), .B2(n20427), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20428) );
  NAND2_X1 U23377 ( .A1(n20428), .A2(n20481), .ZN(n20438) );
  AND2_X1 U23378 ( .A1(n20474), .A2(n11447), .ZN(n20435) );
  OR2_X1 U23379 ( .A1(n20430), .A2(n20429), .ZN(n20567) );
  NAND2_X1 U23380 ( .A1(n20567), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20572) );
  OAI21_X1 U23381 ( .B1(n20841), .B2(n20431), .A(n20572), .ZN(n20432) );
  INV_X1 U23382 ( .A(n20432), .ZN(n20434) );
  OAI211_X1 U23383 ( .C1(n20438), .C2(n20435), .A(n20434), .B(n20433), .ZN(
        n20469) );
  INV_X1 U23384 ( .A(n20435), .ZN(n20437) );
  OAI22_X1 U23385 ( .A1(n20438), .A2(n20437), .B1(n20436), .B2(n20567), .ZN(
        n20468) );
  AOI22_X1 U23386 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20469), .B1(
        n20619), .B2(n20468), .ZN(n20439) );
  OAI211_X1 U23387 ( .C1(n20578), .C2(n20499), .A(n20440), .B(n20439), .ZN(
        P1_U3113) );
  OAI22_X1 U23388 ( .A1(n20472), .A2(n20634), .B1(n20441), .B2(n20465), .ZN(
        n20442) );
  INV_X1 U23389 ( .A(n20442), .ZN(n20444) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20469), .B1(
        n20630), .B2(n20468), .ZN(n20443) );
  OAI211_X1 U23391 ( .C1(n20582), .C2(n20499), .A(n20444), .B(n20443), .ZN(
        P1_U3114) );
  OAI22_X1 U23392 ( .A1(n20499), .A2(n20586), .B1(n20445), .B2(n20465), .ZN(
        n20446) );
  INV_X1 U23393 ( .A(n20446), .ZN(n20448) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20469), .B1(
        n20636), .B2(n20468), .ZN(n20447) );
  OAI211_X1 U23395 ( .C1(n20640), .C2(n20472), .A(n20448), .B(n20447), .ZN(
        P1_U3115) );
  OAI22_X1 U23396 ( .A1(n20499), .A2(n20590), .B1(n20449), .B2(n20465), .ZN(
        n20450) );
  INV_X1 U23397 ( .A(n20450), .ZN(n20452) );
  AOI22_X1 U23398 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20469), .B1(
        n20642), .B2(n20468), .ZN(n20451) );
  OAI211_X1 U23399 ( .C1(n20646), .C2(n20472), .A(n20452), .B(n20451), .ZN(
        P1_U3116) );
  OAI22_X1 U23400 ( .A1(n20472), .A2(n20652), .B1(n20453), .B2(n20465), .ZN(
        n20454) );
  INV_X1 U23401 ( .A(n20454), .ZN(n20456) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20469), .B1(
        n20648), .B2(n20468), .ZN(n20455) );
  OAI211_X1 U23403 ( .C1(n20594), .C2(n20499), .A(n20456), .B(n20455), .ZN(
        P1_U3117) );
  OAI22_X1 U23404 ( .A1(n20499), .A2(n20598), .B1(n20457), .B2(n20465), .ZN(
        n20458) );
  INV_X1 U23405 ( .A(n20458), .ZN(n20460) );
  AOI22_X1 U23406 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20469), .B1(
        n20654), .B2(n20468), .ZN(n20459) );
  OAI211_X1 U23407 ( .C1(n20658), .C2(n20472), .A(n20460), .B(n20459), .ZN(
        P1_U3118) );
  OAI22_X1 U23408 ( .A1(n20472), .A2(n20664), .B1(n20461), .B2(n20465), .ZN(
        n20462) );
  INV_X1 U23409 ( .A(n20462), .ZN(n20464) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20469), .B1(
        n20660), .B2(n20468), .ZN(n20463) );
  OAI211_X1 U23411 ( .C1(n20602), .C2(n20499), .A(n20464), .B(n20463), .ZN(
        P1_U3119) );
  OAI22_X1 U23412 ( .A1(n20499), .A2(n20610), .B1(n20466), .B2(n20465), .ZN(
        n20467) );
  INV_X1 U23413 ( .A(n20467), .ZN(n20471) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20469), .B1(
        n20668), .B2(n20468), .ZN(n20470) );
  OAI211_X1 U23415 ( .C1(n20675), .C2(n20472), .A(n20471), .B(n20470), .ZN(
        P1_U3120) );
  NOR2_X1 U23416 ( .A1(n20611), .A2(n20473), .ZN(n20500) );
  AOI21_X1 U23417 ( .B1(n20474), .B2(n20612), .A(n20500), .ZN(n20476) );
  OAI22_X1 U23418 ( .A1(n20476), .A2(n20620), .B1(n20475), .B2(n20679), .ZN(
        n20501) );
  AOI22_X1 U23419 ( .A1(n20619), .A2(n20501), .B1(n20618), .B2(n20500), .ZN(
        n20485) );
  OAI211_X1 U23420 ( .C1(n20478), .C2(n20477), .A(n20481), .B(n20476), .ZN(
        n20479) );
  OAI211_X1 U23421 ( .C1(n20481), .C2(n20480), .A(n20622), .B(n20479), .ZN(
        n20503) );
  INV_X1 U23422 ( .A(n20534), .ZN(n20496) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20503), .B1(
        n20496), .B2(n20625), .ZN(n20484) );
  OAI211_X1 U23424 ( .C1(n20628), .C2(n20499), .A(n20485), .B(n20484), .ZN(
        P1_U3121) );
  AOI22_X1 U23425 ( .A1(n20630), .A2(n20501), .B1(n20629), .B2(n20500), .ZN(
        n20487) );
  AOI22_X1 U23426 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20503), .B1(
        n20496), .B2(n20631), .ZN(n20486) );
  OAI211_X1 U23427 ( .C1(n20634), .C2(n20499), .A(n20487), .B(n20486), .ZN(
        P1_U3122) );
  AOI22_X1 U23428 ( .A1(n20636), .A2(n20501), .B1(n20635), .B2(n20500), .ZN(
        n20489) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20583), .ZN(n20488) );
  OAI211_X1 U23430 ( .C1(n20586), .C2(n20534), .A(n20489), .B(n20488), .ZN(
        P1_U3123) );
  AOI22_X1 U23431 ( .A1(n20642), .A2(n20501), .B1(n20641), .B2(n20500), .ZN(
        n20491) );
  AOI22_X1 U23432 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20503), .B1(
        n20496), .B2(n20643), .ZN(n20490) );
  OAI211_X1 U23433 ( .C1(n20646), .C2(n20499), .A(n20491), .B(n20490), .ZN(
        P1_U3124) );
  AOI22_X1 U23434 ( .A1(n20648), .A2(n20501), .B1(n20647), .B2(n20500), .ZN(
        n20493) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20591), .ZN(n20492) );
  OAI211_X1 U23436 ( .C1(n20594), .C2(n20534), .A(n20493), .B(n20492), .ZN(
        P1_U3125) );
  AOI22_X1 U23437 ( .A1(n20654), .A2(n20501), .B1(n20653), .B2(n20500), .ZN(
        n20495) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20503), .B1(
        n20496), .B2(n20655), .ZN(n20494) );
  OAI211_X1 U23439 ( .C1(n20658), .C2(n20499), .A(n20495), .B(n20494), .ZN(
        P1_U3126) );
  AOI22_X1 U23440 ( .A1(n20660), .A2(n20501), .B1(n20659), .B2(n20500), .ZN(
        n20498) );
  AOI22_X1 U23441 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20503), .B1(
        n20496), .B2(n20661), .ZN(n20497) );
  OAI211_X1 U23442 ( .C1(n20664), .C2(n20499), .A(n20498), .B(n20497), .ZN(
        P1_U3127) );
  AOI22_X1 U23443 ( .A1(n20668), .A2(n20501), .B1(n20666), .B2(n20500), .ZN(
        n20505) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20605), .ZN(n20504) );
  OAI211_X1 U23445 ( .C1(n20610), .C2(n20534), .A(n20505), .B(n20504), .ZN(
        P1_U3128) );
  NAND2_X1 U23446 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20614) );
  AOI22_X1 U23447 ( .A1(n20559), .A2(n20625), .B1(n20618), .B2(n9683), .ZN(
        n20517) );
  INV_X1 U23448 ( .A(n20559), .ZN(n20508) );
  NAND2_X1 U23449 ( .A1(n20534), .A2(n20508), .ZN(n20509) );
  AOI21_X1 U23450 ( .B1(n20509), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20620), 
        .ZN(n20512) );
  OR2_X1 U23451 ( .A1(n13572), .A2(n20510), .ZN(n20565) );
  OR2_X1 U23452 ( .A1(n20565), .A2(n11447), .ZN(n20514) );
  AOI22_X1 U23453 ( .A1(n20512), .A2(n20514), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20513), .ZN(n20511) );
  OAI211_X1 U23454 ( .C1(n9683), .C2(n20841), .A(n20573), .B(n20511), .ZN(
        n20531) );
  INV_X1 U23455 ( .A(n20512), .ZN(n20515) );
  OAI22_X1 U23456 ( .A1(n20515), .A2(n20514), .B1(n20566), .B2(n20513), .ZN(
        n20530) );
  AOI22_X1 U23457 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20531), .B1(
        n20619), .B2(n20530), .ZN(n20516) );
  OAI211_X1 U23458 ( .C1(n20628), .C2(n20534), .A(n20517), .B(n20516), .ZN(
        P1_U3129) );
  AOI22_X1 U23459 ( .A1(n20559), .A2(n20631), .B1(n20629), .B2(n9683), .ZN(
        n20519) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20531), .B1(
        n20630), .B2(n20530), .ZN(n20518) );
  OAI211_X1 U23461 ( .C1(n20634), .C2(n20534), .A(n20519), .B(n20518), .ZN(
        P1_U3130) );
  AOI22_X1 U23462 ( .A1(n20559), .A2(n20637), .B1(n20635), .B2(n9683), .ZN(
        n20521) );
  AOI22_X1 U23463 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20531), .B1(
        n20636), .B2(n20530), .ZN(n20520) );
  OAI211_X1 U23464 ( .C1(n20640), .C2(n20534), .A(n20521), .B(n20520), .ZN(
        P1_U3131) );
  AOI22_X1 U23465 ( .A1(n20559), .A2(n20643), .B1(n20641), .B2(n9683), .ZN(
        n20523) );
  AOI22_X1 U23466 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20531), .B1(
        n20642), .B2(n20530), .ZN(n20522) );
  OAI211_X1 U23467 ( .C1(n20646), .C2(n20534), .A(n20523), .B(n20522), .ZN(
        P1_U3132) );
  AOI22_X1 U23468 ( .A1(n20559), .A2(n20649), .B1(n20647), .B2(n9683), .ZN(
        n20525) );
  AOI22_X1 U23469 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20531), .B1(
        n20648), .B2(n20530), .ZN(n20524) );
  OAI211_X1 U23470 ( .C1(n20652), .C2(n20534), .A(n20525), .B(n20524), .ZN(
        P1_U3133) );
  AOI22_X1 U23471 ( .A1(n20559), .A2(n20655), .B1(n20653), .B2(n9683), .ZN(
        n20527) );
  AOI22_X1 U23472 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20531), .B1(
        n20654), .B2(n20530), .ZN(n20526) );
  OAI211_X1 U23473 ( .C1(n20658), .C2(n20534), .A(n20527), .B(n20526), .ZN(
        P1_U3134) );
  AOI22_X1 U23474 ( .A1(n20559), .A2(n20661), .B1(n20659), .B2(n9683), .ZN(
        n20529) );
  AOI22_X1 U23475 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20531), .B1(
        n20660), .B2(n20530), .ZN(n20528) );
  OAI211_X1 U23476 ( .C1(n20664), .C2(n20534), .A(n20529), .B(n20528), .ZN(
        P1_U3135) );
  AOI22_X1 U23477 ( .A1(n20559), .A2(n20669), .B1(n20666), .B2(n9683), .ZN(
        n20533) );
  AOI22_X1 U23478 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20531), .B1(
        n20668), .B2(n20530), .ZN(n20532) );
  OAI211_X1 U23479 ( .C1(n20675), .C2(n20534), .A(n20533), .B(n20532), .ZN(
        P1_U3136) );
  NOR2_X1 U23480 ( .A1(n20614), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20541) );
  INV_X1 U23481 ( .A(n20541), .ZN(n20537) );
  NOR2_X1 U23482 ( .A1(n20536), .A2(n20537), .ZN(n20557) );
  INV_X1 U23483 ( .A(n20557), .ZN(n20538) );
  OAI222_X1 U23484 ( .A1(n20565), .A2(n20539), .B1(n20538), .B2(n20620), .C1(
        n20679), .C2(n20537), .ZN(n20558) );
  AOI22_X1 U23485 ( .A1(n20619), .A2(n20558), .B1(n20618), .B2(n20557), .ZN(
        n20544) );
  INV_X1 U23486 ( .A(n20540), .ZN(n20542) );
  OAI21_X1 U23487 ( .B1(n20542), .B2(n20541), .A(n20622), .ZN(n20560) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20560), .B1(
        n20559), .B2(n20575), .ZN(n20543) );
  OAI211_X1 U23489 ( .C1(n20578), .C2(n20568), .A(n20544), .B(n20543), .ZN(
        P1_U3137) );
  AOI22_X1 U23490 ( .A1(n20630), .A2(n20558), .B1(n20629), .B2(n20557), .ZN(
        n20546) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20560), .B1(
        n20559), .B2(n20579), .ZN(n20545) );
  OAI211_X1 U23492 ( .C1(n20582), .C2(n20568), .A(n20546), .B(n20545), .ZN(
        P1_U3138) );
  AOI22_X1 U23493 ( .A1(n20636), .A2(n20558), .B1(n20635), .B2(n20557), .ZN(
        n20548) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20560), .B1(
        n20559), .B2(n20583), .ZN(n20547) );
  OAI211_X1 U23495 ( .C1(n20586), .C2(n20568), .A(n20548), .B(n20547), .ZN(
        P1_U3139) );
  AOI22_X1 U23496 ( .A1(n20642), .A2(n20558), .B1(n20641), .B2(n20557), .ZN(
        n20550) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20560), .B1(
        n20559), .B2(n20587), .ZN(n20549) );
  OAI211_X1 U23498 ( .C1(n20590), .C2(n20568), .A(n20550), .B(n20549), .ZN(
        P1_U3140) );
  AOI22_X1 U23499 ( .A1(n20648), .A2(n20558), .B1(n20647), .B2(n20557), .ZN(
        n20552) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20560), .B1(
        n20559), .B2(n20591), .ZN(n20551) );
  OAI211_X1 U23501 ( .C1(n20594), .C2(n20568), .A(n20552), .B(n20551), .ZN(
        P1_U3141) );
  AOI22_X1 U23502 ( .A1(n20654), .A2(n20558), .B1(n20653), .B2(n20557), .ZN(
        n20554) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20560), .B1(
        n20559), .B2(n20595), .ZN(n20553) );
  OAI211_X1 U23504 ( .C1(n20598), .C2(n20568), .A(n20554), .B(n20553), .ZN(
        P1_U3142) );
  AOI22_X1 U23505 ( .A1(n20660), .A2(n20558), .B1(n20659), .B2(n20557), .ZN(
        n20556) );
  AOI22_X1 U23506 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20560), .B1(
        n20559), .B2(n20599), .ZN(n20555) );
  OAI211_X1 U23507 ( .C1(n20602), .C2(n20568), .A(n20556), .B(n20555), .ZN(
        P1_U3143) );
  AOI22_X1 U23508 ( .A1(n20668), .A2(n20558), .B1(n20666), .B2(n20557), .ZN(
        n20562) );
  AOI22_X1 U23509 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20560), .B1(
        n20559), .B2(n20605), .ZN(n20561) );
  OAI211_X1 U23510 ( .C1(n20610), .C2(n20568), .A(n20562), .B(n20561), .ZN(
        P1_U3144) );
  INV_X1 U23511 ( .A(n20565), .ZN(n20613) );
  NAND2_X1 U23512 ( .A1(n20613), .A2(n11447), .ZN(n20570) );
  OAI22_X1 U23513 ( .A1(n20570), .A2(n20620), .B1(n20567), .B2(n20566), .ZN(
        n20604) );
  AOI22_X1 U23514 ( .A1(n20619), .A2(n20604), .B1(n20618), .B2(n20603), .ZN(
        n20577) );
  INV_X1 U23515 ( .A(n20674), .ZN(n20569) );
  OAI21_X1 U23516 ( .B1(n20606), .B2(n20569), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20571) );
  AOI21_X1 U23517 ( .B1(n20571), .B2(n20570), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20574) );
  OAI211_X1 U23518 ( .C1(n20603), .C2(n20574), .A(n20573), .B(n20572), .ZN(
        n20607) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20607), .B1(
        n20606), .B2(n20575), .ZN(n20576) );
  OAI211_X1 U23520 ( .C1(n20578), .C2(n20674), .A(n20577), .B(n20576), .ZN(
        P1_U3145) );
  AOI22_X1 U23521 ( .A1(n20630), .A2(n20604), .B1(n20629), .B2(n20603), .ZN(
        n20581) );
  AOI22_X1 U23522 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20607), .B1(
        n20606), .B2(n20579), .ZN(n20580) );
  OAI211_X1 U23523 ( .C1(n20582), .C2(n20674), .A(n20581), .B(n20580), .ZN(
        P1_U3146) );
  AOI22_X1 U23524 ( .A1(n20636), .A2(n20604), .B1(n20635), .B2(n20603), .ZN(
        n20585) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20607), .B1(
        n20606), .B2(n20583), .ZN(n20584) );
  OAI211_X1 U23526 ( .C1(n20586), .C2(n20674), .A(n20585), .B(n20584), .ZN(
        P1_U3147) );
  AOI22_X1 U23527 ( .A1(n20642), .A2(n20604), .B1(n20641), .B2(n20603), .ZN(
        n20589) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20607), .B1(
        n20606), .B2(n20587), .ZN(n20588) );
  OAI211_X1 U23529 ( .C1(n20590), .C2(n20674), .A(n20589), .B(n20588), .ZN(
        P1_U3148) );
  AOI22_X1 U23530 ( .A1(n20648), .A2(n20604), .B1(n20647), .B2(n20603), .ZN(
        n20593) );
  AOI22_X1 U23531 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20607), .B1(
        n20606), .B2(n20591), .ZN(n20592) );
  OAI211_X1 U23532 ( .C1(n20594), .C2(n20674), .A(n20593), .B(n20592), .ZN(
        P1_U3149) );
  AOI22_X1 U23533 ( .A1(n20654), .A2(n20604), .B1(n20653), .B2(n20603), .ZN(
        n20597) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20607), .B1(
        n20606), .B2(n20595), .ZN(n20596) );
  OAI211_X1 U23535 ( .C1(n20598), .C2(n20674), .A(n20597), .B(n20596), .ZN(
        P1_U3150) );
  AOI22_X1 U23536 ( .A1(n20660), .A2(n20604), .B1(n20659), .B2(n20603), .ZN(
        n20601) );
  AOI22_X1 U23537 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20607), .B1(
        n20606), .B2(n20599), .ZN(n20600) );
  OAI211_X1 U23538 ( .C1(n20602), .C2(n20674), .A(n20601), .B(n20600), .ZN(
        P1_U3151) );
  AOI22_X1 U23539 ( .A1(n20668), .A2(n20604), .B1(n20666), .B2(n20603), .ZN(
        n20609) );
  AOI22_X1 U23540 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20607), .B1(
        n20606), .B2(n20605), .ZN(n20608) );
  OAI211_X1 U23541 ( .C1(n20610), .C2(n20674), .A(n20609), .B(n20608), .ZN(
        P1_U3152) );
  NOR2_X1 U23542 ( .A1(n20611), .A2(n20614), .ZN(n20665) );
  AOI21_X1 U23543 ( .B1(n20613), .B2(n20612), .A(n20665), .ZN(n20617) );
  NOR2_X1 U23544 ( .A1(n20615), .A2(n20614), .ZN(n20623) );
  INV_X1 U23545 ( .A(n20623), .ZN(n20616) );
  OAI22_X1 U23546 ( .A1(n20617), .A2(n20620), .B1(n20616), .B2(n20679), .ZN(
        n20667) );
  AOI22_X1 U23547 ( .A1(n20619), .A2(n20667), .B1(n20618), .B2(n20665), .ZN(
        n20627) );
  NOR3_X1 U23548 ( .A1(n11720), .A2(n20621), .A3(n20620), .ZN(n20624) );
  OAI21_X1 U23549 ( .B1(n20624), .B2(n20623), .A(n20622), .ZN(n20671) );
  AOI22_X1 U23550 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20625), .ZN(n20626) );
  OAI211_X1 U23551 ( .C1(n20628), .C2(n20674), .A(n20627), .B(n20626), .ZN(
        P1_U3153) );
  AOI22_X1 U23552 ( .A1(n20630), .A2(n20667), .B1(n20629), .B2(n20665), .ZN(
        n20633) );
  AOI22_X1 U23553 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20631), .ZN(n20632) );
  OAI211_X1 U23554 ( .C1(n20634), .C2(n20674), .A(n20633), .B(n20632), .ZN(
        P1_U3154) );
  AOI22_X1 U23555 ( .A1(n20636), .A2(n20667), .B1(n20635), .B2(n20665), .ZN(
        n20639) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20637), .ZN(n20638) );
  OAI211_X1 U23557 ( .C1(n20640), .C2(n20674), .A(n20639), .B(n20638), .ZN(
        P1_U3155) );
  AOI22_X1 U23558 ( .A1(n20642), .A2(n20667), .B1(n20641), .B2(n20665), .ZN(
        n20645) );
  AOI22_X1 U23559 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20643), .ZN(n20644) );
  OAI211_X1 U23560 ( .C1(n20646), .C2(n20674), .A(n20645), .B(n20644), .ZN(
        P1_U3156) );
  AOI22_X1 U23561 ( .A1(n20648), .A2(n20667), .B1(n20647), .B2(n20665), .ZN(
        n20651) );
  AOI22_X1 U23562 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20649), .ZN(n20650) );
  OAI211_X1 U23563 ( .C1(n20652), .C2(n20674), .A(n20651), .B(n20650), .ZN(
        P1_U3157) );
  AOI22_X1 U23564 ( .A1(n20654), .A2(n20667), .B1(n20653), .B2(n20665), .ZN(
        n20657) );
  AOI22_X1 U23565 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20655), .ZN(n20656) );
  OAI211_X1 U23566 ( .C1(n20658), .C2(n20674), .A(n20657), .B(n20656), .ZN(
        P1_U3158) );
  AOI22_X1 U23567 ( .A1(n20660), .A2(n20667), .B1(n20659), .B2(n20665), .ZN(
        n20663) );
  AOI22_X1 U23568 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20661), .ZN(n20662) );
  OAI211_X1 U23569 ( .C1(n20664), .C2(n20674), .A(n20663), .B(n20662), .ZN(
        P1_U3159) );
  AOI22_X1 U23570 ( .A1(n20668), .A2(n20667), .B1(n20666), .B2(n20665), .ZN(
        n20673) );
  AOI22_X1 U23571 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20669), .ZN(n20672) );
  OAI211_X1 U23572 ( .C1(n20675), .C2(n20674), .A(n20673), .B(n20672), .ZN(
        P1_U3160) );
  NOR2_X1 U23573 ( .A1(n20677), .A2(n20676), .ZN(n20680) );
  OAI21_X1 U23574 ( .B1(n20680), .B2(n20679), .A(n20678), .ZN(P1_U3163) );
  AND2_X1 U23575 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20681), .ZN(
        P1_U3164) );
  INV_X1 U23576 ( .A(n20748), .ZN(n20682) );
  AND2_X1 U23577 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20682), .ZN(
        P1_U3165) );
  AND2_X1 U23578 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20681), .ZN(
        P1_U3166) );
  AND2_X1 U23579 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20682), .ZN(
        P1_U3167) );
  AND2_X1 U23580 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20681), .ZN(
        P1_U3168) );
  AND2_X1 U23581 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20682), .ZN(
        P1_U3169) );
  AND2_X1 U23582 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20681), .ZN(
        P1_U3170) );
  AND2_X1 U23583 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20682), .ZN(
        P1_U3171) );
  AND2_X1 U23584 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20681), .ZN(
        P1_U3172) );
  AND2_X1 U23585 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20681), .ZN(
        P1_U3173) );
  AND2_X1 U23586 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20681), .ZN(
        P1_U3174) );
  AND2_X1 U23587 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20682), .ZN(
        P1_U3175) );
  AND2_X1 U23588 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20682), .ZN(
        P1_U3176) );
  AND2_X1 U23589 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20682), .ZN(
        P1_U3177) );
  AND2_X1 U23590 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20682), .ZN(
        P1_U3178) );
  AND2_X1 U23591 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20681), .ZN(
        P1_U3179) );
  AND2_X1 U23592 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20681), .ZN(
        P1_U3180) );
  AND2_X1 U23593 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20681), .ZN(
        P1_U3181) );
  AND2_X1 U23594 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20681), .ZN(
        P1_U3182) );
  AND2_X1 U23595 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20681), .ZN(
        P1_U3183) );
  AND2_X1 U23596 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20681), .ZN(
        P1_U3184) );
  AND2_X1 U23597 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20681), .ZN(
        P1_U3185) );
  AND2_X1 U23598 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20682), .ZN(P1_U3186) );
  AND2_X1 U23599 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20682), .ZN(P1_U3187) );
  INV_X1 U23600 ( .A(P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20880) );
  NOR2_X1 U23601 ( .A1(n20748), .A2(n20880), .ZN(P1_U3188) );
  AND2_X1 U23602 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20682), .ZN(P1_U3189) );
  AND2_X1 U23603 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20682), .ZN(P1_U3190) );
  AND2_X1 U23604 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20682), .ZN(P1_U3191) );
  AND2_X1 U23605 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20682), .ZN(P1_U3192) );
  AND2_X1 U23606 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20682), .ZN(P1_U3193) );
  INV_X1 U23607 ( .A(n20683), .ZN(n20688) );
  NOR2_X1 U23608 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20685) );
  OAI22_X1 U23609 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20694), .B1(n20685), 
        .B2(n20684), .ZN(n20686) );
  OAI21_X1 U23610 ( .B1(n20769), .B2(n20686), .A(n20771), .ZN(n20687) );
  OAI211_X1 U23611 ( .C1(n20689), .C2(n20691), .A(n20688), .B(n20687), .ZN(
        P1_U3194) );
  OAI221_X1 U23612 ( .B1(n20689), .B2(n20762), .C1(n20689), .C2(n20694), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n20699) );
  OAI21_X1 U23613 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20769), .A(HOLD), .ZN(
        n20698) );
  NOR2_X1 U23614 ( .A1(n20695), .A2(n20769), .ZN(n20690) );
  AOI21_X1 U23615 ( .B1(n20690), .B2(n20694), .A(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20697) );
  NOR2_X1 U23616 ( .A1(n20692), .A2(n20691), .ZN(n20693) );
  AOI211_X1 U23617 ( .C1(n20695), .C2(n20694), .A(n20757), .B(n20693), .ZN(
        n20696) );
  OAI22_X1 U23618 ( .A1(n20699), .A2(n20698), .B1(n20697), .B2(n20696), .ZN(
        P1_U3196) );
  NAND2_X1 U23619 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20757), .ZN(n20740) );
  AOI22_X1 U23620 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n20771), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20731), .ZN(n20700) );
  OAI21_X1 U23621 ( .B1(n20749), .B2(n20740), .A(n20700), .ZN(P1_U3197) );
  AOI22_X1 U23622 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20771), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n20731), .ZN(n20701) );
  OAI21_X1 U23623 ( .B1(n13504), .B2(n20740), .A(n20701), .ZN(P1_U3198) );
  INV_X1 U23624 ( .A(n20740), .ZN(n20734) );
  AOI222_X1 U23625 ( .A1(n20734), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20771), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20731), .ZN(n20702) );
  INV_X1 U23626 ( .A(n20702), .ZN(P1_U3199) );
  INV_X1 U23627 ( .A(n20731), .ZN(n20737) );
  INV_X1 U23628 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20774) );
  OAI222_X1 U23629 ( .A1(n20737), .A2(n13781), .B1(n20774), .B2(n20757), .C1(
        n20840), .C2(n20740), .ZN(P1_U3200) );
  AOI222_X1 U23630 ( .A1(n20734), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20771), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20731), .ZN(n20703) );
  INV_X1 U23631 ( .A(n20703), .ZN(P1_U3201) );
  AOI222_X1 U23632 ( .A1(n20734), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20771), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20731), .ZN(n20704) );
  INV_X1 U23633 ( .A(n20704), .ZN(P1_U3202) );
  AOI222_X1 U23634 ( .A1(n20734), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20771), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20731), .ZN(n20705) );
  INV_X1 U23635 ( .A(n20705), .ZN(P1_U3203) );
  AOI222_X1 U23636 ( .A1(n20734), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20771), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n20731), .ZN(n20706) );
  INV_X1 U23637 ( .A(n20706), .ZN(P1_U3204) );
  AOI222_X1 U23638 ( .A1(n20734), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20771), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20731), .ZN(n20707) );
  INV_X1 U23639 ( .A(n20707), .ZN(P1_U3205) );
  AOI222_X1 U23640 ( .A1(n20734), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20771), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20731), .ZN(n20708) );
  INV_X1 U23641 ( .A(n20708), .ZN(P1_U3206) );
  AOI222_X1 U23642 ( .A1(n20734), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20771), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20731), .ZN(n20709) );
  INV_X1 U23643 ( .A(n20709), .ZN(P1_U3207) );
  AOI222_X1 U23644 ( .A1(n20731), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20771), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20734), .ZN(n20710) );
  INV_X1 U23645 ( .A(n20710), .ZN(P1_U3208) );
  AOI22_X1 U23646 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20771), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20731), .ZN(n20711) );
  OAI21_X1 U23647 ( .B1(n20712), .B2(n20740), .A(n20711), .ZN(P1_U3209) );
  AOI22_X1 U23648 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20771), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20734), .ZN(n20713) );
  OAI21_X1 U23649 ( .B1(n20714), .B2(n20737), .A(n20713), .ZN(P1_U3210) );
  AOI222_X1 U23650 ( .A1(n20734), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20771), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20731), .ZN(n20715) );
  INV_X1 U23651 ( .A(n20715), .ZN(P1_U3211) );
  AOI222_X1 U23652 ( .A1(n20734), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20771), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20731), .ZN(n20716) );
  INV_X1 U23653 ( .A(n20716), .ZN(P1_U3212) );
  AOI222_X1 U23654 ( .A1(n20731), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20771), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20734), .ZN(n20717) );
  INV_X1 U23655 ( .A(n20717), .ZN(P1_U3213) );
  AOI222_X1 U23656 ( .A1(n20734), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20771), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20731), .ZN(n20718) );
  INV_X1 U23657 ( .A(n20718), .ZN(P1_U3214) );
  AOI22_X1 U23658 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20771), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20731), .ZN(n20719) );
  OAI21_X1 U23659 ( .B1(n20720), .B2(n20740), .A(n20719), .ZN(P1_U3215) );
  AOI22_X1 U23660 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20771), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20734), .ZN(n20721) );
  OAI21_X1 U23661 ( .B1(n20723), .B2(n20737), .A(n20721), .ZN(P1_U3216) );
  AOI22_X1 U23662 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(n20771), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n20731), .ZN(n20722) );
  OAI21_X1 U23663 ( .B1(n20723), .B2(n20740), .A(n20722), .ZN(P1_U3217) );
  AOI22_X1 U23664 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20771), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n20734), .ZN(n20724) );
  OAI21_X1 U23665 ( .B1(n20726), .B2(n20737), .A(n20724), .ZN(P1_U3218) );
  AOI22_X1 U23666 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n20731), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20771), .ZN(n20725) );
  OAI21_X1 U23667 ( .B1(n20726), .B2(n20740), .A(n20725), .ZN(P1_U3219) );
  INV_X1 U23668 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20728) );
  AOI22_X1 U23669 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n20734), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20771), .ZN(n20727) );
  OAI21_X1 U23670 ( .B1(n20728), .B2(n20737), .A(n20727), .ZN(P1_U3220) );
  AOI222_X1 U23671 ( .A1(n20734), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20771), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20731), .ZN(n20729) );
  INV_X1 U23672 ( .A(n20729), .ZN(P1_U3221) );
  AOI222_X1 U23673 ( .A1(n20734), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20771), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20731), .ZN(n20730) );
  INV_X1 U23674 ( .A(n20730), .ZN(P1_U3222) );
  AOI22_X1 U23675 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20731), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20771), .ZN(n20732) );
  OAI21_X1 U23676 ( .B1(n20733), .B2(n20740), .A(n20732), .ZN(P1_U3223) );
  AOI22_X1 U23677 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20734), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20771), .ZN(n20735) );
  OAI21_X1 U23678 ( .B1(n20736), .B2(n20737), .A(n20735), .ZN(P1_U3224) );
  INV_X1 U23679 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20782) );
  OAI222_X1 U23680 ( .A1(n20737), .A2(n14550), .B1(n20782), .B2(n20757), .C1(
        n20736), .C2(n20740), .ZN(P1_U3225) );
  INV_X1 U23681 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20739) );
  INV_X1 U23682 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20738) );
  OAI222_X1 U23683 ( .A1(n20740), .A2(n14550), .B1(n20739), .B2(n20757), .C1(
        n20738), .C2(n20737), .ZN(P1_U3226) );
  OAI22_X1 U23684 ( .A1(n20771), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20757), .ZN(n20741) );
  INV_X1 U23685 ( .A(n20741), .ZN(P1_U3458) );
  OAI22_X1 U23686 ( .A1(n20771), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20757), .ZN(n20742) );
  INV_X1 U23687 ( .A(n20742), .ZN(P1_U3459) );
  OAI22_X1 U23688 ( .A1(n20771), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20757), .ZN(n20743) );
  INV_X1 U23689 ( .A(n20743), .ZN(P1_U3460) );
  OAI22_X1 U23690 ( .A1(n20771), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20757), .ZN(n20744) );
  INV_X1 U23691 ( .A(n20744), .ZN(P1_U3461) );
  OAI21_X1 U23692 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20748), .A(n20746), 
        .ZN(n20745) );
  INV_X1 U23693 ( .A(n20745), .ZN(P1_U3464) );
  OAI21_X1 U23694 ( .B1(n20748), .B2(n20747), .A(n20746), .ZN(P1_U3465) );
  AOI21_X1 U23695 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20750) );
  AOI22_X1 U23696 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20750), .B2(n20749), .ZN(n20753) );
  INV_X1 U23697 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20752) );
  AOI22_X1 U23698 ( .A1(n20756), .A2(n20753), .B1(n20752), .B2(n20751), .ZN(
        P1_U3481) );
  INV_X1 U23699 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20755) );
  OAI21_X1 U23700 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20756), .ZN(n20754) );
  OAI21_X1 U23701 ( .B1(n20756), .B2(n20755), .A(n20754), .ZN(P1_U3482) );
  AOI22_X1 U23702 ( .A1(n20757), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20792), 
        .B2(n20771), .ZN(P1_U3483) );
  INV_X1 U23703 ( .A(n20758), .ZN(n20759) );
  OAI211_X1 U23704 ( .C1(n20762), .C2(n20761), .A(n20760), .B(n20759), .ZN(
        n20770) );
  NOR2_X1 U23705 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20763), .ZN(n20768) );
  OAI211_X1 U23706 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20765), .A(n20764), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20766) );
  NAND2_X1 U23707 ( .A1(n20770), .A2(n20766), .ZN(n20767) );
  OAI22_X1 U23708 ( .A1(n20770), .A2(n20769), .B1(n20768), .B2(n20767), .ZN(
        P1_U3485) );
  MUX2_X1 U23709 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n20771), .Z(P1_U3486) );
  AOI22_X1 U23710 ( .A1(n20774), .A2(keyinput62), .B1(keyinput12), .B2(n20773), 
        .ZN(n20772) );
  OAI221_X1 U23711 ( .B1(n20774), .B2(keyinput62), .C1(n20773), .C2(keyinput12), .A(n20772), .ZN(n20787) );
  AOI22_X1 U23712 ( .A1(n20777), .A2(keyinput61), .B1(keyinput21), .B2(n20776), 
        .ZN(n20775) );
  OAI221_X1 U23713 ( .B1(n20777), .B2(keyinput61), .C1(n20776), .C2(keyinput21), .A(n20775), .ZN(n20786) );
  AOI22_X1 U23714 ( .A1(n20780), .A2(keyinput55), .B1(n20779), .B2(keyinput35), 
        .ZN(n20778) );
  OAI221_X1 U23715 ( .B1(n20780), .B2(keyinput55), .C1(n20779), .C2(keyinput35), .A(n20778), .ZN(n20785) );
  AOI22_X1 U23716 ( .A1(n20783), .A2(keyinput9), .B1(keyinput37), .B2(n20782), 
        .ZN(n20781) );
  OAI221_X1 U23717 ( .B1(n20783), .B2(keyinput9), .C1(n20782), .C2(keyinput37), 
        .A(n20781), .ZN(n20784) );
  NOR4_X1 U23718 ( .A1(n20787), .A2(n20786), .A3(n20785), .A4(n20784), .ZN(
        n20835) );
  INV_X1 U23719 ( .A(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n20789) );
  AOI22_X1 U23720 ( .A1(n20790), .A2(keyinput60), .B1(n20789), .B2(keyinput3), 
        .ZN(n20788) );
  OAI221_X1 U23721 ( .B1(n20790), .B2(keyinput60), .C1(n20789), .C2(keyinput3), 
        .A(n20788), .ZN(n20802) );
  AOI22_X1 U23722 ( .A1(n20793), .A2(keyinput18), .B1(keyinput0), .B2(n20792), 
        .ZN(n20791) );
  OAI221_X1 U23723 ( .B1(n20793), .B2(keyinput18), .C1(n20792), .C2(keyinput0), 
        .A(n20791), .ZN(n20801) );
  AOI22_X1 U23724 ( .A1(n20796), .A2(keyinput4), .B1(n20795), .B2(keyinput8), 
        .ZN(n20794) );
  OAI221_X1 U23725 ( .B1(n20796), .B2(keyinput4), .C1(n20795), .C2(keyinput8), 
        .A(n20794), .ZN(n20800) );
  INV_X1 U23726 ( .A(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n20798) );
  AOI22_X1 U23727 ( .A1(n12384), .A2(keyinput42), .B1(keyinput11), .B2(n20798), 
        .ZN(n20797) );
  OAI221_X1 U23728 ( .B1(n12384), .B2(keyinput42), .C1(n20798), .C2(keyinput11), .A(n20797), .ZN(n20799) );
  NOR4_X1 U23729 ( .A1(n20802), .A2(n20801), .A3(n20800), .A4(n20799), .ZN(
        n20834) );
  INV_X1 U23730 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n20804) );
  AOI22_X1 U23731 ( .A1(n20804), .A2(keyinput38), .B1(n14983), .B2(keyinput22), 
        .ZN(n20803) );
  OAI221_X1 U23732 ( .B1(n20804), .B2(keyinput38), .C1(n14983), .C2(keyinput22), .A(n20803), .ZN(n20817) );
  AOI22_X1 U23733 ( .A1(n20807), .A2(keyinput57), .B1(keyinput32), .B2(n20806), 
        .ZN(n20805) );
  OAI221_X1 U23734 ( .B1(n20807), .B2(keyinput57), .C1(n20806), .C2(keyinput32), .A(n20805), .ZN(n20816) );
  AOI22_X1 U23735 ( .A1(n20810), .A2(keyinput39), .B1(keyinput58), .B2(n20809), 
        .ZN(n20808) );
  OAI221_X1 U23736 ( .B1(n20810), .B2(keyinput39), .C1(n20809), .C2(keyinput58), .A(n20808), .ZN(n20815) );
  INV_X1 U23737 ( .A(P1_LWORD_REG_4__SCAN_IN), .ZN(n20813) );
  AOI22_X1 U23738 ( .A1(n20813), .A2(keyinput19), .B1(keyinput36), .B2(n20812), 
        .ZN(n20811) );
  OAI221_X1 U23739 ( .B1(n20813), .B2(keyinput19), .C1(n20812), .C2(keyinput36), .A(n20811), .ZN(n20814) );
  NOR4_X1 U23740 ( .A1(n20817), .A2(n20816), .A3(n20815), .A4(n20814), .ZN(
        n20833) );
  AOI22_X1 U23741 ( .A1(n14665), .A2(keyinput52), .B1(n14877), .B2(keyinput45), 
        .ZN(n20818) );
  OAI221_X1 U23742 ( .B1(n14665), .B2(keyinput52), .C1(n14877), .C2(keyinput45), .A(n20818), .ZN(n20831) );
  INV_X1 U23743 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n20821) );
  AOI22_X1 U23744 ( .A1(n20821), .A2(keyinput13), .B1(keyinput24), .B2(n20820), 
        .ZN(n20819) );
  OAI221_X1 U23745 ( .B1(n20821), .B2(keyinput13), .C1(n20820), .C2(keyinput24), .A(n20819), .ZN(n20830) );
  AOI22_X1 U23746 ( .A1(n20824), .A2(keyinput27), .B1(n20823), .B2(keyinput40), 
        .ZN(n20822) );
  OAI221_X1 U23747 ( .B1(n20824), .B2(keyinput27), .C1(n20823), .C2(keyinput40), .A(n20822), .ZN(n20829) );
  XOR2_X1 U23748 ( .A(n20825), .B(keyinput50), .Z(n20827) );
  XNOR2_X1 U23749 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B(keyinput26), .ZN(
        n20826) );
  NAND2_X1 U23750 ( .A1(n20827), .A2(n20826), .ZN(n20828) );
  NOR4_X1 U23751 ( .A1(n20831), .A2(n20830), .A3(n20829), .A4(n20828), .ZN(
        n20832) );
  NAND4_X1 U23752 ( .A1(n20835), .A2(n20834), .A3(n20833), .A4(n20832), .ZN(
        n20900) );
  AOI22_X1 U23753 ( .A1(n15432), .A2(keyinput16), .B1(keyinput44), .B2(n14456), 
        .ZN(n20836) );
  OAI221_X1 U23754 ( .B1(n15432), .B2(keyinput16), .C1(n14456), .C2(keyinput44), .A(n20836), .ZN(n20848) );
  AOI22_X1 U23755 ( .A1(n10900), .A2(keyinput41), .B1(keyinput33), .B2(n20838), 
        .ZN(n20837) );
  OAI221_X1 U23756 ( .B1(n10900), .B2(keyinput41), .C1(n20838), .C2(keyinput33), .A(n20837), .ZN(n20847) );
  AOI22_X1 U23757 ( .A1(n20841), .A2(keyinput15), .B1(keyinput17), .B2(n20840), 
        .ZN(n20839) );
  OAI221_X1 U23758 ( .B1(n20841), .B2(keyinput15), .C1(n20840), .C2(keyinput17), .A(n20839), .ZN(n20846) );
  AOI22_X1 U23759 ( .A1(n20844), .A2(keyinput30), .B1(keyinput28), .B2(n20843), 
        .ZN(n20842) );
  OAI221_X1 U23760 ( .B1(n20844), .B2(keyinput30), .C1(n20843), .C2(keyinput28), .A(n20842), .ZN(n20845) );
  NOR4_X1 U23761 ( .A1(n20848), .A2(n20847), .A3(n20846), .A4(n20845), .ZN(
        n20898) );
  AOI22_X1 U23762 ( .A1(n20850), .A2(keyinput14), .B1(n12365), .B2(keyinput25), 
        .ZN(n20849) );
  OAI221_X1 U23763 ( .B1(n20850), .B2(keyinput14), .C1(n12365), .C2(keyinput25), .A(n20849), .ZN(n20854) );
  XOR2_X1 U23764 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B(keyinput31), .Z(
        n20853) );
  XNOR2_X1 U23765 ( .A(n20851), .B(keyinput54), .ZN(n20852) );
  OR3_X1 U23766 ( .A1(n20854), .A2(n20853), .A3(n20852), .ZN(n20862) );
  AOI22_X1 U23767 ( .A1(n20856), .A2(keyinput47), .B1(n20905), .B2(keyinput5), 
        .ZN(n20855) );
  OAI221_X1 U23768 ( .B1(n20856), .B2(keyinput47), .C1(n20905), .C2(keyinput5), 
        .A(n20855), .ZN(n20861) );
  AOI22_X1 U23769 ( .A1(n20859), .A2(keyinput43), .B1(keyinput53), .B2(n20858), 
        .ZN(n20857) );
  OAI221_X1 U23770 ( .B1(n20859), .B2(keyinput43), .C1(n20858), .C2(keyinput53), .A(n20857), .ZN(n20860) );
  NOR3_X1 U23771 ( .A1(n20862), .A2(n20861), .A3(n20860), .ZN(n20897) );
  AOI22_X1 U23772 ( .A1(n20865), .A2(keyinput63), .B1(keyinput51), .B2(n20864), 
        .ZN(n20863) );
  OAI221_X1 U23773 ( .B1(n20865), .B2(keyinput63), .C1(n20864), .C2(keyinput51), .A(n20863), .ZN(n20878) );
  AOI22_X1 U23774 ( .A1(n20868), .A2(keyinput20), .B1(keyinput1), .B2(n20867), 
        .ZN(n20866) );
  OAI221_X1 U23775 ( .B1(n20868), .B2(keyinput20), .C1(n20867), .C2(keyinput1), 
        .A(n20866), .ZN(n20877) );
  AOI22_X1 U23776 ( .A1(n20871), .A2(keyinput49), .B1(n20870), .B2(keyinput46), 
        .ZN(n20869) );
  OAI221_X1 U23777 ( .B1(n20871), .B2(keyinput49), .C1(n20870), .C2(keyinput46), .A(n20869), .ZN(n20876) );
  AOI22_X1 U23778 ( .A1(n20874), .A2(keyinput34), .B1(n20873), .B2(keyinput10), 
        .ZN(n20872) );
  OAI221_X1 U23779 ( .B1(n20874), .B2(keyinput34), .C1(n20873), .C2(keyinput10), .A(n20872), .ZN(n20875) );
  NOR4_X1 U23780 ( .A1(n20878), .A2(n20877), .A3(n20876), .A4(n20875), .ZN(
        n20896) );
  AOI22_X1 U23781 ( .A1(n20881), .A2(keyinput56), .B1(keyinput29), .B2(n20880), 
        .ZN(n20879) );
  OAI221_X1 U23782 ( .B1(n20881), .B2(keyinput56), .C1(n20880), .C2(keyinput29), .A(n20879), .ZN(n20894) );
  AOI22_X1 U23783 ( .A1(n20916), .A2(keyinput48), .B1(n20883), .B2(keyinput59), 
        .ZN(n20882) );
  OAI221_X1 U23784 ( .B1(n20916), .B2(keyinput48), .C1(n20883), .C2(keyinput59), .A(n20882), .ZN(n20893) );
  AOI22_X1 U23785 ( .A1(n20886), .A2(keyinput6), .B1(keyinput2), .B2(n20885), 
        .ZN(n20884) );
  OAI221_X1 U23786 ( .B1(n20886), .B2(keyinput6), .C1(n20885), .C2(keyinput2), 
        .A(n20884), .ZN(n20891) );
  XNOR2_X1 U23787 ( .A(n20887), .B(keyinput7), .ZN(n20890) );
  XNOR2_X1 U23788 ( .A(n20888), .B(keyinput23), .ZN(n20889) );
  OR3_X1 U23789 ( .A1(n20891), .A2(n20890), .A3(n20889), .ZN(n20892) );
  NOR3_X1 U23790 ( .A1(n20894), .A2(n20893), .A3(n20892), .ZN(n20895) );
  NAND4_X1 U23791 ( .A1(n20898), .A2(n20897), .A3(n20896), .A4(n20895), .ZN(
        n20899) );
  NOR2_X1 U23792 ( .A1(n20900), .A2(n20899), .ZN(n20929) );
  NAND4_X1 U23793 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_4__4__SCAN_IN), .A3(P3_PHYADDRPOINTER_REG_0__SCAN_IN), 
        .A4(P3_EAX_REG_21__SCAN_IN), .ZN(n20904) );
  NAND4_X1 U23794 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A4(
        P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n20903) );
  NAND4_X1 U23795 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(
        P2_EBX_REG_24__SCAN_IN), .A3(P2_EAX_REG_28__SCAN_IN), .A4(
        P2_EAX_REG_24__SCAN_IN), .ZN(n20902) );
  NAND4_X1 U23796 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(
        P2_EBX_REG_28__SCAN_IN), .A3(P1_EBX_REG_16__SCAN_IN), .A4(
        P1_REIP_REG_10__SCAN_IN), .ZN(n20901) );
  NOR4_X1 U23797 ( .A1(n20904), .A2(n20903), .A3(n20902), .A4(n20901), .ZN(
        n20923) );
  NAND3_X1 U23798 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_9__7__SCAN_IN), .A3(P1_INSTQUEUE_REG_13__7__SCAN_IN), 
        .ZN(n20915) );
  NOR4_X1 U23799 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_9__2__SCAN_IN), .A3(P1_INSTQUEUE_REG_2__2__SCAN_IN), 
        .A4(n20905), .ZN(n20908) );
  NOR4_X1 U23800 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_STATEBS16_REG_SCAN_IN), .A3(BUF1_REG_5__SCAN_IN), .A4(
        P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20907) );
  NOR4_X1 U23801 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(BUF2_REG_31__SCAN_IN), 
        .A3(P2_LWORD_REG_2__SCAN_IN), .A4(P2_DATAO_REG_23__SCAN_IN), .ZN(
        n20906) );
  NAND3_X1 U23802 ( .A1(n20908), .A2(n20907), .A3(n20906), .ZN(n20914) );
  NOR4_X1 U23803 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_UWORD_REG_8__SCAN_IN), .A4(
        P3_DATAO_REG_26__SCAN_IN), .ZN(n20912) );
  NOR4_X1 U23804 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(
        P3_REIP_REG_1__SCAN_IN), .A3(P3_EAX_REG_29__SCAN_IN), .A4(
        P2_DATAO_REG_6__SCAN_IN), .ZN(n20911) );
  NOR4_X1 U23805 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(BUF2_REG_22__SCAN_IN), .A4(
        BUF2_REG_20__SCAN_IN), .ZN(n20910) );
  NOR4_X1 U23806 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A4(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n20909) );
  NAND4_X1 U23807 ( .A1(n20912), .A2(n20911), .A3(n20910), .A4(n20909), .ZN(
        n20913) );
  NOR4_X1 U23808 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n20915), .A3(n20914), 
        .A4(n20913), .ZN(n20922) );
  NAND4_X1 U23809 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_DATAO_REG_3__SCAN_IN), .A3(P1_W_R_N_REG_SCAN_IN), .A4(n20916), .ZN(
        n20920) );
  NAND4_X1 U23810 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_4__SCAN_IN), .A3(P1_ADDRESS_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20919) );
  NAND4_X1 U23811 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P1_STATE2_REG_3__SCAN_IN), .A4(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n20918) );
  NAND4_X1 U23812 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(P3_EAX_REG_23__SCAN_IN), .A4(
        P2_CODEFETCH_REG_SCAN_IN), .ZN(n20917) );
  NOR4_X1 U23813 ( .A1(n20920), .A2(n20919), .A3(n20918), .A4(n20917), .ZN(
        n20921) );
  NAND3_X1 U23814 ( .A1(n20923), .A2(n20922), .A3(n20921), .ZN(n20927) );
  AOI222_X1 U23815 ( .A1(P1_EAX_REG_8__SCAN_IN), .A2(n20925), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20021), .C1(n20924), .C2(
        P1_DATAO_REG_8__SCAN_IN), .ZN(n20926) );
  XNOR2_X1 U23816 ( .A(n20927), .B(n20926), .ZN(n20928) );
  XNOR2_X1 U23817 ( .A(n20929), .B(n20928), .ZN(P1_U2928) );
  CLKBUF_X2 U11325 ( .A(n10191), .Z(n9583) );
  AND2_X2 U11089 ( .A1(n14441), .A2(n11922), .ZN(n14352) );
  CLKBUF_X3 U11080 ( .A(n12685), .Z(n9565) );
  INV_X2 U11102 ( .A(n12685), .ZN(n17156) );
  INV_X2 U11016 ( .A(n20931), .ZN(n20932) );
  CLKBUF_X1 U11034 ( .A(n11384), .Z(n11333) );
  AND2_X1 U11039 ( .A1(n10886), .A2(n10181), .ZN(n10219) );
  CLKBUF_X1 U11054 ( .A(n10318), .Z(n9567) );
  NAND2_X1 U11056 ( .A1(n10274), .A2(n19178), .ZN(n10278) );
  AND4_X1 U11093 ( .A1(n11201), .A2(n11200), .A3(n11199), .A4(n11198), .ZN(
        n11208) );
  CLKBUF_X2 U11094 ( .A(n10222), .Z(n9569) );
  CLKBUF_X1 U11120 ( .A(n11157), .Z(n11159) );
  AND2_X1 U11124 ( .A1(n10130), .A2(n10129), .ZN(n10190) );
  CLKBUF_X1 U11303 ( .A(n11324), .Z(n20107) );
  CLKBUF_X1 U11356 ( .A(n11696), .Z(n9587) );
  CLKBUF_X1 U11506 ( .A(n18747), .Z(n18739) );
  CLKBUF_X1 U12291 ( .A(n16488), .Z(n16490) );
  OR2_X1 U12294 ( .A1(n9573), .A2(n19205), .ZN(n20930) );
  INV_X1 U12316 ( .A(n11428), .ZN(n20931) );
  CLKBUF_X1 U12671 ( .A(n11462), .Z(n11428) );
endmodule

