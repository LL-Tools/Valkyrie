
module b15_C_2inp_gates_syn ( 
    DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
    DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
    DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
    DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
    DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
    DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
    READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
    M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
    STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
    W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
    BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
    BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
    REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
    REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
    REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
    REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
    REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
    BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
    ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
    ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
    ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
    ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
    ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
    ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
    ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
    ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
    ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
    ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
    ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN,
    ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
    ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN,
    ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN,
    STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
    DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
    DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
    DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
    DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
    DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
    DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
    DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
    DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
    DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
    DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
    DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
    DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
    DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
    DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
    DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
    DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
    STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
    INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
    INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
    INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
    INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
    INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
    INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
    INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
    INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
    INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
    INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
    INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
    INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
    INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
    INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
    INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
    INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
    INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
    INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
    INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
    INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
    INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
    INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
    INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
    INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
    INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
    INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
    INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
    INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
    INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
    INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
    INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
    INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
    INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
    INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
    INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
    INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
    INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
    INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
    INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
    INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
    INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
    INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
    INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
    INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
    INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
    INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
    INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
    INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
    INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
    INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
    INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
    INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
    INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
    INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
    INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
    INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
    INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
    INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
    INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
    INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
    INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
    INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
    INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
    INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
    INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
    INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
    INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
    INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
    INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
    INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
    INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
    INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
    INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
    INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
    INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
    INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
    INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
    INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
    INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
    INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
    INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
    INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
    INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
    INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
    INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
    PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
    PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
    PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
    PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
    PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
    PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
    PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
    PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
    PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
    PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
    PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
    PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
    PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
    PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
    PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
    PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
    LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
    LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
    LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
    LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
    LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
    LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
    UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
    UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
    UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
    UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
    UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
    DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
    DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
    DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
    DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
    DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
    DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
    DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
    DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
    DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
    DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
    EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
    EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
    EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
    EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
    EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
    EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
    EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
    EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
    EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
    EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
    EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
    EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
    EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
    EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
    EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
    EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
    EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
    EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
    EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
    EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
    EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
    EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
    REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
    REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
    REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
    REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
    REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN,
    U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
    U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
    U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
    U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
    U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
    U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
    U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
    U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
    U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
    U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
    U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
    U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
    U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
    U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
    U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
    U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
    U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
    U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
    U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
    U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
    U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
    U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
    U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
    U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
    U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
    U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
    U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
    U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
    U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
    U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
    U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
    U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
    U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
    U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
    U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
    U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
    U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
    U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
    U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
    U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
    U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
    U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
    U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
    U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
    U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788  );
  input  DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_,
    DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_,
    DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_,
    DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_,
    DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_,
    DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N,
    HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN,
    CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN,
    REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN,
    FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
    BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
    BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
    REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
    REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
    REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
    REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
    REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
    BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
    ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
    ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
    ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
    ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
    ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
    ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
    ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
    ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
    ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
    ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
    ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN,
    ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
    ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN,
    ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN,
    STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
    DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
    DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
    DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
    DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
    DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
    DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
    DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
    DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
    DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
    DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
    DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
    DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
    DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
    DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
    DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
    DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
    STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
    INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
    INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
    INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
    INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
    INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
    INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
    INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
    INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
    INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
    INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
    INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
    INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
    INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
    INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
    INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
    INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
    INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
    INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
    INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
    INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
    INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
    INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
    INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
    INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
    INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
    INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
    INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
    INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
    INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
    INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
    INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
    INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
    INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
    INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
    INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
    INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
    INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
    INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
    INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
    INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
    INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
    INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
    INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
    INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
    INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
    INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
    INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
    INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
    INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
    INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
    INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
    INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
    INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
    INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
    INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
    INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
    INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
    INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
    INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
    INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
    INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
    INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
    INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
    INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
    INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
    INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
    INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
    INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
    INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
    INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
    INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
    INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
    INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
    INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
    INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
    INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
    INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
    INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
    INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
    INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
    INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
    INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
    INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
    INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
    INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
    PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
    PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
    PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
    PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
    PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
    PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
    PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
    PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
    PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
    PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
    PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
    PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
    PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
    PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
    PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
    PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
    LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
    LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
    LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
    LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
    LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
    LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
    UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
    UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
    UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
    UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
    UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
    DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
    DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
    DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
    DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
    DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
    DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
    DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
    DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
    DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
    DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
    EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
    EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
    EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
    EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
    EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
    EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
    EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
    EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
    EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
    EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
    EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
    EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
    EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
    EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
    EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
    EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
    EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
    EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
    EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
    EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
    EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
    EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
    REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
    REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
    REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
    REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
    REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
    U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
    U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
    U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
    U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
    U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
    U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
    U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
    U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
    U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
    U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
    U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
    U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
    U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
    U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
    U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
    U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
    U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
    U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
    U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
    U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
    U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
    U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
    U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
    U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
    U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
    U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
    U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
    U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
    U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
    U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
    U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
    U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
    U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
    U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
    U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
    U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
    U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
    U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
    U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
    U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
    U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
    U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
    U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
    U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire n10200, n9085, n8946, n7515, n7363, n7829, n6998, n9029, n10830,
    n9041, n8985, n11821, n7848, n13693, n9129, n10896, n11536, n11772,
    n10735, n11577, n13177, n9926, n6993, n7541, n9201, n7006, n11826,
    n7988, n7004, n11865, n7774, n11462, n11812, n11519, n10089, n10390,
    n11796, n7956, n6994, n10809, n11401, n9115, n9113, n9126, n9286,
    n8310, n9408, n7253, n7257, n7254, n11813, n9955, n9948, n10146, n9987,
    n8843, n9588, n8676, n8478, n13375, n8309, n7098, n7131, n7201, n10240,
    n10270, n7204, n7162, n10056, n10641, n7208, n7074, n7211, n9794,
    n10174, n11420, n10004, n9002, n9162, n13290, n8227, n10871, n9001,
    n11419, n13367, n10400, n10206, n10848, n11732, n13192, n10837, n11537,
    n11884, n11131, n12242, n11880, n6995, n9199, n11013, n11581, n7783,
    n13764, n7600, n13325, n10841, n10855, n8939, n10862, n7068, n7123,
    n7560, n10864, n7550, n7180, n7673, n9088, n9320, n9298, n9435, n7207,
    n7428, n10481, n8940, n7492, n9304, n9017, n9230, n9847, n11948,
    n13328, n7773, n11908, n9210, n7176, n7531, n7390, n7389, n7324, n7325,
    n7358, n7264, n7265, n8154, n7652, n6996, n8642, n7639, n7326, n7248,
    n6997, n11820, n7245, n6999, n7151, n7000, n7001, n7002, n7003, n11477,
    n7198, n7518, n7065, n8993, n7005, n11809, n7138, n7007, n7546, n7504,
    n9214, n7009, n7010, n7469, n7374, n9218, n7011, n10908, n10869,
    n10770, n7167, n7086, n7087, n7595, n7487, n7154, n7166, n7070, n7113,
    n7185, n7533, n7217, n9786, n9788, n7122, n7147, n7106, n7105, n7164,
    n11806, n9130, n9131, n10360, n10790, n7117, n7195, n7171, n7544,
    n7063, n7062, n7060, n9123, n9122, n7216, n8308, n7967, n7149, n7160,
    n7130, n7135, n7132, n7165, n7134, n7076, n9081, n7727, n7855, n7222,
    n7218, n7188, n7189, n8188, n7209, n8060, n7220, n7223, n8600, n8944,
    n7190, n7191, n7193, n7140, n7104, n7103, n7108, n7109, n7110, n9136,
    n9389, n13342, n7675, n8938, n12929, n7357, n9146, n7877, n9626, n9647,
    n7181, n7182, n10379, n10836, n7178, n10451, n11548, n7096, n7097,
    n7094, n7095, n7093, n9957, n7078, n7139, n10116, n11016, n11092,
    n9456, n9452, n9462, n11739, n9377, n7119, n11803, n13661, n9431,
    n9006, n8973, n8958, n7720, n7672, n7603, n7236, n7258, n7289, n9060,
    n7733, n7129, n8888, n7153, n7143, n7194, n7146, n9161, n7169, n7168,
    n8989, n7059, n7061, n7424, n7373, n7341, n7352, n9155, n9125, n10614,
    n10782, n7875, n7116, n7183, n7184, n10685, n9395, n8839, n8756, n8711,
    n8672, n9703, n8557, n7214, n10079, n10104, n10121, n8306, n8268,
    n7210, n8266, n8179, n8180, n8103, n8061, n10705, n8062, n10718, n8020,
    n8022, n7975, n8955, n9303, n9015, n9611, n7111, n7186, n7187, n7085,
    n7107, n7081, n7159, n11431, n8954, n10443, n11819, n7767, n10456,
    n7730, n7859, n12765, n7319, n7488, n7532, n13315, n11873, n13100,
    n13102, n9446, n7219, n8391, n8351, n8343, n9527, n7982, n10822, n7950,
    n10795, n8887, n8842, n9482, n8716, n9723, n7212, n10647, n11253,
    n9147, n9145, n13741, n11259, n9550, n9566, n11488, n11570, n10921,
    n10167, n9391, n9568, n7192, n7172, n7102, n10239, n7200, n10074,
    n7082, n7084, n7083, n10091, n10115, n10144, n13703, n11867, n13355,
    n13701, n12598, n13203, n12845, n12246, n12841, n13354, n11938, n11967,
    n13652, n9135, n13402, n13655, n11983, n9627, n9988, n10325, n10377,
    n10788, n11017, n11020, n9857, n9864, n11097, n11121, n11123, n11252,
    n11405, n7126, n11530, n10158, n9468, n7092, n7079, n7077, n10102,
    n13662, n13121, n13130, n13139, n13148, n13166, n13176, n13390, n7118,
    n7012, n8906, n10704, n13308, n7013, n7014, n10134, n9764, n8453,
    n7015, n9683, n7016, n9493, n7017, n7018, n10912, n7404, n10821, n8562,
    n7019, n7020, n7021, n7022, n7023, n9480, n7024, n7025, n11454, n7026,
    n10029, n7027, n7028, n10744, n9766, n7029, n10078, n7030, n7031,
    n7032, n7033, n7034, n7035, n7206, n7114, n7115, n7036, n7037, n7141,
    n7142, n7155, n7038, n7039, n7202, n7040, n7041, n7042, n7043, n7044,
    n7045, n7046, n7221, n7047, n7048, n7049, n7050, n7051, n7052, n7173,
    n7174, n8587, n9438, n8880, n8854, n10674, n10644, n7053, n7957, n7054,
    n7055, n13683, n9307, n7144, n11928, n7837, n8384, n13400, n8221,
    n7056, n7057, n7161, n7066, n13597, n13757, n7075, n7965, n7058, n7080,
    n11496, n7064, n11719, n7067, n7936, n7552, n10879, n7069, n10120,
    n9543, n7529, n7071, n9024, n9464, n7158, n9032, n9035, n7072, n7073,
    n9004, n11484, n9005, n7145, n10058, n7150, n10057, n7375, n7088,
    n7136, n11499, n7089, n7090, n10173, n7091, n9466, n9947, n7099,
    n13343, n7148, n9479, n11663, n9120, n10203, n9119, n9128, n7170,
    n7175, n10745, n11421, n9943, n9173, n9012, n9013, n7100, n7101, n7137,
    n9239, n9232, n9235, n9242, n9245, n9251, n9330, n9284, n9292, n9295,
    n9211, n9372, n13760, n9360, n9369, n9363, n9366, n9378, n11775, n9685,
    n7112, n9725, n7196, n7120, n7121, n7601, n10684, n7124, n7125, n7127,
    n7128, n7771, n7769, n7561, n11483, n7133, n9026, n11461, n8994,
    n10213, n7966, n9168, n7156, n7152, n10068, n9034, n7157, n7205, n7163,
    n11418, n9985, n7246, n13310, n7177, n9220, n7179, n10410, n9570,
    n9503, n7197, n10803, n7716, n7861, n7511, n9191, n7501, n9315, n7199,
    n9997, n7203, n7486, n7213, n10147, n10148, n10092, n7215, n10103,
    n9743, n9605, n9481, n9540, n9587, n10927, n9511, n9093, n10018, n7847,
    n7845, n9848, n9747, n9705, n7495, n10457, n8305, n8019, n7224, n7225,
    n11881, n7226, n7227, n7228, n9728, n7229, n7432, n7911, n8899, n11828,
    n9105, n7530, n7232, n9007, n8981, n7635, n9107, n8801, n11829, n8142,
    n7558, n7844, n8877, n8666, n9182, n9451, n8350, n8996, n9225, n13345,
    n7457, n7387, n7537, n8675, n8477, n9688, n7987, n9109, n9778, n10576,
    n9514, n9291, n9471, n8760, n8515, n8229, n10732, n12757, n12759,
    n13110, n13321, n8437, n9501, n10907, n10793, n8222, n11576, n13634,
    n11898, n11980, n12249, n12329, n13665, n12673, n12933, n13669, n9494,
    n10484, n9502, n8392, n10914, n10893, n11046, n11186, n11523, n11529,
    n11559, n11792, n11773, n11808, n12052, n12150, n12235, n12324, n12399,
    n12483, n12550, n12575, n12659, n12748, n12830, n12923, n13007, n13082,
    n13093, n13157, n13227, n13263, n13299, n13742, n9143, n13433, n13404,
    n11010, n11001, n11256, n11503, n11578, n11784, n11901, n12154, n12662,
    n10477, n11263, n11567, n11245, n13710, n13414, n13415, n8586, n7231,
    n13344, n8029, n7230, n7235, n7233, n7612, n7234, n7244, n7472, n7238,
    n7237, n7242, n7240, n8279, n7239, n7241, n7243, n7247, n7252, n7250,
    n7249, n7251, n7263, n7256, n7255, n7261, n7336, n7259, n7260, n7262,
    n7267, n7266, n7271, n7269, n7268, n7270, n7279, n7273, n7272, n7277,
    n7275, n7274, n7276, n7278, n7295, n7281, n7280, n7285, n7283, n7282,
    n7284, n7293, n7287, n7286, n7291, n7288, n7290, n7292, n7294, n7516,
    n7297, n7296, n7301, n7299, n7298, n7300, n7309, n7303, n7302, n7307,
    n7305, n7304, n7306, n7308, n7311, n7310, n7315, n7313, n7312, n7314,
    n7323, n7317, n7316, n7321, n7318, n7320, n7322, n7391, n7328, n7327,
    n7333, n7331, n7330, n7332, n7342, n7335, n7334, n7340, n7338, n7337,
    n7339, n7344, n7343, n7348, n7346, n7345, n7347, n7356, n7350, n7349,
    n7354, n7351, n7353, n7355, n7360, n7359, n7365, n7361, n7362, n7364,
    n7367, n7366, n7371, n7369, n7368, n7370, n7372, n7376, n7380, n7378,
    n7377, n7379, n7388, n7382, n7381, n7386, n7384, n7383, n7385, n7496,
    n7395, n7392, n7393, n7394, n7429, n7397, n7396, n7401, n7399, n7398,
    n7400, n7410, n7403, n7402, n7408, n7406, n7405, n7407, n7409, n7426,
    n7412, n7411, n7416, n7414, n7413, n7415, n7418, n7417, n7422, n7420,
    n7419, n7421, n7423, n7425, n7427, n9849, n7431, n7430, n7436, n7434,
    n8693, n7433, n7435, n7444, n7438, n7437, n7442, n7440, n7439, n7441,
    n7443, n7460, n7446, n7445, n7450, n7448, n7447, n7449, n7458, n7452,
    n7451, n7456, n7454, n7453, n7455, n7459, n7461, n7463, n7462, n7467,
    n7465, n7464, n7466, n7468, n7471, n7470, n7476, n7474, n7473, n7475,
    n7484, n7478, n7477, n7482, n7480, n7479, n7481, n7483, n7485, n7490,
    n7489, n9132, n7491, n9302, n7493, n7494, n9187, n13311, n7497, n7538,
    n7499, n7498, n7500, n7502, n7503, n7508, n7506, n7505, n7507, n7674,
    n7509, n7510, n7513, n9454, n7514, n7527, n7517, n9322, n7520, n7519,
    n7525, n7521, n7523, n13653, n7522, n7524, n7526, n13743, n7528, n7534,
    n7535, n9156, n7536, n9174, n9142, n7539, n7540, n7542, n7549, n7545,
    n7543, n7547, n7551, n7548, n7559, n7557, n13353, n11903, n7553, n7555,
    n7554, n7556, n7724, n7562, n7594, n7880, n7564, n8892, n7563, n7568,
    n8567, n7566, n9401, n7565, n7567, n7576, n7734, n7570, n7569, n7574,
    n7572, n8537, n7571, n7573, n7575, n7592, n7578, n7798, n7577, n7582,
    n7580, n7579, n7581, n7590, n8915, n7584, n7920, n7583, n7588, n7692,
    n7586, n8399, n7807, n7585, n7587, n7589, n7591, n7593, n7596, n7598,
    n7597, n7599, n7602, n7636, n7605, n7604, n7609, n7607, n7606, n7608,
    n7618, n7611, n7610, n7616, n7614, n7613, n7615, n7617, n7634, n7620,
    n7619, n7624, n7622, n7621, n7623, n7632, n7626, n7625, n7630, n7628,
    n7627, n7629, n7631, n7633, n7846, n7638, n7637, n7643, n7641, n7640,
    n7642, n7651, n7645, n7644, n7649, n7647, n7646, n7648, n7650, n7668,
    n7654, n7653, n7658, n7656, n7655, n7657, n7666, n7660, n7659, n7664,
    n7662, n7661, n7663, n7665, n7667, n7670, n7669, n7671, n7719, n7710,
    n7677, n7676, n7681, n7679, n7678, n7680, n7689, n7683, n7682, n7687,
    n7685, n7684, n7686, n7688, n7706, n7691, n7690, n7696, n9398, n7694,
    n7693, n7695, n7704, n7698, n7697, n7702, n7700, n7699, n7701, n7703,
    n7705, n7709, n7969, n7707, n7708, n7713, n7711, n7712, n7715, n7714,
    n7856, n7717, n7718, n7723, n7721, n7722, n7830, n7731, n7725, n12240,
    n12508, n12500, n7726, n12928, n13205, n13197, n12589, n7729, n7728,
    n7732, n7768, n7766, n8130, n7736, n7735, n7740, n7738, n7737, n7739,
    n7748, n7742, n7741, n7746, n7744, n7743, n7745, n7747, n7764, n7750,
    n7927, n7749, n7754, n7752, n7751, n7753, n7762, n7756, n7755, n7760,
    n7758, n7757, n7759, n7761, n7763, n7765, n7770, n7772, n7782, n7863,
    n7778, n7864, n7776, n7775, n7777, n7780, n7824, n11528, n7779, n7781,
    n7817, n7785, n7784, n7789, n7787, n7786, n7788, n7797, n7791, n7790,
    n7795, n7793, n7792, n7794, n7796, n7815, n7800, n7799, n7804, n7802,
    n7801, n7803, n7813, n7806, n7805, n7811, n7809, n7808, n7810, n7812,
    n7814, n7816, n8980, n7818, n7828, n7823, n7821, n8929, n7819, n7820,
    n7822, n7826, n11522, n7825, n7827, n7832, n7831, n7833, n7835, n7834,
    n7843, n7841, n11547, n7836, n7839, n7838, n7840, n7842, n7874, n7873,
    n7854, n7852, n7850, n7849, n7851, n7853, n10887, n7858, n7857, n7860,
    n7862, n10923, n7870, n7868, n7866, n7865, n7867, n7869, n7872, n7871,
    n10886, n10889, n7876, n10766, n7910, n7879, n7878, n7884, n7882,
    n7881, n7883, n7892, n7886, n7885, n7890, n7888, n7887, n7889, n7891,
    n7908, n7894, n7893, n7898, n7896, n7895, n7897, n7906, n7900, n7899,
    n7904, n7902, n7901, n7903, n7905, n7907, n7909, n7958, n7946, n7913,
    n7912, n7917, n7915, n7914, n7916, n7926, n7919, n7918, n7924, n8910,
    n7922, n7921, n7923, n7925, n7944, n7929, n7928, n7933, n7931, n7930,
    n7932, n7942, n7935, n7934, n7940, n7938, n7937, n7939, n7941, n7943,
    n7945, n7955, n7949, n7947, n7948, n7953, n7959, n7951, n11493, n7952,
    n7954, n10765, n7963, n11509, n7961, n7960, n7962, n7964, n10767,
    n7968, n7972, n7970, n7971, n7973, n7974, n7981, n11487, n7979, n7977,
    n7976, n7978, n7980, n11471, n7986, n7984, n7983, n7985, n8021, n8143,
    n7990, n7989, n7994, n7992, n7991, n7993, n8002, n7996, n7995, n8000,
    n7998, n7997, n7999, n8001, n8018, n8004, n8003, n8008, n8006, n8005,
    n8007, n8016, n8010, n8009, n8014, n8012, n8011, n8013, n8015, n8017,
    n11463, n8026, n8024, n8023, n8025, n8059, n8028, n8027, n8033, n8031,
    n8030, n8032, n8049, n8035, n8034, n8039, n8037, n8036, n8038, n8047,
    n8041, n8040, n8045, n8043, n8526, n8042, n8044, n8046, n8048, n8057,
    n8051, n8050, n8055, n8053, n8052, n8054, n8056, n8058, n11446, n8066,
    n8064, n8063, n8065, n8102, n8067, n8070, n8068, n8069, n8075, n8073,
    n8071, n8072, n8074, n8091, n8077, n8076, n8081, n8151, n8079, n8078,
    n8080, n8089, n8083, n8082, n8087, n8085, n8084, n8086, n8088, n8090,
    n8099, n8093, n8092, n8097, n8095, n8094, n8096, n8098, n8100, n8101,
    n8107, n11430, n8105, n8104, n8106, n8141, n8109, n8108, n8113, n8111,
    n8110, n8112, n8129, n8115, n8114, n8119, n8117, n8116, n8118, n8127,
    n8121, n8120, n8125, n8123, n8122, n8124, n8126, n8128, n8138, n8132,
    n8131, n8136, n8134, n8133, n8135, n8137, n8139, n8140, n10662, n8144,
    n8146, n8145, n8150, n8148, n8147, n8149, n8168, n8153, n8152, n8158,
    n8156, n8155, n8157, n8166, n8160, n8159, n8164, n8162, n8161, n8163,
    n8165, n8167, n8176, n8170, n8169, n8174, n8172, n8171, n8173, n8175,
    n8177, n8178, n11412, n8181, n8186, n8184, n8182, n8183, n8185, n8187,
    n8189, n8191, n8190, n8195, n8193, n8192, n8194, n8211, n8197, n8196,
    n8201, n8199, n8198, n8200, n8209, n8203, n8202, n8207, n8205, n8204,
    n8206, n8208, n8210, n8219, n8213, n8212, n8217, n8215, n8214, n8216,
    n8218, n8220, n10624, n8226, n8224, n8223, n8225, n10149, n8228,
    n10605, n8234, n8232, n8230, n8231, n8233, n8267, n8236, n8235, n8240,
    n8238, n8237, n8239, n8256, n8242, n8241, n8246, n8244, n8243, n8245,
    n8254, n8248, n8247, n8252, n8250, n8249, n8251, n8253, n8255, n8264,
    n8258, n8257, n8262, n8260, n8259, n8261, n8263, n8265, n10135, n10590,
    n8272, n8270, n8269, n8271, n8307, n8274, n8273, n8278, n8276, n8275,
    n8277, n8295, n8281, n8280, n8285, n8283, n8282, n8284, n8293, n8287,
    n8286, n8291, n8289, n8288, n8290, n8292, n8294, n8303, n8297, n8296,
    n8301, n8299, n8298, n8300, n8302, n8304, n8311, n8313, n8312, n8317,
    n8315, n8314, n8316, n8325, n8319, n8318, n8323, n8321, n8320, n8322,
    n8324, n8341, n8327, n8326, n8331, n8329, n8328, n8330, n8339, n8333,
    n8332, n8337, n8335, n8334, n8336, n8338, n8340, n8342, n8349, n8347,
    n8345, n10559, n10571, n8344, n8346, n8348, n10555, n8390, n8353,
    n8352, n8357, n8355, n8354, n8356, n8365, n8359, n8358, n8363, n8361,
    n8360, n8362, n8364, n8381, n8367, n8366, n8371, n8369, n8368, n8370,
    n8379, n8373, n8372, n8377, n8375, n8374, n8376, n8378, n8380, n8382,
    n8386, n8383, n8385, n8388, n8387, n8389, n10093, n10537, n8393, n8436,
    n8394, n8396, n8395, n8403, n8397, n8401, n8398, n8400, n8402, n8419,
    n8405, n8404, n8409, n8407, n8406, n8408, n8417, n8411, n8410, n8415,
    n8413, n8412, n8414, n8416, n8418, n8428, n8422, n8420, n8421, n8426,
    n8424, n8423, n8425, n8427, n8429, n8434, n8432, n8430, n8431, n8433,
    n8435, n10061, n8476, n8438, n8472, n8440, n8439, n8444, n8442, n8441,
    n8443, n8452, n8446, n8445, n8450, n8448, n8447, n8449, n8451, n8469,
    n8455, n8454, n8459, n8457, n8456, n8458, n8467, n8461, n8460, n8465,
    n8463, n8462, n8464, n8466, n8468, n8470, n8471, n8474, n8473, n8475,
    n9765, n8480, n8479, n8484, n8482, n8481, n8483, n8500, n8486, n8485,
    n8490, n8488, n8487, n8489, n8498, n8492, n8491, n8496, n8494, n8493,
    n8495, n8497, n8499, n8508, n8502, n8501, n8506, n8504, n8503, n8505,
    n8507, n8509, n8514, n8512, n8510, n8511, n8513, n8518, n8516, n10048,
    n8517, n9744, n8519, n8554, n8521, n8520, n8525, n8523, n8522, n8524,
    n8534, n8528, n8527, n8532, n8530, n8529, n8531, n8533, n8551, n8536,
    n8535, n8541, n8539, n8907, n8538, n8540, n8549, n8543, n8542, n8547,
    n8545, n8544, n8546, n8548, n8550, n8552, n8553, n8556, n8555, n8559,
    n10034, n8558, n8561, n8560, n8566, n8564, n8563, n8565, n8583, n8569,
    n8568, n8573, n8571, n8570, n8572, n8581, n8575, n8574, n8579, n8577,
    n8576, n8578, n8580, n8582, n8593, n8585, n8584, n8591, n8589, n8588,
    n8590, n8592, n8594, n8599, n8597, n8595, n8596, n8598, n8603, n8601,
    n10022, n8602, n8605, n8604, n8609, n8607, n8606, n8608, n8617, n8611,
    n8610, n8615, n8613, n8612, n8614, n8616, n8633, n8619, n8618, n8623,
    n8621, n8620, n8622, n8631, n8625, n8624, n8629, n8627, n8626, n8628,
    n8630, n8632, n8677, n8635, n8634, n8639, n8637, n8636, n8638, n8648,
    n8641, n8640, n8646, n8644, n8643, n8645, n8647, n8664, n8650, n8649,
    n8654, n8652, n8651, n8653, n8662, n8656, n8655, n8660, n8658, n8657,
    n8659, n8661, n8663, n8678, n8665, n8670, n8668, n8667, n8669, n8671,
    n8674, n10010, n8673, n9684, n8718, n8680, n8679, n8684, n8682, n8681,
    n8683, n8692, n8686, n8685, n8690, n8688, n8687, n8689, n8691, n8709,
    n8695, n8694, n8699, n8697, n8696, n8698, n8707, n8701, n8700, n8705,
    n8703, n8702, n8704, n8706, n8708, n8719, n8710, n8717, n8715, n8713,
    n9669, n8712, n8714, n8791, n8721, n8720, n8725, n8723, n8722, n8724,
    n8733, n8727, n8726, n8731, n8729, n8728, n8730, n8732, n8749, n8735,
    n8734, n8739, n8737, n8736, n8738, n8747, n8741, n8740, n8745, n8743,
    n8742, n8744, n8746, n8748, n8792, n8750, n8755, n8752, n8751, n8753,
    n8754, n8758, n9990, n8757, n8759, n9636, n9977, n8800, n8762, n8761,
    n8766, n8764, n8763, n8765, n8774, n8768, n8767, n8772, n8770, n8769,
    n8771, n8773, n8790, n8776, n8775, n8780, n8778, n8777, n8779, n8788,
    n8782, n8781, n8786, n8784, n8783, n8785, n8787, n8789, n8802, n8793,
    n8798, n8796, n8794, n8795, n8797, n8799, n8804, n8803, n8808, n8806,
    n8805, n8807, n8816, n8810, n8809, n8814, n8812, n8811, n8813, n8815,
    n8832, n8818, n8817, n8822, n8820, n8819, n8821, n8830, n8824, n8823,
    n8828, n8826, n8825, n8827, n8829, n8831, n8878, n8833, n8838, n8835,
    n8834, n8836, n8837, n8841, n8845, n9965, n8840, n9607, n8844, n8933,
    n9949, n8847, n8846, n8851, n8849, n8848, n8850, n8860, n8853, n8852,
    n8858, n8856, n8855, n8857, n8859, n8876, n8862, n8861, n8866, n8864,
    n8863, n8865, n8874, n8868, n8867, n8872, n8870, n8869, n8871, n8873,
    n8875, n8889, n8879, n8885, n8883, n8881, n8882, n8884, n8886, n9586,
    n8891, n8890, n8896, n8894, n8893, n8895, n8905, n8898, n8897, n8903,
    n8901, n8900, n8902, n8904, n8925, n8909, n8908, n8914, n8912, n8911,
    n8913, n8923, n8917, n8916, n8921, n8919, n8918, n8920, n8922, n8924,
    n9432, n8926, n8932, n8928, n8927, n8930, n8931, n8935, n9397, n9573,
    n8934, n8936, n8937, n11563, n8943, n8941, n8962, n8942, n9326, n8949,
    n8945, n8948, n8947, n11562, n8950, n8953, n11564, n8951, n8952,
    n11555, n11535, n8965, n8959, n8957, n8956, n8960, n8982, n8961, n8963,
    n8964, n8967, n8974, n11747, n8966, n8972, n8971, n8968, n8969, n8970,
    n11540, n8979, n8977, n8975, n8976, n8978, n11518, n8984, n8988, n8983,
    n9529, n8987, n8986, n11508, n8990, n8995, n8991, n8992, n11497, n8997,
    n9009, n8998, n8999, n9003, n9000, n9008, n9019, n9010, n9011, n11678,
    n9014, n9016, n9018, n9020, n9022, n9021, n11476, n9023, n9025, n9027,
    n11452, n11616, n9028, n11433, n9030, n9031, n9033, n10143, n10397,
    n10114, n10117, n9036, n10370, n9037, n10071, n10070, n10337, n10321,
    n9038, n9039, n9040, n10280, n9042, n10268, n9165, n9044, n9043, n9164,
    n9045, n9169, n9046, n9047, n9049, n9335, n9048, n9050, n9347, n9051,
    n9052, n9054, n10228, n9053, n9984, n9055, n9056, n9972, n10201, n9959,
    n10193, n9973, n9960, n9945, n9057, n9357, n9059, n9058, n9063, n9069,
    n9076, n9079, n9061, n9070, n9062, n9108, n9065, n9064, n9150, n9066,
    n9117, n9068, n9067, n9116, n9121, n9089, n9149, n9071, n9073, n9072,
    n9075, n9074, n9104, n9078, n9077, n9080, n9153, n9082, n9084, n9083,
    n9086, n9087, n9102, n9100, n9091, n9090, n9098, n9092, n9094, n9096,
    n9095, n9097, n9099, n9101, n9103, n9106, n9111, n9148, n9110, n9112,
    n9114, n9118, n9124, n9127, n9134, n9133, n13331, n10176, n13736,
    n9137, n9138, n9141, n9139, n9496, n11580, n9140, n9144, n13304,
    n13735, n13762, n9151, n9152, n9154, n13320, n9157, n9158, n9159,
    n9160, n9163, n10042, n10041, n9166, n10030, n9998, n10256, n10003,
    n9167, n9171, n9170, n9172, n13739, n10434, n9175, n9176, n9180, n9177,
    n9178, n9308, n9179, n9181, n9185, n9183, n9184, n9186, n9190, n9188,
    n9189, n9316, n9193, n9203, n9192, n9194, n9195, n9196, n9197, n9198,
    n9200, n9331, n9204, n9202, n13318, n9208, n9206, n9205, n9207, n9209,
    n9353, n9212, n9215, n9213, n9359, n9217, n9216, n9219, n9227, n9226,
    n9221, n9224, n9222, n9223, n10911, n9229, n9507, n9228, n9231, n10863,
    n9233, n9234, n9236, n9237, n10802, n9238, n9240, n9241, n10787, n9243,
    n9244, n10762, n9246, n9247, n10734, n10725, n9249, n9248, n9250,
    n10724, n9252, n9253, n10694, n9255, n9254, n9256, n10675, n10666,
    n9258, n9257, n9259, n10665, n9261, n9260, n9262, n10645, n9264, n9263,
    n9265, n10422, n9267, n9266, n9268, n10408, n9270, n9269, n9271,
    n10376, n9273, n9272, n9274, n10358, n9276, n9275, n9277, n10341,
    n9279, n9278, n9280, n10324, n9282, n9281, n9283, n9767, n9285, n9287,
    n9745, n9289, n9288, n9290, n9726, n9293, n9294, n9704, n9296, n9297,
    n9686, n9820, n9299, n13380, n9300, n9301, n9486, n9351, n11795, n9306,
    n9305, n9324, n9312, n9310, n9309, n9311, n9314, n9313, n9318, n9317,
    n9319, n11834, n9321, n11847, n9323, n9325, n11794, n9334, n9329,
    n10399, n10387, n9333, n9332, n11731, n11713, n11728, n9327, n11659,
    n11665, n11630, n11599, n9328, n10353, n10278, n10314, n10286, n9344,
    n13324, n11818, n9337, n11752, n11662, n11627, n11602, n10349, n10394,
    n10355, n10315, n10283, n9343, n9336, n9338, n10269, n10259, n11689,
    n9339, n9341, n11778, n11765, n11625, n9340, n9342, n10229, n9346,
    n9345, n9348, n9349, n9350, n9352, n9383, n9354, n9355, n9356, n9358,
    n9934, n9394, n9361, n9362, n9648, n9629, n9364, n9365, n9630, n9609,
    n9367, n9368, n9608, n9370, n9371, n9589, n9373, n9374, n9567, n9505,
    n9375, n9376, n9380, n9379, n9504, n9381, n9938, n9384, n9382, n10230,
    n9385, n9387, n10179, n10159, n9392, n11780, n9386, n9388, n10178,
    n9390, n9393, n9396, n9936, n9445, n9400, n9399, n9405, n9403, n9402,
    n9404, n9414, n9407, n9406, n9412, n9410, n9409, n9411, n9413, n9430,
    n9416, n9415, n9420, n9418, n9417, n9419, n9428, n9422, n9421, n9426,
    n9424, n9423, n9425, n9427, n9429, n9434, n9433, n9436, n9443, n9437,
    n9441, n9439, n9440, n9442, n9444, n9541, n9448, n9447, n9457, n10448,
    n10439, n9449, n9787, n9450, n9453, n13431, n9455, n9459, n9458, n9461,
    n11037, n9460, n10165, n9463, n9465, n9467, n9469, n9478, n9476,
    n10161, n9470, n9474, n9472, n9473, n9475, n9477, n9492, n9484, n9483,
    n9819, n9490, n9485, n9488, n9487, n9489, n9491, n9495, n13409, n9497,
    n13398, n9498, n9499, n13392, n9500, n9539, n9506, n9509, n9508, n9510,
    n9526, n9553, n9512, n9537, n13568, n9513, n10851, n13563, n13558,
    n13548, n13539, n13529, n13519, n13509, n13499, n13489, n13479, n13469,
    n13722, n9515, n10812, n10778, n10760, n10739, n10722, n10693, n10680,
    n10659, n10612, n10619, n10597, n10582, n10563, n10542, n10527, n9773,
    n9756, n9736, n9707, n9695, n9657, n9668, n9517, n9650, n9633, n9613,
    n9521, n9571, n9523, n9516, n9535, n9518, n9519, n9520, n9632, n9522,
    n9572, n9524, n9544, n9533, n9525, n9531, n13379, n9528, n9530, n9532,
    n9534, n9536, n9538, n9542, n9935, n9565, n9563, n9546, n9545, n9549,
    n9547, n9548, n9561, n9551, n9559, n9556, n9552, n9554, n9555, n9557,
    n10904, n9558, n9560, n9562, n9564, n9585, n9569, n9583, n13589, n9581,
    n9592, n9579, n9577, n9575, n9574, n9576, n9578, n9580, n9582, n9584,
    n9604, n10188, n9590, n9602, n9591, n9600, n9598, n9596, n9594, n9593,
    n9595, n9597, n9599, n9601, n9603, n9606, n9963, n9871, n9625, n9610,
    n9612, n9623, n9619, n9615, n9614, n9617, n9616, n9618, n9621, n9620,
    n9622, n9624, n9628, n9975, n9878, n9646, n10214, n9631, n9644, n9635,
    n9634, n9642, n9638, n9637, n9640, n9639, n9641, n9643, n9645, n9885,
    n9665, n10225, n9649, n9663, n9656, n9652, n9651, n9654, n9653, n9655,
    n9661, n9667, n9658, n10831, n9676, n9698, n9659, n9660, n9662, n9664,
    n9892, n9682, n9666, n9680, n9675, n9673, n9671, n9670, n9672, n9674,
    n9678, n9677, n9679, n9681, n10007, n9899, n9702, n10243, n9694, n9687,
    n9690, n9689, n9692, n9691, n9693, n9700, n9696, n9697, n9699, n9701,
    n10019, n9906, n9722, n10251, n9716, n9706, n9714, n9708, n9712, n9710,
    n9709, n9711, n9713, n9715, n9720, n9717, n9759, n9735, n9718, n9719,
    n9721, n9724, n10031, n9913, n9742, n10265, n9734, n9727, n9732, n9730,
    n9729, n9731, n9733, n9738, n9737, n9740, n9739, n9741, n10044, n9763,
    n9746, n10291, n9748, n9755, n9749, n9837, n9753, n9751, n9750, n9752,
    n9754, n9761, n9757, n9758, n9760, n9762, n10059, n9927, n9785, n10303,
    n9771, n9769, n9768, n9770, n9775, n9772, n9774, n9783, n13534, n10525,
    n9776, n10545, n9777, n9781, n10814, n10784, n9779, n9780, n9782,
    n9784, n9790, n9789, n9792, n9791, n9793, n9798, n9796, n9795, n9797,
    n9802, n9800, n9799, n9801, n9806, n9804, n9803, n9805, n9810, n9808,
    n9807, n9809, n9814, n9812, n9811, n9813, n9818, n9816, n9815, n9817,
    n9824, n9822, n9821, n9823, n9828, n9826, n9825, n9827, n9832, n9830,
    n9829, n9831, n9836, n9834, n9833, n9835, n9841, n9839, n9838, n9840,
    n9846, n9842, n9844, n9843, n9845, n11049, n9856, n9850, n11043, n9852,
    n9851, n9854, n9853, n9855, n9863, n9859, n9858, n9861, n9860, n9862,
    n9870, n9866, n9865, n9868, n9867, n9869, n9877, n9873, n9872, n9875,
    n9874, n9876, n9884, n9880, n9879, n9882, n9881, n9883, n9891, n9887,
    n9886, n9889, n9888, n9890, n9898, n9894, n9893, n9896, n9895, n9897,
    n9905, n9901, n9900, n9903, n9902, n9904, n9912, n9908, n9907, n9910,
    n9909, n9911, n9919, n9915, n9914, n9917, n9916, n9918, n9925, n9921,
    n9920, n9923, n9922, n9924, n9933, n9929, n9928, n9931, n9930, n9932,
    n9944, n9942, n9940, n9937, n9939, n9941, n9946, n10187, n9956, n9953,
    n13584, n10190, n9951, n9950, n9952, n9954, n9958, n9962, n9961,
    n10199, n9971, n9969, n10207, n9964, n9967, n9966, n9968, n9970, n9974,
    n9983, n9981, n10215, n9976, n9979, n9978, n9980, n9982, n9986, n10224,
    n9996, n9994, n10226, n9989, n9992, n9991, n9993, n9995, n10001, n9999,
    n10000, n10002, n10005, n10017, n10006, n10238, n10016, n10014, n10244,
    n10009, n10008, n10012, n10011, n10013, n10015, n10250, n10028, n10026,
    n13553, n10252, n10021, n10020, n10024, n10023, n10025, n10027, n10264,
    n10040, n10038, n10266, n10033, n10032, n10036, n10035, n10037, n10039,
    n10043, n10277, n10055, n10053, n10045, n10296, n10047, n10046, n10051,
    n10049, n10050, n10052, n10054, n10302, n10067, n10065, n10305, n10060,
    n10063, n10062, n10064, n10066, n10069, n10101, n10072, n10076, n10073,
    n10075, n10077, n10313, n10088, n10080, n10534, n10086, n10327, n10082,
    n10081, n10084, n10083, n10085, n10087, n10090, n10335, n10100, n11032,
    n10098, n10342, n10094, n10096, n10095, n10097, n10099, n10348, n10113,
    n10105, n11040, n10111, n10362, n10107, n10106, n10109, n10108, n10110,
    n10112, n10131, n10130, n10129, n10119, n10118, n10369, n10122, n10587,
    n10128, n10381, n10124, n10123, n10126, n10125, n10127, n10133, n10132,
    n10386, n10142, n11052, n10140, n10412, n10136, n10138, n10137, n10139,
    n10141, n10145, n10417, n10157, n10150, n10961, n11057, n10155, n10423,
    n10151, n10153, n10152, n10154, n10156, n10172, n10164, n10160, n10162,
    n10163, n10170, n10166, n10168, n10169, n10171, n10186, n10175, n10177,
    n10184, n10182, n10180, n10181, n10183, n10185, n10198, n10192, n10189,
    n10191, n10196, n10194, n10195, n10197, n10212, n10202, n10205, n10204,
    n10210, n10208, n10209, n10211, n10223, n10216, n10219, n10217, n10218,
    n10221, n10220, n10222, n10237, n10227, n10235, n10233, n10231, n10232,
    n10234, n10236, n10249, n10242, n10241, n10247, n10245, n10246, n10248,
    n10263, n10253, n10255, n10254, n10261, n10257, n10258, n10260, n10262,
    n10276, n10267, n10274, n10272, n10271, n10273, n10275, n10301, n10319,
    n10279, n10336, n10292, n10310, n11771, n10281, n10282, n10285, n10284,
    n10288, n10287, n10304, n10289, n10290, n10299, n10295, n10293, n10294,
    n10297, n10298, n10300, n10312, n10308, n10306, n10307, n10309, n10311,
    n10334, n10317, n10316, n10318, n10338, n10320, n10322, n10332, n10323,
    n10330, n10326, n10931, n10328, n10329, n10331, n10333, n10347, n10340,
    n10339, n10345, n10936, n10343, n10344, n10346, n10368, n11598, n10398,
    n11612, n10350, n10351, n10371, n10352, n10366, n11629, n10354, n10357,
    n10356, n10372, n10364, n10359, n10942, n10361, n10363, n10365, n10367,
    n10385, n10375, n10373, n10374, n10383, n10378, n10947, n10380, n10382,
    n10384, n10416, n10388, n10407, n10389, n10393, n10425, n10401, n10391,
    n10392, n10396, n10395, n10426, n10418, n10405, n10403, n10402, n10419,
    n10404, n10406, n10414, n10409, n10952, n10411, n10413, n10415, n10432,
    n10421, n10420, n10430, n10958, n10424, n10428, n10427, n10429, n10431,
    n10433, n10435, n10437, n10436, n10438, n10441, n10440, n10442, n10447,
    n10445, n10444, n10446, n10449, n10450, n13350, n10454, n11810, n10452,
    n13618, n10453, n10462, n10455, n10464, n10458, n11868, n10460, n10459,
    n10461, n10463, n13439, n10465, n10466, n10473, n10470, n10467, n10468,
    n10469, n10471, n10472, n10478, n10474, n10476, n13756, n10475, n13610,
    n10479, n13615, n13613, n10480, n10482, n10483, n13307, n13731, n10485,
    n13713, n13723, n10519, n10516, n10487, n10486, n10491, n10489, n10488,
    n10490, n10499, n10493, n10492, n10497, n10495, n10494, n10496, n10498,
    n10515, n10501, n10500, n10505, n10503, n10502, n10504, n10513, n10507,
    n10506, n10511, n10509, n10508, n10510, n10512, n10514, n13724, n10518,
    n13726, n10517, n10523, n10520, n10521, n10522, n10524, n10529, n10526,
    n10528, n10531, n10530, n10533, n10532, n10536, n11025, n10535, n10541,
    n10539, n10538, n10540, n10543, n10544, n10549, n10547, n10546, n10548,
    n10550, n10554, n10939, n10552, n10551, n10553, n10557, n10556, n10596,
    n10578, n10581, n10558, n10568, n10560, n10562, n10561, n10566, n10564,
    n10565, n10567, n10570, n10569, n10575, n10573, n10572, n10574, n10577,
    n10586, n10580, n10598, n10579, n10584, n10583, n10585, n10589, n10588,
    n10594, n10592, n10591, n10593, n10595, n10602, n10600, n10599, n10601,
    n10604, n10603, n10609, n10955, n10607, n10606, n10608, n10611, n10610,
    n13504, n10632, n10633, n10658, n10653, n10613, n10617, n10615, n10616,
    n10621, n10618, n10620, n10623, n10622, n10628, n10626, n10625, n10627,
    n10630, n10629, n10631, n10635, n10634, n10637, n10636, n10639, n10638,
    n10651, n10640, n11062, n11415, n10643, n10642, n10649, n10646, n11589,
    n10648, n10650, n10652, n10655, n10654, n10657, n10656, n10661, n10660,
    n10671, n11067, n11443, n10664, n10663, n10669, n10667, n11609, n10668,
    n10670, n10692, n10723, n10714, n10672, n10691, n10673, n10677, n11622,
    n10676, n10679, n10678, n10683, n10681, n10682, n10687, n11072, n11449,
    n10686, n10689, n10688, n10690, n10698, n10696, n10695, n11640, n10697,
    n10711, n10700, n10699, n10702, n10701, n10703, n10709, n11077, n11468,
    n10707, n10706, n10708, n10710, n10713, n10712, n10716, n13484, n10715,
    n10717, n10721, n10719, n11474, n11082, n10720, n10731, n10727, n11653,
    n10726, n10729, n10728, n10730, n10733, n10743, n11672, n10737, n10736,
    n10741, n10738, n10740, n10742, n10748, n10746, n10747, n10754, n10910,
    n10749, n10777, n10761, n10750, n10752, n10751, n10753, n10756, n10755,
    n10759, n10757, n10758, n10776, n10764, n11685, n10763, n10774, n10768,
    n10769, n11091, n10772, n10771, n10773, n10775, n10781, n10779, n10780,
    n10799, n10783, n10786, n10785, n10792, n10789, n11707, n10791, n10797,
    n11098, n11514, n10794, n10924, n10796, n10798, n10801, n10800, n11722,
    n10805, n10804, n10808, n10806, n10807, n10818, n10881, n10903, n10811,
    n10810, n10816, n10833, n10838, n10813, n10815, n10817, n10820, n10819,
    n10827, n10824, n10823, n10825, n10996, n10826, n10829, n10828, n10835,
    n10895, n10832, n10854, n10834, n10845, n11738, n10840, n10839, n10843,
    n10842, n10844, n10847, n10846, n10850, n11107, n11533, n10849, n13454,
    n10852, n10853, n10861, n10856, n12248, n10859, n10857, n10858, n10860,
    n10878, n10866, n10865, n11758, n10868, n10867, n10876, n10874, n10870,
    n10872, n11551, n10873, n10875, n10877, n10880, n10883, n10882, n10885,
    n10884, n10892, n10890, n10888, n11571, n10891, n10902, n10894, n10898,
    n10897, n10900, n10899, n10901, n10906, n10905, n10920, n10909, n10918,
    n10916, n10913, n11791, n10915, n10917, n10919, n10926, n10922, n11586,
    n10925, n10928, n10930, n10929, n10933, n10932, n10935, n10934, n10938,
    n10937, n10941, n10940, n10944, n10943, n10946, n10945, n10949, n10948,
    n10951, n10950, n10954, n10953, n10957, n10956, n10960, n10959, n10963,
    n10962, n10965, n10964, n10967, n10966, n10969, n10968, n10971, n10970,
    n10973, n10972, n10975, n10974, n10977, n10976, n10979, n10978, n10981,
    n10980, n10983, n10982, n10985, n10984, n10987, n10986, n10989, n10988,
    n10991, n10990, n10993, n10992, n10995, n10994, n10998, n10997, n11000,
    n10999, n11003, n11002, n11005, n11004, n11007, n11112, n11006, n11009,
    n11008, n11012, n11011, n11015, n11014, n11019, n11018, n11022, n11021,
    n11024, n11023, n11027, n11026, n11029, n11028, n11031, n11030, n11034,
    n11033, n11036, n11035, n11039, n11038, n11042, n11041, n11045, n11044,
    n11048, n11406, n11047, n11051, n11050, n11054, n11398, n11053, n11056,
    n11055, n11059, n11393, n11058, n11061, n11060, n11064, n11388, n11063,
    n11066, n11065, n11069, n11383, n11068, n11071, n11070, n11074, n11378,
    n11073, n11076, n11075, n11079, n11373, n11078, n11081, n11080, n11084,
    n11368, n11083, n11086, n11085, n11088, n11363, n11087, n11090, n11089,
    n11094, n11358, n11093, n11096, n11095, n11951, n11100, n11099, n11102,
    n11101, n11941, n11104, n11103, n11106, n11105, n11931, n11109, n11108,
    n11111, n11110, n11921, n11114, n11113, n11116, n11115, n11911, n11118,
    n11117, n11120, n11119, n11902, n11125, n11122, n11124, n11127, n11126,
    n11129, n11128, n11133, n11130, n11132, n11135, n11134, n11137, n11136,
    n11139, n11138, n11141, n11140, n11143, n11142, n11145, n11144, n11147,
    n11146, n11149, n11148, n11151, n11150, n11153, n11152, n11155, n11154,
    n11157, n11156, n11159, n11158, n11161, n11160, n11163, n11162, n11165,
    n11164, n11167, n11166, n11169, n11168, n11171, n11170, n11173, n11172,
    n11175, n11174, n11177, n11176, n11179, n11178, n11181, n11180, n11183,
    n11182, n11185, n11184, n11188, n11187, n11190, n11189, n11192, n11191,
    n11194, n11193, n11196, n11195, n11198, n11197, n11200, n11199, n11202,
    n11201, n11204, n11203, n11206, n11205, n11208, n11207, n11210, n11209,
    n11212, n11211, n11214, n11213, n11216, n11215, n11218, n11217, n11220,
    n11219, n11222, n11221, n11224, n11223, n11226, n11225, n11228, n11227,
    n11230, n11229, n11232, n11231, n11234, n11233, n11236, n11235, n11238,
    n11237, n11240, n11239, n11242, n11241, n11244, n11243, n11247, n11246,
    n11249, n11248, n11251, n11250, n11255, n11254, n11258, n11257, n11330,
    n11407, n11260, n11261, n11265, n11262, n11264, n11335, n11266, n11267,
    n11269, n11268, n11340, n11270, n11271, n11273, n11272, n11345, n11274,
    n11275, n11277, n11276, n11350, n11278, n11279, n11281, n11280, n11355,
    n11282, n11283, n11285, n11284, n11960, n11360, n11286, n11287, n11289,
    n11288, n11972, n11365, n11290, n11291, n11293, n11292, n11294, n11370,
    n11295, n11296, n11298, n11297, n11299, n11375, n11300, n11301, n11303,
    n11302, n11304, n11380, n11305, n11306, n11308, n11307, n11309, n11385,
    n11310, n11311, n11313, n11312, n11314, n11390, n11315, n11316, n11318,
    n11317, n11319, n11395, n11320, n11321, n11323, n11322, n11324, n11400,
    n11325, n11327, n11326, n11328, n11329, n11332, n11331, n11333, n11334,
    n11337, n11336, n11338, n11339, n11342, n11341, n11343, n11344, n11347,
    n11346, n11348, n11349, n11352, n11351, n11353, n11354, n11357, n11356,
    n11359, n11362, n11361, n11364, n11367, n11366, n11369, n11372, n11371,
    n11374, n11377, n11376, n11379, n11382, n11381, n11384, n11387, n11386,
    n11389, n11392, n11391, n11394, n11397, n11396, n11399, n11403, n11402,
    n11404, n11409, n11408, n11411, n11410, n11414, n11413, n11427, n11591,
    n11417, n11416, n11425, n11453, n11436, n11432, n11423, n11422, n11595,
    n11424, n11426, n11610, n11429, n11428, n11442, n11440, n11434, n11438,
    n11435, n11437, n11613, n11439, n11441, n11445, n11444, n11448, n11447,
    n11459, n13494, n11624, n11451, n11450, n11457, n11455, n11635, n11456,
    n11458, n11641, n11460, n11467, n11643, n11465, n11464, n11466, n11470,
    n11469, n11473, n11472, n11481, n11654, n11475, n11479, n11656, n11478,
    n11480, n11674, n11482, n11486, n11675, n11485, n11492, n11490, n11489,
    n11491, n11495, n11494, n11502, n11686, n11498, n11696, n11500, n11501,
    n11505, n11504, n11708, n11507, n11506, n11513, n11511, n11510, n11512,
    n11516, n11515, n11723, n11517, n11521, n11725, n11520, n11527, n11525,
    n11524, n11526, n11532, n11531, n11546, n11740, n11534, n11544, n11556,
    n11539, n11538, n11542, n11541, n11742, n11543, n11545, n11550, n11549,
    n11554, n11756, n11552, n11553, n11558, n11761, n11557, n11776, n11561,
    n11560, n11569, n11566, n11565, n11783, n11568, n11575, n11573, n11572,
    n11574, n11789, n11802, n11579, n11585, n11583, n11582, n11584, n11588,
    n11587, n11590, n11594, n11592, n11593, n11597, n11596, n11608, n11605,
    n11600, n11601, n11604, n11603, n11617, n11606, n11607, n11611, n11621,
    n11615, n11614, n11619, n11618, n11620, n11623, n11639, n11649, n11626,
    n11694, n11702, n11650, n11634, n11628, n11632, n11631, n11644, n11633,
    n11637, n11636, n11638, n11642, n11648, n11646, n11645, n11647, n11652,
    n11651, n11655, n11658, n11657, n11671, n11660, n11746, n11680, n11661,
    n11669, n11664, n11667, n11666, n11679, n11668, n11670, n11673, n11677,
    n11676, n11684, n11682, n11681, n11683, n11687, n11700, n11688, n11762,
    n11712, n11701, n11691, n11690, n11692, n11716, n11693, n11710, n11695,
    n11698, n11697, n11699, n11706, n11704, n11703, n11705, n11709, n11711,
    n11718, n11714, n11715, n11717, n11721, n11720, n11724, n11727, n11726,
    n11737, n11730, n11729, n11735, n11753, n11733, n11745, n11734, n11736,
    n11741, n11744, n11743, n11751, n11749, n11748, n11750, n11754, n11755,
    n11757, n11760, n11759, n11770, n11764, n11763, n11768, n11766, n11767,
    n11769, n11790, n11774, n11788, n11777, n11782, n11779, n11781, n11786,
    n11785, n11787, n11801, n11793, n11799, n11797, n11798, n11800, n11805,
    n11804, n13749, n11807, n11872, n11859, n11811, n11864, n11845, n11848,
    n11822, n11815, n11814, n11816, n11817, n11843, n11850, n11824, n11823,
    n11825, n11827, n11836, n11832, n11830, n11831, n11833, n13341, n11835,
    n11841, n11837, n11838, n13620, n11839, n11840, n11842, n13622, n11844,
    n11846, n11858, n11857, n11851, n11855, n11849, n11853, n11852, n11854,
    n11856, n13630, n11861, n11860, n13362, n11862, n11863, n13372, n11866,
    n11877, n11870, n11869, n11871, n11875, n11874, n13334, n11876, n13305,
    n11878, n11879, n13188, n12063, n11984, n11968, n11883, n13210, n11882,
    n11897, n12259, n12764, n11891, n13695, n12596, n11889, n11885, n11886,
    n11887, n11888, n11890, n11892, n11895, n11893, n12588, n12260, n11894,
    n12257, n11971, n11896, n11900, n13189, n11899, n11907, n13207, n13675,
    n12429, n12675, n11905, n12064, n12774, n11904, n11973, n11906, n13215,
    n11910, n13216, n11909, n11917, n11913, n13219, n11912, n11915, n13222,
    n11914, n11916, n11920, n13228, n11919, n11927, n11923, n13231, n11922,
    n11925, n13234, n11924, n11926, n13239, n11930, n13246, n11929, n11937,
    n11933, n13243, n11932, n11935, n13240, n11934, n11936, n13251, n11940,
    n13258, n11939, n11947, n11943, n13255, n11942, n11945, n13252, n11944,
    n11946, n11950, n13264, n11949, n11957, n11953, n13267, n11952, n11955,
    n13270, n11954, n11956, n13275, n11959, n13282, n11958, n11966, n11962,
    n13279, n11961, n11964, n13276, n11963, n11965, n13288, n11970, n13298,
    n11969, n11979, n11975, n13295, n11974, n11977, n13289, n11976, n11978,
    n12051, n11982, n11981, n11993, n11985, n11991, n12499, n11996, n12850,
    n11986, n11987, n11998, n11988, n13674, n11989, n11990, n12055, n11992,
    n11995, n11994, n12002, n11997, n12000, n12162, n11999, n12056, n12001,
    n12004, n12003, n12010, n12006, n12005, n12008, n12007, n12009, n12012,
    n12011, n12018, n12014, n12013, n12016, n12015, n12017, n12020, n12019,
    n12026, n12022, n12021, n12024, n12023, n12025, n12028, n12027, n12034,
    n12030, n12029, n12032, n12031, n12033, n12036, n12035, n12042, n12038,
    n12037, n12040, n12039, n12041, n12044, n12043, n12050, n12046, n12045,
    n12048, n12047, n12049, n12054, n12053, n12062, n12058, n12057, n12060,
    n12059, n12061, n12174, n12144, n12069, n12067, n12427, n12066, n12756,
    n12071, n12065, n12143, n12068, n12078, n12167, n12070, n13193, n12072,
    n12073, n12074, n12076, n12421, n12075, n12147, n12077, n12080, n12079,
    n12083, n12081, n12082, n12084, n12086, n12085, n12088, n12087, n12090,
    n12089, n12093, n12091, n12092, n12094, n12096, n12095, n12098, n12097,
    n12100, n12099, n12103, n12101, n12102, n12104, n12106, n12105, n12108,
    n12107, n12110, n12109, n12112, n12536, n12111, n12113, n12115, n12114,
    n12117, n12116, n12119, n12118, n12121, n12545, n12120, n12122, n12124,
    n12123, n12126, n12125, n12128, n12127, n12131, n12129, n12130, n12132,
    n12134, n12133, n12136, n12135, n12138, n12137, n12141, n12139, n12140,
    n12142, n12146, n12145, n12149, n12148, n12152, n12151, n12156, n12153,
    n12155, n12228, n12158, n12157, n12166, n13684, n12159, n13685, n12160,
    n12171, n12161, n12173, n12164, n12163, n12232, n12165, n12169, n12168,
    n12179, n12170, n12172, n12176, n12175, n12177, n12231, n12178, n12181,
    n12180, n12187, n12183, n12182, n12185, n12184, n12186, n12189, n12188,
    n12195, n12191, n12190, n12193, n12192, n12194, n12197, n12196, n12203,
    n12199, n12198, n12201, n12200, n12202, n12205, n12204, n12211, n12207,
    n12206, n12209, n12208, n12210, n12213, n12212, n12219, n12215, n12214,
    n12217, n12216, n12218, n12221, n12220, n12227, n12223, n12222, n12225,
    n12224, n12226, n12230, n12229, n12239, n12234, n12233, n12237, n12236,
    n12238, n12241, n12344, n12317, n12245, n12243, n12244, n12268, n12247,
    n12256, n12932, n12254, n12250, n12251, n12252, n12253, n12255, n12258,
    n12320, n12264, n13112, n12262, n12261, n12321, n12263, n12266, n12265,
    n12267, n12270, n12269, n12276, n12272, n12271, n12274, n12273, n12275,
    n12278, n12277, n12284, n12280, n12279, n12282, n12281, n12283, n12286,
    n12285, n12292, n12288, n12287, n12290, n12289, n12291, n12294, n12293,
    n12300, n12296, n12295, n12298, n12297, n12299, n12302, n12301, n12308,
    n12304, n12303, n12306, n12305, n12307, n12310, n12309, n12316, n12312,
    n12311, n12314, n12313, n12315, n12319, n12318, n12328, n12323, n12322,
    n12326, n12325, n12327, n12398, n12331, n12330, n12338, n12332, n12342,
    n12333, n12334, n12341, n12336, n12335, n12403, n12337, n12340, n12339,
    n12349, n12343, n12346, n12345, n12347, n12402, n12348, n12351, n12350,
    n12357, n12353, n12352, n12355, n12354, n12356, n12359, n12358, n12365,
    n12361, n12360, n12363, n12362, n12364, n12367, n12366, n12373, n12369,
    n12368, n12371, n12370, n12372, n12375, n12374, n12381, n12377, n12376,
    n12379, n12378, n12380, n12383, n12382, n12389, n12385, n12384, n12387,
    n12386, n12388, n12391, n12390, n12397, n12393, n12392, n12395, n12394,
    n12396, n12401, n12400, n12409, n12405, n12404, n12407, n12406, n12408,
    n12482, n12412, n12410, n12411, n12424, n13096, n12417, n12413, n12414,
    n12415, n12416, n12419, n12418, n12420, n12422, n12486, n12423, n12426,
    n12425, n12433, n12428, n12431, n13195, n12430, n12487, n12432, n12435,
    n12434, n12441, n12437, n12436, n12439, n12438, n12440, n12443, n12442,
    n12449, n12445, n12444, n12447, n12446, n12448, n12451, n12450, n12457,
    n12453, n12452, n12455, n12454, n12456, n12459, n12458, n12465, n12461,
    n12460, n12463, n12462, n12464, n12467, n12466, n12473, n12469, n12468,
    n12471, n12470, n12472, n12475, n12474, n12481, n12477, n12476, n12479,
    n12478, n12480, n12485, n12484, n12493, n12489, n12488, n12491, n12490,
    n12492, n12573, n12496, n12494, n12495, n12517, n12497, n12498, n12505,
    n12501, n12506, n12503, n12502, n12504, n12578, n12512, n12507, n12510,
    n12509, n12579, n12511, n12515, n12513, n12514, n12516, n12520, n12518,
    n12519, n12526, n12522, n12521, n12524, n12523, n12525, n12529, n12527,
    n12528, n12535, n12531, n12530, n12533, n12532, n12534, n12538, n12537,
    n12544, n12540, n12539, n12542, n12541, n12543, n12547, n12546, n12554,
    n12549, n12548, n12552, n12551, n12553, n12557, n12555, n12556, n12563,
    n12559, n12558, n12561, n12560, n12562, n12566, n12564, n12565, n12572,
    n12568, n12567, n12570, n12569, n12571, n12577, n12574, n12576, n12585,
    n12581, n12580, n12583, n12582, n12584, n12587, n12753, n12687, n12658,
    n12586, n12593, n12943, n12591, n12590, n12663, n12592, n12595, n12760,
    n12594, n12609, n12604, n12602, n12597, n12599, n12600, n12601, n12603,
    n12605, n12607, n12606, n12939, n12608, n12611, n12610, n12617, n12613,
    n12612, n12615, n12614, n12616, n12619, n12618, n12625, n12621, n12620,
    n12623, n12622, n12624, n12627, n12626, n12633, n12629, n12628, n12631,
    n12630, n12632, n12635, n12634, n12641, n12637, n12636, n12639, n12638,
    n12640, n12643, n12642, n12649, n12645, n12644, n12647, n12646, n12648,
    n12651, n12650, n12657, n12653, n12652, n12655, n12654, n12656, n12661,
    n12660, n12669, n12665, n12664, n12667, n12666, n12668, n12741, n12671,
    n12844, n12670, n12681, n12672, n12674, n12684, n13335, n12676, n12677,
    n12685, n12679, n12859, n12678, n12745, n12680, n12683, n12682, n12692,
    n12686, n12689, n12688, n12690, n12744, n12691, n12694, n12693, n12700,
    n12696, n12695, n12698, n12697, n12699, n12702, n12701, n12708, n12704,
    n12703, n12706, n12705, n12707, n12710, n12709, n12716, n12712, n12711,
    n12714, n12713, n12715, n12718, n12717, n12724, n12720, n12719, n12722,
    n12721, n12723, n12726, n12725, n12732, n12728, n12727, n12730, n12729,
    n12731, n12734, n12733, n12740, n12736, n12735, n12738, n12737, n12739,
    n12743, n12742, n12752, n12747, n12746, n12750, n12749, n12751, n12853,
    n12829, n12755, n12754, n12770, n12758, n12848, n12761, n12762, n12775,
    n12763, n12768, n12773, n13108, n12766, n12767, n12833, n12769, n12772,
    n12771, n12780, n13111, n12778, n12776, n12777, n12834, n12779, n12782,
    n12781, n12788, n12784, n12783, n12786, n12785, n12787, n12790, n12789,
    n12796, n12792, n12791, n12794, n12793, n12795, n12798, n12797, n12804,
    n12800, n12799, n12802, n12801, n12803, n12806, n12805, n12812, n12808,
    n12807, n12810, n12809, n12811, n12814, n12813, n12820, n12816, n12815,
    n12818, n12817, n12819, n12822, n12821, n12828, n12824, n12823, n12826,
    n12825, n12827, n12832, n12831, n12840, n12836, n12835, n12838, n12837,
    n12839, n12843, n12842, n12916, n12847, n12846, n12867, n12849, n12857,
    n12851, n12858, n12852, n12855, n12854, n12856, n12919, n12863, n12861,
    n12860, n12920, n12862, n12865, n12864, n12866, n12869, n12868, n12875,
    n12871, n12870, n12873, n12872, n12874, n12877, n12876, n12883, n12879,
    n12878, n12881, n12880, n12882, n12885, n12884, n12891, n12887, n12886,
    n12889, n12888, n12890, n12893, n12892, n12899, n12895, n12894, n12897,
    n12896, n12898, n12901, n12900, n12907, n12903, n12902, n12905, n12904,
    n12906, n12909, n12908, n12915, n12911, n12910, n12913, n12912, n12914,
    n12918, n12917, n12927, n12922, n12921, n12925, n12924, n12926, n13024,
    n13000, n12931, n12930, n12951, n13014, n12934, n12935, n12936, n12937,
    n12941, n12938, n12940, n12942, n13003, n12947, n12945, n12944, n13004,
    n12946, n12949, n12948, n12950, n12953, n12952, n12959, n12955, n12954,
    n12957, n12956, n12958, n12961, n12960, n12967, n12963, n12962, n12965,
    n12964, n12966, n12969, n12968, n12975, n12971, n12970, n12973, n12972,
    n12974, n12977, n12976, n12983, n12979, n12978, n12981, n12980, n12982,
    n12985, n12984, n12991, n12987, n12986, n12989, n12988, n12990, n12993,
    n12992, n12999, n12995, n12994, n12997, n12996, n12998, n13002, n13001,
    n13011, n13006, n13005, n13009, n13008, n13010, n13081, n13013, n13012,
    n13032, n13015, n13022, n13016, n13017, n13023, n13018, n13020, n13019,
    n13021, n13085, n13028, n13026, n13025, n13086, n13027, n13030, n13029,
    n13031, n13034, n13033, n13040, n13036, n13035, n13038, n13037, n13039,
    n13042, n13041, n13048, n13044, n13043, n13046, n13045, n13047, n13050,
    n13049, n13056, n13052, n13051, n13054, n13053, n13055, n13058, n13057,
    n13064, n13060, n13059, n13062, n13061, n13063, n13066, n13065, n13072,
    n13068, n13067, n13070, n13069, n13071, n13074, n13073, n13080, n13076,
    n13075, n13078, n13077, n13079, n13084, n13083, n13092, n13088, n13087,
    n13090, n13089, n13091, n13175, n13095, n13094, n13120, n13118, n13106,
    n13104, n13098, n13097, n13099, n13101, n13103, n13105, n13107, n13109,
    n13180, n13116, n13114, n13113, n13181, n13115, n13117, n13119, n13123,
    n13122, n13129, n13125, n13124, n13127, n13126, n13128, n13132, n13131,
    n13138, n13134, n13133, n13136, n13135, n13137, n13141, n13140, n13147,
    n13143, n13142, n13145, n13144, n13146, n13150, n13149, n13156, n13152,
    n13151, n13154, n13153, n13155, n13159, n13158, n13165, n13161, n13160,
    n13163, n13162, n13164, n13168, n13167, n13174, n13170, n13169, n13172,
    n13171, n13173, n13179, n13178, n13187, n13183, n13182, n13185, n13184,
    n13186, n13287, n13191, n13190, n13214, n13194, n13673, n13199, n13196,
    n13198, n13204, n13201, n13200, n13202, n13293, n13209, n13206, n13294,
    n13208, n13212, n13211, n13213, n13218, n13217, n13226, n13221, n13220,
    n13224, n13223, n13225, n13230, n13229, n13238, n13233, n13232, n13236,
    n13235, n13237, n13242, n13241, n13250, n13245, n13244, n13248, n13247,
    n13249, n13254, n13253, n13262, n13257, n13256, n13260, n13259, n13261,
    n13266, n13265, n13274, n13269, n13268, n13272, n13271, n13273, n13278,
    n13277, n13286, n13281, n13280, n13284, n13283, n13285, n13292, n13291,
    n13303, n13297, n13296, n13301, n13300, n13302, n13707, n13306, n13330,
    n13309, n13313, n13312, n13314, n13316, n13317, n13319, n13323, n13322,
    n13327, n13326, n13329, n13332, n13333, n13374, n13361, n13340, n13338,
    n13337, n13339, n13654, n13349, n13347, n13646, n13346, n13348, n13641,
    n13352, n13351, n13359, n13357, n13356, n13358, n13360, n13366, n13364,
    n13363, n13365, n13369, n13368, n13370, n13371, n13373, n13391, n13378,
    n13376, n13377, n13382, n13381, n13383, n13616, n13408, n13397, n13384,
    n13389, n13385, n13386, n13387, n13388, n13395, n13393, n13394, n13396,
    n13399, n13407, n13401, n13403, n13405, n13406, n13412, n13410, n13411,
    n13413, n13449, n13416, n13417, n13441, n13429, n13418, n13437, n13424,
    n13446, n13430, n13419, n13422, n13423, n13420, n13421, n13444, n13426,
    n13425, n13428, n13427, n13443, n13432, n13434, n13435, n13436, n13438,
    n13440, n13442, n13448, n13445, n13447, n13451, n13594, n13569, n13450,
    n13453, n13452, n13459, n13456, n13455, n13458, n13457, n13464, n13461,
    n13460, n13463, n13462, n13466, n13465, n13468, n13467, n13474, n13471,
    n13470, n13473, n13472, n13476, n13475, n13478, n13477, n13481, n13480,
    n13483, n13482, n13486, n13485, n13488, n13487, n13491, n13490, n13493,
    n13492, n13496, n13495, n13498, n13497, n13501, n13500, n13503, n13502,
    n13506, n13505, n13508, n13507, n13514, n13511, n13510, n13513, n13512,
    n13516, n13515, n13518, n13517, n13524, n13521, n13520, n13523, n13522,
    n13526, n13525, n13528, n13527, n13531, n13530, n13533, n13532, n13536,
    n13535, n13538, n13537, n13541, n13540, n13543, n13542, n13545, n13544,
    n13547, n13546, n13550, n13549, n13552, n13551, n13555, n13554, n13557,
    n13556, n13560, n13559, n13562, n13561, n13565, n13564, n13567, n13566,
    n13574, n13571, n13570, n13573, n13572, n13576, n13579, n13575, n13578,
    n13577, n13581, n13580, n13583, n13582, n13586, n13585, n13588, n13587,
    n13591, n13595, n13590, n13593, n13592, n13599, n13596, n13598, n13601,
    n13600, n13603, n13602, n13605, n13604, n13607, n13606, n13609, n13608,
    n13612, n13611, n13614, n13617, n13619, n13621, n13624, n13623, n13625,
    n13627, n13626, n13628, n13629, n13640, n13633, n13643, n13631, n13642,
    n13632, n13637, n13635, n13636, n13638, n13639, n13645, n13644, n13648,
    n13647, n13649, n13651, n13650, n13659, n13657, n13656, n13658, n13660,
    n13664, n13663, n13709, n13666, n13668, n13667, n13670, n13672, n13671,
    n13679, n13677, n13702, n13676, n13678, n13680, n13682, n13681, n13686,
    n13687, n13689, n13688, n13690, n13692, n13691, n13694, n13697, n13696,
    n13698, n13700, n13699, n13705, n13704, n13706, n13708, n13712, n13711,
    n13721, n13715, n13714, n13716, n13718, n13717, n13719, n13720, n13725,
    n13728, n13727, n13730, n13729, n13734, n13732, n13733, n13738, n13761,
    n13737, n13753, n13752, n13740, n13745, n13744, n13746, n13747, n13748,
    n13750, n13751, n13755, n13754, n13759, n13758, n13766, n13763, n13765,
    n11918, n7512, n13336;
  assign n10200 = ~n10229 & ~n9386;
  assign n9085 = ~n9454 | ~n13308;
  assign n8946 = ~n9210 | ~n11918;
  assign n7515 = n9302 & n7494;
  assign n7363 = n6997 | n7361;
  assign n7829 = n7600 ^ ~n7599;
  assign n6998 = ~n11826;
  assign n9029 = n9024 | n8178;
  assign n10830 = ~n10851;
  assign n9041 = ~n9464;
  assign n8985 = ~n7067 | ~n7027;
  assign n11821 = ~n11820;
  assign n7848 = ~n13693;
  assign n13693 = n8938;
  assign n9129 = ~n7595 & ~n9085;
  assign n10896 = ~n10907;
  assign n11536 = n8953 & n8952;
  assign n11772 = ~n11732;
  assign n10735 = ~n10790 & ~n10762;
  assign n11577 = n8943 | n8942;
  assign n13177 = ~n13669 | ~n13701;
  assign n9926 = ~n11123;
  assign n6993 = n7675 & n7068;
  assign n7541 = ~n9298 & ~n9201;
  assign n9201 = n9156 & n10793;
  assign n7006 = n7248 & n7253;
  assign n11826 = ~INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n7988 = ~n13310 | ~STATE2_REG_0__SCAN_IN;
  assign n7004 = ~n13310;
  assign n11865 = ~INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n7774 = n13328 | n7773;
  assign n11462 = INSTADDRPOINTER_REG_9__SCAN_IN ^ n9035;
  assign n11812 = ~INSTQUEUERD_ADDR_REG_3__SCAN_IN & ~INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n11519 = n8985 ^ ~n7066;
  assign n10089 = ~n9041;
  assign n10390 = ~n9331 | ~n9325;
  assign n11796 = n9331 & n13342;
  assign n7956 = ~n7771 | ~n7783;
  assign n6994 = ~n11092;
  assign n10809 = n10893 & STATE2_REG_2__SCAN_IN;
  assign n11401 = n11263 | n11262;
  assign n9115 = n9113 | n9112;
  assign n9113 = n9104 & n9103;
  assign n9126 = ~n7733 | ~n7988;
  assign n9286 = n9230;
  assign n8310 = ~n7531 | ~n7516;
  assign n9408 = ~n7880;
  assign n7253 = ~n13344;
  assign n7257 = n13336 & INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n7254 = n7245 & INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n11813 = ~INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n9955 = ~n7126 & ~n9954;
  assign n9948 = ~n7128 | ~n7127;
  assign n10146 = ~n7121 | ~n7205;
  assign n9987 = ~n7172 | ~n7170;
  assign n8843 = ~n9605;
  assign n9588 = ~n9605 & ~n7221;
  assign n8676 = ~n9683;
  assign n8478 = n8309 & n7054;
  assign n13375 = n13391 | STATE2_REG_1__SCAN_IN;
  assign n8309 = n10134 & n10135;
  assign n7098 = n7029 & n9041;
  assign n7131 = n7133 & n7165;
  assign n7201 = ~n10041 & ~n7202;
  assign n10240 = n10270 & n10259;
  assign n10270 = ~n9346 | ~n9345;
  assign n7204 = n7205 & n7206;
  assign n7162 = n10143 | n7163;
  assign n10056 = ~n9162 & ~n9161;
  assign n10641 = ~n8188 | ~n8187;
  assign n7208 = n10745 & n7209;
  assign n7074 = n11484 & n9004;
  assign n7211 = n8228 | n10149;
  assign n9794 = n9380 ^ ~n9504;
  assign n10174 = n9570 | n9569;
  assign n11420 = ~n9029 & ~n9028;
  assign n10004 = ~n9041;
  assign n9002 = n9001 ^ ~INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n9162 = ~n9041 & ~INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n13290 = ~n13192 | ~n13701;
  assign n8227 = n9032 | n8221;
  assign n10871 = n7875 | n7874;
  assign n9001 = ~n7089 | ~n8999;
  assign n11419 = n9035 & INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n13367 = ~n11845 & ~n11844;
  assign n10400 = ~n10390;
  assign n10206 = n9611 & n9610;
  assign n10848 = ~n7782 | ~n7781;
  assign n11732 = ~n9331 | ~n11818;
  assign n13192 = ~n12929 & ~n13693;
  assign n10837 = ~n9512 & ~n9215;
  assign n11537 = ~n8965 | ~n8964;
  assign n11884 = ~n12242 | ~n7772;
  assign n11131 = ~n11130 & ~n13310;
  assign n12242 = ~n7769 | ~n7783;
  assign n11880 = n7832 ^ ~n7831;
  assign n6995 = ~n7956;
  assign n9199 = ~n9185 & ~n9184;
  assign n11013 = ~n11017;
  assign n11581 = ~n11530;
  assign n7783 = ~n7768 | ~n7767;
  assign n13764 = n11263 & n9495;
  assign n7600 = ~n7594 | ~n7593;
  assign n13325 = ~n11806;
  assign n10841 = n10457 ^ ~n10456;
  assign n10855 = n7724 & n7562;
  assign n8939 = n7861 & n7860;
  assign n10862 = ~n10864 & ~n10863;
  assign n7068 = ~n7674 | ~n7673;
  assign n7123 = ~n7545 | ~n7224;
  assign n7560 = n7557 & n7556;
  assign n10864 = ~n7180 | ~n7178;
  assign n7550 = n7549 & n7548;
  assign n7180 = ~n9226 | ~n9225;
  assign n7673 = ~n7530 | ~n9320;
  assign n9088 = ~n9084 & ~n9083;
  assign n9320 = n7529 & n7528;
  assign n9298 = n9303 & n7534;
  assign n9435 = ~n9182 & ~n13400;
  assign n7207 = n7428 & n11908;
  assign n7428 = n7427 & n9849;
  assign n10481 = ~n11908 | ~n13310;
  assign n8940 = ~n13310 & ~n7512;
  assign n7492 = n7495 & n11938;
  assign n9304 = n7516;
  assign n9017 = n7668 | n7667;
  assign n9230 = n7512 & n9210;
  assign n9847 = ~n7488 | ~n7531;
  assign n11948 = ~n7531;
  assign n13328 = ~n7532;
  assign n7773 = n7488;
  assign n11908 = ~n7512;
  assign n9210 = n7426 | n7425;
  assign n7176 = ~n7177 & ~n7080;
  assign n7531 = ~n7358 | ~n7357;
  assign n7390 = n7373 & n7372;
  assign n7389 = n7388 & n7387;
  assign n7324 = n7323 & n7322;
  assign n7325 = n7309 & n7308;
  assign n7358 = n7342 & n7341;
  assign n7264 = n7263 & n7262;
  assign n7265 = n7244 & n7243;
  assign n8154 = n7014;
  assign n7652 = n7253 & n7254;
  assign n6996 = ~n11881;
  assign n8642 = n7257 & n11812;
  assign n7639 = n7254 & n11820;
  assign n7326 = n7254 & n7257;
  assign n7248 = n11809 & INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n6997 = ~n7404;
  assign n11820 = INSTQUEUERD_ADDR_REG_0__SCAN_IN & INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n7245 = ~INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n6999 = ~n11477 | ~n7002;
  assign n7151 = n6999 & n7000;
  assign n7000 = n7001 | n7131;
  assign n7001 = ~n7164;
  assign n7002 = n7130 & n7164;
  assign n7003 = ~n6993 | ~n13400;
  assign n11477 = ~n7073 | ~n9014;
  assign n7198 = ~n6993 | ~n13400;
  assign n7518 = ~n7176 | ~n7484;
  assign n7065 = n8993 ^ ~INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n8993 = ~n7075 | ~n8992;
  assign n7005 = ~n7432;
  assign n11809 = ~INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n7138 = ~n7151 | ~n7154;
  assign n7007 = ~n10434 & ~n9514;
  assign n7546 = ~n7504 | ~n7503;
  assign n7504 = n7490 & n7489;
  assign n9214 = ~n9220 | ~n9218;
  assign n7009 = ~n7374;
  assign n7010 = ~n7009;
  assign n7469 = ~n7374;
  assign n7374 = ~n7257 | ~n6998;
  assign n9218 = ~n9230;
  assign n7011 = ~n10869;
  assign n10908 = ~n10869;
  assign n10869 = n10893 & n9551;
  assign n10770 = n10893 & n9502;
  assign n7167 = ~n7087 | ~n7086;
  assign n7086 = ~n11420;
  assign n7087 = ~n11419 & ~n7088;
  assign n7595 = ~n7487 | ~n13311;
  assign n7487 = ~n9093;
  assign n7154 = n7204 & n7155;
  assign n7166 = ~n9025;
  assign n7070 = n7033 & n7208;
  assign n7113 = ~n7185 & ~n7115;
  assign n7185 = n7186 | n9745;
  assign n7533 = n9210 | n11918;
  assign n7217 = n7031 & n9626;
  assign n9786 = ~n9215;
  assign n9788 = ~n7144 | ~n11948;
  assign n7122 = ~n7967;
  assign n7147 = n7148 & n9998;
  assign n7106 = n7032 & n7013;
  assign n7105 = ~n9040 | ~n7013;
  assign n7164 = ~n7038 | ~n7168;
  assign n11806 = ~n9131 | ~n9130;
  assign n9130 = ~n9155 | ~n9129;
  assign n9131 = ~n9128 | ~n9127;
  assign n10360 = ~n10410 | ~n7114;
  assign n10790 = ~n7117 | ~n10862;
  assign n7117 = ~n7196 & ~n10787;
  assign n7195 = ~n9609 & ~n9608;
  assign n7171 = ~n9984;
  assign n7544 = n12765 | n9136;
  assign n7063 = ~n7326 | ~INSTQUEUE_REG_10__0__SCAN_IN;
  assign n7062 = ~n7652 | ~INSTQUEUE_REG_9__0__SCAN_IN;
  assign n7060 = n7336 & INSTQUEUE_REG_13__0__SCAN_IN;
  assign n9123 = ~n9065 | ~n9064;
  assign n9122 = ~n9123 & ~INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n7216 = n8350 & n8308;
  assign n8308 = ~n10121;
  assign n7967 = ~n7946 | ~n7945;
  assign n7149 = ~n7200;
  assign n7160 = n7055 & n8144;
  assign n7130 = ~n7132 & ~n7135;
  assign n7135 = ~n11462;
  assign n7132 = ~n11476;
  assign n7165 = ~n7167 & ~n7166;
  assign n7134 = ~n9023;
  assign n7076 = ~n6995 | ~n7911;
  assign n9081 = ~n7595;
  assign n7727 = ~n9135;
  assign n7855 = n7709 & n7708;
  assign n7222 = ~n9586;
  assign n7218 = ~n9482 & ~n9684;
  assign n7188 = ~n7189 | ~n10324;
  assign n7189 = ~n10341;
  assign n8188 = ~n7153 | ~n7987;
  assign n7209 = n8060 & n10718;
  assign n8060 = ~n10705;
  assign n7220 = ~n7223 & ~n7221;
  assign n7223 = ~n9395;
  assign n8600 = ~n8557 | ~PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n8944 = ~n8954;
  assign n7190 = ~n7193 | ~n7191;
  assign n7191 = ~n9608;
  assign n7193 = ~n9589 & ~n7194;
  assign n7140 = n7024 & n9055;
  assign n7104 = n7106 & n7020;
  assign n7103 = ~n7105;
  assign n7108 = ~n7110 | ~n7109;
  assign n7109 = ~n9359;
  assign n7110 = ~n7111;
  assign n9136 = ~n13402 | ~n13400;
  assign n9389 = ~n11772 & ~n11689;
  assign n13342 = n9156 & n13743;
  assign n7675 = n7674 | n7673;
  assign n8938 = n7847 ^ ~n7846;
  assign n12929 = n13683 | n12242;
  assign n7357 = n7356 & n7355;
  assign n9146 = STATE_REG_1__SCAN_IN ^ ~STATE_REG_2__SCAN_IN;
  assign n7877 = n10848 & n10822;
  assign n9626 = n8800 & n8799;
  assign n9647 = n8758 & n8757;
  assign n7181 = n7183 & n7182;
  assign n7182 = ~n10422;
  assign n10379 = ~n10410 | ~n7025;
  assign n10836 = n9234 ^ ~n9218;
  assign n7178 = ~n7179 | ~n9786;
  assign n10451 = ~n11806 & ~n13324;
  assign n11548 = n11530 & n11580;
  assign n7096 = n9987 | n7097;
  assign n7097 = ~n7098;
  assign n7094 = n7095 & n9465;
  assign n7095 = ~n7098 | ~n7142;
  assign n7093 = ~n9987 | ~n7140;
  assign n9957 = n9987 & n9055;
  assign n7078 = ~n7138 | ~n7139;
  assign n7139 = ~n7101 | ~n7105;
  assign n10116 = ~n7081 | ~n10370;
  assign n11016 = ~n11017 | ~n13328;
  assign n11092 = ~n9456 | ~n11405;
  assign n9456 = ~n9453 | ~n13390;
  assign n9452 = n9451 & n9450;
  assign n9462 = n7099 & n7029;
  assign n11739 = n9331 & n9300;
  assign n9377 = ~n7195 | ~n9376;
  assign n7119 = ~n9393 & ~n7120;
  assign n11803 = n9331 & n9209;
  assign n13661 = ~n13662;
  assign n9431 = n8889 | n8888;
  assign n9006 = n7072 ^ ~n7973;
  assign n8973 = ~n11555 | ~n11535;
  assign n8958 = n7592 & n7591;
  assign n7720 = ~n7672 | ~n7671;
  assign n7672 = n7670 & n7669;
  assign n7603 = ~n7254 | ~n11865;
  assign n7236 = ~n7248;
  assign n7258 = ~n8642 | ~INSTQUEUE_REG_2__6__SCAN_IN;
  assign n7289 = ~n8642 | ~INSTQUEUE_REG_2__7__SCAN_IN;
  assign n9060 = INSTQUEUERD_ADDR_REG_0__SCAN_IN & n9076;
  assign n7733 = ~n11938 | ~STATE2_REG_0__SCAN_IN;
  assign n7129 = ~n7550 | ~n7551;
  assign n8888 = n8878 | n8877;
  assign n7153 = ~n9029;
  assign n7143 = ~n7911 | ~n7958;
  assign n7194 = ~n9567;
  assign n7146 = n7201 & n10030;
  assign n9161 = ~n10089 & ~n9042;
  assign n7169 = ~n11452;
  assign n7168 = ~n7167;
  assign n8989 = n7815 | n7814;
  assign n7059 = ~n7061 & ~n7060;
  assign n7061 = ~n7063 | ~n7062;
  assign n7424 = ~n7416 & ~n7415;
  assign n7373 = ~n7365 & ~n7364;
  assign n7341 = ~n7340 & ~n7339;
  assign n7352 = ~n8642 | ~INSTQUEUE_REG_2__5__SCAN_IN;
  assign n9155 = ~n9125 | ~n9124;
  assign n9125 = n9122 | INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign n10614 = ~PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n10782 = ~PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n7875 = ~n7835 | ~n7834;
  assign n7116 = ~n10358;
  assign n7183 = n7184 & n10665;
  assign n7184 = ~n10645;
  assign n10685 = n8102 & n8101;
  assign n9395 = ~n8935 & ~n8934;
  assign n8839 = ~n8760 & ~n8759;
  assign n8756 = ~n8711 & ~n9688;
  assign n8711 = ~n8672 | ~PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n8672 = ~n8600 & ~n9728;
  assign n9703 = n8603 & n8602;
  assign n8557 = ~n8515 & ~n9778;
  assign n7214 = n7216 & n7215;
  assign n10079 = n8436 & n8435;
  assign n10104 = n8349 & n8348;
  assign n10121 = n8307 & n8306;
  assign n8306 = n8305 | n8304;
  assign n8268 = ~n8229 & ~n10614;
  assign n7210 = ~n10149;
  assign n8266 = n8305 | n8265;
  assign n8179 = ~PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n8180 = ~n8103 | ~PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n8103 = ~n8062 & ~n8061;
  assign n8061 = ~PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n10705 = n8059 & n8058;
  assign n8062 = ~n8022 | ~PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n10718 = ~n8021 | ~n8020;
  assign n8020 = ~n8019 | ~n7053;
  assign n8022 = ~n7982 & ~n10732;
  assign n7975 = ~n7959 & ~n10782;
  assign n8955 = n7634 & n7633;
  assign n9303 = ~n9788 & ~n10481;
  assign n9015 = ~n7710 & ~n13400;
  assign n9611 = ~n7195;
  assign n7111 = ~n7112 | ~n9686;
  assign n7186 = n7188 | n7187;
  assign n7187 = ~n9767;
  assign n7085 = ~n10101;
  assign n7107 = n8144 & n9109;
  assign n7081 = ~n9035;
  assign n7159 = n7160 & n9109;
  assign n11431 = ~n9035 & ~INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n8954 = n7706 & n7705;
  assign n10443 = n9194 & n13320;
  assign n11819 = ~n9203 & ~n9202;
  assign n7767 = n7766 & n7765;
  assign n10456 = n7731 & n7730;
  assign n7730 = n7729 & n7728;
  assign n7859 = ~n7855;
  assign n12765 = INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n7319 = ~n7639 | ~INSTQUEUE_REG_11__2__SCAN_IN;
  assign n7488 = n7265 & n7264;
  assign n7532 = n7295 | n7294;
  assign n13315 = n9134 & n9133;
  assign n11873 = ~INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n13100 = ~STATEBS16_REG_SCAN_IN;
  assign n13102 = ~n8937;
  assign n9446 = n11983 & STATEBS16_REG_SCAN_IN;
  assign n7219 = ~n9541;
  assign n8391 = ~PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n8351 = ~n8343 & ~n10576;
  assign n8343 = ~n8268 | ~PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n9527 = EBX_REG_31__SCAN_IN & n10809;
  assign n7982 = ~n7975 | ~PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n10822 = ~n7828 | ~n7827;
  assign n7950 = ~n7824 & ~n11529;
  assign n10795 = ~n10770;
  assign n8887 = n9949 | n8384;
  assign n8842 = ~n9607;
  assign n9482 = n8717 & n8716;
  assign n8716 = n8715 & n8714;
  assign n9723 = n8559 & n8558;
  assign n7212 = ~n7213;
  assign n10647 = ~n10666 | ~n7183;
  assign n11253 = ~n9147 & ~n13742;
  assign n9147 = ~n11259 & ~n9145;
  assign n9145 = ~n13325 & ~n9144;
  assign n13741 = n8940;
  assign n11259 = ~n11263 & ~n9454;
  assign n9550 = PHYADDRPOINTER_REG_31__SCAN_IN ^ ~n9472;
  assign n9566 = n9588 ^ ~n9395;
  assign n11488 = n7030 | n10746;
  assign n11570 = ~n11548;
  assign n10921 = n7870 & n7869;
  assign n10167 = ~n10178 & ~n9390;
  assign n9391 = n10167 & INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n9568 = n7195 & n7192;
  assign n7192 = ~n9589;
  assign n7172 = ~n7137 | ~n7138;
  assign n7102 = ~n7103 | ~n7020;
  assign n10239 = ~n10269 & ~n9339;
  assign n7200 = ~n9164 | ~n7037;
  assign n10074 = ~n7084 | ~n7082;
  assign n7082 = n7083 & n10071;
  assign n7084 = ~n10068 | ~n7085;
  assign n7083 = ~n7085 | ~n10069;
  assign n10091 = ~n10074;
  assign n10115 = ~n7081 | ~n10397;
  assign n10144 = ~n7151 & ~n11421;
  assign n13703 = n6993;
  assign n11867 = n9201;
  assign n13355 = ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n13701 = ~n8939;
  assign n12598 = ~n13665 & ~n12513;
  assign n13203 = ~n12246 & ~n12170;
  assign n12845 = ~n12759;
  assign n12246 = ~n11901;
  assign n12841 = ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n13354 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n11938 = ~n7496;
  assign n11967 = ~n11901 | ~STATE2_REG_3__SCAN_IN;
  assign n13652 = n11806 & STATE2_REG_3__SCAN_IN;
  assign n9135 = n13655 & STATE2_REG_2__SCAN_IN;
  assign n13402 = ~STATE2_REG_1__SCAN_IN & ~STATE2_REG_3__SCAN_IN;
  assign n13655 = ~STATE2_REG_1__SCAN_IN;
  assign n11983 = ~STATE2_REG_2__SCAN_IN;
  assign n9627 = n8676 & n7031;
  assign n9988 = n9480 ^ ~n9647;
  assign n10325 = ~n10360 & ~n10341;
  assign n10377 = n10410 & n10408;
  assign n10788 = ~n10862 | ~n7197;
  assign n11017 = n9793 & n13390;
  assign n11020 = n11017 & n9849;
  assign n9857 = ~n9566;
  assign n9864 = ~n9948;
  assign n11097 = ~n6994 & ~n11049;
  assign n11121 = ~n11097;
  assign n11123 = ~n11092 | ~n11049;
  assign n11252 = ~n13735;
  assign n11405 = n11263 | n9455;
  assign n7126 = ~n9948 & ~n11881;
  assign n11530 = ~n11567 | ~n9137;
  assign n10158 = n9469 ^ ~INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n9468 = ~n7096 | ~n7094;
  assign n7092 = ~n9945;
  assign n7079 = ~n7077;
  assign n7077 = n7078;
  assign n10102 = ~n10068 & ~n10069;
  assign n13662 = ~n10462 & ~n10455;
  assign n13121 = ~n13215;
  assign n13130 = ~n13227;
  assign n13139 = ~n13239;
  assign n13148 = ~n13251;
  assign n13166 = ~n13275;
  assign n13176 = ~n13288;
  assign n13390 = ~n13404;
  assign n7118 = ~n9381 | ~n11739;
  assign n7012 = n7017 & n7054;
  assign n8906 = ~n8130;
  assign n10704 = ~n7030 | ~n10718;
  assign n13308 = n7531;
  assign n7013 = n9041 | n10280;
  assign n7014 = n6998 & n11865;
  assign n10134 = ~n7152 | ~n7045;
  assign n9764 = ~n8478;
  assign n8453 = ~n7603;
  assign n7015 = n10369 | n11567;
  assign n9683 = ~n8309 | ~n7012;
  assign n7016 = n7041 & n9723;
  assign n9493 = n9543 ^ ~n7056;
  assign n7017 = n7016 & n9703;
  assign n7018 = n7162 & n7046;
  assign n10912 = ~n9214;
  assign n7404 = n11812 & n11820;
  assign n10821 = n7876 & n10871;
  assign n8562 = ~n7336;
  assign n7019 = n9705 | n7108;
  assign n7020 = n9049 & n9048;
  assign n7021 = n10725 | n10724;
  assign n7022 = ~n10766 & ~n10685;
  assign n7023 = ~n13329 & ~n13328;
  assign n9480 = n8676 & n7218;
  assign n7024 = n9972 & n9959;
  assign n7025 = n10376 & n10408;
  assign n11454 = ~n9026 | ~n9025;
  assign n7026 = n9041 | n9355;
  assign n10029 = ~n7150 | ~n7200;
  assign n7027 = n8983 | n9529;
  assign n7028 = n10089 | n9052;
  assign n10744 = ~n10766 & ~n7125;
  assign n9766 = ~n10360 & ~n7188;
  assign n7029 = n9357 & n9356;
  assign n10078 = n8309 & n7214;
  assign n7030 = n10744 & n10745;
  assign n7031 = n7218 & n9647;
  assign n7032 = n10116 & n10071;
  assign n7033 = n7124 & n7211;
  assign n7034 = n7022 & n7070;
  assign n7035 = n9394 & n7119;
  assign n7206 = ~n9036;
  assign n7114 = ~n7115;
  assign n7115 = ~n7025 | ~n7116;
  assign n7036 = ~n9464 | ~n10193;
  assign n7037 = ~n7203 | ~n9163;
  assign n7141 = ~n7142;
  assign n7142 = ~n7026 | ~n9055;
  assign n7155 = ~n9040;
  assign n7038 = n11431 | n7169;
  assign n7039 = ~n9141 & ~n9140;
  assign n7202 = ~n10056;
  assign n7040 = n7022 & n7069;
  assign n7041 = ~n9744 & ~n9765;
  assign n7042 = ~n7143 & ~n7122;
  assign n7043 = n9705 | n7111;
  assign n7044 = n10128 & n10127;
  assign n7045 = n8227 | n7210;
  assign n7046 = n7157 & n10115;
  assign n7221 = ~n7222 | ~n8842;
  assign n7047 = n8478 & n7041;
  assign n7048 = n7220 & n7219;
  assign n7049 = n7018 | n9036;
  assign n7050 = n10360 | n7186;
  assign n7051 = n7140 & n7036;
  assign n7052 = n8478 & n7016;
  assign n7173 = ~n7174;
  assign n7174 = n7175 & n7028;
  assign n8587 = n8586;
  assign n9438 = ~n7864;
  assign n8880 = ~n9438;
  assign n8854 = ~n7603;
  assign n10674 = ~n7021 & ~n10694;
  assign n10644 = ~n10666 | ~n10665;
  assign n7053 = n8018 | n8017;
  assign n7957 = n7817 & n7816;
  assign n7054 = n7214 & n10079;
  assign n7055 = n8220 | n9015;
  assign n13683 = n11880;
  assign n9307 = ~n11928 | ~n11918;
  assign n7144 = ~n9307;
  assign n11928 = ~n9210;
  assign n7837 = ~STATE2_REG_2__SCAN_IN & ~STATEBS16_REG_SCAN_IN;
  assign n8384 = ~n7837;
  assign n13400 = ~STATE2_REG_0__SCAN_IN;
  assign n8221 = ~n7773 | ~STATE2_REG_2__SCAN_IN;
  assign n7056 = ~n9448 | ~n9447;
  assign n7057 = n7180 & n7179;
  assign n7161 = ~INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n7066 = ~INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n13597 = ~n13757 | ~n13449;
  assign n13757 = ~STATE_REG_0__SCAN_IN & ~n13433;
  assign n7075 = ~n7058 | ~n9109;
  assign n7965 = ~n7058 | ~n7987;
  assign n7058 = n7076 ^ ~n7958;
  assign n7080 = ~n7059 | ~n7461;
  assign n11496 = ~n11508 | ~n7064;
  assign n7064 = ~n7065;
  assign n11719 = n11508 ^ ~n7065;
  assign n7067 = ~n8984;
  assign n7936 = n11812 & n11865;
  assign n7552 = ~n7123 | ~n7068;
  assign n10879 = n7601 ^ ~n7068;
  assign n7069 = n7208 & n7124;
  assign n10120 = ~n8309;
  assign n9543 = ~n8843 | ~n7048;
  assign n7529 = ~n10793 | ~n7071;
  assign n7071 = ~n7429 | ~n7428;
  assign n9024 = ~n7072 | ~n8144;
  assign n9464 = ~n7072 | ~n9016;
  assign n7158 = ~n7072 | ~n7159;
  assign n9032 = ~n7072 | ~n7160;
  assign n9035 = n7072 & n7107;
  assign n7072 = ~n6995 | ~n7042;
  assign n7073 = ~n9005 | ~n7074;
  assign n9004 = ~n9002 | ~n9003;
  assign n11484 = n9013 ^ ~n11678;
  assign n9005 = ~n11496 | ~n9000;
  assign n7145 = ~n7078 | ~n7146;
  assign n10058 = ~n7078 | ~n10056;
  assign n7150 = ~n7078 | ~n7201;
  assign n10057 = ~n7079 | ~n7202;
  assign n7375 = ~n8642 | ~INSTQUEUE_REG_2__4__SCAN_IN;
  assign n7088 = ~n11433;
  assign n7136 = ~n11477 | ~n11476;
  assign n11499 = ~n9002;
  assign n7089 = ~n8994 | ~n9109;
  assign U2957 = ~n7091 | ~n7090;
  assign n7090 = ~n10173 | ~n11578;
  assign n10173 = n9059 ^ ~n9058;
  assign n7091 = n7225 & n7039;
  assign n9466 = ~n9987 | ~n7051;
  assign n9947 = n7093 & n7092;
  assign n7099 = ~n9987 | ~n7141;
  assign n13343 = ~n7257;
  assign n7148 = ~n7149 | ~n10030;
  assign n9479 = n9173 ^ ~n9172;
  assign n11663 = ~n10400 & ~n11796;
  assign n9120 = ~n9119 & ~n9118;
  assign n10203 = ~n10230 & ~n9385;
  assign n9119 = ~n9115 | ~n9114;
  assign n9128 = ~n9121 & ~n9120;
  assign n7170 = ~n7173 & ~n7171;
  assign n7175 = ~n9045 | ~n7020;
  assign n10745 = ~n7981 | ~n7980;
  assign n11421 = ~n9030 & ~INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n9943 = ~n9942 & ~n9941;
  assign n9173 = ~n9171 & ~n9170;
  assign n9012 = n9006 | n9085;
  assign n9013 = ~n9012 | ~n9011;
  assign n7100 = ~n7049 | ~n7104;
  assign n7101 = ~n7049 | ~n7106;
  assign n7137 = ~n7100 | ~n7102;
  assign n9239 = ~n9215 | ~INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n9232 = ~n9215 | ~INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n9235 = ~n9215 | ~INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n9242 = ~n9215 | ~INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n9245 = ~n9215 | ~INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n9251 = ~n9215 | ~INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n9330 = n9786 & n9210;
  assign n9284 = ~n9215 | ~INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n9292 = ~n9507 | ~INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n9295 = ~n9507 | ~INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n9211 = ~n9507 | ~INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n9372 = ~n9215 | ~INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n13760 = ~n9215 | ~n10481;
  assign n9360 = ~n9215 | ~INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n9369 = ~n9215 | ~INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n9363 = ~n9215 | ~INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n9366 = ~n9215 | ~INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n9378 = ~n9215 | ~INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n11775 = n7057 ^ ~n9215;
  assign n9685 = ~n9705 & ~n9704;
  assign n7112 = ~n9704;
  assign n9725 = n10410 & n7113;
  assign n7196 = ~n9238 | ~n10836;
  assign U2988 = ~n7035 | ~n7118;
  assign n7120 = ~n9938;
  assign U2971 = ~n7015 | ~n7044;
  assign n7121 = ~n10144;
  assign n7601 = ~n7129 | ~n7123;
  assign n10684 = ~n10744 | ~n7208;
  assign n7124 = ~n7125;
  assign n7125 = ~n10765 | ~n10767;
  assign n7127 = ~n9588;
  assign n7128 = ~n9587 | ~n9586;
  assign n7771 = n7830 & n7829;
  assign n7769 = ~n7771;
  assign n7561 = ~n7552 | ~n7129;
  assign n11483 = n9005 & n9004;
  assign n7133 = ~n11462 | ~n7134;
  assign n9026 = ~n11461 | ~n11462;
  assign n11461 = ~n7136 | ~n9023;
  assign n8994 = n7966 ^ ~n7967;
  assign n10213 = n9957 ^ ~n9974;
  assign n7966 = n7956 | n7143;
  assign n9168 = ~n7145 | ~n7147;
  assign n7156 = ~n7151 | ~n7204;
  assign n7152 = ~n7034 | ~n8189;
  assign n10068 = ~n7156 | ~n7049;
  assign n9034 = ~n7157;
  assign n7157 = ~n7158 | ~n7161;
  assign n7205 = ~n10143;
  assign n7163 = ~n11421;
  assign n11418 = ~n11454 | ~n11452;
  assign n9985 = n7172 & n7174;
  assign n7246 = ~n8453 | ~INSTQUEUE_REG_8__6__SCAN_IN;
  assign n13310 = ~n7518;
  assign n7177 = ~n7483 | ~n7468;
  assign n9220 = ~n7004 | ~n11928;
  assign n7179 = ~n9227 | ~n10911;
  assign n10410 = n10666 & n7181;
  assign n9570 = ~n9609 & ~n7190;
  assign n9503 = ~n9570;
  assign n7197 = ~n7196;
  assign n10803 = ~n10862 | ~n10836;
  assign n7716 = ~n7198 | ~n7855;
  assign n7861 = ~n7003 | ~n7857;
  assign n7511 = ~n7199;
  assign n9191 = ~n7199 & ~n8946;
  assign n7501 = ~n7199 & ~n7500;
  assign n9315 = ~n7199 | ~n9286;
  assign n7199 = ~n7497 | ~n9187;
  assign n9997 = ~n10058 | ~n9163;
  assign n7203 = ~n10042;
  assign n7486 = ~n7207 | ~n7429;
  assign n7213 = ~n7040 | ~n8189;
  assign n10147 = ~n7213 | ~n8227;
  assign n10148 = ~n7212 | ~n8228;
  assign n10092 = ~n8309 | ~n7216;
  assign n7215 = ~n10093;
  assign n10103 = ~n8309 | ~n8308;
  assign n9743 = ~n8478 | ~n8477;
  assign n9605 = ~n8676 | ~n7217;
  assign n9481 = ~n8676 | ~n8675;
  assign n9540 = ~n8843 | ~n7220;
  assign n9587 = ~n8843 | ~n8842;
  assign n10927 = n9511 ^ ~n9510;
  assign n9511 = ~n9506 | ~n9505;
  assign n9093 = ~n7518 | ~STATE2_REG_0__SCAN_IN;
  assign n10018 = n9168;
  assign n7847 = n7845 ^ ~n7844;
  assign n7845 = ~n7717 | ~n8142;
  assign n9848 = ~n9935;
  assign n9747 = ~n9725;
  assign n9705 = ~n9725 | ~n9291;
  assign n7495 = n7531 | n7488;
  assign n10457 = n7724;
  assign n8305 = n8221 | n8143;
  assign n8019 = ~n8305;
  assign n7224 = n7547 | INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n7225 = n9566 | n11881;
  assign n11881 = ~n13414 | ~n8937;
  assign n7226 = n11846 & n13655;
  assign n7227 = ~n13204 | ~n8937;
  assign n7228 = ~n12757 & ~n13102;
  assign n9728 = ~PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n7229 = ~n8057 | ~n8056;
  assign n7432 = ~n7404;
  assign n7911 = ~n7957;
  assign n8899 = n9401;
  assign n11828 = n9174;
  assign n9105 = n10481 & n9074;
  assign n7530 = ~n7527 & ~n7526;
  assign n7232 = ~n7612 | ~INSTQUEUE_REG_4__6__SCAN_IN;
  assign n9007 = n7944 | n7943;
  assign n8981 = n7764 | n7763;
  assign n7635 = n7733 | n8955;
  assign n9107 = INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n8801 = n8792 | n8791;
  assign n11829 = n9303;
  assign n8142 = ~n9015;
  assign n7558 = ~n7560;
  assign n7844 = ~n7720;
  assign n8877 = n8802 | n8801;
  assign n8666 = ~n9435;
  assign n9182 = n8310 | n8311;
  assign n9451 = n10439 | READY_N;
  assign n8350 = ~n10104;
  assign n8996 = n7908 | n7907;
  assign n9225 = ~n10911;
  assign n13345 = ~n9182;
  assign n7457 = ~n7456 & ~n7455;
  assign n7387 = ~n7386 & ~n7385;
  assign n7537 = ~n8946 & ~n7536;
  assign n8675 = ~n9684;
  assign n8477 = ~n9765;
  assign n9688 = ~PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n7987 = ~n8221;
  assign n9109 = ~n9085;
  assign n9778 = ~PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n10576 = ~PHYADDRPOINTER_REG_15__SCAN_IN;
  assign n9514 = n13310 | n9513;
  assign n9291 = ~n9726;
  assign n9471 = ~n9397 & ~n9396;
  assign n8760 = ~n8756 | ~PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n8515 = ~n8437 | ~PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n8229 = ~n8222 | ~PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n10732 = ~PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n12757 = n10841;
  assign n12759 = n13683 & n7848;
  assign n13110 = ~n12246 & ~n12774;
  assign n13321 = ~n9155 & ~n9154;
  assign n8437 = ~n8392 & ~n8391;
  assign n9501 = n9500 & n11559;
  assign n10907 = ~n10893 | ~STATE2_REG_3__SCAN_IN;
  assign n10793 = ~n10481;
  assign n8222 = ~n8180 & ~n8179;
  assign n11576 = ~n11559;
  assign n13634 = n11821;
  assign n11898 = n11980 & n8939;
  assign n11980 = ~n12673 & ~n11884;
  assign n12249 = ~n12167 & ~n8939;
  assign n12329 = ~n13665 & ~n7848;
  assign n13665 = n12243 | n13683;
  assign n12673 = ~n13683 | ~n13693;
  assign n12933 = ~n12845 & ~n12844;
  assign n13669 = ~n12929 & ~n7848;
  assign n9494 = n13321 & n9157;
  assign n10484 = n10470 & n10469;
  assign n9502 = n9550 & STATE2_REG_1__SCAN_IN;
  assign n8392 = ~n8351 | ~PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n10914 = ~n10837;
  assign n10893 = ~n13764 | ~n9501;
  assign n11046 = ~n10587;
  assign n11186 = ~n13304 & ~STATE2_REG_0__SCAN_IN;
  assign n11523 = ~n10996;
  assign n11529 = ~PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n11559 = n9136 | STATE2_REG_2__SCAN_IN;
  assign n11792 = ~n11739;
  assign n11773 = ~n11795 & ~n11794;
  assign n11808 = n13652 | n11807;
  assign n12052 = ~n11898;
  assign n12150 = ~n11980 | ~n13701;
  assign n12235 = n12167 | n13701;
  assign n12324 = ~n12249;
  assign n12399 = ~n12329 | ~n8939;
  assign n12483 = ~n12329 | ~n13701;
  assign n12550 = ~n12575;
  assign n12575 = ~n13665 & ~n12410;
  assign n12659 = ~n12598;
  assign n12748 = n12673 | n12760;
  assign n12830 = n12673 | n12844;
  assign n12923 = n12845 | n12760;
  assign n13007 = ~n12933;
  assign n13082 = ~n13669 | ~n8939;
  assign n13093 = ~n13188;
  assign n13157 = ~n13263;
  assign n13227 = ~n11967 & ~n11918;
  assign n13263 = ~n11967 & ~n11948;
  assign n13299 = ~n13192 | ~n8939;
  assign n13742 = n9146 | STATE_REG_0__SCAN_IN;
  assign n9143 = ~n9142 & ~n13404;
  assign n13433 = ~STATE_REG_1__SCAN_IN;
  assign n13404 = ~n9135 | ~STATE2_REG_0__SCAN_IN;
  assign n11010 = ~n11020;
  assign n11001 = ~n11016;
  assign n11256 = ~n11253 & ~n11252;
  assign n11503 = ~n11091;
  assign n11578 = ~n11567;
  assign n11784 = ~n11803;
  assign n11901 = n11808 & n13400;
  assign n12154 = ~n12235;
  assign n12662 = ~n12607 | ~n12939;
  assign n10477 = n13439 | n10465;
  assign n11263 = ~n11806 | ~n9143;
  assign n11567 = n13331 | n13404;
  assign n11245 = n11256;
  assign n13710 = ~n11901 & ~n11879;
  assign n13414 = ~n8936 & ~n13655;
  assign n13415 = ~n13756 | ~n10477;
  assign n8586 = n7257 & n7248;
  assign n7231 = ~n8586 | ~INSTQUEUE_REG_6__6__SCAN_IN;
  assign n13344 = ~n11813 | ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n8029 = n7253 & n11812;
  assign n7230 = ~n8029 | ~INSTQUEUE_REG_1__6__SCAN_IN;
  assign n7235 = ~n7231 | ~n7230;
  assign n7233 = ~n7798 | ~INSTQUEUE_REG_14__6__SCAN_IN;
  assign n7612 = n7248 & n11865;
  assign n7234 = ~n7233 | ~n7232;
  assign n7244 = ~n7235 & ~n7234;
  assign n7472 = ~n7236 & ~n11821;
  assign n7238 = ~n7472 | ~INSTQUEUE_REG_7__6__SCAN_IN;
  assign n7237 = ~n7936 | ~INSTQUEUE_REG_0__6__SCAN_IN;
  assign n7242 = ~n7238 | ~n7237;
  assign n7240 = ~n7404 | ~INSTQUEUE_REG_3__6__SCAN_IN;
  assign n8279 = n6998 & n11820;
  assign n7239 = ~n8279 | ~INSTQUEUE_REG_15__6__SCAN_IN;
  assign n7241 = ~n7240 | ~n7239;
  assign n7243 = ~n7242 & ~n7241;
  assign n7247 = ~n7326 | ~INSTQUEUE_REG_10__6__SCAN_IN;
  assign n7252 = ~n7247 | ~n7246;
  assign n7250 = ~n7006 | ~INSTQUEUE_REG_5__6__SCAN_IN;
  assign n7249 = ~n7014 | ~INSTQUEUE_REG_12__6__SCAN_IN;
  assign n7251 = ~n7250 | ~n7249;
  assign n7263 = ~n7252 & ~n7251;
  assign n7256 = ~n7652 | ~INSTQUEUE_REG_9__6__SCAN_IN;
  assign n7255 = ~n7639 | ~INSTQUEUE_REG_11__6__SCAN_IN;
  assign n7261 = ~n7256 | ~n7255;
  assign n7336 = ~n13344 & ~n11826;
  assign n7259 = ~n7336 | ~INSTQUEUE_REG_13__6__SCAN_IN;
  assign n7260 = ~n7259 | ~n7258;
  assign n7262 = ~n7261 & ~n7260;
  assign n7267 = ~n7326 | ~INSTQUEUE_REG_10__7__SCAN_IN;
  assign n7266 = ~n7652 | ~INSTQUEUE_REG_9__7__SCAN_IN;
  assign n7271 = ~n7267 | ~n7266;
  assign n7269 = ~n7639 | ~INSTQUEUE_REG_11__7__SCAN_IN;
  assign n7268 = ~n7404 | ~INSTQUEUE_REG_3__7__SCAN_IN;
  assign n7270 = ~n7269 | ~n7268;
  assign n7279 = ~n7271 & ~n7270;
  assign n7273 = ~n8586 | ~INSTQUEUE_REG_6__7__SCAN_IN;
  assign n7272 = ~n7612 | ~INSTQUEUE_REG_4__7__SCAN_IN;
  assign n7277 = ~n7273 | ~n7272;
  assign n7275 = ~n7336 | ~INSTQUEUE_REG_13__7__SCAN_IN;
  assign n7274 = ~n7014 | ~INSTQUEUE_REG_12__7__SCAN_IN;
  assign n7276 = ~n7275 | ~n7274;
  assign n7278 = ~n7277 & ~n7276;
  assign n7295 = ~n7279 | ~n7278;
  assign n7281 = ~n7798 | ~INSTQUEUE_REG_14__7__SCAN_IN;
  assign n7280 = ~n8453 | ~INSTQUEUE_REG_8__7__SCAN_IN;
  assign n7285 = ~n7281 | ~n7280;
  assign n7283 = ~n7472 | ~INSTQUEUE_REG_7__7__SCAN_IN;
  assign n7282 = ~n8279 | ~INSTQUEUE_REG_15__7__SCAN_IN;
  assign n7284 = ~n7283 | ~n7282;
  assign n7293 = ~n7285 & ~n7284;
  assign n7287 = ~n7006 | ~INSTQUEUE_REG_5__7__SCAN_IN;
  assign n7286 = ~n8029 | ~INSTQUEUE_REG_1__7__SCAN_IN;
  assign n7291 = ~n7287 | ~n7286;
  assign n7288 = ~n7936 | ~INSTQUEUE_REG_0__7__SCAN_IN;
  assign n7290 = ~n7289 | ~n7288;
  assign n7292 = ~n7291 & ~n7290;
  assign n7294 = ~n7293 | ~n7292;
  assign n7516 = n7488 & n7532;
  assign n7297 = ~n7469 | ~INSTQUEUE_REG_14__2__SCAN_IN;
  assign n7296 = ~n8642 | ~INSTQUEUE_REG_2__2__SCAN_IN;
  assign n7301 = ~n7297 | ~n7296;
  assign n7299 = ~n7472 | ~INSTQUEUE_REG_7__2__SCAN_IN;
  assign n7298 = ~n7014 | ~INSTQUEUE_REG_12__2__SCAN_IN;
  assign n7300 = ~n7299 | ~n7298;
  assign n7309 = ~n7301 & ~n7300;
  assign n7303 = ~n7612 | ~INSTQUEUE_REG_4__2__SCAN_IN;
  assign n7302 = ~n8029 | ~INSTQUEUE_REG_1__2__SCAN_IN;
  assign n7307 = ~n7303 | ~n7302;
  assign n7305 = ~n8453 | ~INSTQUEUE_REG_8__2__SCAN_IN;
  assign n7304 = ~n7936 | ~INSTQUEUE_REG_0__2__SCAN_IN;
  assign n7306 = ~n7305 | ~n7304;
  assign n7308 = ~n7307 & ~n7306;
  assign n7311 = ~n7326 | ~INSTQUEUE_REG_10__2__SCAN_IN;
  assign n7310 = ~n7336 | ~INSTQUEUE_REG_13__2__SCAN_IN;
  assign n7315 = ~n7311 | ~n7310;
  assign n7313 = ~n7652 | ~INSTQUEUE_REG_9__2__SCAN_IN;
  assign n7312 = ~n7404 | ~INSTQUEUE_REG_3__2__SCAN_IN;
  assign n7314 = ~n7313 | ~n7312;
  assign n7323 = ~n7315 & ~n7314;
  assign n7317 = ~n8586 | ~INSTQUEUE_REG_6__2__SCAN_IN;
  assign n7316 = ~n7006 | ~INSTQUEUE_REG_5__2__SCAN_IN;
  assign n7321 = ~n7317 | ~n7316;
  assign n7318 = ~n8279 | ~INSTQUEUE_REG_15__2__SCAN_IN;
  assign n7320 = ~n7319 | ~n7318;
  assign n7322 = ~n7321 & ~n7320;
  assign n7391 = ~n7516 & ~n11918;
  assign n7328 = ~n7326 | ~INSTQUEUE_REG_10__5__SCAN_IN;
  assign n7327 = ~n7404 | ~INSTQUEUE_REG_3__5__SCAN_IN;
  assign n7333 = ~n7328 | ~n7327;
  assign n7331 = ~n7798 | ~INSTQUEUE_REG_14__5__SCAN_IN;
  assign n7330 = ~n7472 | ~INSTQUEUE_REG_7__5__SCAN_IN;
  assign n7332 = ~n7331 | ~n7330;
  assign n7342 = ~n7333 & ~n7332;
  assign n7335 = ~n7652 | ~INSTQUEUE_REG_9__5__SCAN_IN;
  assign n7334 = ~n7612 | ~INSTQUEUE_REG_4__5__SCAN_IN;
  assign n7340 = ~n7335 | ~n7334;
  assign n7338 = ~n7336 | ~INSTQUEUE_REG_13__5__SCAN_IN;
  assign n7337 = ~n7936 | ~INSTQUEUE_REG_0__5__SCAN_IN;
  assign n7339 = ~n7338 | ~n7337;
  assign n7344 = ~n7006 | ~INSTQUEUE_REG_5__5__SCAN_IN;
  assign n7343 = ~n8453 | ~INSTQUEUE_REG_8__5__SCAN_IN;
  assign n7348 = ~n7344 | ~n7343;
  assign n7346 = ~n8029 | ~INSTQUEUE_REG_1__5__SCAN_IN;
  assign n7345 = ~n7014 | ~INSTQUEUE_REG_12__5__SCAN_IN;
  assign n7347 = ~n7346 | ~n7345;
  assign n7356 = ~n7348 & ~n7347;
  assign n7350 = ~n8586 | ~INSTQUEUE_REG_6__5__SCAN_IN;
  assign n7349 = ~n7639 | ~INSTQUEUE_REG_11__5__SCAN_IN;
  assign n7354 = ~n7350 | ~n7349;
  assign n7351 = ~n8279 | ~INSTQUEUE_REG_15__5__SCAN_IN;
  assign n7353 = ~n7352 | ~n7351;
  assign n7355 = ~n7354 & ~n7353;
  assign n7360 = ~n7326 | ~INSTQUEUE_REG_10__4__SCAN_IN;
  assign n7359 = ~n7336 | ~INSTQUEUE_REG_13__4__SCAN_IN;
  assign n7365 = ~n7360 | ~n7359;
  assign n7361 = ~INSTQUEUE_REG_3__4__SCAN_IN;
  assign n7362 = ~n7652 | ~INSTQUEUE_REG_9__4__SCAN_IN;
  assign n7364 = ~n7363 | ~n7362;
  assign n7367 = ~n8586 | ~INSTQUEUE_REG_6__4__SCAN_IN;
  assign n7366 = ~n7006 | ~INSTQUEUE_REG_5__4__SCAN_IN;
  assign n7371 = ~n7367 | ~n7366;
  assign n7369 = ~n7639 | ~INSTQUEUE_REG_11__4__SCAN_IN;
  assign n7368 = ~n8279 | ~INSTQUEUE_REG_15__4__SCAN_IN;
  assign n7370 = ~n7369 | ~n7368;
  assign n7372 = ~n7371 & ~n7370;
  assign n7376 = ~n7469 | ~INSTQUEUE_REG_14__4__SCAN_IN;
  assign n7380 = ~n7376 | ~n7375;
  assign n7378 = ~n7472 | ~INSTQUEUE_REG_7__4__SCAN_IN;
  assign n7377 = ~n7014 | ~INSTQUEUE_REG_12__4__SCAN_IN;
  assign n7379 = ~n7378 | ~n7377;
  assign n7388 = ~n7380 & ~n7379;
  assign n7382 = ~n7612 | ~INSTQUEUE_REG_4__4__SCAN_IN;
  assign n7381 = ~n8029 | ~INSTQUEUE_REG_1__4__SCAN_IN;
  assign n7386 = ~n7382 | ~n7381;
  assign n7384 = ~n8453 | ~INSTQUEUE_REG_8__4__SCAN_IN;
  assign n7383 = ~n7936 | ~INSTQUEUE_REG_0__4__SCAN_IN;
  assign n7385 = ~n7384 | ~n7383;
  assign n7496 = ~n7390 | ~n7389;
  assign n7395 = ~n7391 | ~n7492;
  assign n7392 = ~n7496 | ~n7773;
  assign n7393 = ~n7392 | ~n7495;
  assign n7394 = ~n7393 | ~n11918;
  assign n7429 = ~n7395 | ~n7394;
  assign n7397 = ~n7639 | ~INSTQUEUE_REG_11__3__SCAN_IN;
  assign n7396 = ~n7798 | ~INSTQUEUE_REG_14__3__SCAN_IN;
  assign n7401 = ~n7397 | ~n7396;
  assign n7399 = ~n7006 | ~INSTQUEUE_REG_5__3__SCAN_IN;
  assign n7398 = ~n8642 | ~INSTQUEUE_REG_2__3__SCAN_IN;
  assign n7400 = ~n7399 | ~n7398;
  assign n7410 = ~n7401 & ~n7400;
  assign n7403 = ~n8586 | ~INSTQUEUE_REG_6__3__SCAN_IN;
  assign n7402 = ~n8453 | ~INSTQUEUE_REG_8__3__SCAN_IN;
  assign n7408 = ~n7403 | ~n7402;
  assign n7406 = ~n7336 | ~INSTQUEUE_REG_13__3__SCAN_IN;
  assign n7405 = ~n7404 | ~INSTQUEUE_REG_3__3__SCAN_IN;
  assign n7407 = ~n7406 | ~n7405;
  assign n7409 = ~n7408 & ~n7407;
  assign n7426 = ~n7410 | ~n7409;
  assign n7412 = ~n7326 | ~INSTQUEUE_REG_10__3__SCAN_IN;
  assign n7411 = ~n7652 | ~INSTQUEUE_REG_9__3__SCAN_IN;
  assign n7416 = ~n7412 | ~n7411;
  assign n7414 = ~n8029 | ~INSTQUEUE_REG_1__3__SCAN_IN;
  assign n7413 = ~n7014 | ~INSTQUEUE_REG_12__3__SCAN_IN;
  assign n7415 = ~n7414 | ~n7413;
  assign n7418 = ~n7472 | ~INSTQUEUE_REG_7__3__SCAN_IN;
  assign n7417 = ~n7612 | ~INSTQUEUE_REG_4__3__SCAN_IN;
  assign n7422 = ~n7418 | ~n7417;
  assign n7420 = ~n7936 | ~INSTQUEUE_REG_0__3__SCAN_IN;
  assign n7419 = ~n8279 | ~INSTQUEUE_REG_15__3__SCAN_IN;
  assign n7421 = ~n7420 | ~n7419;
  assign n7423 = ~n7422 & ~n7421;
  assign n7425 = ~n7424 | ~n7423;
  assign n7427 = ~n8310 | ~n9210;
  assign n9849 = n7532;
  assign n7431 = ~n7326 | ~INSTQUEUE_REG_10__1__SCAN_IN;
  assign n7430 = ~n7336 | ~INSTQUEUE_REG_13__1__SCAN_IN;
  assign n7436 = ~n7431 | ~n7430;
  assign n7434 = ~n7652 | ~INSTQUEUE_REG_9__1__SCAN_IN;
  assign n8693 = ~n7432;
  assign n7433 = ~n7005 | ~INSTQUEUE_REG_3__1__SCAN_IN;
  assign n7435 = ~n7434 | ~n7433;
  assign n7444 = ~n7436 & ~n7435;
  assign n7438 = ~n8586 | ~INSTQUEUE_REG_6__1__SCAN_IN;
  assign n7437 = ~n7006 | ~INSTQUEUE_REG_5__1__SCAN_IN;
  assign n7442 = ~n7438 | ~n7437;
  assign n7440 = ~n7639 | ~INSTQUEUE_REG_11__1__SCAN_IN;
  assign n7439 = ~n8279 | ~INSTQUEUE_REG_15__1__SCAN_IN;
  assign n7441 = ~n7440 | ~n7439;
  assign n7443 = ~n7442 & ~n7441;
  assign n7460 = ~n7444 | ~n7443;
  assign n7446 = ~n7798 | ~INSTQUEUE_REG_14__1__SCAN_IN;
  assign n7445 = ~n8642 | ~INSTQUEUE_REG_2__1__SCAN_IN;
  assign n7450 = ~n7446 | ~n7445;
  assign n7448 = ~n7472 | ~INSTQUEUE_REG_7__1__SCAN_IN;
  assign n7447 = ~n7014 | ~INSTQUEUE_REG_12__1__SCAN_IN;
  assign n7449 = ~n7448 | ~n7447;
  assign n7458 = ~n7450 & ~n7449;
  assign n7452 = ~n7612 | ~INSTQUEUE_REG_4__1__SCAN_IN;
  assign n7451 = ~n8029 | ~INSTQUEUE_REG_1__1__SCAN_IN;
  assign n7456 = ~n7452 | ~n7451;
  assign n7454 = ~n8453 | ~INSTQUEUE_REG_8__1__SCAN_IN;
  assign n7453 = ~n7936 | ~INSTQUEUE_REG_0__1__SCAN_IN;
  assign n7455 = ~n7454 | ~n7453;
  assign n7459 = ~n7458 | ~n7457;
  assign n7461 = ~n7404 | ~INSTQUEUE_REG_3__0__SCAN_IN;
  assign n7463 = ~n8586 | ~INSTQUEUE_REG_6__0__SCAN_IN;
  assign n7462 = ~n7006 | ~INSTQUEUE_REG_5__0__SCAN_IN;
  assign n7467 = ~n7463 | ~n7462;
  assign n7465 = ~n7639 | ~INSTQUEUE_REG_11__0__SCAN_IN;
  assign n7464 = ~n8279 | ~INSTQUEUE_REG_15__0__SCAN_IN;
  assign n7466 = ~n7465 | ~n7464;
  assign n7468 = ~n7467 & ~n7466;
  assign n7471 = ~n7469 | ~INSTQUEUE_REG_14__0__SCAN_IN;
  assign n7470 = ~n8642 | ~INSTQUEUE_REG_2__0__SCAN_IN;
  assign n7476 = ~n7471 | ~n7470;
  assign n7474 = ~n7472 | ~INSTQUEUE_REG_7__0__SCAN_IN;
  assign n7473 = ~n7014 | ~INSTQUEUE_REG_12__0__SCAN_IN;
  assign n7475 = ~n7474 | ~n7473;
  assign n7484 = ~n7476 & ~n7475;
  assign n7478 = ~n7612 | ~INSTQUEUE_REG_4__0__SCAN_IN;
  assign n7477 = ~n8029 | ~INSTQUEUE_REG_1__0__SCAN_IN;
  assign n7482 = ~n7478 | ~n7477;
  assign n7480 = ~n8453 | ~INSTQUEUE_REG_8__0__SCAN_IN;
  assign n7479 = ~n7936 | ~INSTQUEUE_REG_0__0__SCAN_IN;
  assign n7481 = ~n7480 | ~n7479;
  assign n7483 = ~n7482 & ~n7481;
  assign n7485 = ~n7988;
  assign n7490 = ~n7486 | ~n7485;
  assign n7489 = ~n9081 | ~n9847;
  assign n9132 = ~n11938 | ~n7531;
  assign n7491 = ~n9132;
  assign n9302 = ~n7491 | ~n9230;
  assign n7493 = ~n7492 | ~n9849;
  assign n7494 = ~n7493 | ~n8940;
  assign n9187 = n7495 & n9849;
  assign n13311 = n7496;
  assign n7497 = n9847 | n13311;
  assign n7538 = ~n11908 | ~n9146;
  assign n7499 = ~n7538 | ~n11948;
  assign n7498 = ~n8946;
  assign n7500 = ~n7499 | ~n7498;
  assign n7502 = ~n7515 | ~n7501;
  assign n7503 = ~n7502 | ~STATE2_REG_0__SCAN_IN;
  assign n7508 = ~n7546 | ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n7506 = ~n9136 | ~n13354;
  assign n7505 = ~n9135 | ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n7507 = ~n7506 | ~n7505;
  assign n7674 = ~n7508 | ~n7507;
  assign n7509 = ~n9847 | ~n13311;
  assign n7510 = n9210 & n7509;
  assign n7513 = ~n7511 | ~n7510;
  assign n9454 = n7512;
  assign n7514 = ~n7513 | ~n9454;
  assign n7527 = ~n7515 | ~n7514;
  assign n7517 = ~n9307 & ~n11938;
  assign n9322 = ~n7517 | ~n9304;
  assign n7520 = ~n9322 | ~n13310;
  assign n7519 = ~n7004 | ~n11918;
  assign n7525 = ~n7520 | ~n7519;
  assign n7521 = ~n9847 | ~n9210;
  assign n7523 = ~n8940 | ~n7521;
  assign n13653 = ~n13402;
  assign n7522 = ~n13653 & ~n13400;
  assign n7524 = n7523 & n7522;
  assign n7526 = ~n7525 | ~n7524;
  assign n13743 = n13310 & n9454;
  assign n7528 = ~n13743 | ~n9132;
  assign n7534 = ~n7774;
  assign n7535 = ~n9132 & ~n7533;
  assign n9156 = n7535 & n7534;
  assign n7536 = ~n11948 | ~n11938;
  assign n9174 = ~n7537 | ~n9304;
  assign n9142 = n9174 | n13310;
  assign n7539 = ~n9142;
  assign n7540 = ~n7539 | ~n7538;
  assign n7542 = ~n7541 | ~n7540;
  assign n7549 = ~n7542 | ~STATE2_REG_0__SCAN_IN;
  assign n7545 = ~n7549;
  assign n7543 = ~n7727 | ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n7547 = ~n7544 | ~n7543;
  assign n7551 = ~n7546 | ~INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n7548 = ~n7547;
  assign n7559 = ~n7561;
  assign n7557 = ~n7546 | ~INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n13353 = ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n11903 = n13353 ^ ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n7553 = ~n9136;
  assign n7555 = ~n11903 | ~n7553;
  assign n7554 = ~n7727 | ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n7556 = n7555 & n7554;
  assign n7724 = ~n7559 | ~n7558;
  assign n7562 = ~n7561 | ~n7560;
  assign n7594 = ~n10855 | ~n13400;
  assign n7880 = ~n7006;
  assign n7564 = ~n9408 | ~INSTQUEUE_REG_6__2__SCAN_IN;
  assign n8892 = n7612;
  assign n7563 = ~n8892 | ~INSTQUEUE_REG_5__2__SCAN_IN;
  assign n7568 = ~n7564 | ~n7563;
  assign n8567 = ~n7927;
  assign n7566 = ~n8567 | ~INSTQUEUE_REG_3__2__SCAN_IN;
  assign n9401 = n8029;
  assign n7565 = ~n9401 | ~INSTQUEUE_REG_2__2__SCAN_IN;
  assign n7567 = ~n7566 | ~n7565;
  assign n7576 = ~n7568 & ~n7567;
  assign n7734 = ~n8562;
  assign n7570 = ~n7734 | ~INSTQUEUE_REG_14__2__SCAN_IN;
  assign n7569 = ~n8854 | ~INSTQUEUE_REG_9__2__SCAN_IN;
  assign n7574 = ~n7570 | ~n7569;
  assign n7572 = ~n8154 | ~INSTQUEUE_REG_13__2__SCAN_IN;
  assign n8537 = ~n8279;
  assign n7571 = ~n8279 | ~INSTQUEUE_REG_0__2__SCAN_IN;
  assign n7573 = ~n7572 | ~n7571;
  assign n7575 = ~n7574 & ~n7573;
  assign n7592 = n7576 & n7575;
  assign n7578 = ~n8587 | ~INSTQUEUE_REG_7__2__SCAN_IN;
  assign n7798 = ~n7374;
  assign n7577 = ~n7009 | ~INSTQUEUE_REG_15__2__SCAN_IN;
  assign n7582 = ~n7578 | ~n7577;
  assign n7580 = ~n8906 | ~INSTQUEUE_REG_11__2__SCAN_IN;
  assign n7579 = ~n8420 | ~INSTQUEUE_REG_4__2__SCAN_IN;
  assign n7581 = ~n7580 | ~n7579;
  assign n7590 = ~n7582 & ~n7581;
  assign n8915 = n7652;
  assign n7584 = ~n8915 | ~INSTQUEUE_REG_10__2__SCAN_IN;
  assign n7920 = ~n7639;
  assign n7583 = ~n8910 | ~INSTQUEUE_REG_12__2__SCAN_IN;
  assign n7588 = ~n7584 | ~n7583;
  assign n7692 = ~n7472;
  assign n7586 = ~n9398 | ~INSTQUEUE_REG_8__2__SCAN_IN;
  assign n8399 = ~n7936;
  assign n7807 = ~n8399;
  assign n7585 = ~n7807 | ~INSTQUEUE_REG_1__2__SCAN_IN;
  assign n7587 = ~n7586 | ~n7585;
  assign n7589 = ~n7588 & ~n7587;
  assign n7591 = n7590 & n7589;
  assign n7593 = n7733 | n8958;
  assign n7596 = ~INSTQUEUE_REG_0__2__SCAN_IN;
  assign n7598 = ~n7595 & ~n7596;
  assign n7597 = ~n7988 & ~n8958;
  assign n7599 = ~n7598 & ~n7597;
  assign n7602 = ~n10879;
  assign n7636 = ~n7602 | ~n13400;
  assign n7605 = ~n7734 | ~INSTQUEUE_REG_14__1__SCAN_IN;
  assign n7604 = ~n8854 | ~INSTQUEUE_REG_9__1__SCAN_IN;
  assign n7609 = ~n7605 | ~n7604;
  assign n7607 = ~n8587 | ~INSTQUEUE_REG_7__1__SCAN_IN;
  assign n7606 = ~n9401 | ~INSTQUEUE_REG_2__1__SCAN_IN;
  assign n7608 = ~n7607 | ~n7606;
  assign n7618 = ~n7609 & ~n7608;
  assign n7611 = ~n8910 | ~INSTQUEUE_REG_12__1__SCAN_IN;
  assign n7610 = ~n9398 | ~INSTQUEUE_REG_8__1__SCAN_IN;
  assign n7616 = ~n7611 | ~n7610;
  assign n7614 = ~n8892 | ~INSTQUEUE_REG_5__1__SCAN_IN;
  assign n7613 = ~n7014 | ~INSTQUEUE_REG_13__1__SCAN_IN;
  assign n7615 = ~n7614 | ~n7613;
  assign n7617 = ~n7616 & ~n7615;
  assign n7634 = n7618 & n7617;
  assign n7620 = ~n9408 | ~INSTQUEUE_REG_6__1__SCAN_IN;
  assign n7619 = ~n8151 | ~INSTQUEUE_REG_3__1__SCAN_IN;
  assign n7624 = ~n7620 | ~n7619;
  assign n7622 = ~n8915 | ~INSTQUEUE_REG_10__1__SCAN_IN;
  assign n7621 = ~n8420 | ~INSTQUEUE_REG_4__1__SCAN_IN;
  assign n7623 = ~n7622 | ~n7621;
  assign n7632 = ~n7624 & ~n7623;
  assign n7626 = ~n8906 | ~INSTQUEUE_REG_11__1__SCAN_IN;
  assign n7625 = ~n8279 | ~INSTQUEUE_REG_0__1__SCAN_IN;
  assign n7630 = ~n7626 | ~n7625;
  assign n7628 = ~n7009 | ~INSTQUEUE_REG_15__1__SCAN_IN;
  assign n7627 = ~n7807 | ~INSTQUEUE_REG_1__1__SCAN_IN;
  assign n7629 = ~n7628 | ~n7627;
  assign n7631 = ~n7630 & ~n7629;
  assign n7633 = n7632 & n7631;
  assign n7846 = ~n7636 | ~n7635;
  assign n7638 = ~n8587 | ~INSTQUEUE_REG_7__7__SCAN_IN;
  assign n7637 = ~n7009 | ~INSTQUEUE_REG_15__7__SCAN_IN;
  assign n7643 = ~n7638 | ~n7637;
  assign n7641 = ~n7639 | ~INSTQUEUE_REG_12__7__SCAN_IN;
  assign n7640 = ~n9401 | ~INSTQUEUE_REG_2__7__SCAN_IN;
  assign n7642 = ~n7641 | ~n7640;
  assign n7651 = ~n7643 & ~n7642;
  assign n7645 = ~n9408 | ~INSTQUEUE_REG_6__7__SCAN_IN;
  assign n7644 = ~n8854 | ~INSTQUEUE_REG_9__7__SCAN_IN;
  assign n7649 = ~n7645 | ~n7644;
  assign n7647 = ~n7807 | ~INSTQUEUE_REG_1__7__SCAN_IN;
  assign n7646 = ~n7014 | ~INSTQUEUE_REG_13__7__SCAN_IN;
  assign n7648 = ~n7647 | ~n7646;
  assign n7650 = ~n7649 & ~n7648;
  assign n7668 = ~n7651 | ~n7650;
  assign n7654 = ~n7326 | ~INSTQUEUE_REG_11__7__SCAN_IN;
  assign n7653 = ~n8915 | ~INSTQUEUE_REG_10__7__SCAN_IN;
  assign n7658 = ~n7654 | ~n7653;
  assign n7656 = ~n7734 | ~INSTQUEUE_REG_14__7__SCAN_IN;
  assign n7655 = ~n8892 | ~INSTQUEUE_REG_5__7__SCAN_IN;
  assign n7657 = ~n7656 | ~n7655;
  assign n7666 = ~n7658 & ~n7657;
  assign n7660 = ~n9398 | ~INSTQUEUE_REG_8__7__SCAN_IN;
  assign n7659 = ~n8279 | ~INSTQUEUE_REG_0__7__SCAN_IN;
  assign n7664 = ~n7660 | ~n7659;
  assign n7662 = ~n8567 | ~INSTQUEUE_REG_3__7__SCAN_IN;
  assign n7661 = ~n8693 | ~INSTQUEUE_REG_4__7__SCAN_IN;
  assign n7663 = ~n7662 | ~n7661;
  assign n7665 = ~n7664 & ~n7663;
  assign n7667 = ~n7666 | ~n7665;
  assign n7670 = n7733 | n9017;
  assign n7669 = n7988 | n8955;
  assign n7671 = ~n9081 | ~INSTQUEUE_REG_0__1__SCAN_IN;
  assign n7719 = ~n7846 | ~n7720;
  assign n7710 = ~n11938 | ~n9017;
  assign n7677 = ~n7326 | ~INSTQUEUE_REG_11__0__SCAN_IN;
  assign n7676 = ~n7734 | ~INSTQUEUE_REG_14__0__SCAN_IN;
  assign n7681 = ~n7677 | ~n7676;
  assign n7679 = ~n8915 | ~INSTQUEUE_REG_10__0__SCAN_IN;
  assign n7678 = ~n8420 | ~INSTQUEUE_REG_4__0__SCAN_IN;
  assign n7680 = ~n7679 | ~n7678;
  assign n7689 = ~n7681 & ~n7680;
  assign n7683 = ~n8587 | ~INSTQUEUE_REG_7__0__SCAN_IN;
  assign n7682 = ~n9408 | ~INSTQUEUE_REG_6__0__SCAN_IN;
  assign n7687 = ~n7683 | ~n7682;
  assign n7685 = ~n8910 | ~INSTQUEUE_REG_12__0__SCAN_IN;
  assign n7684 = ~n8279 | ~INSTQUEUE_REG_0__0__SCAN_IN;
  assign n7686 = ~n7685 | ~n7684;
  assign n7688 = ~n7687 & ~n7686;
  assign n7706 = n7689 & n7688;
  assign n7691 = ~n7009 | ~INSTQUEUE_REG_15__0__SCAN_IN;
  assign n7690 = ~n8567 | ~INSTQUEUE_REG_3__0__SCAN_IN;
  assign n7696 = ~n7691 | ~n7690;
  assign n9398 = ~n7692;
  assign n7694 = ~n9398 | ~INSTQUEUE_REG_8__0__SCAN_IN;
  assign n7693 = ~n7014 | ~INSTQUEUE_REG_13__0__SCAN_IN;
  assign n7695 = ~n7694 | ~n7693;
  assign n7704 = ~n7696 & ~n7695;
  assign n7698 = ~n8892 | ~INSTQUEUE_REG_5__0__SCAN_IN;
  assign n7697 = ~n9401 | ~INSTQUEUE_REG_2__0__SCAN_IN;
  assign n7702 = ~n7698 | ~n7697;
  assign n7700 = ~n8854 | ~INSTQUEUE_REG_9__0__SCAN_IN;
  assign n7699 = ~n7807 | ~INSTQUEUE_REG_1__0__SCAN_IN;
  assign n7701 = ~n7700 | ~n7699;
  assign n7703 = ~n7702 & ~n7701;
  assign n7705 = n7704 & n7703;
  assign n7709 = ~n9015 | ~n8954;
  assign n7969 = ~n9017;
  assign n7707 = ~n7969 | ~n8944;
  assign n7708 = n7733 | n7707;
  assign n7713 = ~n7710;
  assign n7711 = ~n13310 | ~n8944;
  assign n7712 = ~n7711 | ~STATE2_REG_0__SCAN_IN;
  assign n7715 = ~n7713 & ~n7712;
  assign n7714 = ~n9081 | ~INSTQUEUE_REG_0__0__SCAN_IN;
  assign n7856 = ~n7715 | ~n7714;
  assign n7717 = ~n7716 | ~n7856;
  assign n7718 = ~n7845;
  assign n7723 = ~n7719 | ~n7718;
  assign n7721 = ~n7846;
  assign n7722 = ~n7721 | ~n7844;
  assign n7830 = n7723 & n7722;
  assign n7731 = ~n7546 | ~INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n7725 = ~n12841 | ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n12240 = ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n12508 = ~n7725 & ~n12240;
  assign n12500 = ~n12508 | ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n7726 = ~n12500 | ~n12841;
  assign n12928 = ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n13205 = ~n12928 & ~n13355;
  assign n13197 = ~n13205 | ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n12589 = ~n7726 | ~n13197;
  assign n7729 = n12589 | n9136;
  assign n7728 = ~n7727 | ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n7732 = ~n10841;
  assign n7768 = ~n7732 | ~n13400;
  assign n7766 = ~n9081 | ~INSTQUEUE_REG_0__3__SCAN_IN;
  assign n8130 = ~n7326;
  assign n7736 = ~n8906 | ~INSTQUEUE_REG_11__3__SCAN_IN;
  assign n7735 = ~n7734 | ~INSTQUEUE_REG_14__3__SCAN_IN;
  assign n7740 = ~n7736 | ~n7735;
  assign n7738 = ~n8915 | ~INSTQUEUE_REG_10__3__SCAN_IN;
  assign n7737 = ~n8420 | ~INSTQUEUE_REG_4__3__SCAN_IN;
  assign n7739 = ~n7738 | ~n7737;
  assign n7748 = ~n7740 & ~n7739;
  assign n7742 = ~n8587 | ~INSTQUEUE_REG_7__3__SCAN_IN;
  assign n7741 = ~n9408 | ~INSTQUEUE_REG_6__3__SCAN_IN;
  assign n7746 = ~n7742 | ~n7741;
  assign n7744 = ~n8910 | ~INSTQUEUE_REG_12__3__SCAN_IN;
  assign n7743 = ~n8907 | ~INSTQUEUE_REG_0__3__SCAN_IN;
  assign n7745 = ~n7744 | ~n7743;
  assign n7747 = ~n7746 & ~n7745;
  assign n7764 = ~n7748 | ~n7747;
  assign n7750 = ~n7009 | ~INSTQUEUE_REG_15__3__SCAN_IN;
  assign n7927 = ~n8642;
  assign n7749 = ~n8151 | ~INSTQUEUE_REG_3__3__SCAN_IN;
  assign n7754 = ~n7750 | ~n7749;
  assign n7752 = ~n9398 | ~INSTQUEUE_REG_8__3__SCAN_IN;
  assign n7751 = ~n7014 | ~INSTQUEUE_REG_13__3__SCAN_IN;
  assign n7753 = ~n7752 | ~n7751;
  assign n7762 = ~n7754 & ~n7753;
  assign n7756 = ~n8892 | ~INSTQUEUE_REG_5__3__SCAN_IN;
  assign n7755 = ~n9401 | ~INSTQUEUE_REG_2__3__SCAN_IN;
  assign n7760 = ~n7756 | ~n7755;
  assign n7758 = ~n8854 | ~INSTQUEUE_REG_9__3__SCAN_IN;
  assign n7757 = ~n7807 | ~INSTQUEUE_REG_1__3__SCAN_IN;
  assign n7759 = ~n7758 | ~n7757;
  assign n7761 = ~n7760 & ~n7759;
  assign n7763 = ~n7762 | ~n7761;
  assign n7765 = ~n9126 | ~n8981;
  assign n7770 = ~n7783;
  assign n7772 = ~n7771 | ~n7770;
  assign n7782 = ~n11884 | ~n7987;
  assign n7863 = ~n7774 & ~n11983;
  assign n7778 = ~n7863 | ~INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n7864 = ~n9849 & ~n11983;
  assign n7776 = ~n8880 | ~EAX_REG_3__SCAN_IN;
  assign n7775 = ~n9446 | ~PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n7777 = n7776 & n7775;
  assign n7780 = ~n7778 | ~n7777;
  assign n7824 = ~PHYADDRPOINTER_REG_1__SCAN_IN | ~PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n11528 = PHYADDRPOINTER_REG_3__SCAN_IN ^ n7824;
  assign n7779 = n11528 & n8929;
  assign n7781 = ~n7780 & ~n7779;
  assign n7817 = ~n9081 | ~INSTQUEUE_REG_0__4__SCAN_IN;
  assign n7785 = ~n8906 | ~INSTQUEUE_REG_11__4__SCAN_IN;
  assign n7784 = ~n8526 | ~INSTQUEUE_REG_14__4__SCAN_IN;
  assign n7789 = ~n7785 | ~n7784;
  assign n7787 = ~n8915 | ~INSTQUEUE_REG_10__4__SCAN_IN;
  assign n7786 = ~n8693 | ~INSTQUEUE_REG_4__4__SCAN_IN;
  assign n7788 = ~n7787 | ~n7786;
  assign n7797 = ~n7789 & ~n7788;
  assign n7791 = ~n8587 | ~INSTQUEUE_REG_7__4__SCAN_IN;
  assign n7790 = ~n9408 | ~INSTQUEUE_REG_6__4__SCAN_IN;
  assign n7795 = ~n7791 | ~n7790;
  assign n7793 = ~n8910 | ~INSTQUEUE_REG_12__4__SCAN_IN;
  assign n7792 = ~n8907 | ~INSTQUEUE_REG_0__4__SCAN_IN;
  assign n7794 = ~n7793 | ~n7792;
  assign n7796 = ~n7795 & ~n7794;
  assign n7815 = ~n7797 | ~n7796;
  assign n7800 = ~n7009 | ~INSTQUEUE_REG_15__4__SCAN_IN;
  assign n7799 = ~n8151 | ~INSTQUEUE_REG_3__4__SCAN_IN;
  assign n7804 = ~n7800 | ~n7799;
  assign n7802 = ~n9398 | ~INSTQUEUE_REG_8__4__SCAN_IN;
  assign n7801 = ~n8154 | ~INSTQUEUE_REG_13__4__SCAN_IN;
  assign n7803 = ~n7802 | ~n7801;
  assign n7813 = ~n7804 & ~n7803;
  assign n7806 = ~n8892 | ~INSTQUEUE_REG_5__4__SCAN_IN;
  assign n7805 = ~n9401 | ~INSTQUEUE_REG_2__4__SCAN_IN;
  assign n7811 = ~n7806 | ~n7805;
  assign n7809 = ~n8854 | ~INSTQUEUE_REG_9__4__SCAN_IN;
  assign n7808 = ~n7807 | ~INSTQUEUE_REG_1__4__SCAN_IN;
  assign n7810 = ~n7809 | ~n7808;
  assign n7812 = ~n7811 & ~n7810;
  assign n7814 = ~n7813 | ~n7812;
  assign n7816 = ~n9126 | ~n8989;
  assign n8980 = n7956 ^ ~n7957;
  assign n7818 = ~n8980;
  assign n7828 = ~n7818 | ~n7987;
  assign n7823 = ~n7863 | ~INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n7821 = ~n8880 | ~EAX_REG_4__SCAN_IN;
  assign n8929 = ~n8384;
  assign n7819 = n9446 & PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n7820 = ~n8929 & ~n7819;
  assign n7822 = n7821 & n7820;
  assign n7826 = ~n7823 | ~n7822;
  assign n11522 = n7950 ^ ~PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n7825 = n11522 | n8384;
  assign n7827 = ~n7826 | ~n7825;
  assign n7832 = ~n7829;
  assign n7831 = ~n7830;
  assign n7833 = ~n11880;
  assign n7835 = ~n7833 | ~n7987;
  assign n7834 = ~n9446;
  assign n7843 = ~n7863 | ~INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n7841 = ~n8880 | ~EAX_REG_2__SCAN_IN;
  assign n11547 = PHYADDRPOINTER_REG_1__SCAN_IN ^ PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n7836 = ~n11547;
  assign n7839 = ~n7837 | ~n7836;
  assign n7838 = ~n9446 | ~PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n7840 = n7839 & n7838;
  assign n7842 = n7841 & n7840;
  assign n7874 = ~n7843 | ~n7842;
  assign n7873 = ~n7875 | ~n7874;
  assign n7854 = ~n7848 | ~n7987;
  assign n7852 = ~n7863 | ~INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n7850 = ~n8880 | ~EAX_REG_1__SCAN_IN;
  assign n7849 = ~n11983 | ~PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n7851 = n7850 & n7849;
  assign n7853 = n7852 & n7851;
  assign n10887 = ~n7854 | ~n7853;
  assign n7858 = ~n7856;
  assign n7857 = ~n7859 & ~n7858;
  assign n7860 = ~n7859 | ~n7858;
  assign n7862 = ~n8939 | ~n9304;
  assign n10923 = ~n7862 | ~STATE2_REG_2__SCAN_IN;
  assign n7870 = ~n13703 | ~n7987;
  assign n7868 = ~n7863 | ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n7866 = ~n7864 | ~EAX_REG_0__SCAN_IN;
  assign n7865 = ~n11983 | ~PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n7867 = n7866 & n7865;
  assign n7869 = n7868 & n7867;
  assign n7872 = n10923 | n10921;
  assign n7871 = ~n10921 | ~n7837;
  assign n10886 = ~n7872 | ~n7871;
  assign n10889 = ~n10887 | ~n10886;
  assign n7876 = ~n7873 | ~n10889;
  assign n10766 = ~n7877 | ~n10821;
  assign n7910 = ~n9081 | ~INSTQUEUE_REG_0__5__SCAN_IN;
  assign n7879 = ~n8906 | ~INSTQUEUE_REG_11__5__SCAN_IN;
  assign n7878 = ~n8915 | ~INSTQUEUE_REG_10__5__SCAN_IN;
  assign n7884 = ~n7879 | ~n7878;
  assign n7882 = ~n9408 | ~INSTQUEUE_REG_6__5__SCAN_IN;
  assign n7881 = ~n8892 | ~INSTQUEUE_REG_5__5__SCAN_IN;
  assign n7883 = ~n7882 | ~n7881;
  assign n7892 = ~n7884 & ~n7883;
  assign n7886 = ~n7009 | ~INSTQUEUE_REG_15__5__SCAN_IN;
  assign n7885 = ~n8151 | ~INSTQUEUE_REG_3__5__SCAN_IN;
  assign n7890 = ~n7886 | ~n7885;
  assign n7888 = ~n8587 | ~INSTQUEUE_REG_7__5__SCAN_IN;
  assign n7887 = ~n8154 | ~INSTQUEUE_REG_13__5__SCAN_IN;
  assign n7889 = ~n7888 | ~n7887;
  assign n7891 = ~n7890 & ~n7889;
  assign n7908 = ~n7892 | ~n7891;
  assign n7894 = ~n8526 | ~INSTQUEUE_REG_14__5__SCAN_IN;
  assign n7893 = ~n8854 | ~INSTQUEUE_REG_9__5__SCAN_IN;
  assign n7898 = ~n7894 | ~n7893;
  assign n7896 = ~n9401 | ~INSTQUEUE_REG_2__5__SCAN_IN;
  assign n7895 = ~n7807 | ~INSTQUEUE_REG_1__5__SCAN_IN;
  assign n7897 = ~n7896 | ~n7895;
  assign n7906 = ~n7898 & ~n7897;
  assign n7900 = ~n8910 | ~INSTQUEUE_REG_12__5__SCAN_IN;
  assign n7899 = ~n9398 | ~INSTQUEUE_REG_8__5__SCAN_IN;
  assign n7904 = ~n7900 | ~n7899;
  assign n7902 = ~n8420 | ~INSTQUEUE_REG_4__5__SCAN_IN;
  assign n7901 = ~n8907 | ~INSTQUEUE_REG_0__5__SCAN_IN;
  assign n7903 = ~n7902 | ~n7901;
  assign n7905 = ~n7904 & ~n7903;
  assign n7907 = ~n7906 | ~n7905;
  assign n7909 = ~n9126 | ~n8996;
  assign n7958 = ~n7910 | ~n7909;
  assign n7946 = ~n9081 | ~INSTQUEUE_REG_0__6__SCAN_IN;
  assign n7913 = ~n8906 | ~INSTQUEUE_REG_11__6__SCAN_IN;
  assign n7912 = ~n8526 | ~INSTQUEUE_REG_14__6__SCAN_IN;
  assign n7917 = ~n7913 | ~n7912;
  assign n7915 = ~n8915 | ~INSTQUEUE_REG_10__6__SCAN_IN;
  assign n7914 = ~n8693 | ~INSTQUEUE_REG_4__6__SCAN_IN;
  assign n7916 = ~n7915 | ~n7914;
  assign n7926 = ~n7917 & ~n7916;
  assign n7919 = ~n8587 | ~INSTQUEUE_REG_7__6__SCAN_IN;
  assign n7918 = ~n9408 | ~INSTQUEUE_REG_6__6__SCAN_IN;
  assign n7924 = ~n7919 | ~n7918;
  assign n8910 = ~n7920;
  assign n7922 = ~n8910 | ~INSTQUEUE_REG_12__6__SCAN_IN;
  assign n7921 = ~n8907 | ~INSTQUEUE_REG_0__6__SCAN_IN;
  assign n7923 = ~n7922 | ~n7921;
  assign n7925 = ~n7924 & ~n7923;
  assign n7944 = ~n7926 | ~n7925;
  assign n7929 = ~n7009 | ~INSTQUEUE_REG_15__6__SCAN_IN;
  assign n7928 = ~n8151 | ~INSTQUEUE_REG_3__6__SCAN_IN;
  assign n7933 = ~n7929 | ~n7928;
  assign n7931 = ~n9398 | ~INSTQUEUE_REG_8__6__SCAN_IN;
  assign n7930 = ~n8154 | ~INSTQUEUE_REG_13__6__SCAN_IN;
  assign n7932 = ~n7931 | ~n7930;
  assign n7942 = ~n7933 & ~n7932;
  assign n7935 = ~n8892 | ~INSTQUEUE_REG_5__6__SCAN_IN;
  assign n7934 = ~n9401 | ~INSTQUEUE_REG_2__6__SCAN_IN;
  assign n7940 = ~n7935 | ~n7934;
  assign n7938 = ~n8854 | ~INSTQUEUE_REG_9__6__SCAN_IN;
  assign n7937 = ~n7807 | ~INSTQUEUE_REG_1__6__SCAN_IN;
  assign n7939 = ~n7938 | ~n7937;
  assign n7941 = ~n7940 & ~n7939;
  assign n7943 = ~n7942 | ~n7941;
  assign n7945 = ~n9126 | ~n9007;
  assign n7955 = ~n8994 | ~n7987;
  assign n7949 = ~n8880 | ~EAX_REG_6__SCAN_IN;
  assign n7947 = PHYADDRPOINTER_REG_6__SCAN_IN & n11983;
  assign n7948 = ~n8929 & ~n7947;
  assign n7953 = ~n7949 | ~n7948;
  assign n7959 = ~n7950 | ~PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n7951 = ~n7975;
  assign n11493 = PHYADDRPOINTER_REG_6__SCAN_IN ^ ~n7951;
  assign n7952 = ~n11493 | ~n8929;
  assign n7954 = ~n7953 | ~n7952;
  assign n10765 = ~n7955 | ~n7954;
  assign n7963 = ~n8880 | ~EAX_REG_5__SCAN_IN;
  assign n11509 = PHYADDRPOINTER_REG_5__SCAN_IN ^ ~n7959;
  assign n7961 = n11509 | n8384;
  assign n7960 = ~n9446 | ~PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n7962 = n7961 & n7960;
  assign n7964 = n7963 & n7962;
  assign n10767 = ~n7965 | ~n7964;
  assign n7968 = ~INSTQUEUE_REG_0__7__SCAN_IN;
  assign n7972 = ~n7595 & ~n7968;
  assign n7970 = n7988 | n7969;
  assign n7971 = ~n8142 | ~n7970;
  assign n7973 = ~n7972 & ~n7971;
  assign n7974 = ~n9006;
  assign n7981 = ~n7974 | ~n7987;
  assign n11487 = PHYADDRPOINTER_REG_7__SCAN_IN ^ n7982;
  assign n7979 = n11487 & n8929;
  assign n7977 = ~n7864 | ~EAX_REG_7__SCAN_IN;
  assign n7976 = ~n9446 | ~PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n7978 = ~n7977 | ~n7976;
  assign n7980 = ~n7979 & ~n7978;
  assign n11471 = PHYADDRPOINTER_REG_8__SCAN_IN ^ ~n8022;
  assign n7986 = n11471 & n8929;
  assign n7984 = ~n8880 | ~EAX_REG_8__SCAN_IN;
  assign n7983 = ~n9446 | ~PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n7985 = ~n7984 | ~n7983;
  assign n8021 = ~n7986 & ~n7985;
  assign n8143 = n7595 & n7988;
  assign n7990 = ~n8906 | ~INSTQUEUE_REG_12__0__SCAN_IN;
  assign n7989 = ~n8892 | ~INSTQUEUE_REG_6__0__SCAN_IN;
  assign n7994 = ~n7990 | ~n7989;
  assign n7992 = ~n9398 | ~INSTQUEUE_REG_9__0__SCAN_IN;
  assign n7991 = ~n9401 | ~INSTQUEUE_REG_3__0__SCAN_IN;
  assign n7993 = ~n7992 | ~n7991;
  assign n8002 = ~n7994 & ~n7993;
  assign n7996 = ~n8910 | ~INSTQUEUE_REG_13__0__SCAN_IN;
  assign n7995 = ~n7469 | ~INSTQUEUE_REG_0__0__SCAN_IN;
  assign n8000 = ~n7996 | ~n7995;
  assign n7998 = ~n8587 | ~INSTQUEUE_REG_8__0__SCAN_IN;
  assign n7997 = ~n8693 | ~INSTQUEUE_REG_5__0__SCAN_IN;
  assign n7999 = ~n7998 | ~n7997;
  assign n8001 = ~n8000 & ~n7999;
  assign n8018 = ~n8002 | ~n8001;
  assign n8004 = ~n7734 | ~INSTQUEUE_REG_15__0__SCAN_IN;
  assign n8003 = ~n8854 | ~INSTQUEUE_REG_10__0__SCAN_IN;
  assign n8008 = ~n8004 | ~n8003;
  assign n8006 = ~n8915 | ~INSTQUEUE_REG_11__0__SCAN_IN;
  assign n8005 = ~n8154 | ~INSTQUEUE_REG_14__0__SCAN_IN;
  assign n8007 = ~n8006 | ~n8005;
  assign n8016 = ~n8008 & ~n8007;
  assign n8010 = ~n9408 | ~INSTQUEUE_REG_7__0__SCAN_IN;
  assign n8009 = ~n8907 | ~INSTQUEUE_REG_1__0__SCAN_IN;
  assign n8014 = ~n8010 | ~n8009;
  assign n8012 = ~n8151 | ~INSTQUEUE_REG_4__0__SCAN_IN;
  assign n8011 = ~n7807 | ~INSTQUEUE_REG_2__0__SCAN_IN;
  assign n8013 = ~n8012 | ~n8011;
  assign n8015 = ~n8014 & ~n8013;
  assign n8017 = ~n8016 | ~n8015;
  assign n11463 = PHYADDRPOINTER_REG_9__SCAN_IN ^ ~n8062;
  assign n8026 = ~n11463 & ~n8384;
  assign n8024 = ~n8880 | ~EAX_REG_9__SCAN_IN;
  assign n8023 = ~n9446 | ~PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n8025 = ~n8024 | ~n8023;
  assign n8059 = ~n8026 & ~n8025;
  assign n8028 = ~n9408 | ~INSTQUEUE_REG_7__1__SCAN_IN;
  assign n8027 = ~n7469 | ~INSTQUEUE_REG_0__1__SCAN_IN;
  assign n8033 = ~n8028 | ~n8027;
  assign n8031 = ~n8892 | ~INSTQUEUE_REG_6__1__SCAN_IN;
  assign n8030 = ~n8899 | ~INSTQUEUE_REG_3__1__SCAN_IN;
  assign n8032 = ~n8031 | ~n8030;
  assign n8049 = n8033 | n8032;
  assign n8035 = ~n9398 | ~INSTQUEUE_REG_9__1__SCAN_IN;
  assign n8034 = ~n8420 | ~INSTQUEUE_REG_5__1__SCAN_IN;
  assign n8039 = ~n8035 | ~n8034;
  assign n8037 = ~n8906 | ~INSTQUEUE_REG_12__1__SCAN_IN;
  assign n8036 = ~n8154 | ~INSTQUEUE_REG_14__1__SCAN_IN;
  assign n8038 = ~n8037 | ~n8036;
  assign n8047 = ~n8039 & ~n8038;
  assign n8041 = ~n8910 | ~INSTQUEUE_REG_13__1__SCAN_IN;
  assign n8040 = ~n8907 | ~INSTQUEUE_REG_1__1__SCAN_IN;
  assign n8045 = ~n8041 | ~n8040;
  assign n8043 = ~n8587 | ~INSTQUEUE_REG_8__1__SCAN_IN;
  assign n8526 = ~n8562;
  assign n8042 = ~n8526 | ~INSTQUEUE_REG_15__1__SCAN_IN;
  assign n8044 = ~n8043 | ~n8042;
  assign n8046 = ~n8045 & ~n8044;
  assign n8048 = ~n8047 | ~n8046;
  assign n8057 = ~n8049 & ~n8048;
  assign n8051 = ~n8915 | ~INSTQUEUE_REG_11__1__SCAN_IN;
  assign n8050 = ~n7807 | ~INSTQUEUE_REG_2__1__SCAN_IN;
  assign n8055 = ~n8051 | ~n8050;
  assign n8053 = ~n8854 | ~INSTQUEUE_REG_10__1__SCAN_IN;
  assign n8052 = ~n8151 | ~INSTQUEUE_REG_4__1__SCAN_IN;
  assign n8054 = ~n8053 | ~n8052;
  assign n8056 = ~n8055 & ~n8054;
  assign n8058 = ~n8019 | ~n7229;
  assign n11446 = n8103 ^ ~PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n8066 = ~n11446 | ~n7837;
  assign n8064 = ~n7864 | ~EAX_REG_10__SCAN_IN;
  assign n8063 = ~n9446 | ~PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n8065 = n8064 & n8063;
  assign n8102 = n8066 & n8065;
  assign n8067 = ~INSTQUEUE_REG_13__2__SCAN_IN;
  assign n8070 = ~n7920 & ~n8067;
  assign n8068 = ~INSTQUEUE_REG_9__2__SCAN_IN;
  assign n8069 = ~n7692 & ~n8068;
  assign n8075 = ~n8070 & ~n8069;
  assign n8073 = ~n7010 & ~n7596;
  assign n8071 = ~INSTQUEUE_REG_2__2__SCAN_IN;
  assign n8072 = ~n8399 & ~n8071;
  assign n8074 = ~n8073 & ~n8072;
  assign n8091 = ~n8075 | ~n8074;
  assign n8077 = ~n8906 | ~INSTQUEUE_REG_12__2__SCAN_IN;
  assign n8076 = ~n9408 | ~INSTQUEUE_REG_7__2__SCAN_IN;
  assign n8081 = ~n8077 | ~n8076;
  assign n8151 = ~n7927;
  assign n8079 = ~n8151 | ~INSTQUEUE_REG_4__2__SCAN_IN;
  assign n8078 = ~n8154 | ~INSTQUEUE_REG_14__2__SCAN_IN;
  assign n8080 = ~n8079 | ~n8078;
  assign n8089 = ~n8081 & ~n8080;
  assign n8083 = ~n8915 | ~INSTQUEUE_REG_11__2__SCAN_IN;
  assign n8082 = ~n8892 | ~INSTQUEUE_REG_6__2__SCAN_IN;
  assign n8087 = ~n8083 | ~n8082;
  assign n8085 = ~n8526 | ~INSTQUEUE_REG_15__2__SCAN_IN;
  assign n8084 = ~n8907 | ~INSTQUEUE_REG_1__2__SCAN_IN;
  assign n8086 = ~n8085 | ~n8084;
  assign n8088 = ~n8087 & ~n8086;
  assign n8090 = ~n8089 | ~n8088;
  assign n8099 = ~n8091 & ~n8090;
  assign n8093 = ~n8587 | ~INSTQUEUE_REG_8__2__SCAN_IN;
  assign n8092 = ~n8854 | ~INSTQUEUE_REG_10__2__SCAN_IN;
  assign n8097 = ~n8093 | ~n8092;
  assign n8095 = ~n8899 | ~INSTQUEUE_REG_3__2__SCAN_IN;
  assign n8094 = ~n8420 | ~INSTQUEUE_REG_5__2__SCAN_IN;
  assign n8096 = ~n8095 | ~n8094;
  assign n8098 = ~n8097 & ~n8096;
  assign n8100 = n8099 & n8098;
  assign n8101 = n8305 | n8100;
  assign n8107 = ~n7864 | ~EAX_REG_11__SCAN_IN;
  assign n11430 = PHYADDRPOINTER_REG_11__SCAN_IN ^ ~n8180;
  assign n8105 = n11430 | n8384;
  assign n8104 = ~n9446 | ~PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n8106 = n8105 & n8104;
  assign n8141 = n8107 & n8106;
  assign n8109 = ~n7469 | ~INSTQUEUE_REG_0__3__SCAN_IN;
  assign n8108 = ~n8892 | ~INSTQUEUE_REG_6__3__SCAN_IN;
  assign n8113 = ~n8109 | ~n8108;
  assign n8111 = ~n8567 | ~INSTQUEUE_REG_4__3__SCAN_IN;
  assign n8110 = ~n8693 | ~INSTQUEUE_REG_5__3__SCAN_IN;
  assign n8112 = ~n8111 | ~n8110;
  assign n8129 = n8113 | n8112;
  assign n8115 = ~n8526 | ~INSTQUEUE_REG_15__3__SCAN_IN;
  assign n8114 = ~n8910 | ~INSTQUEUE_REG_13__3__SCAN_IN;
  assign n8119 = ~n8115 | ~n8114;
  assign n8117 = ~n9398 | ~INSTQUEUE_REG_9__3__SCAN_IN;
  assign n8116 = ~n7807 | ~INSTQUEUE_REG_2__3__SCAN_IN;
  assign n8118 = ~n8117 | ~n8116;
  assign n8127 = ~n8119 & ~n8118;
  assign n8121 = ~n8899 | ~INSTQUEUE_REG_3__3__SCAN_IN;
  assign n8120 = ~n8907 | ~INSTQUEUE_REG_1__3__SCAN_IN;
  assign n8125 = ~n8121 | ~n8120;
  assign n8123 = ~n9408 | ~INSTQUEUE_REG_7__3__SCAN_IN;
  assign n8122 = ~n8586 | ~INSTQUEUE_REG_8__3__SCAN_IN;
  assign n8124 = ~n8123 | ~n8122;
  assign n8126 = ~n8125 & ~n8124;
  assign n8128 = ~n8127 | ~n8126;
  assign n8138 = ~n8129 & ~n8128;
  assign n8132 = ~n8906 | ~INSTQUEUE_REG_12__3__SCAN_IN;
  assign n8131 = ~n8154 | ~INSTQUEUE_REG_14__3__SCAN_IN;
  assign n8136 = ~n8132 | ~n8131;
  assign n8134 = ~n8915 | ~INSTQUEUE_REG_11__3__SCAN_IN;
  assign n8133 = ~n8854 | ~INSTQUEUE_REG_10__3__SCAN_IN;
  assign n8135 = ~n8134 | ~n8133;
  assign n8137 = ~n8136 & ~n8135;
  assign n8139 = n8138 & n8137;
  assign n8140 = n8305 | n8139;
  assign n10662 = ~n8141 | ~n8140;
  assign n8144 = ~n8143 | ~n8142;
  assign n8146 = ~n8915 | ~INSTQUEUE_REG_11__4__SCAN_IN;
  assign n8145 = ~n8526 | ~INSTQUEUE_REG_15__4__SCAN_IN;
  assign n8150 = ~n8146 | ~n8145;
  assign n8148 = ~n7469 | ~INSTQUEUE_REG_0__4__SCAN_IN;
  assign n8147 = ~n8899 | ~INSTQUEUE_REG_3__4__SCAN_IN;
  assign n8149 = ~n8148 | ~n8147;
  assign n8168 = n8150 | n8149;
  assign n8153 = ~n8587 | ~INSTQUEUE_REG_8__4__SCAN_IN;
  assign n8152 = ~n8151 | ~INSTQUEUE_REG_4__4__SCAN_IN;
  assign n8158 = ~n8153 | ~n8152;
  assign n8156 = ~n9408 | ~INSTQUEUE_REG_7__4__SCAN_IN;
  assign n8155 = ~n8154 | ~INSTQUEUE_REG_14__4__SCAN_IN;
  assign n8157 = ~n8156 | ~n8155;
  assign n8166 = ~n8158 & ~n8157;
  assign n8160 = ~n8906 | ~INSTQUEUE_REG_12__4__SCAN_IN;
  assign n8159 = ~n8892 | ~INSTQUEUE_REG_6__4__SCAN_IN;
  assign n8164 = ~n8160 | ~n8159;
  assign n8162 = ~n8693 | ~INSTQUEUE_REG_5__4__SCAN_IN;
  assign n8161 = ~n8907 | ~INSTQUEUE_REG_1__4__SCAN_IN;
  assign n8163 = ~n8162 | ~n8161;
  assign n8165 = ~n8164 & ~n8163;
  assign n8167 = ~n8166 | ~n8165;
  assign n8176 = ~n8168 & ~n8167;
  assign n8170 = ~n9398 | ~INSTQUEUE_REG_9__4__SCAN_IN;
  assign n8169 = ~n7807 | ~INSTQUEUE_REG_2__4__SCAN_IN;
  assign n8174 = ~n8170 | ~n8169;
  assign n8172 = ~n8910 | ~INSTQUEUE_REG_13__4__SCAN_IN;
  assign n8171 = ~n8854 | ~INSTQUEUE_REG_10__4__SCAN_IN;
  assign n8173 = ~n8172 | ~n8171;
  assign n8175 = ~n8174 & ~n8173;
  assign n8177 = ~n8176 | ~n8175;
  assign n8178 = ~n8177 & ~n9015;
  assign n11412 = PHYADDRPOINTER_REG_12__SCAN_IN ^ ~n8222;
  assign n8181 = ~n11412;
  assign n8186 = ~n8181 | ~n8929;
  assign n8184 = ~n7864 | ~EAX_REG_12__SCAN_IN;
  assign n8182 = ~PHYADDRPOINTER_REG_12__SCAN_IN & ~n13100;
  assign n8183 = STATE2_REG_2__SCAN_IN | n8182;
  assign n8185 = ~n8184 | ~n8183;
  assign n8187 = ~n8186 | ~n8185;
  assign n8189 = n10662 & n10641;
  assign n8191 = ~n8906 | ~INSTQUEUE_REG_12__5__SCAN_IN;
  assign n8190 = ~n8907 | ~INSTQUEUE_REG_1__5__SCAN_IN;
  assign n8195 = ~n8191 | ~n8190;
  assign n8193 = ~n9398 | ~INSTQUEUE_REG_9__5__SCAN_IN;
  assign n8192 = ~n7009 | ~INSTQUEUE_REG_0__5__SCAN_IN;
  assign n8194 = ~n8193 | ~n8192;
  assign n8211 = n8195 | n8194;
  assign n8197 = ~n8910 | ~INSTQUEUE_REG_13__5__SCAN_IN;
  assign n8196 = ~n8151 | ~INSTQUEUE_REG_4__5__SCAN_IN;
  assign n8201 = ~n8197 | ~n8196;
  assign n8199 = ~n9408 | ~INSTQUEUE_REG_7__5__SCAN_IN;
  assign n8198 = ~n8587 | ~INSTQUEUE_REG_8__5__SCAN_IN;
  assign n8200 = ~n8199 | ~n8198;
  assign n8209 = ~n8201 & ~n8200;
  assign n8203 = ~n8526 | ~INSTQUEUE_REG_15__5__SCAN_IN;
  assign n8202 = ~n8154 | ~INSTQUEUE_REG_14__5__SCAN_IN;
  assign n8207 = ~n8203 | ~n8202;
  assign n8205 = ~n8892 | ~INSTQUEUE_REG_6__5__SCAN_IN;
  assign n8204 = ~n8693 | ~INSTQUEUE_REG_5__5__SCAN_IN;
  assign n8206 = ~n8205 | ~n8204;
  assign n8208 = ~n8207 & ~n8206;
  assign n8210 = ~n8209 | ~n8208;
  assign n8219 = ~n8211 & ~n8210;
  assign n8213 = ~n8915 | ~INSTQUEUE_REG_11__5__SCAN_IN;
  assign n8212 = ~n8854 | ~INSTQUEUE_REG_10__5__SCAN_IN;
  assign n8217 = ~n8213 | ~n8212;
  assign n8215 = ~n8899 | ~INSTQUEUE_REG_3__5__SCAN_IN;
  assign n8214 = ~n7807 | ~INSTQUEUE_REG_2__5__SCAN_IN;
  assign n8216 = ~n8215 | ~n8214;
  assign n8218 = ~n8217 & ~n8216;
  assign n8220 = ~n8219 | ~n8218;
  assign n10624 = n8229 ^ ~PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n8226 = n10624 | n8384;
  assign n8224 = ~n8880 | ~EAX_REG_13__SCAN_IN;
  assign n8223 = ~n9446 | ~PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n8225 = n8224 & n8223;
  assign n10149 = ~n8226 | ~n8225;
  assign n8228 = ~n8227;
  assign n10605 = PHYADDRPOINTER_REG_14__SCAN_IN ^ n8268;
  assign n8234 = ~n10605 | ~n7837;
  assign n8232 = ~n7864 | ~EAX_REG_14__SCAN_IN;
  assign n8230 = PHYADDRPOINTER_REG_14__SCAN_IN | n13100;
  assign n8231 = ~n8230 | ~n11983;
  assign n8233 = ~n8232 | ~n8231;
  assign n8267 = ~n8234 | ~n8233;
  assign n8236 = ~n8906 | ~INSTQUEUE_REG_12__6__SCAN_IN;
  assign n8235 = ~n7469 | ~INSTQUEUE_REG_0__6__SCAN_IN;
  assign n8240 = ~n8236 | ~n8235;
  assign n8238 = ~n8854 | ~INSTQUEUE_REG_10__6__SCAN_IN;
  assign n8237 = ~n8892 | ~INSTQUEUE_REG_6__6__SCAN_IN;
  assign n8239 = ~n8238 | ~n8237;
  assign n8256 = n8240 | n8239;
  assign n8242 = ~n9398 | ~INSTQUEUE_REG_9__6__SCAN_IN;
  assign n8241 = ~n8899 | ~INSTQUEUE_REG_3__6__SCAN_IN;
  assign n8246 = ~n8242 | ~n8241;
  assign n8244 = ~n8526 | ~INSTQUEUE_REG_15__6__SCAN_IN;
  assign n8243 = ~n8910 | ~INSTQUEUE_REG_13__6__SCAN_IN;
  assign n8245 = ~n8244 | ~n8243;
  assign n8254 = ~n8246 & ~n8245;
  assign n8248 = ~n8915 | ~INSTQUEUE_REG_11__6__SCAN_IN;
  assign n8247 = ~n8154 | ~INSTQUEUE_REG_14__6__SCAN_IN;
  assign n8252 = ~n8248 | ~n8247;
  assign n8250 = ~n7006 | ~INSTQUEUE_REG_7__6__SCAN_IN;
  assign n8249 = ~n8420 | ~INSTQUEUE_REG_5__6__SCAN_IN;
  assign n8251 = ~n8250 | ~n8249;
  assign n8253 = ~n8252 & ~n8251;
  assign n8255 = ~n8254 | ~n8253;
  assign n8264 = ~n8256 & ~n8255;
  assign n8258 = ~n8586 | ~INSTQUEUE_REG_8__6__SCAN_IN;
  assign n8257 = ~n8279 | ~INSTQUEUE_REG_1__6__SCAN_IN;
  assign n8262 = ~n8258 | ~n8257;
  assign n8260 = ~n8151 | ~INSTQUEUE_REG_4__6__SCAN_IN;
  assign n8259 = ~n7807 | ~INSTQUEUE_REG_2__6__SCAN_IN;
  assign n8261 = ~n8260 | ~n8259;
  assign n8263 = ~n8262 & ~n8261;
  assign n8265 = n8264 & n8263;
  assign n10135 = ~n8267 | ~n8266;
  assign n10590 = PHYADDRPOINTER_REG_15__SCAN_IN ^ n8343;
  assign n8272 = n10590 & n7837;
  assign n8270 = ~n7864 | ~EAX_REG_15__SCAN_IN;
  assign n8269 = ~n9446 | ~PHYADDRPOINTER_REG_15__SCAN_IN;
  assign n8271 = ~n8270 | ~n8269;
  assign n8307 = ~n8272 & ~n8271;
  assign n8274 = ~n8587 | ~INSTQUEUE_REG_8__7__SCAN_IN;
  assign n8273 = ~n8526 | ~INSTQUEUE_REG_15__7__SCAN_IN;
  assign n8278 = ~n8274 | ~n8273;
  assign n8276 = ~n7009 | ~INSTQUEUE_REG_0__7__SCAN_IN;
  assign n8275 = ~n8892 | ~INSTQUEUE_REG_6__7__SCAN_IN;
  assign n8277 = ~n8276 | ~n8275;
  assign n8295 = n8278 | n8277;
  assign n8281 = ~n8854 | ~INSTQUEUE_REG_10__7__SCAN_IN;
  assign n8280 = ~n8279 | ~INSTQUEUE_REG_1__7__SCAN_IN;
  assign n8285 = ~n8281 | ~n8280;
  assign n8283 = ~n8906 | ~INSTQUEUE_REG_12__7__SCAN_IN;
  assign n8282 = ~n8420 | ~INSTQUEUE_REG_5__7__SCAN_IN;
  assign n8284 = ~n8283 | ~n8282;
  assign n8293 = ~n8285 & ~n8284;
  assign n8287 = ~n8915 | ~INSTQUEUE_REG_11__7__SCAN_IN;
  assign n8286 = ~n8151 | ~INSTQUEUE_REG_4__7__SCAN_IN;
  assign n8291 = ~n8287 | ~n8286;
  assign n8289 = ~n8910 | ~INSTQUEUE_REG_13__7__SCAN_IN;
  assign n8288 = ~n8154 | ~INSTQUEUE_REG_14__7__SCAN_IN;
  assign n8290 = ~n8289 | ~n8288;
  assign n8292 = ~n8291 & ~n8290;
  assign n8294 = ~n8293 | ~n8292;
  assign n8303 = ~n8295 & ~n8294;
  assign n8297 = ~n9398 | ~INSTQUEUE_REG_9__7__SCAN_IN;
  assign n8296 = ~n7807 | ~INSTQUEUE_REG_2__7__SCAN_IN;
  assign n8301 = ~n8297 | ~n8296;
  assign n8299 = ~n9408 | ~INSTQUEUE_REG_7__7__SCAN_IN;
  assign n8298 = ~n8899 | ~INSTQUEUE_REG_3__7__SCAN_IN;
  assign n8300 = ~n8299 | ~n8298;
  assign n8302 = ~n8301 & ~n8300;
  assign n8304 = n8303 & n8302;
  assign n8311 = ~n13311 | ~n11918;
  assign n8313 = ~n7009 | ~INSTQUEUE_REG_1__0__SCAN_IN;
  assign n8312 = ~n8907 | ~INSTQUEUE_REG_2__0__SCAN_IN;
  assign n8317 = ~n8313 | ~n8312;
  assign n8315 = ~n9408 | ~INSTQUEUE_REG_8__0__SCAN_IN;
  assign n8314 = ~n8910 | ~INSTQUEUE_REG_14__0__SCAN_IN;
  assign n8316 = ~n8315 | ~n8314;
  assign n8325 = ~n8317 & ~n8316;
  assign n8319 = ~n8526 | ~INSTQUEUE_REG_0__0__SCAN_IN;
  assign n8318 = ~n8899 | ~INSTQUEUE_REG_4__0__SCAN_IN;
  assign n8323 = ~n8319 | ~n8318;
  assign n8321 = ~n8154 | ~INSTQUEUE_REG_15__0__SCAN_IN;
  assign n8320 = ~n8693 | ~INSTQUEUE_REG_6__0__SCAN_IN;
  assign n8322 = ~n8321 | ~n8320;
  assign n8324 = ~n8323 & ~n8322;
  assign n8341 = ~n8325 | ~n8324;
  assign n8327 = ~n8586 | ~INSTQUEUE_REG_9__0__SCAN_IN;
  assign n8326 = ~n8892 | ~INSTQUEUE_REG_7__0__SCAN_IN;
  assign n8331 = ~n8327 | ~n8326;
  assign n8329 = ~n8642 | ~INSTQUEUE_REG_5__0__SCAN_IN;
  assign n8328 = ~n7807 | ~INSTQUEUE_REG_3__0__SCAN_IN;
  assign n8330 = ~n8329 | ~n8328;
  assign n8339 = ~n8331 & ~n8330;
  assign n8333 = ~n8915 | ~INSTQUEUE_REG_12__0__SCAN_IN;
  assign n8332 = ~n8906 | ~INSTQUEUE_REG_13__0__SCAN_IN;
  assign n8337 = ~n8333 | ~n8332;
  assign n8335 = ~n9398 | ~INSTQUEUE_REG_10__0__SCAN_IN;
  assign n8334 = ~n8854 | ~INSTQUEUE_REG_11__0__SCAN_IN;
  assign n8336 = ~n8335 | ~n8334;
  assign n8338 = ~n8337 & ~n8336;
  assign n8340 = ~n8339 | ~n8338;
  assign n8342 = n8341 | n8340;
  assign n8349 = ~n9435 | ~n8342;
  assign n8347 = ~n7864 | ~EAX_REG_16__SCAN_IN;
  assign n8345 = ~n9446 | ~PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n10559 = ~PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n10571 = n10559 ^ n8351;
  assign n8344 = ~n8929 | ~n10571;
  assign n8346 = n8345 & n8344;
  assign n8348 = n8347 & n8346;
  assign n10555 = PHYADDRPOINTER_REG_17__SCAN_IN ^ ~n8392;
  assign n8390 = ~n10555 | ~n8929;
  assign n8353 = ~n9398 | ~INSTQUEUE_REG_10__1__SCAN_IN;
  assign n8352 = ~n8642 | ~INSTQUEUE_REG_5__1__SCAN_IN;
  assign n8357 = ~n8353 | ~n8352;
  assign n8355 = ~n8906 | ~INSTQUEUE_REG_13__1__SCAN_IN;
  assign n8354 = ~n8899 | ~INSTQUEUE_REG_4__1__SCAN_IN;
  assign n8356 = ~n8355 | ~n8354;
  assign n8365 = ~n8357 & ~n8356;
  assign n8359 = ~n8892 | ~INSTQUEUE_REG_7__1__SCAN_IN;
  assign n8358 = ~n8154 | ~INSTQUEUE_REG_15__1__SCAN_IN;
  assign n8363 = ~n8359 | ~n8358;
  assign n8361 = ~n8587 | ~INSTQUEUE_REG_9__1__SCAN_IN;
  assign n8360 = ~n7807 | ~INSTQUEUE_REG_3__1__SCAN_IN;
  assign n8362 = ~n8361 | ~n8360;
  assign n8364 = ~n8363 & ~n8362;
  assign n8381 = ~n8365 | ~n8364;
  assign n8367 = ~n9408 | ~INSTQUEUE_REG_8__1__SCAN_IN;
  assign n8366 = ~n8907 | ~INSTQUEUE_REG_2__1__SCAN_IN;
  assign n8371 = ~n8367 | ~n8366;
  assign n8369 = ~n8854 | ~INSTQUEUE_REG_11__1__SCAN_IN;
  assign n8368 = ~n8693 | ~INSTQUEUE_REG_6__1__SCAN_IN;
  assign n8370 = ~n8369 | ~n8368;
  assign n8379 = ~n8371 & ~n8370;
  assign n8373 = ~n7469 | ~INSTQUEUE_REG_1__1__SCAN_IN;
  assign n8372 = ~n8910 | ~INSTQUEUE_REG_14__1__SCAN_IN;
  assign n8377 = ~n8373 | ~n8372;
  assign n8375 = ~n8915 | ~INSTQUEUE_REG_12__1__SCAN_IN;
  assign n8374 = ~n8526 | ~INSTQUEUE_REG_0__1__SCAN_IN;
  assign n8376 = ~n8375 | ~n8374;
  assign n8378 = ~n8377 & ~n8376;
  assign n8380 = ~n8379 | ~n8378;
  assign n8382 = ~n8381 & ~n8380;
  assign n8386 = ~n8666 & ~n8382;
  assign n8383 = ~n8880 | ~EAX_REG_17__SCAN_IN;
  assign n8385 = ~n8384 | ~n8383;
  assign n8388 = ~n8386 & ~n8385;
  assign n8387 = ~n11983 | ~PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n8389 = ~n8388 | ~n8387;
  assign n10093 = ~n8390 | ~n8389;
  assign n10537 = PHYADDRPOINTER_REG_18__SCAN_IN ^ ~n8437;
  assign n8393 = ~n10537;
  assign n8436 = ~n8393 | ~n8929;
  assign n8394 = ~INSTQUEUE_REG_8__2__SCAN_IN;
  assign n8396 = ~n7880 & ~n8394;
  assign n8395 = ~n8562 & ~n7596;
  assign n8403 = ~n8396 & ~n8395;
  assign n8397 = ~INSTQUEUE_REG_10__2__SCAN_IN;
  assign n8401 = ~n7692 & ~n8397;
  assign n8398 = ~INSTQUEUE_REG_3__2__SCAN_IN;
  assign n8400 = ~n8399 & ~n8398;
  assign n8402 = ~n8401 & ~n8400;
  assign n8419 = ~n8403 | ~n8402;
  assign n8405 = ~n8899 | ~INSTQUEUE_REG_4__2__SCAN_IN;
  assign n8404 = ~n8907 | ~INSTQUEUE_REG_2__2__SCAN_IN;
  assign n8409 = ~n8405 | ~n8404;
  assign n8407 = ~n8906 | ~INSTQUEUE_REG_13__2__SCAN_IN;
  assign n8406 = ~n8587 | ~INSTQUEUE_REG_9__2__SCAN_IN;
  assign n8408 = ~n8407 | ~n8406;
  assign n8417 = ~n8409 & ~n8408;
  assign n8411 = ~n8910 | ~INSTQUEUE_REG_14__2__SCAN_IN;
  assign n8410 = ~n8854 | ~INSTQUEUE_REG_11__2__SCAN_IN;
  assign n8415 = ~n8411 | ~n8410;
  assign n8413 = ~n7009 | ~INSTQUEUE_REG_1__2__SCAN_IN;
  assign n8412 = ~n8892 | ~INSTQUEUE_REG_7__2__SCAN_IN;
  assign n8414 = ~n8413 | ~n8412;
  assign n8416 = ~n8415 & ~n8414;
  assign n8418 = ~n8417 | ~n8416;
  assign n8428 = ~n8419 & ~n8418;
  assign n8422 = ~n8567 | ~INSTQUEUE_REG_5__2__SCAN_IN;
  assign n8420 = ~n6997;
  assign n8421 = ~n8693 | ~INSTQUEUE_REG_6__2__SCAN_IN;
  assign n8426 = ~n8422 | ~n8421;
  assign n8424 = ~n8915 | ~INSTQUEUE_REG_12__2__SCAN_IN;
  assign n8423 = ~n8154 | ~INSTQUEUE_REG_15__2__SCAN_IN;
  assign n8425 = ~n8424 | ~n8423;
  assign n8427 = ~n8426 & ~n8425;
  assign n8429 = ~n8428 | ~n8427;
  assign n8434 = ~n9435 | ~n8429;
  assign n8432 = ~n7864 | ~EAX_REG_18__SCAN_IN;
  assign n8430 = ~PHYADDRPOINTER_REG_18__SCAN_IN & ~n13100;
  assign n8431 = STATE2_REG_2__SCAN_IN | n8430;
  assign n8433 = n8432 & n8431;
  assign n8435 = ~n8434 | ~n8433;
  assign n10061 = n8515 ^ ~PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n8476 = ~n10061 | ~n8929;
  assign n8438 = ~PHYADDRPOINTER_REG_19__SCAN_IN | ~n11983;
  assign n8472 = ~n8384 | ~n8438;
  assign n8440 = ~n8906 | ~INSTQUEUE_REG_13__3__SCAN_IN;
  assign n8439 = ~n8154 | ~INSTQUEUE_REG_15__3__SCAN_IN;
  assign n8444 = ~n8440 | ~n8439;
  assign n8442 = ~n9408 | ~INSTQUEUE_REG_8__3__SCAN_IN;
  assign n8441 = ~n8910 | ~INSTQUEUE_REG_14__3__SCAN_IN;
  assign n8443 = ~n8442 | ~n8441;
  assign n8452 = ~n8444 & ~n8443;
  assign n8446 = ~n8899 | ~INSTQUEUE_REG_4__3__SCAN_IN;
  assign n8445 = ~n8151 | ~INSTQUEUE_REG_5__3__SCAN_IN;
  assign n8450 = ~n8446 | ~n8445;
  assign n8448 = ~n8526 | ~INSTQUEUE_REG_0__3__SCAN_IN;
  assign n8447 = ~n8892 | ~INSTQUEUE_REG_7__3__SCAN_IN;
  assign n8449 = ~n8448 | ~n8447;
  assign n8451 = ~n8450 & ~n8449;
  assign n8469 = ~n8452 | ~n8451;
  assign n8455 = ~n8453 | ~INSTQUEUE_REG_11__3__SCAN_IN;
  assign n8454 = ~n7807 | ~INSTQUEUE_REG_3__3__SCAN_IN;
  assign n8459 = ~n8455 | ~n8454;
  assign n8457 = ~n8587 | ~INSTQUEUE_REG_9__3__SCAN_IN;
  assign n8456 = ~n8907 | ~INSTQUEUE_REG_2__3__SCAN_IN;
  assign n8458 = ~n8457 | ~n8456;
  assign n8467 = ~n8459 & ~n8458;
  assign n8461 = ~n8915 | ~INSTQUEUE_REG_12__3__SCAN_IN;
  assign n8460 = ~n9398 | ~INSTQUEUE_REG_10__3__SCAN_IN;
  assign n8465 = ~n8461 | ~n8460;
  assign n8463 = ~n7009 | ~INSTQUEUE_REG_1__3__SCAN_IN;
  assign n8462 = ~n8420 | ~INSTQUEUE_REG_6__3__SCAN_IN;
  assign n8464 = ~n8463 | ~n8462;
  assign n8466 = ~n8465 & ~n8464;
  assign n8468 = ~n8467 | ~n8466;
  assign n8470 = ~n8469 & ~n8468;
  assign n8471 = ~n8666 & ~n8470;
  assign n8474 = ~n8472 & ~n8471;
  assign n8473 = ~n8880 | ~EAX_REG_19__SCAN_IN;
  assign n8475 = ~n8474 | ~n8473;
  assign n9765 = ~n8476 | ~n8475;
  assign n8480 = ~n8915 | ~INSTQUEUE_REG_12__4__SCAN_IN;
  assign n8479 = ~n8151 | ~INSTQUEUE_REG_5__4__SCAN_IN;
  assign n8484 = ~n8480 | ~n8479;
  assign n8482 = ~n8906 | ~INSTQUEUE_REG_13__4__SCAN_IN;
  assign n8481 = ~n8526 | ~INSTQUEUE_REG_0__4__SCAN_IN;
  assign n8483 = ~n8482 | ~n8481;
  assign n8500 = n8484 | n8483;
  assign n8486 = ~n9398 | ~INSTQUEUE_REG_10__4__SCAN_IN;
  assign n8485 = ~n7807 | ~INSTQUEUE_REG_3__4__SCAN_IN;
  assign n8490 = ~n8486 | ~n8485;
  assign n8488 = ~n7469 | ~INSTQUEUE_REG_1__4__SCAN_IN;
  assign n8487 = ~n8907 | ~INSTQUEUE_REG_2__4__SCAN_IN;
  assign n8489 = ~n8488 | ~n8487;
  assign n8498 = ~n8490 & ~n8489;
  assign n8492 = ~n8910 | ~INSTQUEUE_REG_14__4__SCAN_IN;
  assign n8491 = ~n8854 | ~INSTQUEUE_REG_11__4__SCAN_IN;
  assign n8496 = ~n8492 | ~n8491;
  assign n8494 = ~n8899 | ~INSTQUEUE_REG_4__4__SCAN_IN;
  assign n8493 = ~n8420 | ~INSTQUEUE_REG_6__4__SCAN_IN;
  assign n8495 = ~n8494 | ~n8493;
  assign n8497 = ~n8496 & ~n8495;
  assign n8499 = ~n8498 | ~n8497;
  assign n8508 = ~n8500 & ~n8499;
  assign n8502 = ~n9408 | ~INSTQUEUE_REG_8__4__SCAN_IN;
  assign n8501 = ~n8586 | ~INSTQUEUE_REG_9__4__SCAN_IN;
  assign n8506 = ~n8502 | ~n8501;
  assign n8504 = ~n8892 | ~INSTQUEUE_REG_7__4__SCAN_IN;
  assign n8503 = ~n7014 | ~INSTQUEUE_REG_15__4__SCAN_IN;
  assign n8505 = ~n8504 | ~n8503;
  assign n8507 = ~n8506 & ~n8505;
  assign n8509 = ~n8508 | ~n8507;
  assign n8514 = ~n9435 | ~n8509;
  assign n8512 = ~n8880 | ~EAX_REG_20__SCAN_IN;
  assign n8510 = ~PHYADDRPOINTER_REG_20__SCAN_IN & ~n13100;
  assign n8511 = STATE2_REG_2__SCAN_IN | n8510;
  assign n8513 = n8512 & n8511;
  assign n8518 = ~n8514 | ~n8513;
  assign n8516 = ~n8557;
  assign n10048 = PHYADDRPOINTER_REG_20__SCAN_IN ^ ~n8516;
  assign n8517 = ~n10048 | ~n7837;
  assign n9744 = ~n8518 | ~n8517;
  assign n8519 = ~PHYADDRPOINTER_REG_21__SCAN_IN | ~n11983;
  assign n8554 = ~n8384 | ~n8519;
  assign n8521 = ~n7807 | ~INSTQUEUE_REG_3__5__SCAN_IN;
  assign n8520 = ~n7014 | ~INSTQUEUE_REG_15__5__SCAN_IN;
  assign n8525 = ~n8521 | ~n8520;
  assign n8523 = ~n8587 | ~INSTQUEUE_REG_9__5__SCAN_IN;
  assign n8522 = ~n8892 | ~INSTQUEUE_REG_7__5__SCAN_IN;
  assign n8524 = ~n8523 | ~n8522;
  assign n8534 = ~n8525 & ~n8524;
  assign n8528 = ~n8526 | ~INSTQUEUE_REG_0__5__SCAN_IN;
  assign n8527 = ~n8899 | ~INSTQUEUE_REG_4__5__SCAN_IN;
  assign n8532 = ~n8528 | ~n8527;
  assign n8530 = ~n8906 | ~INSTQUEUE_REG_13__5__SCAN_IN;
  assign n8529 = ~n7009 | ~INSTQUEUE_REG_1__5__SCAN_IN;
  assign n8531 = ~n8530 | ~n8529;
  assign n8533 = ~n8532 & ~n8531;
  assign n8551 = ~n8534 | ~n8533;
  assign n8536 = ~n9398 | ~INSTQUEUE_REG_10__5__SCAN_IN;
  assign n8535 = ~n8151 | ~INSTQUEUE_REG_5__5__SCAN_IN;
  assign n8541 = ~n8536 | ~n8535;
  assign n8539 = ~n8915 | ~INSTQUEUE_REG_12__5__SCAN_IN;
  assign n8907 = ~n8537;
  assign n8538 = ~n8907 | ~INSTQUEUE_REG_2__5__SCAN_IN;
  assign n8540 = ~n8539 | ~n8538;
  assign n8549 = ~n8541 & ~n8540;
  assign n8543 = ~n9408 | ~INSTQUEUE_REG_8__5__SCAN_IN;
  assign n8542 = ~n8693 | ~INSTQUEUE_REG_6__5__SCAN_IN;
  assign n8547 = ~n8543 | ~n8542;
  assign n8545 = ~n8910 | ~INSTQUEUE_REG_14__5__SCAN_IN;
  assign n8544 = ~n8854 | ~INSTQUEUE_REG_11__5__SCAN_IN;
  assign n8546 = ~n8545 | ~n8544;
  assign n8548 = ~n8547 & ~n8546;
  assign n8550 = ~n8549 | ~n8548;
  assign n8552 = ~n8551 & ~n8550;
  assign n8553 = ~n8666 & ~n8552;
  assign n8556 = ~n8554 & ~n8553;
  assign n8555 = ~n8880 | ~EAX_REG_21__SCAN_IN;
  assign n8559 = ~n8556 | ~n8555;
  assign n10034 = PHYADDRPOINTER_REG_21__SCAN_IN ^ ~n8600;
  assign n8558 = ~n10034 | ~n7837;
  assign n8561 = ~n8854 | ~INSTQUEUE_REG_11__6__SCAN_IN;
  assign n8560 = ~n8892 | ~INSTQUEUE_REG_7__6__SCAN_IN;
  assign n8566 = ~n8561 | ~n8560;
  assign n8564 = ~n8526 | ~INSTQUEUE_REG_0__6__SCAN_IN;
  assign n8563 = ~n8693 | ~INSTQUEUE_REG_6__6__SCAN_IN;
  assign n8565 = ~n8564 | ~n8563;
  assign n8583 = n8566 | n8565;
  assign n8569 = ~n8567 | ~INSTQUEUE_REG_5__6__SCAN_IN;
  assign n8568 = ~n8907 | ~INSTQUEUE_REG_2__6__SCAN_IN;
  assign n8573 = ~n8569 | ~n8568;
  assign n8571 = ~n8915 | ~INSTQUEUE_REG_12__6__SCAN_IN;
  assign n8570 = ~n8899 | ~INSTQUEUE_REG_4__6__SCAN_IN;
  assign n8572 = ~n8571 | ~n8570;
  assign n8581 = ~n8573 & ~n8572;
  assign n8575 = ~n8906 | ~INSTQUEUE_REG_13__6__SCAN_IN;
  assign n8574 = ~n9398 | ~INSTQUEUE_REG_10__6__SCAN_IN;
  assign n8579 = ~n8575 | ~n8574;
  assign n8577 = ~n7009 | ~INSTQUEUE_REG_1__6__SCAN_IN;
  assign n8576 = ~n8910 | ~INSTQUEUE_REG_14__6__SCAN_IN;
  assign n8578 = ~n8577 | ~n8576;
  assign n8580 = ~n8579 & ~n8578;
  assign n8582 = ~n8581 | ~n8580;
  assign n8593 = ~n8583 & ~n8582;
  assign n8585 = ~n7006 | ~INSTQUEUE_REG_8__6__SCAN_IN;
  assign n8584 = ~n7807 | ~INSTQUEUE_REG_3__6__SCAN_IN;
  assign n8591 = ~n8585 | ~n8584;
  assign n8589 = ~n8587 | ~INSTQUEUE_REG_9__6__SCAN_IN;
  assign n8588 = ~n8154 | ~INSTQUEUE_REG_15__6__SCAN_IN;
  assign n8590 = ~n8589 | ~n8588;
  assign n8592 = ~n8591 & ~n8590;
  assign n8594 = ~n8593 | ~n8592;
  assign n8599 = ~n9435 | ~n8594;
  assign n8597 = ~n8880 | ~EAX_REG_22__SCAN_IN;
  assign n8595 = ~PHYADDRPOINTER_REG_22__SCAN_IN & ~n13100;
  assign n8596 = STATE2_REG_2__SCAN_IN | n8595;
  assign n8598 = n8597 & n8596;
  assign n8603 = ~n8599 | ~n8598;
  assign n8601 = ~n8672;
  assign n10022 = PHYADDRPOINTER_REG_22__SCAN_IN ^ ~n8601;
  assign n8602 = ~n10022 | ~n7837;
  assign n8605 = ~n8526 | ~INSTQUEUE_REG_1__0__SCAN_IN;
  assign n8604 = ~n8151 | ~INSTQUEUE_REG_6__0__SCAN_IN;
  assign n8609 = ~n8605 | ~n8604;
  assign n8607 = ~n8854 | ~INSTQUEUE_REG_12__0__SCAN_IN;
  assign n8606 = ~n8420 | ~INSTQUEUE_REG_7__0__SCAN_IN;
  assign n8608 = ~n8607 | ~n8606;
  assign n8617 = ~n8609 & ~n8608;
  assign n8611 = ~n8915 | ~INSTQUEUE_REG_13__0__SCAN_IN;
  assign n8610 = ~n7009 | ~INSTQUEUE_REG_2__0__SCAN_IN;
  assign n8615 = ~n8611 | ~n8610;
  assign n8613 = ~n9408 | ~INSTQUEUE_REG_9__0__SCAN_IN;
  assign n8612 = ~n8154 | ~INSTQUEUE_REG_0__0__SCAN_IN;
  assign n8614 = ~n8613 | ~n8612;
  assign n8616 = ~n8615 & ~n8614;
  assign n8633 = ~n8617 | ~n8616;
  assign n8619 = ~n8899 | ~INSTQUEUE_REG_5__0__SCAN_IN;
  assign n8618 = ~n8907 | ~INSTQUEUE_REG_3__0__SCAN_IN;
  assign n8623 = ~n8619 | ~n8618;
  assign n8621 = ~n8587 | ~INSTQUEUE_REG_10__0__SCAN_IN;
  assign n8620 = ~n8910 | ~INSTQUEUE_REG_15__0__SCAN_IN;
  assign n8622 = ~n8621 | ~n8620;
  assign n8631 = ~n8623 & ~n8622;
  assign n8625 = ~n8906 | ~INSTQUEUE_REG_14__0__SCAN_IN;
  assign n8624 = ~n8892 | ~INSTQUEUE_REG_8__0__SCAN_IN;
  assign n8629 = ~n8625 | ~n8624;
  assign n8627 = ~n9398 | ~INSTQUEUE_REG_11__0__SCAN_IN;
  assign n8626 = ~n7807 | ~INSTQUEUE_REG_4__0__SCAN_IN;
  assign n8628 = ~n8627 | ~n8626;
  assign n8630 = ~n8629 & ~n8628;
  assign n8632 = ~n8631 | ~n8630;
  assign n8677 = ~n8633 & ~n8632;
  assign n8635 = ~n8906 | ~INSTQUEUE_REG_13__7__SCAN_IN;
  assign n8634 = ~n8154 | ~INSTQUEUE_REG_15__7__SCAN_IN;
  assign n8639 = ~n8635 | ~n8634;
  assign n8637 = ~n8915 | ~INSTQUEUE_REG_12__7__SCAN_IN;
  assign n8636 = ~n8892 | ~INSTQUEUE_REG_7__7__SCAN_IN;
  assign n8638 = ~n8637 | ~n8636;
  assign n8648 = ~n8639 & ~n8638;
  assign n8641 = ~n7009 | ~INSTQUEUE_REG_1__7__SCAN_IN;
  assign n8640 = ~n9398 | ~INSTQUEUE_REG_10__7__SCAN_IN;
  assign n8646 = ~n8641 | ~n8640;
  assign n8644 = ~n8910 | ~INSTQUEUE_REG_14__7__SCAN_IN;
  assign n8643 = ~n8642 | ~INSTQUEUE_REG_5__7__SCAN_IN;
  assign n8645 = ~n8644 | ~n8643;
  assign n8647 = ~n8646 & ~n8645;
  assign n8664 = ~n8648 | ~n8647;
  assign n8650 = ~n8526 | ~INSTQUEUE_REG_0__7__SCAN_IN;
  assign n8649 = ~n8899 | ~INSTQUEUE_REG_4__7__SCAN_IN;
  assign n8654 = ~n8650 | ~n8649;
  assign n8652 = ~n8587 | ~INSTQUEUE_REG_9__7__SCAN_IN;
  assign n8651 = ~n8693 | ~INSTQUEUE_REG_6__7__SCAN_IN;
  assign n8653 = ~n8652 | ~n8651;
  assign n8662 = ~n8654 & ~n8653;
  assign n8656 = ~n9408 | ~INSTQUEUE_REG_8__7__SCAN_IN;
  assign n8655 = ~n8854 | ~INSTQUEUE_REG_11__7__SCAN_IN;
  assign n8660 = ~n8656 | ~n8655;
  assign n8658 = ~n7807 | ~INSTQUEUE_REG_3__7__SCAN_IN;
  assign n8657 = ~n8907 | ~INSTQUEUE_REG_2__7__SCAN_IN;
  assign n8659 = ~n8658 | ~n8657;
  assign n8661 = ~n8660 & ~n8659;
  assign n8663 = ~n8662 | ~n8661;
  assign n8678 = ~n8664 & ~n8663;
  assign n8665 = n8677 ^ ~n8678;
  assign n8670 = ~n8666 & ~n8665;
  assign n8668 = ~n7864 | ~EAX_REG_23__SCAN_IN;
  assign n8667 = ~PHYADDRPOINTER_REG_23__SCAN_IN | ~n11983;
  assign n8669 = ~n8668 | ~n8667;
  assign n8671 = ~n8670 & ~n8669;
  assign n8674 = ~n8671 | ~n8384;
  assign n10010 = PHYADDRPOINTER_REG_23__SCAN_IN ^ ~n8711;
  assign n8673 = ~n10010 | ~n7837;
  assign n9684 = ~n8674 | ~n8673;
  assign n8718 = n8678 | n8677;
  assign n8680 = ~n9398 | ~INSTQUEUE_REG_11__1__SCAN_IN;
  assign n8679 = ~n8154 | ~INSTQUEUE_REG_0__1__SCAN_IN;
  assign n8684 = ~n8680 | ~n8679;
  assign n8682 = ~n8587 | ~INSTQUEUE_REG_10__1__SCAN_IN;
  assign n8681 = ~n8892 | ~INSTQUEUE_REG_8__1__SCAN_IN;
  assign n8683 = ~n8682 | ~n8681;
  assign n8692 = ~n8684 & ~n8683;
  assign n8686 = ~n9408 | ~INSTQUEUE_REG_9__1__SCAN_IN;
  assign n8685 = ~n8899 | ~INSTQUEUE_REG_5__1__SCAN_IN;
  assign n8690 = ~n8686 | ~n8685;
  assign n8688 = ~n8915 | ~INSTQUEUE_REG_13__1__SCAN_IN;
  assign n8687 = ~n8151 | ~INSTQUEUE_REG_6__1__SCAN_IN;
  assign n8689 = ~n8688 | ~n8687;
  assign n8691 = ~n8690 & ~n8689;
  assign n8709 = ~n8692 | ~n8691;
  assign n8695 = ~n7009 | ~INSTQUEUE_REG_2__1__SCAN_IN;
  assign n8694 = ~n8420 | ~INSTQUEUE_REG_7__1__SCAN_IN;
  assign n8699 = ~n8695 | ~n8694;
  assign n8697 = ~n8906 | ~INSTQUEUE_REG_14__1__SCAN_IN;
  assign n8696 = ~n8910 | ~INSTQUEUE_REG_15__1__SCAN_IN;
  assign n8698 = ~n8697 | ~n8696;
  assign n8707 = ~n8699 & ~n8698;
  assign n8701 = ~n8854 | ~INSTQUEUE_REG_12__1__SCAN_IN;
  assign n8700 = ~n7807 | ~INSTQUEUE_REG_4__1__SCAN_IN;
  assign n8705 = ~n8701 | ~n8700;
  assign n8703 = ~n8526 | ~INSTQUEUE_REG_1__1__SCAN_IN;
  assign n8702 = ~n8907 | ~INSTQUEUE_REG_3__1__SCAN_IN;
  assign n8704 = ~n8703 | ~n8702;
  assign n8706 = ~n8705 & ~n8704;
  assign n8708 = ~n8707 | ~n8706;
  assign n8719 = ~n8709 & ~n8708;
  assign n8710 = n8718 ^ n8719;
  assign n8717 = ~n8710 | ~n9435;
  assign n8715 = ~n8880 | ~EAX_REG_24__SCAN_IN;
  assign n8713 = ~n9446 | ~PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n9669 = PHYADDRPOINTER_REG_24__SCAN_IN ^ ~n8756;
  assign n8712 = ~n7837 | ~n9669;
  assign n8714 = n8713 & n8712;
  assign n8791 = n8719 | n8718;
  assign n8721 = ~n8915 | ~INSTQUEUE_REG_13__2__SCAN_IN;
  assign n8720 = ~n8154 | ~INSTQUEUE_REG_0__2__SCAN_IN;
  assign n8725 = ~n8721 | ~n8720;
  assign n8723 = ~n9408 | ~INSTQUEUE_REG_9__2__SCAN_IN;
  assign n8722 = ~n8899 | ~INSTQUEUE_REG_5__2__SCAN_IN;
  assign n8724 = ~n8723 | ~n8722;
  assign n8733 = ~n8725 & ~n8724;
  assign n8727 = ~n8910 | ~INSTQUEUE_REG_15__2__SCAN_IN;
  assign n8726 = ~n8907 | ~INSTQUEUE_REG_3__2__SCAN_IN;
  assign n8731 = ~n8727 | ~n8726;
  assign n8729 = ~n8892 | ~INSTQUEUE_REG_8__2__SCAN_IN;
  assign n8728 = ~n8151 | ~INSTQUEUE_REG_6__2__SCAN_IN;
  assign n8730 = ~n8729 | ~n8728;
  assign n8732 = ~n8731 & ~n8730;
  assign n8749 = ~n8733 | ~n8732;
  assign n8735 = ~n8526 | ~INSTQUEUE_REG_1__2__SCAN_IN;
  assign n8734 = ~n8854 | ~INSTQUEUE_REG_12__2__SCAN_IN;
  assign n8739 = ~n8735 | ~n8734;
  assign n8737 = ~n8906 | ~INSTQUEUE_REG_14__2__SCAN_IN;
  assign n8736 = ~n8587 | ~INSTQUEUE_REG_10__2__SCAN_IN;
  assign n8738 = ~n8737 | ~n8736;
  assign n8747 = ~n8739 & ~n8738;
  assign n8741 = ~n7009 | ~INSTQUEUE_REG_2__2__SCAN_IN;
  assign n8740 = ~n8420 | ~INSTQUEUE_REG_7__2__SCAN_IN;
  assign n8745 = ~n8741 | ~n8740;
  assign n8743 = ~n9398 | ~INSTQUEUE_REG_11__2__SCAN_IN;
  assign n8742 = ~n7807 | ~INSTQUEUE_REG_4__2__SCAN_IN;
  assign n8744 = ~n8743 | ~n8742;
  assign n8746 = ~n8745 & ~n8744;
  assign n8748 = ~n8747 | ~n8746;
  assign n8792 = ~n8749 & ~n8748;
  assign n8750 = n8791 ^ n8792;
  assign n8755 = ~n8750 | ~n9435;
  assign n8752 = ~n8880 | ~EAX_REG_25__SCAN_IN;
  assign n8751 = ~PHYADDRPOINTER_REG_25__SCAN_IN | ~n11983;
  assign n8753 = ~n8752 | ~n8751;
  assign n8754 = ~n8753 & ~n8929;
  assign n8758 = ~n8755 | ~n8754;
  assign n9990 = PHYADDRPOINTER_REG_25__SCAN_IN ^ ~n8760;
  assign n8757 = ~n9990 | ~n7837;
  assign n8759 = ~PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n9636 = ~PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n9977 = n8839 ^ ~n9636;
  assign n8800 = ~n9977 | ~n8929;
  assign n8762 = ~n8910 | ~INSTQUEUE_REG_15__3__SCAN_IN;
  assign n8761 = ~n8854 | ~INSTQUEUE_REG_12__3__SCAN_IN;
  assign n8766 = ~n8762 | ~n8761;
  assign n8764 = ~n9408 | ~INSTQUEUE_REG_9__3__SCAN_IN;
  assign n8763 = ~n7469 | ~INSTQUEUE_REG_2__3__SCAN_IN;
  assign n8765 = ~n8764 | ~n8763;
  assign n8774 = ~n8766 & ~n8765;
  assign n8768 = ~n9398 | ~INSTQUEUE_REG_11__3__SCAN_IN;
  assign n8767 = ~n7807 | ~INSTQUEUE_REG_4__3__SCAN_IN;
  assign n8772 = ~n8768 | ~n8767;
  assign n8770 = ~n8899 | ~INSTQUEUE_REG_5__3__SCAN_IN;
  assign n8769 = ~n8693 | ~INSTQUEUE_REG_7__3__SCAN_IN;
  assign n8771 = ~n8770 | ~n8769;
  assign n8773 = ~n8772 & ~n8771;
  assign n8790 = ~n8774 | ~n8773;
  assign n8776 = ~n8151 | ~INSTQUEUE_REG_6__3__SCAN_IN;
  assign n8775 = ~n8907 | ~INSTQUEUE_REG_3__3__SCAN_IN;
  assign n8780 = ~n8776 | ~n8775;
  assign n8778 = ~n8915 | ~INSTQUEUE_REG_13__3__SCAN_IN;
  assign n8777 = ~n8587 | ~INSTQUEUE_REG_10__3__SCAN_IN;
  assign n8779 = ~n8778 | ~n8777;
  assign n8788 = ~n8780 & ~n8779;
  assign n8782 = ~n8906 | ~INSTQUEUE_REG_14__3__SCAN_IN;
  assign n8781 = ~n8892 | ~INSTQUEUE_REG_8__3__SCAN_IN;
  assign n8786 = ~n8782 | ~n8781;
  assign n8784 = ~n8526 | ~INSTQUEUE_REG_1__3__SCAN_IN;
  assign n8783 = ~n8154 | ~INSTQUEUE_REG_0__3__SCAN_IN;
  assign n8785 = ~n8784 | ~n8783;
  assign n8787 = ~n8786 & ~n8785;
  assign n8789 = ~n8788 | ~n8787;
  assign n8802 = ~n8790 & ~n8789;
  assign n8793 = n8802 ^ n8801;
  assign n8798 = ~n8793 | ~n9435;
  assign n8796 = ~n8880 | ~EAX_REG_26__SCAN_IN;
  assign n8794 = PHYADDRPOINTER_REG_26__SCAN_IN & n11983;
  assign n8795 = ~n8929 & ~n8794;
  assign n8797 = n8796 & n8795;
  assign n8799 = ~n8798 | ~n8797;
  assign n8804 = ~n7807 | ~INSTQUEUE_REG_4__4__SCAN_IN;
  assign n8803 = ~n8420 | ~INSTQUEUE_REG_7__4__SCAN_IN;
  assign n8808 = ~n8804 | ~n8803;
  assign n8806 = ~n8915 | ~INSTQUEUE_REG_13__4__SCAN_IN;
  assign n8805 = ~n8892 | ~INSTQUEUE_REG_8__4__SCAN_IN;
  assign n8807 = ~n8806 | ~n8805;
  assign n8816 = ~n8808 & ~n8807;
  assign n8810 = ~n8906 | ~INSTQUEUE_REG_14__4__SCAN_IN;
  assign n8809 = ~n8151 | ~INSTQUEUE_REG_6__4__SCAN_IN;
  assign n8814 = ~n8810 | ~n8809;
  assign n8812 = ~n8910 | ~INSTQUEUE_REG_15__4__SCAN_IN;
  assign n8811 = ~n8907 | ~INSTQUEUE_REG_3__4__SCAN_IN;
  assign n8813 = ~n8812 | ~n8811;
  assign n8815 = ~n8814 & ~n8813;
  assign n8832 = ~n8816 | ~n8815;
  assign n8818 = ~n7009 | ~INSTQUEUE_REG_2__4__SCAN_IN;
  assign n8817 = ~n8899 | ~INSTQUEUE_REG_5__4__SCAN_IN;
  assign n8822 = ~n8818 | ~n8817;
  assign n8820 = ~n8526 | ~INSTQUEUE_REG_1__4__SCAN_IN;
  assign n8819 = ~n8154 | ~INSTQUEUE_REG_0__4__SCAN_IN;
  assign n8821 = ~n8820 | ~n8819;
  assign n8830 = ~n8822 & ~n8821;
  assign n8824 = ~n9398 | ~INSTQUEUE_REG_11__4__SCAN_IN;
  assign n8823 = ~n8854 | ~INSTQUEUE_REG_12__4__SCAN_IN;
  assign n8828 = ~n8824 | ~n8823;
  assign n8826 = ~n9408 | ~INSTQUEUE_REG_9__4__SCAN_IN;
  assign n8825 = ~n8586 | ~INSTQUEUE_REG_10__4__SCAN_IN;
  assign n8827 = ~n8826 | ~n8825;
  assign n8829 = ~n8828 & ~n8827;
  assign n8831 = ~n8830 | ~n8829;
  assign n8878 = ~n8832 & ~n8831;
  assign n8833 = n8877 ^ n8878;
  assign n8838 = ~n8833 | ~n9435;
  assign n8835 = ~n8880 | ~EAX_REG_27__SCAN_IN;
  assign n8834 = ~PHYADDRPOINTER_REG_27__SCAN_IN | ~n11983;
  assign n8836 = ~n8835 | ~n8834;
  assign n8837 = ~n8836 & ~n8929;
  assign n8841 = ~n8838 | ~n8837;
  assign n8845 = ~n8839 | ~PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n9965 = PHYADDRPOINTER_REG_27__SCAN_IN ^ ~n8845;
  assign n8840 = ~n9965 | ~n8929;
  assign n9607 = ~n8841 | ~n8840;
  assign n8844 = ~PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n8933 = ~n8845 & ~n8844;
  assign n9949 = n8933 ^ ~PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n8847 = ~n8906 | ~INSTQUEUE_REG_14__5__SCAN_IN;
  assign n8846 = ~n8420 | ~INSTQUEUE_REG_7__5__SCAN_IN;
  assign n8851 = ~n8847 | ~n8846;
  assign n8849 = ~n8899 | ~INSTQUEUE_REG_5__5__SCAN_IN;
  assign n8848 = ~n7807 | ~INSTQUEUE_REG_4__5__SCAN_IN;
  assign n8850 = ~n8849 | ~n8848;
  assign n8860 = ~n8851 & ~n8850;
  assign n8853 = ~n9408 | ~INSTQUEUE_REG_9__5__SCAN_IN;
  assign n8852 = ~n8910 | ~INSTQUEUE_REG_15__5__SCAN_IN;
  assign n8858 = ~n8853 | ~n8852;
  assign n8856 = ~n8915 | ~INSTQUEUE_REG_13__5__SCAN_IN;
  assign n8855 = ~n8854 | ~INSTQUEUE_REG_12__5__SCAN_IN;
  assign n8857 = ~n8856 | ~n8855;
  assign n8859 = ~n8858 & ~n8857;
  assign n8876 = ~n8860 | ~n8859;
  assign n8862 = ~n8151 | ~INSTQUEUE_REG_6__5__SCAN_IN;
  assign n8861 = ~n8154 | ~INSTQUEUE_REG_0__5__SCAN_IN;
  assign n8866 = ~n8862 | ~n8861;
  assign n8864 = ~n7469 | ~INSTQUEUE_REG_2__5__SCAN_IN;
  assign n8863 = ~n8907 | ~INSTQUEUE_REG_3__5__SCAN_IN;
  assign n8865 = ~n8864 | ~n8863;
  assign n8874 = ~n8866 & ~n8865;
  assign n8868 = ~n8586 | ~INSTQUEUE_REG_10__5__SCAN_IN;
  assign n8867 = ~n8526 | ~INSTQUEUE_REG_1__5__SCAN_IN;
  assign n8872 = ~n8868 | ~n8867;
  assign n8870 = ~n9398 | ~INSTQUEUE_REG_11__5__SCAN_IN;
  assign n8869 = ~n8892 | ~INSTQUEUE_REG_8__5__SCAN_IN;
  assign n8871 = ~n8870 | ~n8869;
  assign n8873 = ~n8872 & ~n8871;
  assign n8875 = ~n8874 | ~n8873;
  assign n8889 = ~n8876 & ~n8875;
  assign n8879 = n8889 ^ n8888;
  assign n8885 = ~n8879 | ~n9435;
  assign n8883 = ~n8880 | ~EAX_REG_28__SCAN_IN;
  assign n8881 = PHYADDRPOINTER_REG_28__SCAN_IN & n11983;
  assign n8882 = ~n8929 & ~n8881;
  assign n8884 = n8883 & n8882;
  assign n8886 = ~n8885 | ~n8884;
  assign n9586 = ~n8887 | ~n8886;
  assign n8891 = ~n8854 | ~INSTQUEUE_REG_12__6__SCAN_IN;
  assign n8890 = ~n7807 | ~INSTQUEUE_REG_4__6__SCAN_IN;
  assign n8896 = ~n8891 | ~n8890;
  assign n8894 = ~n8892 | ~INSTQUEUE_REG_8__6__SCAN_IN;
  assign n8893 = ~n8567 | ~INSTQUEUE_REG_6__6__SCAN_IN;
  assign n8895 = ~n8894 | ~n8893;
  assign n8905 = ~n8896 & ~n8895;
  assign n8898 = ~n8526 | ~INSTQUEUE_REG_1__6__SCAN_IN;
  assign n8897 = ~n8154 | ~INSTQUEUE_REG_0__6__SCAN_IN;
  assign n8903 = ~n8898 | ~n8897;
  assign n8901 = ~n8586 | ~INSTQUEUE_REG_10__6__SCAN_IN;
  assign n8900 = ~n8899 | ~INSTQUEUE_REG_5__6__SCAN_IN;
  assign n8902 = ~n8901 | ~n8900;
  assign n8904 = ~n8903 & ~n8902;
  assign n8925 = ~n8905 | ~n8904;
  assign n8909 = ~n8906 | ~INSTQUEUE_REG_14__6__SCAN_IN;
  assign n8908 = ~n8907 | ~INSTQUEUE_REG_3__6__SCAN_IN;
  assign n8914 = ~n8909 | ~n8908;
  assign n8912 = ~n9408 | ~INSTQUEUE_REG_9__6__SCAN_IN;
  assign n8911 = ~n8910 | ~INSTQUEUE_REG_15__6__SCAN_IN;
  assign n8913 = ~n8912 | ~n8911;
  assign n8923 = ~n8914 & ~n8913;
  assign n8917 = ~n8915 | ~INSTQUEUE_REG_13__6__SCAN_IN;
  assign n8916 = ~n9398 | ~INSTQUEUE_REG_11__6__SCAN_IN;
  assign n8921 = ~n8917 | ~n8916;
  assign n8919 = ~n7469 | ~INSTQUEUE_REG_2__6__SCAN_IN;
  assign n8918 = ~n8420 | ~INSTQUEUE_REG_7__6__SCAN_IN;
  assign n8920 = ~n8919 | ~n8918;
  assign n8922 = ~n8921 & ~n8920;
  assign n8924 = ~n8923 | ~n8922;
  assign n9432 = ~n8925 & ~n8924;
  assign n8926 = n9431 ^ n9432;
  assign n8932 = ~n8926 | ~n9435;
  assign n8928 = ~n7864 | ~EAX_REG_29__SCAN_IN;
  assign n8927 = ~PHYADDRPOINTER_REG_29__SCAN_IN | ~n11983;
  assign n8930 = ~n8928 | ~n8927;
  assign n8931 = ~n8930 & ~n8929;
  assign n8935 = n8932 & n8931;
  assign n9397 = ~n8933 | ~PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n9573 = n9397 ^ PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n8934 = ~n9573 & ~n8384;
  assign n8936 = ~n13400 | ~STATEBS16_REG_SCAN_IN;
  assign n8937 = ~STATE2_REG_3__SCAN_IN & ~STATE2_REG_2__SCAN_IN;
  assign n11563 = n8938 | n9085;
  assign n8943 = ~n8939 & ~n9085;
  assign n8941 = ~n13741 | ~n8954;
  assign n8962 = ~n13310 | ~n9210;
  assign n8942 = ~n8941 | ~n8962;
  assign n9326 = INSTADDRPOINTER_REG_0__SCAN_IN & INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n8949 = ~n11577 | ~n9326;
  assign n8945 = n8944 ^ ~n8955;
  assign n8948 = ~n8945 | ~n13741;
  assign n8947 = ~n8946 & ~n11948;
  assign n11562 = n8948 & n8947;
  assign n8950 = n8949 & n11562;
  assign n8953 = ~n11563 | ~n8950;
  assign n11564 = ~n11577 | ~INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n8951 = ~INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n8952 = ~n11564 | ~n8951;
  assign n11555 = ~n11536;
  assign n11535 = ~INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n8965 = n11880 | n9085;
  assign n8959 = n8955 | n8954;
  assign n8957 = ~n8959;
  assign n8956 = ~n8958;
  assign n8960 = ~n8957 | ~n8956;
  assign n8982 = ~n8959 | ~n8958;
  assign n8961 = ~n8960 | ~n8982;
  assign n8963 = ~n8961 | ~n13741;
  assign n8964 = n8963 & n8962;
  assign n8967 = ~n8973 | ~n11537;
  assign n8974 = ~n11536 | ~INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n11747 = ~INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n8966 = n8974 & n11747;
  assign n8972 = ~n8967 | ~n8966;
  assign n8971 = ~n11884 | ~n9109;
  assign n8968 = ~n8981;
  assign n8969 = n8982 ^ ~n8968;
  assign n8970 = ~n8969 | ~n13741;
  assign n11540 = ~n8971 | ~n8970;
  assign n8979 = ~n8972 | ~n11540;
  assign n8977 = n8973 & INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n8975 = ~n11537;
  assign n8976 = ~n8975 | ~n8974;
  assign n8978 = ~n8977 | ~n8976;
  assign n11518 = ~n8979 | ~n8978;
  assign n8984 = ~n8980 & ~n9085;
  assign n8988 = ~n8982 | ~n8981;
  assign n8983 = n8989 ^ n8988;
  assign n9529 = ~n13741;
  assign n8987 = ~n11518 | ~n11519;
  assign n8986 = ~n8985 | ~INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n11508 = ~n8987 | ~n8986;
  assign n8990 = ~n8988;
  assign n8995 = ~n8990 | ~n8989;
  assign n8991 = n8995 ^ ~n8996;
  assign n8992 = ~n8991 | ~n13741;
  assign n11497 = ~n8993 | ~INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n8997 = ~n8995;
  assign n9009 = ~n8997 | ~n8996;
  assign n8998 = n9009 ^ ~n9007;
  assign n8999 = ~n8998 | ~n13741;
  assign n9003 = ~n9001 | ~INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n9000 = n11497 & n9003;
  assign n9008 = ~n9007;
  assign n9019 = n9009 | n9008;
  assign n9010 = n9019 ^ ~n9017;
  assign n9011 = ~n9010 | ~n13741;
  assign n11678 = ~INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n9014 = ~n9013 | ~INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n9016 = n9015 & n9109;
  assign n9018 = ~n13741 | ~n9017;
  assign n9020 = n9019 | n9018;
  assign n9022 = ~n9464 | ~n9020;
  assign n9021 = ~INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n11476 = n9022 ^ ~n9021;
  assign n9023 = ~n9022 | ~INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n9025 = ~n9035 | ~INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n9027 = ~INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n11452 = ~n9464 | ~n9027;
  assign n11616 = ~INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n9028 = ~n9109 | ~INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n11433 = ~n9035 | ~INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n9030 = ~n9029 & ~n9085;
  assign n9031 = ~n9109 | ~INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n9033 = ~n9032 & ~n9031;
  assign n10143 = n9034 | n9033;
  assign n10397 = ~INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n10114 = ~n9035 | ~INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n10117 = ~n9035 | ~INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n9036 = ~n10114 | ~n10117;
  assign n10370 = ~INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n9037 = ~INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n10071 = ~n9464 | ~n9037;
  assign n10070 = ~n9041 | ~INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n10337 = ~INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n10321 = ~INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n9038 = ~n10337 | ~n10321;
  assign n9039 = ~n9041 | ~n9038;
  assign n9040 = ~n10070 | ~n9039;
  assign n10280 = INSTADDRPOINTER_REG_17__SCAN_IN & INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n9042 = ~INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n10268 = ~INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n9165 = ~n10089 & ~n10268;
  assign n9044 = ~n9161 & ~n9165;
  assign n9043 = ~INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n9164 = n10004 | n9043;
  assign n9045 = ~n9044 | ~n9164;
  assign n9169 = ~INSTADDRPOINTER_REG_22__SCAN_IN | ~INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n9046 = ~INSTADDRPOINTER_REG_21__SCAN_IN | ~INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n9047 = n9169 | n9046;
  assign n9049 = ~n10089 | ~n9047;
  assign n9335 = ~INSTADDRPOINTER_REG_20__SCAN_IN | ~INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n9048 = ~n10089 | ~n9335;
  assign n9050 = ~INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n9347 = ~INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n9051 = ~n9050 | ~n9347;
  assign n9052 = ~n9051 & ~INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n9054 = ~n9041 & ~INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n10228 = ~INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n9053 = ~n10089 & ~n10228;
  assign n9984 = ~n9054 & ~n9053;
  assign n9055 = ~n9054;
  assign n9056 = ~INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n9972 = ~n10089 | ~n9056;
  assign n10201 = ~INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n9959 = ~n10089 | ~n10201;
  assign n10193 = ~INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n9973 = n10004 | n9056;
  assign n9960 = n10004 | n10201;
  assign n9945 = ~n9973 | ~n9960;
  assign n9057 = ~n10089 & ~n10193;
  assign n9357 = ~n9945 & ~n9057;
  assign n9059 = ~n9466 | ~n9357;
  assign n9058 = INSTADDRPOINTER_REG_29__SCAN_IN ^ n9464;
  assign n9063 = ~INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~n12240;
  assign n9069 = INSTQUEUERD_ADDR_REG_2__SCAN_IN ^ ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n9076 = INSTQUEUERD_ADDR_REG_1__SCAN_IN ^ ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n9079 = ~n9060 | ~n13354;
  assign n9061 = ~n13355 | ~INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n9070 = ~n9079 | ~n9061;
  assign n9062 = ~n9069 | ~n9070;
  assign n9108 = ~n9063 | ~n9062;
  assign n9065 = ~n9108 | ~n9107;
  assign n9064 = ~n12841 | ~INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n9150 = ~INSTQUEUEWR_ADDR_REG_4__SCAN_IN | ~n9122;
  assign n9066 = ~n9126 & ~n9085;
  assign n9117 = ~n9150 & ~n9066;
  assign n9068 = ~n9150 & ~n7595;
  assign n9067 = ~STATE2_REG_0__SCAN_IN & ~n11873;
  assign n9116 = ~n9068 & ~n9067;
  assign n9121 = ~n9117 & ~n9116;
  assign n9089 = ~n9126;
  assign n9149 = n9070 ^ ~n9069;
  assign n9071 = ~n9149;
  assign n9073 = ~n9089 | ~n9071;
  assign n9072 = ~n7595 | ~n9149;
  assign n9075 = ~n9073 | ~n9072;
  assign n9074 = ~n11908 | ~n13308;
  assign n9104 = ~n9075 | ~n9105;
  assign n9078 = ~n13354 | ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n9077 = ~n9076;
  assign n9080 = ~n9078 | ~n9077;
  assign n9153 = ~n9080 | ~n9079;
  assign n9082 = ~n9081 | ~n9153;
  assign n9084 = ~n9082 | ~n13308;
  assign n9083 = n9126 & n9454;
  assign n9086 = ~n9153 & ~n13400;
  assign n9087 = ~n9129 & ~n9086;
  assign n9102 = n9088 | n9087;
  assign n9100 = ~n9088 | ~n9087;
  assign n9091 = INSTQUEUERD_ADDR_REG_0__SCAN_IN ^ INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n9090 = ~n9089 & ~n9091;
  assign n9098 = ~n9090 & ~n9129;
  assign n9092 = ~n9091;
  assign n9094 = n9092 & n9132;
  assign n9096 = ~n9094 & ~n9093;
  assign n9095 = ~n9105;
  assign n9097 = ~n9096 & ~n9095;
  assign n9099 = ~n9098 & ~n9097;
  assign n9101 = ~n9100 | ~n9099;
  assign n9103 = ~n9102 | ~n9101;
  assign n9106 = ~n9105 & ~n9149;
  assign n9111 = ~n9106 | ~n9126;
  assign n9148 = n9108 ^ ~n9107;
  assign n9110 = ~n9148 | ~n9109;
  assign n9112 = ~n9111 | ~n9110;
  assign n9114 = ~n9148 | ~n7595;
  assign n9118 = n9117 & n9116;
  assign n9124 = ~INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~n9123;
  assign n9127 = ~n9155 | ~n9126;
  assign n9134 = ~n7774 & ~n8946;
  assign n9133 = ~n9132 & ~n13310;
  assign n13331 = ~n11806 | ~n13315;
  assign n10176 = ~n11576 | ~REIP_REG_29__SCAN_IN;
  assign n13736 = ~n13102 | ~n9136;
  assign n9137 = ~n13736 | ~n13400;
  assign n9138 = ~n11581 | ~PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n9141 = ~n10176 | ~n9138;
  assign n9139 = ~n13400 | ~STATE2_REG_2__SCAN_IN;
  assign n9496 = ~STATE2_REG_1__SCAN_IN | ~n13100;
  assign n11580 = ~n9139 | ~n9496;
  assign n9140 = ~n11570 & ~n9573;
  assign n9144 = ~n13342 | ~n13390;
  assign n13304 = ~STATE2_REG_2__SCAN_IN | ~STATE2_REG_1__SCAN_IN;
  assign n13735 = ~n11186;
  assign U2892 = n11245 & DATAO_REG_31__SCAN_IN;
  assign n13762 = ~n13102 & ~STATE2_REG_1__SCAN_IN;
  assign n9151 = ~n9149 & ~n9148;
  assign n9152 = ~n9151 | ~n9150;
  assign n9154 = ~n9153 & ~n9152;
  assign n13320 = ~n9156 | ~n13310;
  assign n9157 = ~n13320 & ~n13404;
  assign n9158 = ~MEMORYFETCH_REG_SCAN_IN;
  assign n9159 = ~n9494 & ~n9158;
  assign n9160 = ~n13762 & ~n9159;
  assign U2788 = ~n11263 | ~n9160;
  assign n9163 = ~n9162;
  assign n10042 = ~n9041 & ~INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n10041 = ~n9164;
  assign n9166 = n10004 & n10268;
  assign n10030 = ~n9165 & ~n9166;
  assign n9998 = ~n9166;
  assign n10256 = ~INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n10003 = ~n9168 | ~n10256;
  assign n9167 = ~n10003 & ~INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n9171 = ~n9167 & ~n10089;
  assign n9170 = ~n10018 & ~n9169;
  assign n9172 = n10004 ^ ~INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n13739 = ~n13742;
  assign n10434 = ~n9454 & ~n13739;
  assign n9175 = ~n11828 & ~n10434;
  assign n9176 = ~n11806 | ~n9175;
  assign n9180 = ~n9176 | ~n11918;
  assign n9177 = ~n9454 | ~n13742;
  assign n9178 = ~n13321 | ~n9177;
  assign n9308 = ~n11918;
  assign n9179 = ~n9178 | ~n9308;
  assign n9181 = ~n9180 | ~n9179;
  assign n9185 = ~READY_N & ~n9181;
  assign n9183 = ~n13345 | ~n9454;
  assign n9184 = ~n11806 & ~n9183;
  assign n9186 = n9847 & n11938;
  assign n9190 = ~n9187 | ~n9186;
  assign n9188 = n9847 | n11908;
  assign n9189 = n9188 & n7004;
  assign n9316 = ~n9190 | ~n9189;
  assign n9193 = n9191 & n9316;
  assign n9203 = n8310 | n11938;
  assign n9192 = ~n9203 | ~n13310;
  assign n9194 = ~n9193 | ~n9192;
  assign n9195 = ~n7774 | ~n7004;
  assign n9196 = ~n9195 | ~n11918;
  assign n9197 = ~n13325 & ~n9196;
  assign n9198 = ~n10443 & ~n9197;
  assign n9200 = ~n9199 | ~n9198;
  assign n9331 = n9200 & n13390;
  assign n9204 = ~n11867 & ~n13315;
  assign n9202 = n10481 | n8946;
  assign n13318 = ~n11819;
  assign n9208 = n9204 & n13318;
  assign n9206 = ~n9298 | ~n13311;
  assign n9205 = n9142 | n11908;
  assign n9207 = n9206 & n9205;
  assign n9209 = ~n9208 | ~n9207;
  assign n9353 = ~n9479 | ~n11803;
  assign n9212 = ~n9214 | ~EBX_REG_24__SCAN_IN;
  assign n9215 = n11908 | n13310;
  assign n9213 = ~n9212 | ~n9211;
  assign n9359 = n9213 ^ ~n9286;
  assign n9217 = ~n9214 | ~EBX_REG_1__SCAN_IN;
  assign n9216 = ~n9215 | ~INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n9219 = ~n9217 | ~n9216;
  assign n9227 = n9219 ^ ~n9218;
  assign n9226 = ~n9227;
  assign n9221 = ~n9220;
  assign n9224 = ~n9221 | ~EBX_REG_0__SCAN_IN;
  assign n9222 = ~EBX_REG_0__SCAN_IN;
  assign n9223 = ~n9286 | ~n9222;
  assign n10911 = ~n9224 | ~n9223;
  assign n9229 = ~n9214 | ~EBX_REG_2__SCAN_IN;
  assign n9507 = ~n9786;
  assign n9228 = ~n9507 | ~INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n9231 = ~n9229 | ~n9228;
  assign n10863 = n9231 ^ ~n9286;
  assign n9233 = ~n9214 | ~EBX_REG_3__SCAN_IN;
  assign n9234 = ~n9233 | ~n9232;
  assign n9236 = ~n9214 | ~EBX_REG_4__SCAN_IN;
  assign n9237 = ~n9236 | ~n9235;
  assign n10802 = n9237 ^ ~n9286;
  assign n9238 = ~n10802;
  assign n9240 = ~n9214 | ~EBX_REG_5__SCAN_IN;
  assign n9241 = ~n9240 | ~n9239;
  assign n10787 = n9241 ^ ~n9286;
  assign n9243 = ~n9214 | ~EBX_REG_6__SCAN_IN;
  assign n9244 = ~n9243 | ~n9242;
  assign n10762 = n9244 ^ ~n9286;
  assign n9246 = ~n9214 | ~EBX_REG_7__SCAN_IN;
  assign n9247 = ~n9246 | ~n9245;
  assign n10734 = n9247 ^ ~n9218;
  assign n10725 = ~n10735 | ~n10734;
  assign n9249 = ~n9214 | ~EBX_REG_8__SCAN_IN;
  assign n9248 = ~n9507 | ~INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n9250 = ~n9249 | ~n9248;
  assign n10724 = n9250 ^ ~n9286;
  assign n9252 = ~n9214 | ~EBX_REG_9__SCAN_IN;
  assign n9253 = ~n9252 | ~n9251;
  assign n10694 = n9253 ^ ~n9286;
  assign n9255 = ~n9214 | ~EBX_REG_10__SCAN_IN;
  assign n9254 = ~n9507 | ~INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n9256 = ~n9255 | ~n9254;
  assign n10675 = n9256 ^ ~n9218;
  assign n10666 = n10674 & n10675;
  assign n9258 = ~n9214 | ~EBX_REG_11__SCAN_IN;
  assign n9257 = ~n9507 | ~INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n9259 = ~n9258 | ~n9257;
  assign n10665 = n9259 ^ ~n9218;
  assign n9261 = ~n9214 | ~EBX_REG_12__SCAN_IN;
  assign n9260 = ~n9507 | ~INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n9262 = ~n9261 | ~n9260;
  assign n10645 = n9262 ^ ~n9286;
  assign n9264 = ~n9214 | ~EBX_REG_13__SCAN_IN;
  assign n9263 = ~n9507 | ~INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n9265 = ~n9264 | ~n9263;
  assign n10422 = n9265 ^ ~n9286;
  assign n9267 = ~n9214 | ~EBX_REG_14__SCAN_IN;
  assign n9266 = ~n9507 | ~INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n9268 = ~n9267 | ~n9266;
  assign n10408 = n9268 ^ ~n9218;
  assign n9270 = ~n9214 | ~EBX_REG_15__SCAN_IN;
  assign n9269 = ~n9507 | ~INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n9271 = ~n9270 | ~n9269;
  assign n10376 = n9271 ^ ~n9218;
  assign n9273 = ~n9214 | ~EBX_REG_16__SCAN_IN;
  assign n9272 = ~n9507 | ~INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n9274 = ~n9273 | ~n9272;
  assign n10358 = n9274 ^ ~n9286;
  assign n9276 = ~n9214 | ~EBX_REG_17__SCAN_IN;
  assign n9275 = ~n9507 | ~INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n9277 = ~n9276 | ~n9275;
  assign n10341 = n9277 ^ ~n9286;
  assign n9279 = ~n9214 | ~EBX_REG_18__SCAN_IN;
  assign n9278 = ~n9507 | ~INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n9280 = ~n9279 | ~n9278;
  assign n10324 = n9280 ^ ~n9218;
  assign n9282 = ~n9214 | ~EBX_REG_19__SCAN_IN;
  assign n9281 = ~n9507 | ~INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n9283 = ~n9282 | ~n9281;
  assign n9767 = n9283 ^ ~n9218;
  assign n9285 = ~n9214 | ~EBX_REG_20__SCAN_IN;
  assign n9287 = ~n9285 | ~n9284;
  assign n9745 = n9287 ^ ~n9286;
  assign n9289 = ~n9214 | ~EBX_REG_21__SCAN_IN;
  assign n9288 = ~n9507 | ~INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n9290 = ~n9289 | ~n9288;
  assign n9726 = n9290 ^ ~n9286;
  assign n9293 = ~n9214 | ~EBX_REG_22__SCAN_IN;
  assign n9294 = ~n9293 | ~n9292;
  assign n9704 = n9294 ^ ~n9286;
  assign n9296 = ~n9214 | ~EBX_REG_23__SCAN_IN;
  assign n9297 = ~n9296 | ~n9295;
  assign n9686 = n9297 ^ ~n9218;
  assign n9820 = n9359 ^ n7043;
  assign n9299 = ~n9298 | ~n11938;
  assign n13380 = n9142 | n9454;
  assign n9300 = ~n9299 | ~n13380;
  assign n9301 = ~n9820 | ~n11739;
  assign n9486 = ~n11576 | ~REIP_REG_24__SCAN_IN;
  assign n9351 = ~n9301 | ~n9486;
  assign n11795 = ~n9331 & ~n11576;
  assign n9306 = n9302 | n7004;
  assign n9305 = ~n11829 | ~n9304;
  assign n9324 = n9306 & n9305;
  assign n9312 = n7144 & n13743;
  assign n9310 = ~n7774 | ~n9308;
  assign n9309 = n11918 | n13310;
  assign n9311 = ~n9310 | ~n9309;
  assign n9314 = ~n9312 & ~n9311;
  assign n9313 = ~n9214 | ~n8946;
  assign n9318 = ~n9314 | ~n9313;
  assign n9317 = ~n9316 | ~n9315;
  assign n9319 = ~n9318 & ~n9317;
  assign n11834 = ~n9320 | ~n9319;
  assign n9321 = ~n13310 | ~n13308;
  assign n11847 = ~n9322 & ~n9321;
  assign n9323 = ~n11834 & ~n11847;
  assign n9325 = ~n9324 | ~n9323;
  assign n11794 = ~INSTADDRPOINTER_REG_0__SCAN_IN & ~n10390;
  assign n9334 = ~INSTADDRPOINTER_REG_16__SCAN_IN | ~INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n9329 = ~n9334;
  assign n10399 = INSTADDRPOINTER_REG_12__SCAN_IN & INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n10387 = ~INSTADDRPOINTER_REG_13__SCAN_IN | ~n10399;
  assign n9333 = ~INSTADDRPOINTER_REG_10__SCAN_IN | ~INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n9332 = ~n9021 & ~n11678;
  assign n11731 = ~INSTADDRPOINTER_REG_2__SCAN_IN & ~n9326;
  assign n11713 = ~INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n11728 = ~INSTADDRPOINTER_REG_4__SCAN_IN | ~INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n9327 = ~n11713 & ~n11728;
  assign n11659 = ~INSTADDRPOINTER_REG_6__SCAN_IN | ~n9327;
  assign n11665 = ~n11731 & ~n11659;
  assign n11630 = ~n9332 | ~n11665;
  assign n11599 = ~n9333 & ~n11630;
  assign n9328 = ~INSTADDRPOINTER_REG_14__SCAN_IN | ~n11599;
  assign n10353 = ~n10387 & ~n9328;
  assign n10278 = ~n9329 | ~n10353;
  assign n10314 = ~n10337 & ~n10278;
  assign n10286 = ~INSTADDRPOINTER_REG_18__SCAN_IN | ~n10314;
  assign n9344 = ~n9335 & ~n10286;
  assign n13324 = ~n13345 | ~n9330;
  assign n11818 = ~n13324;
  assign n9337 = ~n9344 & ~n11732;
  assign n11752 = ~INSTADDRPOINTER_REG_2__SCAN_IN | ~INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n11662 = ~n11752 & ~n11659;
  assign n11627 = ~n11662 | ~n9332;
  assign n11602 = ~n11627 & ~n9333;
  assign n10349 = ~n11602;
  assign n10394 = ~n10349 & ~n10387;
  assign n10355 = ~INSTADDRPOINTER_REG_14__SCAN_IN | ~n10394;
  assign n10315 = ~n10355 & ~n9334;
  assign n10283 = ~n10280 | ~n10315;
  assign n9343 = ~n10283 & ~n9335;
  assign n9336 = ~n11663 & ~n9343;
  assign n9338 = ~n9337 & ~n9336;
  assign n10269 = ~n11773 | ~n9338;
  assign n10259 = ~n10256 & ~n10268;
  assign n11689 = ~n11663;
  assign n9339 = ~n10259 & ~n9389;
  assign n9341 = ~INSTADDRPOINTER_REG_24__SCAN_IN | ~INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n11778 = ~INSTADDRPOINTER_REG_0__SCAN_IN & ~n11796;
  assign n11765 = ~n11663 & ~n11778;
  assign n11625 = ~n11765;
  assign n9340 = ~n11625 | ~n11732;
  assign n9342 = ~n9341 | ~n9340;
  assign n10229 = ~n10239 | ~n9342;
  assign n9346 = ~n9343 | ~n11765;
  assign n9345 = ~n9344 | ~n11772;
  assign n9348 = ~n10240 | ~INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n9349 = ~n9348 | ~n9347;
  assign n9350 = n10229 & n9349;
  assign n9352 = ~n9351 & ~n9350;
  assign U2994 = ~n9353 | ~n9352;
  assign n9383 = ~INSTADDRPOINTER_REG_28__SCAN_IN | ~INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n9354 = ~INSTADDRPOINTER_REG_26__SCAN_IN | ~INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n9355 = ~n9383 & ~n9354;
  assign n9356 = ~n9041 | ~INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n9358 = n10004 ^ ~INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n9934 = n9462 ^ ~n9358;
  assign n9394 = ~n9934 | ~n11803;
  assign n9361 = ~n9214 | ~EBX_REG_25__SCAN_IN;
  assign n9362 = ~n9361 | ~n9360;
  assign n9648 = n9362 ^ ~n9286;
  assign n9629 = ~n7019 & ~n9648;
  assign n9364 = ~n9214 | ~EBX_REG_26__SCAN_IN;
  assign n9365 = ~n9364 | ~n9363;
  assign n9630 = n9365 ^ ~n9218;
  assign n9609 = ~n9629 | ~n9630;
  assign n9367 = ~n9214 | ~EBX_REG_27__SCAN_IN;
  assign n9368 = ~n9367 | ~n9366;
  assign n9608 = n9368 ^ ~n9286;
  assign n9370 = ~n9214 | ~EBX_REG_28__SCAN_IN;
  assign n9371 = ~n9370 | ~n9369;
  assign n9589 = n9371 ^ ~n9286;
  assign n9373 = ~n9214 | ~EBX_REG_29__SCAN_IN;
  assign n9374 = ~n9373 | ~n9372;
  assign n9567 = n9374 ^ ~n9218;
  assign n9505 = ~n9503 | ~n9286;
  assign n9375 = ~n9374;
  assign n9376 = ~n9589 & ~n9375;
  assign n9380 = ~n9505 | ~n9377;
  assign n9379 = ~n9214 | ~EBX_REG_30__SCAN_IN;
  assign n9504 = ~n9379 | ~n9378;
  assign n9381 = ~n9794;
  assign n9938 = ~n11576 | ~REIP_REG_30__SCAN_IN;
  assign n9384 = ~INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n9382 = INSTADDRPOINTER_REG_23__SCAN_IN & INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n10230 = ~n10240 | ~n9382;
  assign n9385 = ~INSTADDRPOINTER_REG_26__SCAN_IN | ~INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n9387 = ~n9383;
  assign n10179 = ~n10203 | ~n9387;
  assign n10159 = ~n9384 & ~n10179;
  assign n9392 = ~n10159 & ~INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n11780 = ~n9389;
  assign n9386 = n9385 & n11780;
  assign n9388 = n9387 | n9389;
  assign n10178 = ~n10200 | ~n9388;
  assign n9390 = ~INSTADDRPOINTER_REG_29__SCAN_IN & ~n9389;
  assign n9393 = ~n9392 & ~n9391;
  assign n9396 = ~PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n9936 = PHYADDRPOINTER_REG_30__SCAN_IN ^ n9471;
  assign n9445 = ~n9936 | ~n8929;
  assign n9400 = ~n9398 | ~INSTQUEUE_REG_11__7__SCAN_IN;
  assign n9399 = ~n8567 | ~INSTQUEUE_REG_6__7__SCAN_IN;
  assign n9405 = ~n9400 | ~n9399;
  assign n9403 = ~n9401 | ~INSTQUEUE_REG_5__7__SCAN_IN;
  assign n9402 = ~n8693 | ~INSTQUEUE_REG_7__7__SCAN_IN;
  assign n9404 = ~n9403 | ~n9402;
  assign n9414 = ~n9405 & ~n9404;
  assign n9407 = ~n8526 | ~INSTQUEUE_REG_1__7__SCAN_IN;
  assign n9406 = ~n8279 | ~INSTQUEUE_REG_3__7__SCAN_IN;
  assign n9412 = ~n9407 | ~n9406;
  assign n9410 = ~n7006 | ~INSTQUEUE_REG_9__7__SCAN_IN;
  assign n9409 = ~n8910 | ~INSTQUEUE_REG_15__7__SCAN_IN;
  assign n9411 = ~n9410 | ~n9409;
  assign n9413 = ~n9412 & ~n9411;
  assign n9430 = ~n9414 | ~n9413;
  assign n9416 = ~n8854 | ~INSTQUEUE_REG_12__7__SCAN_IN;
  assign n9415 = ~n7807 | ~INSTQUEUE_REG_4__7__SCAN_IN;
  assign n9420 = ~n9416 | ~n9415;
  assign n9418 = ~n7009 | ~INSTQUEUE_REG_2__7__SCAN_IN;
  assign n9417 = ~n8892 | ~INSTQUEUE_REG_8__7__SCAN_IN;
  assign n9419 = ~n9418 | ~n9417;
  assign n9428 = ~n9420 & ~n9419;
  assign n9422 = ~n8906 | ~INSTQUEUE_REG_14__7__SCAN_IN;
  assign n9421 = ~n8586 | ~INSTQUEUE_REG_10__7__SCAN_IN;
  assign n9426 = ~n9422 | ~n9421;
  assign n9424 = ~n8915 | ~INSTQUEUE_REG_13__7__SCAN_IN;
  assign n9423 = ~n7014 | ~INSTQUEUE_REG_0__7__SCAN_IN;
  assign n9425 = ~n9424 | ~n9423;
  assign n9427 = ~n9426 & ~n9425;
  assign n9429 = ~n9428 | ~n9427;
  assign n9434 = ~n9430 & ~n9429;
  assign n9433 = ~n9432 & ~n9431;
  assign n9436 = n9434 ^ ~n9433;
  assign n9443 = ~n9436 | ~n9435;
  assign n9437 = ~EAX_REG_30__SCAN_IN;
  assign n9441 = ~n9438 & ~n9437;
  assign n9439 = ~PHYADDRPOINTER_REG_30__SCAN_IN | ~n11983;
  assign n9440 = ~n8384 | ~n9439;
  assign n9442 = ~n9441 & ~n9440;
  assign n9444 = ~n9443 | ~n9442;
  assign n9541 = ~n9445 | ~n9444;
  assign n9448 = ~n7864 | ~EAX_REG_31__SCAN_IN;
  assign n9447 = ~n9446 | ~PHYADDRPOINTER_REG_31__SCAN_IN;
  assign n9457 = ~n9493 | ~n13328;
  assign n10448 = ~n11806 | ~n11819;
  assign n10439 = ~n13321 | ~n11867;
  assign n9449 = ~n13328 | ~n11938;
  assign n9787 = ~n9449 & ~n7773;
  assign n9450 = ~n11829 | ~n9787;
  assign n9453 = ~n10448 | ~n9452;
  assign n13431 = ~READY_N;
  assign n9455 = ~n9454 | ~n13431;
  assign n9459 = ~n9457 | ~n11092;
  assign n9458 = n11092 | EAX_REG_31__SCAN_IN;
  assign n9461 = ~n9459 | ~n9458;
  assign n11037 = ~n6994 & ~n7774;
  assign n9460 = ~n11037 | ~DATAI_31_;
  assign U2860 = ~n9461 | ~n9460;
  assign n10165 = ~INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n9463 = ~n10165 & ~n9384;
  assign n9465 = ~n9464 | ~n9463;
  assign n9467 = ~n9466 | ~INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n9469 = ~n9468 | ~n9467;
  assign n9478 = ~n10158 | ~n11578;
  assign n9476 = n9493 & n6996;
  assign n10161 = ~REIP_REG_31__SCAN_IN | ~n11576;
  assign n9470 = ~n11581 | ~PHYADDRPOINTER_REG_31__SCAN_IN;
  assign n9474 = n10161 & n9470;
  assign n9472 = ~n9471 | ~PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n9473 = ~n11548 | ~n9550;
  assign n9475 = ~n9474 | ~n9473;
  assign n9477 = ~n9476 & ~n9475;
  assign U2955 = ~n9478 | ~n9477;
  assign n9492 = ~n9479 | ~n11578;
  assign n9484 = ~n9480;
  assign n9483 = ~n9481 | ~n9482;
  assign n9819 = ~n9484 | ~n9483;
  assign n9490 = ~n9819 & ~n11881;
  assign n9485 = ~n11581 | ~PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n9488 = ~n9486 | ~n9485;
  assign n9487 = ~n11570 & ~n9669;
  assign n9489 = n9488 | n9487;
  assign n9491 = ~n9490 & ~n9489;
  assign U2962 = ~n9492 | ~n9491;
  assign n9495 = ~n9494;
  assign n13409 = ~STATE2_REG_0__SCAN_IN & ~STATE2_REG_2__SCAN_IN;
  assign n9497 = ~n9496;
  assign n13398 = ~n13409 | ~n9497;
  assign n9498 = STATE2_REG_3__SCAN_IN & n11983;
  assign n9499 = STATE2_REG_0__SCAN_IN & n9498;
  assign n13392 = ~n9499 | ~n13655;
  assign n9500 = n13398 & n13392;
  assign n9539 = ~n9493 | ~n10770;
  assign n9506 = ~n9570 | ~n9504;
  assign n9509 = ~n9214 | ~EBX_REG_31__SCAN_IN;
  assign n9508 = ~n9507 | ~INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n9510 = ~n9509 | ~n9508;
  assign n9526 = ~STATEBS16_REG_SCAN_IN & ~READY_N;
  assign n9553 = ~n9526;
  assign n9512 = ~n9553 | ~n9527;
  assign n9537 = ~n10927 & ~n10914;
  assign n13568 = ~REIP_REG_25__SCAN_IN;
  assign n9513 = ~n10809 | ~n9526;
  assign n10851 = ~n10434 & ~n9514;
  assign n13563 = ~REIP_REG_24__SCAN_IN;
  assign n13558 = ~REIP_REG_23__SCAN_IN;
  assign n13548 = ~REIP_REG_21__SCAN_IN;
  assign n13539 = ~REIP_REG_19__SCAN_IN;
  assign n13529 = ~REIP_REG_17__SCAN_IN;
  assign n13519 = ~REIP_REG_15__SCAN_IN;
  assign n13509 = ~REIP_REG_13__SCAN_IN;
  assign n13499 = ~REIP_REG_11__SCAN_IN;
  assign n13489 = ~REIP_REG_9__SCAN_IN;
  assign n13479 = ~REIP_REG_7__SCAN_IN;
  assign n13469 = ~REIP_REG_5__SCAN_IN;
  assign n13722 = ~REIP_REG_1__SCAN_IN;
  assign n9515 = ~REIP_REG_3__SCAN_IN | ~REIP_REG_2__SCAN_IN;
  assign n10812 = ~n13722 & ~n9515;
  assign n10778 = ~REIP_REG_4__SCAN_IN | ~n10812;
  assign n10760 = ~n13469 & ~n10778;
  assign n10739 = ~REIP_REG_6__SCAN_IN | ~n10760;
  assign n10722 = ~n13479 & ~n10739;
  assign n10693 = ~REIP_REG_8__SCAN_IN | ~n10722;
  assign n10680 = ~n13489 & ~n10693;
  assign n10659 = ~REIP_REG_10__SCAN_IN | ~n10680;
  assign n10612 = ~n13499 & ~n10659;
  assign n10619 = ~REIP_REG_12__SCAN_IN | ~n10612;
  assign n10597 = ~n13509 & ~n10619;
  assign n10582 = ~REIP_REG_14__SCAN_IN | ~n10597;
  assign n10563 = ~n13519 & ~n10582;
  assign n10542 = ~REIP_REG_16__SCAN_IN | ~n10563;
  assign n10527 = ~n13529 & ~n10542;
  assign n9773 = ~REIP_REG_18__SCAN_IN | ~n10527;
  assign n9756 = ~n13539 & ~n9773;
  assign n9736 = ~REIP_REG_20__SCAN_IN | ~n9756;
  assign n9707 = ~n13548 & ~n9736;
  assign n9695 = ~REIP_REG_22__SCAN_IN | ~n9707;
  assign n9657 = ~n13558 & ~n9695;
  assign n9668 = ~n9657;
  assign n9517 = ~n13563 & ~n9668;
  assign n9650 = ~n7007 | ~n9517;
  assign n9633 = ~n13568 & ~n9650;
  assign n9613 = ~REIP_REG_26__SCAN_IN | ~n9633;
  assign n9521 = ~REIP_REG_28__SCAN_IN | ~REIP_REG_27__SCAN_IN;
  assign n9571 = ~n9613 & ~n9521;
  assign n9523 = ~REIP_REG_30__SCAN_IN | ~REIP_REG_29__SCAN_IN;
  assign n9516 = ~REIP_REG_31__SCAN_IN & ~n9523;
  assign n9535 = ~n9571 | ~n9516;
  assign n9518 = REIP_REG_25__SCAN_IN & n9517;
  assign n9519 = ~n9518 | ~REIP_REG_26__SCAN_IN;
  assign n9520 = ~n9519 | ~n10851;
  assign n9632 = ~n9520 | ~n10893;
  assign n9522 = n9521 & n10851;
  assign n9572 = ~n9632 & ~n9522;
  assign n9524 = ~n10851 | ~n9523;
  assign n9544 = ~n9572 | ~n9524;
  assign n9533 = ~REIP_REG_31__SCAN_IN | ~n9544;
  assign n9525 = ~PHYADDRPOINTER_REG_31__SCAN_IN;
  assign n9531 = ~n10907 & ~n9525;
  assign n13379 = ~n13739 | ~n9526;
  assign n9528 = ~n13379 | ~n9527;
  assign n9530 = ~n9529 & ~n9528;
  assign n9532 = ~n9531 & ~n9530;
  assign n9534 = n9533 & n9532;
  assign n9536 = ~n9535 | ~n9534;
  assign n9538 = ~n9537 & ~n9536;
  assign U2796 = ~n9539 | ~n9538;
  assign n9542 = ~n9540 | ~n9541;
  assign n9935 = ~n9543 | ~n9542;
  assign n9565 = ~n9848 | ~n10770;
  assign n9563 = ~n9794 & ~n10914;
  assign n9546 = ~n10896 | ~PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n9545 = ~REIP_REG_30__SCAN_IN | ~n9544;
  assign n9549 = ~n9546 | ~n9545;
  assign n9547 = ~n9571 | ~REIP_REG_29__SCAN_IN;
  assign n9548 = ~REIP_REG_30__SCAN_IN & ~n9547;
  assign n9561 = ~n9549 & ~n9548;
  assign n9551 = ~n9550 & ~n13655;
  assign n9559 = ~n9936 | ~n10869;
  assign n9556 = ~n13741 | ~n13379;
  assign n9552 = ~EBX_REG_31__SCAN_IN;
  assign n9554 = ~n9553 | ~n9552;
  assign n9555 = n13310 | n9554;
  assign n9557 = ~n9556 | ~n9555;
  assign n10904 = n10809 & n9557;
  assign n9558 = ~EBX_REG_30__SCAN_IN | ~n10904;
  assign n9560 = n9559 & n9558;
  assign n9562 = ~n9561 | ~n9560;
  assign n9564 = ~n9563 & ~n9562;
  assign U2797 = ~n9565 | ~n9564;
  assign n9585 = ~n9857 | ~n10770;
  assign n9569 = ~n9568 & ~n9567;
  assign n9583 = ~n10174 & ~n10914;
  assign n13589 = ~REIP_REG_29__SCAN_IN;
  assign n9581 = ~n9571 | ~n13589;
  assign n9592 = ~n9572;
  assign n9579 = ~REIP_REG_29__SCAN_IN | ~n9592;
  assign n9577 = ~n10908 & ~n9573;
  assign n9575 = ~n10896 | ~PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n9574 = ~n10904 | ~EBX_REG_29__SCAN_IN;
  assign n9576 = ~n9575 | ~n9574;
  assign n9578 = ~n9577 & ~n9576;
  assign n9580 = n9579 & n9578;
  assign n9582 = ~n9581 | ~n9580;
  assign n9584 = ~n9583 & ~n9582;
  assign U2798 = ~n9585 | ~n9584;
  assign n9604 = ~n9864 | ~n10770;
  assign n10188 = n9589 ^ n9611;
  assign n9590 = ~n10188;
  assign n9602 = ~n9590 & ~n10914;
  assign n9591 = ~REIP_REG_28__SCAN_IN & ~n9613;
  assign n9600 = ~REIP_REG_27__SCAN_IN | ~n9591;
  assign n9598 = ~REIP_REG_28__SCAN_IN | ~n9592;
  assign n9596 = ~n9949 & ~n7011;
  assign n9594 = ~n10896 | ~PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n9593 = ~n10904 | ~EBX_REG_28__SCAN_IN;
  assign n9595 = ~n9594 | ~n9593;
  assign n9597 = ~n9596 & ~n9595;
  assign n9599 = n9598 & n9597;
  assign n9601 = ~n9600 | ~n9599;
  assign n9603 = ~n9602 & ~n9601;
  assign U2799 = ~n9604 | ~n9603;
  assign n9606 = n9605;
  assign n9963 = n9606 ^ ~n9607;
  assign n9871 = ~n9963;
  assign n9625 = ~n9871 | ~n10770;
  assign n9610 = ~n9609 | ~n9608;
  assign n9612 = ~n10206;
  assign n9623 = ~n9612 & ~n10914;
  assign n9619 = n10896 & PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n9615 = n9613 | REIP_REG_27__SCAN_IN;
  assign n9614 = ~n10904 | ~EBX_REG_27__SCAN_IN;
  assign n9617 = n9615 & n9614;
  assign n9616 = ~n9632 | ~REIP_REG_27__SCAN_IN;
  assign n9618 = ~n9617 | ~n9616;
  assign n9621 = ~n9619 & ~n9618;
  assign n9620 = ~n10869 | ~n9965;
  assign n9622 = ~n9621 | ~n9620;
  assign n9624 = ~n9623 & ~n9622;
  assign U2800 = ~n9625 | ~n9624;
  assign n9628 = n9627 | n9626;
  assign n9975 = ~n9606 | ~n9628;
  assign n9878 = ~n9975;
  assign n9646 = ~n9878 | ~n10770;
  assign n10214 = n9630 ^ n9629;
  assign n9631 = ~n10214;
  assign n9644 = ~n9631 & ~n10914;
  assign n9635 = ~n9632;
  assign n9634 = ~REIP_REG_26__SCAN_IN & ~n9633;
  assign n9642 = ~n9635 & ~n9634;
  assign n9638 = ~n10904 | ~EBX_REG_26__SCAN_IN;
  assign n9637 = n10907 | n9636;
  assign n9640 = n9638 & n9637;
  assign n9639 = ~n9977 | ~n10869;
  assign n9641 = ~n9640 | ~n9639;
  assign n9643 = n9642 | n9641;
  assign n9645 = ~n9644 & ~n9643;
  assign U2801 = ~n9646 | ~n9645;
  assign n9885 = ~n9988;
  assign n9665 = ~n9885 | ~n10770;
  assign n10225 = n7019 ^ n9648;
  assign n9649 = ~n10225;
  assign n9663 = ~n9649 & ~n10914;
  assign n9656 = ~REIP_REG_25__SCAN_IN & ~n9650;
  assign n9652 = ~n10896 | ~PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n9651 = ~n10904 | ~EBX_REG_25__SCAN_IN;
  assign n9654 = n9652 & n9651;
  assign n9653 = ~n10869 | ~n9990;
  assign n9655 = ~n9654 | ~n9653;
  assign n9661 = ~n9656 & ~n9655;
  assign n9667 = ~n10851 | ~n13563;
  assign n9658 = ~n9657 & ~n10830;
  assign n10831 = ~n10893;
  assign n9676 = n9658 | n10831;
  assign n9698 = ~n9676;
  assign n9659 = ~n9667 | ~n9698;
  assign n9660 = ~n9659 | ~REIP_REG_25__SCAN_IN;
  assign n9662 = ~n9661 | ~n9660;
  assign n9664 = ~n9663 & ~n9662;
  assign U2802 = ~n9665 | ~n9664;
  assign n9892 = ~n9819;
  assign n9682 = ~n9892 | ~n10770;
  assign n9666 = ~n9820;
  assign n9680 = ~n9666 & ~n10914;
  assign n9675 = ~n9668 & ~n9667;
  assign n9673 = ~n7011 & ~n9669;
  assign n9671 = ~n10896 | ~PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n9670 = ~EBX_REG_24__SCAN_IN | ~n10904;
  assign n9672 = ~n9671 | ~n9670;
  assign n9674 = n9673 | n9672;
  assign n9678 = ~n9675 & ~n9674;
  assign n9677 = ~n9676 | ~REIP_REG_24__SCAN_IN;
  assign n9679 = ~n9678 | ~n9677;
  assign n9681 = ~n9680 & ~n9679;
  assign U2803 = ~n9682 | ~n9681;
  assign n10007 = n9683 ^ ~n9684;
  assign n9899 = ~n10007;
  assign n9702 = ~n9899 | ~n10770;
  assign n10243 = n9686 ^ n9685;
  assign n9694 = ~n10243 | ~n10837;
  assign n9687 = ~n10010;
  assign n9690 = ~n7011 & ~n9687;
  assign n9689 = ~n10907 & ~n9688;
  assign n9692 = ~n9690 & ~n9689;
  assign n9691 = ~n10904 | ~EBX_REG_23__SCAN_IN;
  assign n9693 = n9692 & n9691;
  assign n9700 = ~n9694 | ~n9693;
  assign n9696 = ~n9695 & ~n10830;
  assign n9697 = ~REIP_REG_23__SCAN_IN & ~n9696;
  assign n9699 = ~n9698 & ~n9697;
  assign n9701 = ~n9700 & ~n9699;
  assign U2804 = ~n9702 | ~n9701;
  assign n10019 = n7052 ^ ~n9703;
  assign n9906 = ~n10019;
  assign n9722 = ~n9906 | ~n10770;
  assign n10251 = n9705 ^ ~n9704;
  assign n9716 = ~n10251 & ~n10914;
  assign n9706 = ~REIP_REG_22__SCAN_IN & ~n10830;
  assign n9714 = ~n9707 | ~n9706;
  assign n9708 = ~n10022;
  assign n9712 = ~n10908 & ~n9708;
  assign n9710 = ~n10896 | ~PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n9709 = ~n10904 | ~EBX_REG_22__SCAN_IN;
  assign n9711 = ~n9710 | ~n9709;
  assign n9713 = ~n9712 & ~n9711;
  assign n9715 = ~n9714 | ~n9713;
  assign n9720 = ~n9716 & ~n9715;
  assign n9717 = n9736 & n10851;
  assign n9759 = ~n9717 & ~n10831;
  assign n9735 = ~n10851 | ~n13548;
  assign n9718 = ~n9759 | ~n9735;
  assign n9719 = ~REIP_REG_22__SCAN_IN | ~n9718;
  assign n9721 = n9720 & n9719;
  assign U2805 = ~n9722 | ~n9721;
  assign n9724 = ~n7047 & ~n9723;
  assign n10031 = n7052 | n9724;
  assign n9913 = ~n10031;
  assign n9742 = ~n9913 | ~n10770;
  assign n10265 = n9747 ^ n9726;
  assign n9734 = ~n10265 | ~n10837;
  assign n9727 = ~n10034;
  assign n9732 = ~n10908 & ~n9727;
  assign n9730 = n10907 | n9728;
  assign n9729 = ~EBX_REG_21__SCAN_IN | ~n10904;
  assign n9731 = ~n9730 | ~n9729;
  assign n9733 = ~n9732 & ~n9731;
  assign n9738 = ~n9734 | ~n9733;
  assign n9737 = ~n9736 & ~n9735;
  assign n9740 = n9738 | n9737;
  assign n9739 = ~n9759 & ~n13548;
  assign n9741 = ~n9740 & ~n9739;
  assign U2806 = ~n9742 | ~n9741;
  assign n10044 = n9744 ^ n9743;
  assign n9763 = ~n10044 | ~n10770;
  assign n9746 = ~n7050 | ~n9745;
  assign n10291 = ~n9747 | ~n9746;
  assign n9748 = ~n10291;
  assign n9755 = ~n9748 | ~n10837;
  assign n9749 = ~n10904;
  assign n9837 = ~EBX_REG_20__SCAN_IN;
  assign n9753 = ~n9749 & ~n9837;
  assign n9751 = ~n10896 | ~PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n9750 = ~n10869 | ~n10048;
  assign n9752 = ~n9751 | ~n9750;
  assign n9754 = ~n9753 & ~n9752;
  assign n9761 = ~n9755 | ~n9754;
  assign n9757 = n10851 & n9756;
  assign n9758 = ~REIP_REG_20__SCAN_IN & ~n9757;
  assign n9760 = ~n9759 & ~n9758;
  assign n9762 = ~n9761 & ~n9760;
  assign U2807 = ~n9763 | ~n9762;
  assign n10059 = n9764 ^ ~n9765;
  assign n9927 = ~n10059;
  assign n9785 = ~n9927 | ~n10770;
  assign n10303 = n9766 ^ ~n9767;
  assign n9771 = ~n10303 & ~n10914;
  assign n9769 = ~n10904 | ~EBX_REG_19__SCAN_IN;
  assign n9768 = ~n10869 | ~n10061;
  assign n9770 = ~n9769 | ~n9768;
  assign n9775 = n9771 | n9770;
  assign n9772 = ~n10851 | ~n13539;
  assign n9774 = ~n9773 & ~n9772;
  assign n9783 = n9775 | n9774;
  assign n13534 = ~REIP_REG_18__SCAN_IN;
  assign n10525 = ~n10851 | ~n13534;
  assign n9776 = ~n10527 & ~n10830;
  assign n10545 = ~n10831 & ~n9776;
  assign n9777 = ~n10525 | ~n10545;
  assign n9781 = ~n9777 | ~REIP_REG_19__SCAN_IN;
  assign n10814 = ~n10893 | ~n13762;
  assign n10784 = ~n10814;
  assign n9779 = ~n10907 & ~n9778;
  assign n9780 = ~n10784 & ~n9779;
  assign n9782 = ~n9781 | ~n9780;
  assign n9784 = ~n9783 & ~n9782;
  assign U2808 = ~n9785 | ~n9784;
  assign n9790 = n9787 & n9786;
  assign n9789 = ~n9788;
  assign n9792 = ~n9790 | ~n9789;
  assign n9791 = ~n10451;
  assign n9793 = ~n9792 | ~n9791;
  assign n9798 = ~n9848 | ~n11020;
  assign n9796 = ~n9794 & ~n11016;
  assign n9795 = n11013 & EBX_REG_30__SCAN_IN;
  assign n9797 = ~n9796 & ~n9795;
  assign U2829 = ~n9798 | ~n9797;
  assign n9802 = ~n9857 | ~n11020;
  assign n9800 = ~n10174 & ~n11016;
  assign n9799 = n11013 & EBX_REG_29__SCAN_IN;
  assign n9801 = ~n9800 & ~n9799;
  assign U2830 = ~n9802 | ~n9801;
  assign n9806 = ~n9948 & ~n11010;
  assign n9804 = ~n10188 | ~n11001;
  assign n9803 = ~n11013 | ~EBX_REG_28__SCAN_IN;
  assign n9805 = ~n9804 | ~n9803;
  assign U2831 = n9806 | n9805;
  assign n9810 = ~n9963 & ~n11010;
  assign n9808 = ~n10206 | ~n11001;
  assign n9807 = ~n11013 | ~EBX_REG_27__SCAN_IN;
  assign n9809 = ~n9808 | ~n9807;
  assign U2832 = n9810 | n9809;
  assign n9814 = ~n9975 & ~n11010;
  assign n9812 = ~n10214 | ~n11001;
  assign n9811 = ~n11013 | ~EBX_REG_26__SCAN_IN;
  assign n9813 = ~n9812 | ~n9811;
  assign U2833 = n9814 | n9813;
  assign n9818 = ~n9988 & ~n11010;
  assign n9816 = ~n10225 | ~n11001;
  assign n9815 = ~n11013 | ~EBX_REG_25__SCAN_IN;
  assign n9817 = ~n9816 | ~n9815;
  assign U2834 = n9818 | n9817;
  assign n9824 = ~n9819 & ~n11010;
  assign n9822 = ~n9820 | ~n11001;
  assign n9821 = ~n11013 | ~EBX_REG_24__SCAN_IN;
  assign n9823 = ~n9822 | ~n9821;
  assign U2835 = n9824 | n9823;
  assign n9828 = ~n10007 & ~n11010;
  assign n9826 = ~n10243 | ~n11001;
  assign n9825 = ~n11013 | ~EBX_REG_23__SCAN_IN;
  assign n9827 = ~n9826 | ~n9825;
  assign U2836 = n9828 | n9827;
  assign n9832 = ~n9906 | ~n11020;
  assign n9830 = ~n10251 & ~n11016;
  assign n9829 = n11013 & EBX_REG_22__SCAN_IN;
  assign n9831 = ~n9830 & ~n9829;
  assign U2837 = ~n9832 | ~n9831;
  assign n9836 = ~n10031 & ~n11010;
  assign n9834 = ~n10265 | ~n11001;
  assign n9833 = ~n11013 | ~EBX_REG_21__SCAN_IN;
  assign n9835 = ~n9834 | ~n9833;
  assign U2838 = n9836 | n9835;
  assign n9841 = ~n10044 | ~n11020;
  assign n9839 = ~n10291 & ~n11016;
  assign n9838 = ~n11017 & ~n9837;
  assign n9840 = ~n9839 & ~n9838;
  assign U2839 = ~n9841 | ~n9840;
  assign n9846 = ~n10059 & ~n11010;
  assign n9842 = ~n10303;
  assign n9844 = ~n9842 | ~n11001;
  assign n9843 = ~n11013 | ~EBX_REG_19__SCAN_IN;
  assign n9845 = ~n9844 | ~n9843;
  assign U2840 = n9846 | n9845;
  assign n11049 = ~n9847 | ~n9849;
  assign n9856 = ~n9848 | ~n9926;
  assign n9850 = ~n11948 | ~n9849;
  assign n11043 = ~n6994 & ~n9850;
  assign n9852 = ~n11043 | ~DATAI_14_;
  assign n9851 = ~n6994 | ~EAX_REG_30__SCAN_IN;
  assign n9854 = ~n9852 | ~n9851;
  assign n9853 = n11037 & DATAI_30_;
  assign n9855 = ~n9854 & ~n9853;
  assign U2861 = ~n9856 | ~n9855;
  assign n9863 = ~n9857 | ~n9926;
  assign n9859 = ~n11043 | ~DATAI_13_;
  assign n9858 = ~n6994 | ~EAX_REG_29__SCAN_IN;
  assign n9861 = ~n9859 | ~n9858;
  assign n9860 = n11037 & DATAI_29_;
  assign n9862 = ~n9861 & ~n9860;
  assign U2862 = ~n9863 | ~n9862;
  assign n9870 = ~n9864 | ~n9926;
  assign n9866 = ~n11043 | ~DATAI_12_;
  assign n9865 = ~n6994 | ~EAX_REG_28__SCAN_IN;
  assign n9868 = ~n9866 | ~n9865;
  assign n9867 = n11037 & DATAI_28_;
  assign n9869 = ~n9868 & ~n9867;
  assign U2863 = ~n9870 | ~n9869;
  assign n9877 = ~n9871 | ~n9926;
  assign n9873 = ~n11043 | ~DATAI_11_;
  assign n9872 = ~n6994 | ~EAX_REG_27__SCAN_IN;
  assign n9875 = ~n9873 | ~n9872;
  assign n9874 = n11037 & DATAI_27_;
  assign n9876 = ~n9875 & ~n9874;
  assign U2864 = ~n9877 | ~n9876;
  assign n9884 = ~n9878 | ~n9926;
  assign n9880 = ~n11043 | ~DATAI_10_;
  assign n9879 = ~n6994 | ~EAX_REG_26__SCAN_IN;
  assign n9882 = ~n9880 | ~n9879;
  assign n9881 = n11037 & DATAI_26_;
  assign n9883 = ~n9882 & ~n9881;
  assign U2865 = ~n9884 | ~n9883;
  assign n9891 = ~n9885 | ~n9926;
  assign n9887 = ~n11043 | ~DATAI_9_;
  assign n9886 = ~n6994 | ~EAX_REG_25__SCAN_IN;
  assign n9889 = ~n9887 | ~n9886;
  assign n9888 = n11037 & DATAI_25_;
  assign n9890 = ~n9889 & ~n9888;
  assign U2866 = ~n9891 | ~n9890;
  assign n9898 = ~n9892 | ~n9926;
  assign n9894 = ~n11043 | ~DATAI_8_;
  assign n9893 = ~n6994 | ~EAX_REG_24__SCAN_IN;
  assign n9896 = ~n9894 | ~n9893;
  assign n9895 = n11037 & DATAI_24_;
  assign n9897 = ~n9896 & ~n9895;
  assign U2867 = ~n9898 | ~n9897;
  assign n9905 = ~n9899 | ~n9926;
  assign n9901 = ~n11043 | ~DATAI_7_;
  assign n9900 = ~n6994 | ~EAX_REG_23__SCAN_IN;
  assign n9903 = ~n9901 | ~n9900;
  assign n9902 = n11037 & DATAI_23_;
  assign n9904 = ~n9903 & ~n9902;
  assign U2868 = ~n9905 | ~n9904;
  assign n9912 = ~n9906 | ~n9926;
  assign n9908 = ~n11043 | ~DATAI_6_;
  assign n9907 = ~n6994 | ~EAX_REG_22__SCAN_IN;
  assign n9910 = ~n9908 | ~n9907;
  assign n9909 = n11037 & DATAI_22_;
  assign n9911 = ~n9910 & ~n9909;
  assign U2869 = ~n9912 | ~n9911;
  assign n9919 = ~n9913 | ~n9926;
  assign n9915 = ~n11043 | ~DATAI_5_;
  assign n9914 = ~n6994 | ~EAX_REG_21__SCAN_IN;
  assign n9917 = ~n9915 | ~n9914;
  assign n9916 = n11037 & DATAI_21_;
  assign n9918 = ~n9917 & ~n9916;
  assign U2870 = ~n9919 | ~n9918;
  assign n9925 = ~n10044 | ~n9926;
  assign n9921 = ~n11043 | ~DATAI_4_;
  assign n9920 = ~n6994 | ~EAX_REG_20__SCAN_IN;
  assign n9923 = ~n9921 | ~n9920;
  assign n9922 = n11037 & DATAI_20_;
  assign n9924 = ~n9923 & ~n9922;
  assign U2871 = ~n9925 | ~n9924;
  assign n9933 = ~n9927 | ~n9926;
  assign n9929 = ~n11043 | ~DATAI_3_;
  assign n9928 = ~n6994 | ~EAX_REG_19__SCAN_IN;
  assign n9931 = ~n9929 | ~n9928;
  assign n9930 = n11037 & DATAI_19_;
  assign n9932 = ~n9931 & ~n9930;
  assign U2872 = ~n9933 | ~n9932;
  assign n9944 = ~n9934 | ~n11578;
  assign n9942 = ~n9935 & ~n11881;
  assign n9940 = ~n9936 | ~n11548;
  assign n9937 = ~n11581 | ~PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n9939 = n9938 & n9937;
  assign n9941 = ~n9940 | ~n9939;
  assign U2956 = ~n9944 | ~n9943;
  assign n9946 = n10004 ^ ~INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n10187 = n9947 ^ ~n9946;
  assign n9956 = ~n10187 | ~n11578;
  assign n9953 = ~n9949 & ~n11570;
  assign n13584 = ~REIP_REG_28__SCAN_IN;
  assign n10190 = ~n11559 & ~n13584;
  assign n9951 = ~n10190;
  assign n9950 = ~n11581 | ~PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n9952 = ~n9951 | ~n9950;
  assign n9954 = n9953 | n9952;
  assign U2958 = ~n9956 | ~n9955;
  assign n9958 = ~n9957 | ~n9972;
  assign n9962 = ~n9958 | ~n9973;
  assign n9961 = ~n9960 | ~n9959;
  assign n10199 = n9962 ^ ~n9961;
  assign n9971 = ~n10199 | ~n11578;
  assign n9969 = ~n9963 & ~n11881;
  assign n10207 = ~n11576 | ~REIP_REG_27__SCAN_IN;
  assign n9964 = ~n11581 | ~PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n9967 = n10207 & n9964;
  assign n9966 = ~n11548 | ~n9965;
  assign n9968 = ~n9967 | ~n9966;
  assign n9970 = ~n9969 & ~n9968;
  assign U2959 = ~n9971 | ~n9970;
  assign n9974 = ~n9973 | ~n9972;
  assign n9983 = ~n10213 | ~n11578;
  assign n9981 = ~n9975 & ~n11881;
  assign n10215 = ~n11576 | ~REIP_REG_26__SCAN_IN;
  assign n9976 = ~n11581 | ~PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n9979 = n10215 & n9976;
  assign n9978 = ~n9977 | ~n11548;
  assign n9980 = ~n9979 | ~n9978;
  assign n9982 = ~n9981 & ~n9980;
  assign U2960 = ~n9983 | ~n9982;
  assign n9986 = n9985 | n9984;
  assign n10224 = ~n9987 | ~n9986;
  assign n9996 = ~n10224 | ~n11578;
  assign n9994 = ~n9988 & ~n11881;
  assign n10226 = ~n11576 | ~REIP_REG_25__SCAN_IN;
  assign n9989 = ~n11581 | ~PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n9992 = n10226 & n9989;
  assign n9991 = ~n11548 | ~n9990;
  assign n9993 = ~n9992 | ~n9991;
  assign n9995 = ~n9994 & ~n9993;
  assign U2961 = ~n9996 | ~n9995;
  assign n10001 = ~n9997;
  assign n9999 = ~n9998 | ~INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n10000 = ~n9999 & ~n10042;
  assign n10002 = ~n10001 | ~n10000;
  assign n10005 = ~n10003 | ~n10002;
  assign n10017 = n10004 ^ ~INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n10006 = ~n10005 | ~n10017;
  assign n10238 = n10006 ^ ~INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n10016 = ~n10238 | ~n11578;
  assign n10014 = ~n10007 & ~n11881;
  assign n10244 = ~n11576 | ~REIP_REG_23__SCAN_IN;
  assign n10009 = ~n10244;
  assign n10008 = ~n11530 & ~n9688;
  assign n10012 = ~n10009 & ~n10008;
  assign n10011 = ~n11548 | ~n10010;
  assign n10013 = ~n10012 | ~n10011;
  assign n10015 = ~n10014 & ~n10013;
  assign U2963 = ~n10016 | ~n10015;
  assign n10250 = n10018 ^ ~n10017;
  assign n10028 = ~n10250 | ~n11578;
  assign n10026 = ~n10019 & ~n11881;
  assign n13553 = ~REIP_REG_22__SCAN_IN;
  assign n10252 = ~n11559 & ~n13553;
  assign n10021 = ~n10252;
  assign n10020 = ~n11581 | ~PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n10024 = n10021 & n10020;
  assign n10023 = ~n11548 | ~n10022;
  assign n10025 = ~n10024 | ~n10023;
  assign n10027 = ~n10026 & ~n10025;
  assign U2964 = ~n10028 | ~n10027;
  assign n10264 = n10029 ^ ~n10030;
  assign n10040 = ~n10264 | ~n11578;
  assign n10038 = ~n10031 & ~n11881;
  assign n10266 = ~n11576 | ~REIP_REG_21__SCAN_IN;
  assign n10033 = ~n10266;
  assign n10032 = ~n11530 & ~n9728;
  assign n10036 = ~n10033 & ~n10032;
  assign n10035 = ~n11548 | ~n10034;
  assign n10037 = ~n10036 | ~n10035;
  assign n10039 = ~n10038 & ~n10037;
  assign U2965 = ~n10040 | ~n10039;
  assign n10043 = ~n10042 & ~n10041;
  assign n10277 = n10043 ^ n9997;
  assign n10055 = ~n10277 & ~n11567;
  assign n10053 = ~n10044 | ~n6996;
  assign n10045 = ~REIP_REG_20__SCAN_IN;
  assign n10296 = ~n11559 & ~n10045;
  assign n10047 = ~n10296;
  assign n10046 = ~n11581 | ~PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n10051 = ~n10047 | ~n10046;
  assign n10049 = ~n10048;
  assign n10050 = ~n11570 & ~n10049;
  assign n10052 = ~n10051 & ~n10050;
  assign n10054 = ~n10053 | ~n10052;
  assign U2966 = n10055 | n10054;
  assign n10302 = ~n10058 | ~n10057;
  assign n10067 = ~n10302 | ~n11578;
  assign n10065 = ~n10059 & ~n11881;
  assign n10305 = ~n11576 | ~REIP_REG_19__SCAN_IN;
  assign n10060 = ~n11581 | ~PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n10063 = n10305 & n10060;
  assign n10062 = ~n11548 | ~n10061;
  assign n10064 = ~n10063 | ~n10062;
  assign n10066 = ~n10065 & ~n10064;
  assign U2967 = ~n10067 | ~n10066;
  assign n10069 = ~n10116;
  assign n10101 = ~n10070 | ~n10071;
  assign n10072 = ~n9041 & ~n10337;
  assign n10076 = ~n10091 | ~n10072;
  assign n10073 = ~n10089 & ~INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n10075 = ~n10074 | ~n10073;
  assign n10077 = ~n10076 | ~n10075;
  assign n10313 = n10077 ^ ~n10321;
  assign n10088 = ~n10313 | ~n11578;
  assign n10080 = ~n10078 & ~n10079;
  assign n10534 = ~n8478 & ~n10080;
  assign n10086 = ~n10534 | ~n6996;
  assign n10327 = n11576 & REIP_REG_18__SCAN_IN;
  assign n10082 = ~n10327;
  assign n10081 = ~n11581 | ~PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n10084 = ~n10082 | ~n10081;
  assign n10083 = ~n11570 & ~n10537;
  assign n10085 = ~n10084 & ~n10083;
  assign n10087 = n10086 & n10085;
  assign U2968 = ~n10088 | ~n10087;
  assign n10090 = n10089 ^ ~n10337;
  assign n10335 = n10091 ^ ~n10090;
  assign n10100 = ~n10335 | ~n11578;
  assign n11032 = n10092 ^ ~n10093;
  assign n10098 = ~n11032 & ~n11881;
  assign n10342 = ~n11576 | ~REIP_REG_17__SCAN_IN;
  assign n10094 = ~n11581 | ~PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n10096 = n10342 & n10094;
  assign n10095 = ~n11548 | ~n10555;
  assign n10097 = ~n10096 | ~n10095;
  assign n10099 = ~n10098 & ~n10097;
  assign U2969 = ~n10100 | ~n10099;
  assign n10348 = n10102 ^ ~n10101;
  assign n10113 = ~n10348 | ~n11578;
  assign n10105 = ~n10103 | ~n10104;
  assign n11040 = ~n10092 | ~n10105;
  assign n10111 = ~n11040 & ~n11881;
  assign n10362 = n11576 & REIP_REG_16__SCAN_IN;
  assign n10107 = ~n10362;
  assign n10106 = ~n11581 | ~PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n10109 = ~n10107 | ~n10106;
  assign n10108 = ~n11570 & ~n10571;
  assign n10110 = n10109 | n10108;
  assign n10112 = ~n10111 & ~n10110;
  assign U2970 = ~n10113 | ~n10112;
  assign n10131 = ~n10146 | ~n7157;
  assign n10130 = n10114 & n10115;
  assign n10129 = ~n10131 | ~n10130;
  assign n10119 = ~n10129 | ~n10115;
  assign n10118 = ~n10117 | ~n10116;
  assign n10369 = n10119 ^ ~n10118;
  assign n10122 = ~n10120 | ~n10121;
  assign n10587 = n10103 & n10122;
  assign n10128 = ~n10587 | ~n6996;
  assign n10381 = ~n11559 & ~n13519;
  assign n10124 = ~n10381;
  assign n10123 = ~n11581 | ~PHYADDRPOINTER_REG_15__SCAN_IN;
  assign n10126 = ~n10124 | ~n10123;
  assign n10125 = ~n11570 & ~n10590;
  assign n10127 = ~n10126 & ~n10125;
  assign n10133 = ~n10129;
  assign n10132 = ~n10131 & ~n10130;
  assign n10386 = ~n10133 & ~n10132;
  assign n10142 = n10386 | n11567;
  assign n11052 = n10134 ^ ~n10135;
  assign n10140 = ~n11052 & ~n11881;
  assign n10412 = ~n11576 | ~REIP_REG_14__SCAN_IN;
  assign n10136 = ~n11581 | ~PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n10138 = n10412 & n10136;
  assign n10137 = ~n11548 | ~n10605;
  assign n10139 = ~n10138 | ~n10137;
  assign n10141 = ~n10140 & ~n10139;
  assign U2972 = ~n10142 | ~n10141;
  assign n10145 = ~n10144 | ~n10143;
  assign n10417 = ~n10146 | ~n10145;
  assign n10157 = ~n10417 | ~n11578;
  assign n10150 = ~n10148 | ~n10147;
  assign n10961 = n10150 ^ ~n10149;
  assign n11057 = ~n10961;
  assign n10155 = ~n11057 & ~n11881;
  assign n10423 = ~n11576 | ~REIP_REG_13__SCAN_IN;
  assign n10151 = ~n11581 | ~PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n10153 = n10423 & n10151;
  assign n10152 = ~n11548 | ~n10624;
  assign n10154 = ~n10153 | ~n10152;
  assign n10156 = ~n10155 & ~n10154;
  assign U2973 = ~n10157 | ~n10156;
  assign n10172 = ~n10158 | ~n11803;
  assign n10164 = ~n10927 & ~n11792;
  assign n10160 = ~n10159 | ~INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n10162 = INSTADDRPOINTER_REG_31__SCAN_IN | n10160;
  assign n10163 = ~n10162 | ~n10161;
  assign n10170 = ~n10164 & ~n10163;
  assign n10166 = ~n10165 | ~n11780;
  assign n10168 = ~n10167 | ~n10166;
  assign n10169 = ~INSTADDRPOINTER_REG_31__SCAN_IN | ~n10168;
  assign n10171 = n10170 & n10169;
  assign U2987 = ~n10172 | ~n10171;
  assign n10186 = ~n10173 | ~n11803;
  assign n10175 = ~n10174;
  assign n10177 = ~n10175 | ~n11739;
  assign n10184 = ~n10177 | ~n10176;
  assign n10182 = ~n10178 & ~n9384;
  assign n10180 = ~n10179;
  assign n10181 = ~n10180 & ~INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n10183 = ~n10182 & ~n10181;
  assign n10185 = ~n10184 & ~n10183;
  assign U2989 = ~n10186 | ~n10185;
  assign n10198 = ~n10187 | ~n11803;
  assign n10192 = ~n10188 | ~n11739;
  assign n10189 = ~n10200 & ~n10193;
  assign n10191 = ~n10190 & ~n10189;
  assign n10196 = ~n10192 | ~n10191;
  assign n10194 = n10193 ^ ~INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n10195 = n10203 & n10194;
  assign n10197 = ~n10196 & ~n10195;
  assign U2990 = ~n10198 | ~n10197;
  assign n10212 = ~n10199 | ~n11803;
  assign n10202 = ~n10200;
  assign n10205 = ~n10202 & ~n10201;
  assign n10204 = ~n10203 & ~INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n10210 = ~n10205 & ~n10204;
  assign n10208 = ~n10206 | ~n11739;
  assign n10209 = ~n10208 | ~n10207;
  assign n10211 = ~n10210 & ~n10209;
  assign U2991 = ~n10212 | ~n10211;
  assign n10223 = ~n10213 | ~n11803;
  assign n10216 = ~n10214 | ~n11739;
  assign n10219 = ~n10216 | ~n10215;
  assign n10217 = INSTADDRPOINTER_REG_25__SCAN_IN ^ ~INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n10218 = ~n10230 & ~n10217;
  assign n10221 = ~n10219 & ~n10218;
  assign n10220 = ~n10229 | ~INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n10222 = n10221 & n10220;
  assign U2992 = ~n10223 | ~n10222;
  assign n10237 = ~n10224 | ~n11803;
  assign n10227 = ~n10225 | ~n11739;
  assign n10235 = ~n10227 | ~n10226;
  assign n10233 = ~n10229 & ~n10228;
  assign n10231 = ~n10230;
  assign n10232 = ~n10231 & ~INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n10234 = ~n10233 & ~n10232;
  assign n10236 = ~n10235 & ~n10234;
  assign U2993 = ~n10237 | ~n10236;
  assign n10249 = ~n10238 | ~n11803;
  assign n10242 = n10239 & INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n10241 = ~n10240 & ~INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n10247 = ~n10242 & ~n10241;
  assign n10245 = ~n10243 | ~n11739;
  assign n10246 = ~n10245 | ~n10244;
  assign n10248 = ~n10247 & ~n10246;
  assign U2995 = ~n10249 | ~n10248;
  assign n10263 = ~n10250 | ~n11803;
  assign n10253 = ~n10251 & ~n11792;
  assign n10255 = ~n10253 & ~n10252;
  assign n10254 = ~n10269 | ~INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n10261 = ~n10255 | ~n10254;
  assign n10257 = ~n10256 | ~n10268;
  assign n10258 = ~n10270 | ~n10257;
  assign n10260 = ~n10259 & ~n10258;
  assign n10262 = ~n10261 & ~n10260;
  assign U2996 = ~n10263 | ~n10262;
  assign n10276 = ~n10264 | ~n11803;
  assign n10267 = ~n10265 | ~n11739;
  assign n10274 = ~n10267 | ~n10266;
  assign n10272 = ~n10269 & ~n10268;
  assign n10271 = ~n10270 & ~INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n10273 = ~n10272 & ~n10271;
  assign n10275 = ~n10274 & ~n10273;
  assign U2997 = ~n10276 | ~n10275;
  assign n10301 = ~n10277 & ~n11784;
  assign n10319 = ~n11765 | ~n10315;
  assign n10279 = n11732 | n10278;
  assign n10336 = ~n10319 | ~n10279;
  assign n10292 = ~n10336 | ~n10280;
  assign n10310 = n10292 | INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n11771 = ~INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n10281 = ~n11771 & ~n10283;
  assign n10282 = ~n10390 & ~n10281;
  assign n10285 = ~n11795 & ~n10282;
  assign n10284 = ~n10283 | ~n11796;
  assign n10288 = n10285 & n10284;
  assign n10287 = ~n11772 | ~n10286;
  assign n10304 = ~n10288 | ~n10287;
  assign n10289 = ~n10304;
  assign n10290 = ~n10310 | ~n10289;
  assign n10299 = ~n10290 | ~INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n10295 = n10291 | n11792;
  assign n10293 = ~INSTADDRPOINTER_REG_20__SCAN_IN & ~n10292;
  assign n10294 = ~INSTADDRPOINTER_REG_19__SCAN_IN | ~n10293;
  assign n10297 = ~n10295 | ~n10294;
  assign n10298 = ~n10297 & ~n10296;
  assign n10300 = ~n10299 | ~n10298;
  assign U2998 = n10301 | n10300;
  assign n10312 = n10302 & n11803;
  assign n10308 = n10303 | n11792;
  assign n10306 = ~INSTADDRPOINTER_REG_19__SCAN_IN | ~n10304;
  assign n10307 = n10306 & n10305;
  assign n10309 = n10308 & n10307;
  assign n10311 = ~n10310 | ~n10309;
  assign U2999 = n10312 | n10311;
  assign n10334 = ~n10313 | ~n11803;
  assign n10317 = ~n10314 & ~n11732;
  assign n10316 = ~n11663 & ~n10315;
  assign n10318 = ~n10317 & ~n10316;
  assign n10338 = ~n11773 | ~n10318;
  assign n10320 = ~INSTADDRPOINTER_REG_17__SCAN_IN & ~n10319;
  assign n10322 = ~n10338 & ~n10320;
  assign n10332 = ~n10322 & ~n10321;
  assign n10323 = ~INSTADDRPOINTER_REG_18__SCAN_IN & ~n10337;
  assign n10330 = ~n10336 | ~n10323;
  assign n10326 = ~n10325 & ~n10324;
  assign n10931 = n9766 | n10326;
  assign n10328 = ~n10931 & ~n11792;
  assign n10329 = ~n10328 & ~n10327;
  assign n10331 = ~n10330 | ~n10329;
  assign n10333 = ~n10332 & ~n10331;
  assign U3000 = ~n10334 | ~n10333;
  assign n10347 = ~n10335 | ~n11803;
  assign n10340 = ~n10336 & ~INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n10339 = ~n10338 & ~n10337;
  assign n10345 = ~n10340 & ~n10339;
  assign n10936 = n10341 ^ n10360;
  assign n10343 = ~n10936 | ~n11739;
  assign n10344 = ~n10343 | ~n10342;
  assign n10346 = ~n10345 & ~n10344;
  assign U3001 = ~n10347 | ~n10346;
  assign n10368 = ~n10348 | ~n11803;
  assign n11598 = ~n11625 & ~n10349;
  assign n10398 = n11772 & n11599;
  assign n11612 = ~n11598 & ~n10398;
  assign n10350 = ~n10387;
  assign n10351 = ~n10350 | ~INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n10371 = n11612 | n10351;
  assign n10352 = INSTADDRPOINTER_REG_15__SCAN_IN ^ ~INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n10366 = ~n10371 & ~n10352;
  assign n11629 = ~n11773;
  assign n10354 = ~n10353 & ~n11732;
  assign n10357 = ~n11629 & ~n10354;
  assign n10356 = ~n11689 | ~n10355;
  assign n10372 = ~n10357 | ~n10356;
  assign n10364 = ~n10372 | ~INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n10359 = ~n10379 | ~n10358;
  assign n10942 = ~n10360 | ~n10359;
  assign n10361 = ~n10942 & ~n11792;
  assign n10363 = ~n10362 & ~n10361;
  assign n10365 = ~n10364 | ~n10363;
  assign n10367 = ~n10366 & ~n10365;
  assign U3002 = ~n10368 | ~n10367;
  assign n10385 = ~n10369 & ~n11784;
  assign n10375 = ~n10371 | ~n10370;
  assign n10373 = ~n10372;
  assign n10374 = ~n10373 | ~INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n10383 = ~n10375 | ~n10374;
  assign n10378 = n10377 | n10376;
  assign n10947 = ~n10379 | ~n10378;
  assign n10380 = ~n11792 & ~n10947;
  assign n10382 = ~n10381 & ~n10380;
  assign n10384 = ~n10383 | ~n10382;
  assign U3003 = n10385 | n10384;
  assign n10416 = ~n10386 & ~n11784;
  assign n10388 = n11612 | n10387;
  assign n10407 = ~n10388 | ~n10397;
  assign n10389 = ~n11599 | ~n10399;
  assign n10393 = ~n10389 | ~n11772;
  assign n10425 = ~n11602 | ~n10399;
  assign n10401 = ~n11771 & ~n10425;
  assign n10391 = ~n10401 & ~n10390;
  assign n10392 = ~n11795 & ~n10391;
  assign n10396 = n10393 & n10392;
  assign n10395 = ~n10394;
  assign n10426 = ~n11796 | ~n10395;
  assign n10418 = ~n10396 | ~n10426;
  assign n10405 = ~n10418 & ~n10397;
  assign n10403 = ~n10399 | ~n10398;
  assign n10402 = ~n10401 | ~n10400;
  assign n10419 = ~n10403 | ~n10402;
  assign n10404 = ~n10419 | ~n7161;
  assign n10406 = ~n10405 | ~n10404;
  assign n10414 = ~n10407 | ~n10406;
  assign n10409 = ~n10408;
  assign n10952 = n10410 ^ ~n10409;
  assign n10411 = ~n10952 | ~n11739;
  assign n10413 = n10412 & n10411;
  assign n10415 = ~n10414 | ~n10413;
  assign U3004 = n10416 | n10415;
  assign n10432 = ~n10417 | ~n11803;
  assign n10421 = ~n10418 & ~n7161;
  assign n10420 = ~n10419 & ~INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n10430 = ~n10421 & ~n10420;
  assign n10958 = n10422 ^ n10647;
  assign n10424 = ~n11739 | ~n10958;
  assign n10428 = ~n10424 | ~n10423;
  assign n10427 = ~n10426 & ~n10425;
  assign n10429 = n10428 | n10427;
  assign n10431 = ~n10430 & ~n10429;
  assign U3005 = ~n10432 | ~n10431;
  assign n10433 = ~n11828;
  assign n10435 = ~n13342 & ~n10433;
  assign n10437 = ~n10435 & ~n10434;
  assign n10436 = ~n9142 | ~n13742;
  assign n10438 = ~n10437 | ~n10436;
  assign n10441 = ~n13325 & ~n10438;
  assign n10440 = ~n10439;
  assign n10442 = ~n10441 & ~n10440;
  assign n10447 = ~READY_N & ~n10442;
  assign n10445 = ~n10443;
  assign n10444 = ~n13743 | ~n11918;
  assign n10446 = ~n10445 | ~n10444;
  assign n10449 = ~n10447 & ~n10446;
  assign n10450 = ~n10449 | ~n10448;
  assign n13350 = ~n10451 & ~n10450;
  assign n10454 = n13350 | n13404;
  assign n11810 = ~FLUSH_REG_SCAN_IN;
  assign n10452 = ~n13304;
  assign n13618 = ~n10452 | ~STATE2_REG_0__SCAN_IN;
  assign n10453 = n11810 | n13618;
  assign n10462 = ~n10454 | ~n10453;
  assign n10455 = n13400 & STATE2_REG_3__SCAN_IN;
  assign n10464 = ~n13662 | ~INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n10458 = ~n10457 & ~n10456;
  assign n11868 = n10458 ^ ~n11873;
  assign n10460 = ~n11868;
  assign n10459 = ~n11867 | ~n13402;
  assign n10461 = ~n10460 & ~n10459;
  assign n10463 = ~n10462 | ~n10461;
  assign U3455 = ~n10464 | ~n10463;
  assign n13439 = ~STATE_REG_0__SCAN_IN;
  assign n10465 = ~STATE_REG_2__SCAN_IN & ~n13433;
  assign n10466 = ~ADS_N_REG_SCAN_IN & ~n10477;
  assign U2789 = ~n13757 & ~n10466;
  assign n10473 = ~STATE2_REG_0__SCAN_IN | ~n13762;
  assign n10470 = n11806 | n10793;
  assign n10467 = ~n13320;
  assign n10468 = ~n13321 | ~n10467;
  assign n10469 = ~n10468 | ~n9142;
  assign n10471 = ~n10484 | ~n13390;
  assign n10472 = ~CODEFETCH_REG_SCAN_IN | ~n10471;
  assign U2790 = ~n10473 | ~n10472;
  assign n10478 = ~STATE_REG_2__SCAN_IN & ~STATE_REG_0__SCAN_IN;
  assign n10474 = ~n10478 & ~D_C_N_REG_SCAN_IN;
  assign n10476 = ~n13757 & ~n10474;
  assign n13756 = ~n13757;
  assign n10475 = ~CODEFETCH_REG_SCAN_IN & ~n13756;
  assign U2791 = n10476 | n10475;
  assign n13610 = ~n13415;
  assign n10479 = BS16_N | n10478;
  assign n13615 = ~n13610 | ~n10479;
  assign n13613 = ~n13610;
  assign n10480 = ~STATEBS16_REG_SCAN_IN | ~n13613;
  assign U2792 = ~n13615 | ~n10480;
  assign n10482 = n13739 | n13760;
  assign n10483 = ~n13431 | ~n10482;
  assign n13307 = ~n10484 | ~n10483;
  assign n13731 = ~n13307 | ~n13390;
  assign n10485 = ~FLUSH_REG_SCAN_IN | ~n13731;
  assign U2793 = ~n11567 | ~n10485;
  assign n13713 = ~DATAWIDTH_REG_0__SCAN_IN & ~DATAWIDTH_REG_1__SCAN_IN;
  assign n13723 = ~REIP_REG_0__SCAN_IN;
  assign n10519 = ~n13713 | ~n13723;
  assign n10516 = ~n10519 | ~n13722;
  assign n10487 = ~DATAWIDTH_REG_20__SCAN_IN & ~DATAWIDTH_REG_21__SCAN_IN;
  assign n10486 = ~DATAWIDTH_REG_22__SCAN_IN & ~DATAWIDTH_REG_23__SCAN_IN;
  assign n10491 = ~n10487 | ~n10486;
  assign n10489 = ~DATAWIDTH_REG_16__SCAN_IN & ~DATAWIDTH_REG_17__SCAN_IN;
  assign n10488 = ~DATAWIDTH_REG_18__SCAN_IN & ~DATAWIDTH_REG_19__SCAN_IN;
  assign n10490 = ~n10489 | ~n10488;
  assign n10499 = ~n10491 & ~n10490;
  assign n10493 = ~DATAWIDTH_REG_28__SCAN_IN & ~DATAWIDTH_REG_29__SCAN_IN;
  assign n10492 = ~DATAWIDTH_REG_30__SCAN_IN & ~DATAWIDTH_REG_31__SCAN_IN;
  assign n10497 = ~n10493 | ~n10492;
  assign n10495 = ~DATAWIDTH_REG_24__SCAN_IN & ~DATAWIDTH_REG_25__SCAN_IN;
  assign n10494 = ~DATAWIDTH_REG_26__SCAN_IN & ~DATAWIDTH_REG_27__SCAN_IN;
  assign n10496 = ~n10495 | ~n10494;
  assign n10498 = ~n10497 & ~n10496;
  assign n10515 = ~n10499 | ~n10498;
  assign n10501 = ~DATAWIDTH_REG_4__SCAN_IN & ~DATAWIDTH_REG_5__SCAN_IN;
  assign n10500 = ~DATAWIDTH_REG_6__SCAN_IN & ~DATAWIDTH_REG_7__SCAN_IN;
  assign n10505 = ~n10501 | ~n10500;
  assign n10503 = ~DATAWIDTH_REG_2__SCAN_IN & ~DATAWIDTH_REG_3__SCAN_IN;
  assign n10502 = ~DATAWIDTH_REG_0__SCAN_IN | ~DATAWIDTH_REG_1__SCAN_IN;
  assign n10504 = ~n10503 | ~n10502;
  assign n10513 = ~n10505 & ~n10504;
  assign n10507 = ~DATAWIDTH_REG_12__SCAN_IN & ~DATAWIDTH_REG_13__SCAN_IN;
  assign n10506 = ~DATAWIDTH_REG_14__SCAN_IN & ~DATAWIDTH_REG_15__SCAN_IN;
  assign n10511 = ~n10507 | ~n10506;
  assign n10509 = ~DATAWIDTH_REG_8__SCAN_IN & ~DATAWIDTH_REG_9__SCAN_IN;
  assign n10508 = ~DATAWIDTH_REG_10__SCAN_IN & ~DATAWIDTH_REG_11__SCAN_IN;
  assign n10510 = ~n10509 | ~n10508;
  assign n10512 = ~n10511 & ~n10510;
  assign n10514 = ~n10513 | ~n10512;
  assign n13724 = ~n10515 & ~n10514;
  assign n10518 = ~n10516 | ~n13724;
  assign n13726 = ~n13724;
  assign n10517 = ~BYTEENABLE_REG_1__SCAN_IN | ~n13726;
  assign U2794 = ~n10518 | ~n10517;
  assign n10523 = ~BYTEENABLE_REG_3__SCAN_IN | ~n13726;
  assign n10520 = DATAWIDTH_REG_1__SCAN_IN | REIP_REG_1__SCAN_IN;
  assign n10521 = ~n10520 | ~n10519;
  assign n10522 = ~n10521 | ~n13724;
  assign U2795 = ~n10523 | ~n10522;
  assign n10524 = n10896 & PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n10529 = ~n10784 & ~n10524;
  assign n10526 = ~n10525;
  assign n10528 = ~n10527 | ~n10526;
  assign n10531 = ~n10529 | ~n10528;
  assign n10530 = ~n13534 & ~n10545;
  assign n10533 = ~n10531 & ~n10530;
  assign n10532 = ~EBX_REG_18__SCAN_IN | ~n10904;
  assign n10536 = ~n10533 | ~n10532;
  assign n11025 = ~n10534;
  assign n10535 = ~n11025 & ~n10795;
  assign n10541 = ~n10536 & ~n10535;
  assign n10539 = ~n10931 & ~n10914;
  assign n10538 = ~n10908 & ~n10537;
  assign n10540 = ~n10539 & ~n10538;
  assign U2809 = ~n10541 | ~n10540;
  assign n10543 = ~n10830 & ~n10542;
  assign n10544 = ~REIP_REG_17__SCAN_IN & ~n10543;
  assign n10549 = ~n10545 & ~n10544;
  assign n10547 = ~n10904 | ~EBX_REG_17__SCAN_IN;
  assign n10546 = ~n10896 | ~PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n10548 = ~n10547 | ~n10546;
  assign n10550 = ~n10549 & ~n10548;
  assign n10554 = ~n10550 | ~n10814;
  assign n10939 = ~n11032;
  assign n10552 = ~n10939 | ~n10770;
  assign n10551 = ~n10936 | ~n10837;
  assign n10553 = ~n10552 | ~n10551;
  assign n10557 = ~n10554 & ~n10553;
  assign n10556 = ~n10555 | ~n10869;
  assign U2810 = ~n10557 | ~n10556;
  assign n10596 = n10582 & n10851;
  assign n10578 = ~n10831 & ~n10596;
  assign n10581 = ~n10851 | ~n13519;
  assign n10558 = ~n10578 | ~n10581;
  assign n10568 = ~n10558 | ~REIP_REG_16__SCAN_IN;
  assign n10560 = ~n10907 & ~n10559;
  assign n10562 = ~n10784 & ~n10560;
  assign n10561 = ~EBX_REG_16__SCAN_IN | ~n10904;
  assign n10566 = ~n10562 | ~n10561;
  assign n10564 = ~n10563 | ~n10851;
  assign n10565 = ~REIP_REG_16__SCAN_IN & ~n10564;
  assign n10567 = ~n10566 & ~n10565;
  assign n10570 = ~n10568 | ~n10567;
  assign n10569 = ~n11040 & ~n10795;
  assign n10575 = ~n10570 & ~n10569;
  assign n10573 = ~n10914 & ~n10942;
  assign n10572 = ~n7011 & ~n10571;
  assign n10574 = ~n10573 & ~n10572;
  assign U2811 = ~n10575 | ~n10574;
  assign n10577 = ~n10907 & ~n10576;
  assign n10586 = ~n10784 & ~n10577;
  assign n10580 = ~EBX_REG_15__SCAN_IN | ~n10904;
  assign n10598 = ~n10578;
  assign n10579 = ~REIP_REG_15__SCAN_IN | ~n10598;
  assign n10584 = ~n10580 | ~n10579;
  assign n10583 = ~n10582 & ~n10581;
  assign n10585 = ~n10584 & ~n10583;
  assign n10589 = ~n10586 | ~n10585;
  assign n10588 = ~n11046 & ~n10795;
  assign n10594 = ~n10589 & ~n10588;
  assign n10592 = ~n10914 & ~n10947;
  assign n10591 = ~n10908 & ~n10590;
  assign n10593 = ~n10592 & ~n10591;
  assign U2812 = ~n10594 | ~n10593;
  assign n10595 = ~n10896 | ~PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n10602 = ~n10814 | ~n10595;
  assign n10600 = ~n10597 | ~n10596;
  assign n10599 = ~REIP_REG_14__SCAN_IN | ~n10598;
  assign n10601 = ~n10600 | ~n10599;
  assign n10604 = ~n10602 & ~n10601;
  assign n10603 = ~EBX_REG_14__SCAN_IN | ~n10904;
  assign n10609 = ~n10604 | ~n10603;
  assign n10955 = ~n11052;
  assign n10607 = ~n10955 | ~n10770;
  assign n10606 = ~n10869 | ~n10605;
  assign n10608 = ~n10607 | ~n10606;
  assign n10611 = ~n10609 & ~n10608;
  assign n10610 = ~n10837 | ~n10952;
  assign U2813 = ~n10611 | ~n10610;
  assign n13504 = ~REIP_REG_12__SCAN_IN;
  assign n10632 = ~n10851 | ~n13504;
  assign n10633 = ~n10612;
  assign n10658 = ~n10633 | ~n10851;
  assign n10653 = n10893 & n10658;
  assign n10613 = ~n10632 | ~n10653;
  assign n10617 = ~n10613 | ~REIP_REG_13__SCAN_IN;
  assign n10615 = ~n10907 & ~n10614;
  assign n10616 = ~n10784 & ~n10615;
  assign n10621 = ~n10617 | ~n10616;
  assign n10618 = ~n10851 | ~n13509;
  assign n10620 = ~n10619 & ~n10618;
  assign n10623 = ~n10621 & ~n10620;
  assign n10622 = ~EBX_REG_13__SCAN_IN | ~n10904;
  assign n10628 = ~n10623 | ~n10622;
  assign n10626 = ~n10624 | ~n10869;
  assign n10625 = ~n10770 | ~n10961;
  assign n10627 = ~n10626 | ~n10625;
  assign n10630 = ~n10628 & ~n10627;
  assign n10629 = ~n10837 | ~n10958;
  assign U2814 = ~n10630 | ~n10629;
  assign n10631 = ~n10896 | ~PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n10635 = ~n10814 | ~n10631;
  assign n10634 = ~n10633 & ~n10632;
  assign n10637 = ~n10635 & ~n10634;
  assign n10636 = ~EBX_REG_12__SCAN_IN | ~n10904;
  assign n10639 = ~n10637 | ~n10636;
  assign n10638 = ~n10653 & ~n13504;
  assign n10651 = ~n10639 & ~n10638;
  assign n10640 = ~n7040 | ~n10662;
  assign n11062 = n10641 ^ n10640;
  assign n11415 = ~n11062;
  assign n10643 = ~n11415 | ~n10770;
  assign n10642 = n10908 | n11412;
  assign n10649 = ~n10643 | ~n10642;
  assign n10646 = ~n10644 | ~n10645;
  assign n11589 = ~n10647 | ~n10646;
  assign n10648 = ~n10914 & ~n11589;
  assign n10650 = ~n10649 & ~n10648;
  assign U2815 = ~n10651 | ~n10650;
  assign n10652 = ~n10896 | ~PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n10655 = ~n10814 | ~n10652;
  assign n10654 = ~n10653 & ~n13499;
  assign n10657 = ~n10655 & ~n10654;
  assign n10656 = ~EBX_REG_11__SCAN_IN | ~n10904;
  assign n10661 = ~n10657 | ~n10656;
  assign n10660 = ~n10659 & ~n10658;
  assign n10671 = ~n10661 & ~n10660;
  assign n11067 = n7040 ^ ~n10662;
  assign n11443 = ~n11067;
  assign n10664 = ~n11443 | ~n10770;
  assign n10663 = ~n10869 | ~n11430;
  assign n10669 = ~n10664 | ~n10663;
  assign n10667 = n10666 | n10665;
  assign n11609 = ~n10644 | ~n10667;
  assign n10668 = ~n10914 & ~n11609;
  assign n10670 = ~n10669 & ~n10668;
  assign U2816 = ~n10671 | ~n10670;
  assign n10692 = ~n10851 | ~n13489;
  assign n10723 = n10693 & n10851;
  assign n10714 = ~n10831 & ~n10723;
  assign n10672 = ~n10692 | ~n10714;
  assign n10691 = ~n10672 | ~REIP_REG_10__SCAN_IN;
  assign n10673 = ~n10896 | ~PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n10677 = ~n10814 | ~n10673;
  assign n11622 = n10674 ^ ~n10675;
  assign n10676 = ~n10914 & ~n11622;
  assign n10679 = ~n10677 & ~n10676;
  assign n10678 = ~EBX_REG_10__SCAN_IN | ~n10904;
  assign n10683 = ~n10679 | ~n10678;
  assign n10681 = ~n10680 | ~n10851;
  assign n10682 = ~REIP_REG_10__SCAN_IN & ~n10681;
  assign n10687 = ~n10683 & ~n10682;
  assign n11072 = n10684 ^ ~n10685;
  assign n11449 = ~n11072;
  assign n10686 = ~n11449 | ~n10770;
  assign n10689 = ~n10687 | ~n10686;
  assign n10688 = ~n11446 & ~n7011;
  assign n10690 = ~n10689 & ~n10688;
  assign U2817 = ~n10691 | ~n10690;
  assign n10698 = ~n10693 & ~n10692;
  assign n10696 = ~n10674;
  assign n10695 = ~n7021 | ~n10694;
  assign n11640 = ~n10696 | ~n10695;
  assign n10697 = ~n11640 & ~n10914;
  assign n10711 = ~n10698 & ~n10697;
  assign n10700 = ~n10904 | ~EBX_REG_9__SCAN_IN;
  assign n10699 = ~n10896 | ~PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n10702 = ~n10700 | ~n10699;
  assign n10701 = ~n10714 & ~n13489;
  assign n10703 = ~n10702 & ~n10701;
  assign n10709 = ~n10703 | ~n10814;
  assign n11077 = n10705 ^ ~n10704;
  assign n11468 = ~n11077;
  assign n10707 = ~n11468 | ~n10770;
  assign n10706 = ~n10869 | ~n11463;
  assign n10708 = ~n10707 | ~n10706;
  assign n10710 = ~n10709 & ~n10708;
  assign U2818 = ~n10711 | ~n10710;
  assign n10713 = ~n10904 | ~EBX_REG_8__SCAN_IN;
  assign n10712 = ~n10896 | ~PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n10716 = ~n10713 | ~n10712;
  assign n13484 = ~REIP_REG_8__SCAN_IN;
  assign n10715 = ~n10714 & ~n13484;
  assign n10717 = ~n10716 & ~n10715;
  assign n10721 = ~n10717 | ~n10814;
  assign n10719 = n7030 | n10718;
  assign n11474 = n10704 & n10719;
  assign n11082 = ~n11474;
  assign n10720 = ~n11082 & ~n10795;
  assign n10731 = ~n10721 & ~n10720;
  assign n10727 = ~n10723 | ~n10722;
  assign n11653 = n10725 ^ n10724;
  assign n10726 = ~n11653 | ~n10837;
  assign n10729 = ~n10727 | ~n10726;
  assign n10728 = ~n11471 & ~n10908;
  assign n10730 = ~n10729 & ~n10728;
  assign U2819 = ~n10731 | ~n10730;
  assign n10733 = ~n10907 & ~n10732;
  assign n10743 = ~n10784 & ~n10733;
  assign n11672 = n10735 ^ n10734;
  assign n10737 = ~n11672 | ~n10837;
  assign n10736 = ~n10904 | ~EBX_REG_7__SCAN_IN;
  assign n10741 = ~n10737 | ~n10736;
  assign n10738 = ~n10851 | ~n13479;
  assign n10740 = ~n10739 & ~n10738;
  assign n10742 = ~n10741 & ~n10740;
  assign n10748 = ~n10743 | ~n10742;
  assign n10746 = ~n10744 & ~n10745;
  assign n10747 = ~n11488 & ~n10795;
  assign n10754 = ~n10748 & ~n10747;
  assign n10910 = ~n10831 & ~n10851;
  assign n10749 = n10893 & n10760;
  assign n10777 = ~n10910 & ~n10749;
  assign n10761 = ~REIP_REG_6__SCAN_IN & ~n10830;
  assign n10750 = ~n10777 & ~n10761;
  assign n10752 = ~n13479 & ~n10750;
  assign n10751 = ~n10908 & ~n11487;
  assign n10753 = ~n10752 & ~n10751;
  assign U2820 = ~n10754 | ~n10753;
  assign n10756 = ~n10904 | ~EBX_REG_6__SCAN_IN;
  assign n10755 = ~n10896 | ~PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n10759 = ~n10756 | ~n10755;
  assign n10757 = ~REIP_REG_6__SCAN_IN | ~n10777;
  assign n10758 = ~n10814 | ~n10757;
  assign n10776 = ~n10759 & ~n10758;
  assign n10764 = ~n10761 | ~n10760;
  assign n11685 = n10762 ^ n10790;
  assign n10763 = ~n11685 | ~n10837;
  assign n10774 = ~n10764 | ~n10763;
  assign n10768 = ~n10766;
  assign n10769 = ~n10768 | ~n10767;
  assign n11091 = n10765 ^ n10769;
  assign n10772 = ~n11503 | ~n10770;
  assign n10771 = ~n10869 | ~n11493;
  assign n10773 = ~n10772 | ~n10771;
  assign n10775 = ~n10774 & ~n10773;
  assign U2821 = ~n10776 | ~n10775;
  assign n10781 = ~n10777;
  assign n10779 = ~n10830 & ~n10778;
  assign n10780 = ~REIP_REG_5__SCAN_IN & ~n10779;
  assign n10799 = ~n10781 & ~n10780;
  assign n10783 = ~n10907 & ~n10782;
  assign n10786 = ~n10784 & ~n10783;
  assign n10785 = ~EBX_REG_5__SCAN_IN | ~n10904;
  assign n10792 = ~n10786 | ~n10785;
  assign n10789 = ~n10788 | ~n10787;
  assign n11707 = ~n10790 | ~n10789;
  assign n10791 = ~n10914 & ~n11707;
  assign n10797 = ~n10792 & ~n10791;
  assign n11098 = n10767 ^ n10766;
  assign n11514 = ~n11098;
  assign n10794 = ~n10809 | ~n10793;
  assign n10924 = ~n10795 | ~n10794;
  assign n10796 = ~n11514 | ~n10924;
  assign n10798 = ~n10797 | ~n10796;
  assign n10801 = ~n10799 & ~n10798;
  assign n10800 = ~n11509 | ~n10869;
  assign U2822 = ~n10801 | ~n10800;
  assign n11722 = n10803 ^ n10802;
  assign n10805 = ~n11722 | ~n10837;
  assign n10804 = ~n10904 | ~EBX_REG_4__SCAN_IN;
  assign n10808 = ~n10805 | ~n10804;
  assign n10806 = ~n10812 | ~n10851;
  assign n10807 = ~REIP_REG_4__SCAN_IN & ~n10806;
  assign n10818 = ~n10808 & ~n10807;
  assign n10881 = ~n10809 | ~n13743;
  assign n10903 = ~n10881;
  assign n10811 = ~n10903 | ~n11868;
  assign n10810 = ~n10896 | ~PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n10816 = ~n10811 | ~n10810;
  assign n10833 = n10830 | n10812;
  assign n10838 = ~n10893 | ~n10833;
  assign n10813 = ~REIP_REG_4__SCAN_IN | ~n10838;
  assign n10815 = ~n10814 | ~n10813;
  assign n10817 = ~n10816 & ~n10815;
  assign n10820 = ~n10818 | ~n10817;
  assign n10819 = ~n11522 & ~n10908;
  assign n10827 = ~n10820 & ~n10819;
  assign n10824 = ~n10821 | ~n10848;
  assign n10823 = ~n10822;
  assign n10825 = ~n10824 | ~n10823;
  assign n10996 = n10766 & n10825;
  assign n10826 = ~n10996 | ~n10924;
  assign U2823 = ~n10827 | ~n10826;
  assign n10829 = ~n10904 | ~EBX_REG_3__SCAN_IN;
  assign n10828 = ~n10896 | ~PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n10835 = ~n10829 | ~n10828;
  assign n10895 = ~REIP_REG_1__SCAN_IN & ~n10830;
  assign n10832 = ~n10831 & ~n10895;
  assign n10854 = ~REIP_REG_2__SCAN_IN | ~n10832;
  assign n10834 = ~n10833 & ~n10854;
  assign n10845 = ~n10835 & ~n10834;
  assign n11738 = n10862 ^ n10836;
  assign n10840 = ~n10837 | ~n11738;
  assign n10839 = ~REIP_REG_3__SCAN_IN | ~n10838;
  assign n10843 = ~n10840 | ~n10839;
  assign n10842 = ~n10881 & ~n12757;
  assign n10844 = ~n10843 & ~n10842;
  assign n10847 = ~n10845 | ~n10844;
  assign n10846 = ~n11528 & ~n7011;
  assign n10850 = ~n10847 & ~n10846;
  assign n11107 = n10848 ^ ~n10821;
  assign n11533 = ~n11107;
  assign n10849 = ~n11533 | ~n10924;
  assign U2824 = ~n10850 | ~n10849;
  assign n13454 = ~REIP_REG_2__SCAN_IN;
  assign n10852 = ~n10851 | ~REIP_REG_1__SCAN_IN;
  assign n10853 = ~n13454 | ~n10852;
  assign n10861 = ~n10854 | ~n10853;
  assign n10856 = n10855;
  assign n12248 = ~n10856;
  assign n10859 = ~n10881 & ~n12248;
  assign n10857 = ~PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n10858 = ~n10907 & ~n10857;
  assign n10860 = ~n10859 & ~n10858;
  assign n10878 = n10861 & n10860;
  assign n10866 = ~n10862;
  assign n10865 = ~n10864 | ~n10863;
  assign n11758 = ~n10866 | ~n10865;
  assign n10868 = n11758 | n10914;
  assign n10867 = ~n10904 | ~EBX_REG_2__SCAN_IN;
  assign n10876 = ~n10868 | ~n10867;
  assign n10874 = ~n11547 | ~n10869;
  assign n10870 = ~n10889;
  assign n10872 = ~n10871 & ~n10870;
  assign n11551 = ~n10821 & ~n10872;
  assign n10873 = ~n11551 | ~n10924;
  assign n10875 = ~n10874 | ~n10873;
  assign n10877 = ~n10876 & ~n10875;
  assign U2825 = ~n10878 | ~n10877;
  assign n10880 = n10879;
  assign n10883 = ~n10881 & ~n10880;
  assign n10882 = ~n11775 & ~n10914;
  assign n10885 = ~n10883 & ~n10882;
  assign n10884 = ~EBX_REG_1__SCAN_IN | ~n10904;
  assign n10892 = ~n10885 | ~n10884;
  assign n10890 = ~n10924;
  assign n10888 = n10887 | n10886;
  assign n11571 = ~n10889 | ~n10888;
  assign n10891 = ~n10890 & ~n11571;
  assign n10902 = ~n10892 & ~n10891;
  assign n10894 = ~n13722 & ~n10893;
  assign n10898 = ~n10895 & ~n10894;
  assign n10897 = ~n10896 | ~PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n10900 = ~n10898 | ~n10897;
  assign n10899 = ~PHYADDRPOINTER_REG_1__SCAN_IN & ~n7011;
  assign n10901 = ~n10900 & ~n10899;
  assign U2826 = ~n10902 | ~n10901;
  assign n10906 = ~n10903 | ~n13703;
  assign n10905 = ~n10904 | ~EBX_REG_0__SCAN_IN;
  assign n10920 = ~n10906 | ~n10905;
  assign n10909 = ~n10908 | ~n10907;
  assign n10918 = ~n10909 | ~PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n10916 = ~n10910 & ~n13723;
  assign n10913 = ~n10912 | ~n11771;
  assign n11791 = ~n9225 | ~n10913;
  assign n10915 = ~n10914 & ~n11791;
  assign n10917 = ~n10916 & ~n10915;
  assign n10919 = ~n10918 | ~n10917;
  assign n10926 = ~n10920 & ~n10919;
  assign n10922 = ~n10921;
  assign n11586 = n10923 ^ ~n10922;
  assign n10925 = ~n10924 | ~n11586;
  assign U2827 = ~n10926 | ~n10925;
  assign n10928 = ~n10927;
  assign n10930 = ~n10928 | ~n11001;
  assign n10929 = ~EBX_REG_31__SCAN_IN | ~n11013;
  assign U2828 = ~n10930 | ~n10929;
  assign n10933 = ~n10931 & ~n11016;
  assign n10932 = ~n11025 & ~n11010;
  assign n10935 = ~n10933 & ~n10932;
  assign n10934 = ~EBX_REG_18__SCAN_IN | ~n11013;
  assign U2841 = ~n10935 | ~n10934;
  assign n10938 = ~n11013 | ~EBX_REG_17__SCAN_IN;
  assign n10937 = ~n10936 | ~n11001;
  assign n10941 = n10938 & n10937;
  assign n10940 = ~n10939 | ~n11020;
  assign U2842 = ~n10941 | ~n10940;
  assign n10944 = ~n10942 & ~n11016;
  assign n10943 = ~n11040 & ~n11010;
  assign n10946 = ~n10944 & ~n10943;
  assign n10945 = ~EBX_REG_16__SCAN_IN | ~n11013;
  assign U2843 = ~n10946 | ~n10945;
  assign n10949 = ~n10947 & ~n11016;
  assign n10948 = ~n11046 & ~n11010;
  assign n10951 = ~n10949 & ~n10948;
  assign n10950 = ~EBX_REG_15__SCAN_IN | ~n11013;
  assign U2844 = ~n10951 | ~n10950;
  assign n10954 = ~n11013 | ~EBX_REG_14__SCAN_IN;
  assign n10953 = ~n10952 | ~n11001;
  assign n10957 = n10954 & n10953;
  assign n10956 = ~n10955 | ~n11020;
  assign U2845 = ~n10957 | ~n10956;
  assign n10960 = ~n11013 | ~EBX_REG_13__SCAN_IN;
  assign n10959 = ~n10958 | ~n11001;
  assign n10963 = n10960 & n10959;
  assign n10962 = ~n10961 | ~n11020;
  assign U2846 = ~n10963 | ~n10962;
  assign n10965 = ~n11589 & ~n11016;
  assign n10964 = ~n11062 & ~n11010;
  assign n10967 = ~n10965 & ~n10964;
  assign n10966 = ~EBX_REG_12__SCAN_IN | ~n11013;
  assign U2847 = ~n10967 | ~n10966;
  assign n10969 = ~n11609 & ~n11016;
  assign n10968 = ~n11067 & ~n11010;
  assign n10971 = ~n10969 & ~n10968;
  assign n10970 = ~EBX_REG_11__SCAN_IN | ~n11013;
  assign U2848 = ~n10971 | ~n10970;
  assign n10973 = ~n11622 & ~n11016;
  assign n10972 = ~n11072 & ~n11010;
  assign n10975 = ~n10973 & ~n10972;
  assign n10974 = ~EBX_REG_10__SCAN_IN | ~n11013;
  assign U2849 = ~n10975 | ~n10974;
  assign n10977 = ~n11640 & ~n11016;
  assign n10976 = ~n11077 & ~n11010;
  assign n10979 = ~n10977 & ~n10976;
  assign n10978 = ~EBX_REG_9__SCAN_IN | ~n11013;
  assign U2850 = ~n10979 | ~n10978;
  assign n10981 = ~n11082 & ~n11010;
  assign n10980 = n11013 & EBX_REG_8__SCAN_IN;
  assign n10983 = ~n10981 & ~n10980;
  assign n10982 = ~n11653 | ~n11001;
  assign U2851 = ~n10983 | ~n10982;
  assign n10985 = ~n11488 & ~n11010;
  assign n10984 = n11013 & EBX_REG_7__SCAN_IN;
  assign n10987 = ~n10985 & ~n10984;
  assign n10986 = ~n11672 | ~n11001;
  assign U2852 = ~n10987 | ~n10986;
  assign n10989 = ~n11013 | ~EBX_REG_6__SCAN_IN;
  assign n10988 = ~n11685 | ~n11001;
  assign n10991 = n10989 & n10988;
  assign n10990 = ~n11503 | ~n11020;
  assign U2853 = ~n10991 | ~n10990;
  assign n10993 = ~n11707 & ~n11016;
  assign n10992 = ~n11098 & ~n11010;
  assign n10995 = ~n10993 & ~n10992;
  assign n10994 = ~EBX_REG_5__SCAN_IN | ~n11013;
  assign U2854 = ~n10995 | ~n10994;
  assign n10998 = ~n11523 & ~n11010;
  assign n10997 = n11013 & EBX_REG_4__SCAN_IN;
  assign n11000 = ~n10998 & ~n10997;
  assign n10999 = ~n11722 | ~n11001;
  assign U2855 = ~n11000 | ~n10999;
  assign n11003 = ~n11013 | ~EBX_REG_3__SCAN_IN;
  assign n11002 = ~n11738 | ~n11001;
  assign n11005 = n11003 & n11002;
  assign n11004 = ~n11533 | ~n11020;
  assign U2856 = ~n11005 | ~n11004;
  assign n11007 = ~n11758 & ~n11016;
  assign n11112 = ~n11551;
  assign n11006 = ~n11112 & ~n11010;
  assign n11009 = ~n11007 & ~n11006;
  assign n11008 = ~EBX_REG_2__SCAN_IN | ~n11013;
  assign U2857 = ~n11009 | ~n11008;
  assign n11012 = ~n11775 & ~n11016;
  assign n11011 = ~n11571 & ~n11010;
  assign n11015 = ~n11012 & ~n11011;
  assign n11014 = ~EBX_REG_1__SCAN_IN | ~n11013;
  assign U2858 = ~n11015 | ~n11014;
  assign n11019 = ~n11016 & ~n11791;
  assign n11018 = ~n11017 & ~n9222;
  assign n11022 = ~n11019 & ~n11018;
  assign n11021 = ~n11586 | ~n11020;
  assign U2859 = ~n11022 | ~n11021;
  assign n11024 = ~n11043 | ~DATAI_2_;
  assign n11023 = ~n11037 | ~DATAI_18_;
  assign n11027 = ~n11024 | ~n11023;
  assign n11026 = ~n11025 & ~n11123;
  assign n11029 = ~n11027 & ~n11026;
  assign n11028 = ~EAX_REG_18__SCAN_IN | ~n6994;
  assign U2873 = ~n11029 | ~n11028;
  assign n11031 = ~n11043 | ~DATAI_1_;
  assign n11030 = ~n11037 | ~DATAI_17_;
  assign n11034 = ~n11031 | ~n11030;
  assign n11033 = ~n11032 & ~n11123;
  assign n11036 = ~n11034 & ~n11033;
  assign n11035 = ~EAX_REG_17__SCAN_IN | ~n6994;
  assign U2874 = ~n11036 | ~n11035;
  assign n11039 = ~n11037 | ~DATAI_16_;
  assign n11038 = ~n6994 | ~EAX_REG_16__SCAN_IN;
  assign n11042 = ~n11039 | ~n11038;
  assign n11041 = ~n11040 & ~n11123;
  assign n11045 = ~n11042 & ~n11041;
  assign n11044 = ~n11043 | ~DATAI_0_;
  assign U2875 = ~n11045 | ~n11044;
  assign n11048 = ~n11046 & ~n11123;
  assign n11406 = ~EAX_REG_15__SCAN_IN;
  assign n11047 = ~n11092 & ~n11406;
  assign n11051 = ~n11048 & ~n11047;
  assign n11050 = ~DATAI_15_ | ~n11097;
  assign U2876 = ~n11051 | ~n11050;
  assign n11054 = ~n11052 & ~n11123;
  assign n11398 = ~EAX_REG_14__SCAN_IN;
  assign n11053 = ~n11092 & ~n11398;
  assign n11056 = ~n11054 & ~n11053;
  assign n11055 = ~DATAI_14_ | ~n11097;
  assign U2877 = ~n11056 | ~n11055;
  assign n11059 = ~n11057 & ~n11123;
  assign n11393 = ~EAX_REG_13__SCAN_IN;
  assign n11058 = ~n11092 & ~n11393;
  assign n11061 = ~n11059 & ~n11058;
  assign n11060 = ~DATAI_13_ | ~n11097;
  assign U2878 = ~n11061 | ~n11060;
  assign n11064 = ~n11062 & ~n11123;
  assign n11388 = ~EAX_REG_12__SCAN_IN;
  assign n11063 = ~n11092 & ~n11388;
  assign n11066 = ~n11064 & ~n11063;
  assign n11065 = ~DATAI_12_ | ~n11097;
  assign U2879 = ~n11066 | ~n11065;
  assign n11069 = ~n11067 & ~n11123;
  assign n11383 = ~EAX_REG_11__SCAN_IN;
  assign n11068 = ~n11092 & ~n11383;
  assign n11071 = ~n11069 & ~n11068;
  assign n11070 = ~DATAI_11_ | ~n11097;
  assign U2880 = ~n11071 | ~n11070;
  assign n11074 = ~n11072 & ~n11123;
  assign n11378 = ~EAX_REG_10__SCAN_IN;
  assign n11073 = ~n11092 & ~n11378;
  assign n11076 = ~n11074 & ~n11073;
  assign n11075 = ~DATAI_10_ | ~n11097;
  assign U2881 = ~n11076 | ~n11075;
  assign n11079 = ~n11077 & ~n11123;
  assign n11373 = ~EAX_REG_9__SCAN_IN;
  assign n11078 = ~n11092 & ~n11373;
  assign n11081 = ~n11079 & ~n11078;
  assign n11080 = ~DATAI_9_ | ~n11097;
  assign U2882 = ~n11081 | ~n11080;
  assign n11084 = ~n11082 & ~n11123;
  assign n11368 = ~EAX_REG_8__SCAN_IN;
  assign n11083 = ~n11092 & ~n11368;
  assign n11086 = ~n11084 & ~n11083;
  assign n11085 = ~DATAI_8_ | ~n11097;
  assign U2883 = ~n11086 | ~n11085;
  assign n11088 = ~n11488 & ~n11123;
  assign n11363 = ~EAX_REG_7__SCAN_IN;
  assign n11087 = ~n11092 & ~n11363;
  assign n11090 = ~n11088 & ~n11087;
  assign n11089 = ~DATAI_7_ | ~n11097;
  assign U2884 = ~n11090 | ~n11089;
  assign n11094 = ~n11091 & ~n11123;
  assign n11358 = ~EAX_REG_6__SCAN_IN;
  assign n11093 = ~n11092 & ~n11358;
  assign n11096 = ~n11094 & ~n11093;
  assign n11095 = ~DATAI_6_ | ~n11097;
  assign U2885 = ~n11096 | ~n11095;
  assign n11951 = ~DATAI_5_;
  assign n11100 = ~n11951 & ~n11121;
  assign n11099 = ~n11098 & ~n11123;
  assign n11102 = ~n11100 & ~n11099;
  assign n11101 = ~EAX_REG_5__SCAN_IN | ~n6994;
  assign U2886 = ~n11102 | ~n11101;
  assign n11941 = ~DATAI_4_;
  assign n11104 = ~n11941 & ~n11121;
  assign n11103 = ~n11523 & ~n11123;
  assign n11106 = ~n11104 & ~n11103;
  assign n11105 = ~EAX_REG_4__SCAN_IN | ~n6994;
  assign U2887 = ~n11106 | ~n11105;
  assign n11931 = ~DATAI_3_;
  assign n11109 = ~n11931 & ~n11121;
  assign n11108 = ~n11107 & ~n11123;
  assign n11111 = ~n11109 & ~n11108;
  assign n11110 = ~EAX_REG_3__SCAN_IN | ~n6994;
  assign U2888 = ~n11111 | ~n11110;
  assign n11921 = ~DATAI_2_;
  assign n11114 = ~n11921 & ~n11121;
  assign n11113 = ~n11112 & ~n11123;
  assign n11116 = ~n11114 & ~n11113;
  assign n11115 = ~EAX_REG_2__SCAN_IN | ~n6994;
  assign U2889 = ~n11116 | ~n11115;
  assign n11911 = ~DATAI_1_;
  assign n11118 = ~n11911 & ~n11121;
  assign n11117 = ~n11123 & ~n11571;
  assign n11120 = ~n11118 & ~n11117;
  assign n11119 = ~EAX_REG_1__SCAN_IN | ~n6994;
  assign U2890 = ~n11120 | ~n11119;
  assign n11902 = ~DATAI_0_;
  assign n11125 = ~n11902 & ~n11121;
  assign n11122 = ~n11586;
  assign n11124 = ~n11123 & ~n11122;
  assign n11127 = ~n11125 & ~n11124;
  assign n11126 = ~EAX_REG_0__SCAN_IN | ~n6994;
  assign U2891 = ~n11127 | ~n11126;
  assign n11129 = ~DATAO_REG_30__SCAN_IN | ~n11245;
  assign n11128 = ~n11252 | ~UWORD_REG_14__SCAN_IN;
  assign n11133 = n11129 & n11128;
  assign n11130 = ~n11253;
  assign n11132 = ~n11131 | ~EAX_REG_30__SCAN_IN;
  assign U2893 = ~n11133 | ~n11132;
  assign n11135 = ~n11245 | ~DATAO_REG_29__SCAN_IN;
  assign n11134 = ~n11252 | ~UWORD_REG_13__SCAN_IN;
  assign n11137 = n11135 & n11134;
  assign n11136 = ~n11131 | ~EAX_REG_29__SCAN_IN;
  assign U2894 = ~n11137 | ~n11136;
  assign n11139 = ~n11245 | ~DATAO_REG_28__SCAN_IN;
  assign n11138 = ~n11252 | ~UWORD_REG_12__SCAN_IN;
  assign n11141 = n11139 & n11138;
  assign n11140 = ~n11131 | ~EAX_REG_28__SCAN_IN;
  assign U2895 = ~n11141 | ~n11140;
  assign n11143 = ~n11256 | ~DATAO_REG_27__SCAN_IN;
  assign n11142 = ~n11252 | ~UWORD_REG_11__SCAN_IN;
  assign n11145 = n11143 & n11142;
  assign n11144 = ~n11131 | ~EAX_REG_27__SCAN_IN;
  assign U2896 = ~n11145 | ~n11144;
  assign n11147 = ~n11256 | ~DATAO_REG_26__SCAN_IN;
  assign n11146 = ~n11186 | ~UWORD_REG_10__SCAN_IN;
  assign n11149 = n11147 & n11146;
  assign n11148 = ~n11131 | ~EAX_REG_26__SCAN_IN;
  assign U2897 = ~n11149 | ~n11148;
  assign n11151 = ~n11245 | ~DATAO_REG_25__SCAN_IN;
  assign n11150 = ~n11186 | ~UWORD_REG_9__SCAN_IN;
  assign n11153 = n11151 & n11150;
  assign n11152 = ~n11131 | ~EAX_REG_25__SCAN_IN;
  assign U2898 = ~n11153 | ~n11152;
  assign n11155 = ~n11245 | ~DATAO_REG_24__SCAN_IN;
  assign n11154 = ~n11186 | ~UWORD_REG_8__SCAN_IN;
  assign n11157 = n11155 & n11154;
  assign n11156 = ~n11131 | ~EAX_REG_24__SCAN_IN;
  assign U2899 = ~n11157 | ~n11156;
  assign n11159 = ~n11245 | ~DATAO_REG_23__SCAN_IN;
  assign n11158 = ~n11186 | ~UWORD_REG_7__SCAN_IN;
  assign n11161 = n11159 & n11158;
  assign n11160 = ~n11131 | ~EAX_REG_23__SCAN_IN;
  assign U2900 = ~n11161 | ~n11160;
  assign n11163 = ~DATAO_REG_22__SCAN_IN | ~n11245;
  assign n11162 = ~n11186 | ~UWORD_REG_6__SCAN_IN;
  assign n11165 = n11163 & n11162;
  assign n11164 = ~n11131 | ~EAX_REG_22__SCAN_IN;
  assign U2901 = ~n11165 | ~n11164;
  assign n11167 = ~DATAO_REG_21__SCAN_IN | ~n11245;
  assign n11166 = ~n11186 | ~UWORD_REG_5__SCAN_IN;
  assign n11169 = n11167 & n11166;
  assign n11168 = ~n11131 | ~EAX_REG_21__SCAN_IN;
  assign U2902 = ~n11169 | ~n11168;
  assign n11171 = ~n11256 | ~DATAO_REG_20__SCAN_IN;
  assign n11170 = ~n11252 | ~UWORD_REG_4__SCAN_IN;
  assign n11173 = n11171 & n11170;
  assign n11172 = ~n11131 | ~EAX_REG_20__SCAN_IN;
  assign U2903 = ~n11173 | ~n11172;
  assign n11175 = ~n11245 | ~DATAO_REG_19__SCAN_IN;
  assign n11174 = ~n11186 | ~UWORD_REG_3__SCAN_IN;
  assign n11177 = n11175 & n11174;
  assign n11176 = ~n11131 | ~EAX_REG_19__SCAN_IN;
  assign U2904 = ~n11177 | ~n11176;
  assign n11179 = ~n11256 | ~DATAO_REG_18__SCAN_IN;
  assign n11178 = ~n11186 | ~UWORD_REG_2__SCAN_IN;
  assign n11181 = n11179 & n11178;
  assign n11180 = ~n11131 | ~EAX_REG_18__SCAN_IN;
  assign U2905 = ~n11181 | ~n11180;
  assign n11183 = ~n11245 | ~DATAO_REG_17__SCAN_IN;
  assign n11182 = ~n11186 | ~UWORD_REG_1__SCAN_IN;
  assign n11185 = n11183 & n11182;
  assign n11184 = ~n11131 | ~EAX_REG_17__SCAN_IN;
  assign U2906 = ~n11185 | ~n11184;
  assign n11188 = ~n11256 | ~DATAO_REG_16__SCAN_IN;
  assign n11187 = ~n11186 | ~UWORD_REG_0__SCAN_IN;
  assign n11190 = n11188 & n11187;
  assign n11189 = ~n11131 | ~EAX_REG_16__SCAN_IN;
  assign U2907 = ~n11190 | ~n11189;
  assign n11192 = ~n11252 | ~LWORD_REG_15__SCAN_IN;
  assign n11191 = ~n11253 | ~EAX_REG_15__SCAN_IN;
  assign n11194 = n11192 & n11191;
  assign n11193 = ~n11245 | ~DATAO_REG_15__SCAN_IN;
  assign U2908 = ~n11194 | ~n11193;
  assign n11196 = ~n11252 | ~LWORD_REG_14__SCAN_IN;
  assign n11195 = ~n11253 | ~EAX_REG_14__SCAN_IN;
  assign n11198 = n11196 & n11195;
  assign n11197 = ~n11256 | ~DATAO_REG_14__SCAN_IN;
  assign U2909 = ~n11198 | ~n11197;
  assign n11200 = ~n11252 | ~LWORD_REG_13__SCAN_IN;
  assign n11199 = ~n11253 | ~EAX_REG_13__SCAN_IN;
  assign n11202 = n11200 & n11199;
  assign n11201 = ~n11245 | ~DATAO_REG_13__SCAN_IN;
  assign U2910 = ~n11202 | ~n11201;
  assign n11204 = ~n11252 | ~LWORD_REG_12__SCAN_IN;
  assign n11203 = ~n11253 | ~EAX_REG_12__SCAN_IN;
  assign n11206 = n11204 & n11203;
  assign n11205 = ~n11245 | ~DATAO_REG_12__SCAN_IN;
  assign U2911 = ~n11206 | ~n11205;
  assign n11208 = ~n11252 | ~LWORD_REG_11__SCAN_IN;
  assign n11207 = ~n11253 | ~EAX_REG_11__SCAN_IN;
  assign n11210 = n11208 & n11207;
  assign n11209 = ~n11245 | ~DATAO_REG_11__SCAN_IN;
  assign U2912 = ~n11210 | ~n11209;
  assign n11212 = ~n11252 | ~LWORD_REG_10__SCAN_IN;
  assign n11211 = ~n11253 | ~EAX_REG_10__SCAN_IN;
  assign n11214 = n11212 & n11211;
  assign n11213 = ~n11256 | ~DATAO_REG_10__SCAN_IN;
  assign U2913 = ~n11214 | ~n11213;
  assign n11216 = ~n11252 | ~LWORD_REG_9__SCAN_IN;
  assign n11215 = ~n11253 | ~EAX_REG_9__SCAN_IN;
  assign n11218 = n11216 & n11215;
  assign n11217 = ~n11256 | ~DATAO_REG_9__SCAN_IN;
  assign U2914 = ~n11218 | ~n11217;
  assign n11220 = ~n11252 | ~LWORD_REG_8__SCAN_IN;
  assign n11219 = ~n11253 | ~EAX_REG_8__SCAN_IN;
  assign n11222 = n11220 & n11219;
  assign n11221 = ~n11245 | ~DATAO_REG_8__SCAN_IN;
  assign U2915 = ~n11222 | ~n11221;
  assign n11224 = ~n11252 | ~LWORD_REG_7__SCAN_IN;
  assign n11223 = ~n11253 | ~EAX_REG_7__SCAN_IN;
  assign n11226 = n11224 & n11223;
  assign n11225 = ~n11245 | ~DATAO_REG_7__SCAN_IN;
  assign U2916 = ~n11226 | ~n11225;
  assign n11228 = ~n11252 | ~LWORD_REG_6__SCAN_IN;
  assign n11227 = ~n11253 | ~EAX_REG_6__SCAN_IN;
  assign n11230 = n11228 & n11227;
  assign n11229 = ~n11245 | ~DATAO_REG_6__SCAN_IN;
  assign U2917 = ~n11230 | ~n11229;
  assign n11232 = ~n11252 | ~LWORD_REG_5__SCAN_IN;
  assign n11231 = ~n11253 | ~EAX_REG_5__SCAN_IN;
  assign n11234 = n11232 & n11231;
  assign n11233 = ~n11256 | ~DATAO_REG_5__SCAN_IN;
  assign U2918 = ~n11234 | ~n11233;
  assign n11236 = ~n11252 | ~LWORD_REG_4__SCAN_IN;
  assign n11235 = ~n11253 | ~EAX_REG_4__SCAN_IN;
  assign n11238 = n11236 & n11235;
  assign n11237 = ~n11245 | ~DATAO_REG_4__SCAN_IN;
  assign U2919 = ~n11238 | ~n11237;
  assign n11240 = ~n11252 | ~LWORD_REG_3__SCAN_IN;
  assign n11239 = ~n11253 | ~EAX_REG_3__SCAN_IN;
  assign n11242 = n11240 & n11239;
  assign n11241 = ~n11245 | ~DATAO_REG_3__SCAN_IN;
  assign U2920 = ~n11242 | ~n11241;
  assign n11244 = ~n11252 | ~LWORD_REG_2__SCAN_IN;
  assign n11243 = ~n11253 | ~EAX_REG_2__SCAN_IN;
  assign n11247 = n11244 & n11243;
  assign n11246 = ~n11245 | ~DATAO_REG_2__SCAN_IN;
  assign U2921 = ~n11247 | ~n11246;
  assign n11249 = ~n11252 | ~LWORD_REG_1__SCAN_IN;
  assign n11248 = ~n11253 | ~EAX_REG_1__SCAN_IN;
  assign n11251 = n11249 & n11248;
  assign n11250 = ~n11256 | ~DATAO_REG_1__SCAN_IN;
  assign U2922 = ~n11251 | ~n11250;
  assign n11255 = ~n11252 | ~LWORD_REG_0__SCAN_IN;
  assign n11254 = ~n11253 | ~EAX_REG_0__SCAN_IN;
  assign n11258 = n11255 & n11254;
  assign n11257 = ~n11256 | ~DATAO_REG_0__SCAN_IN;
  assign U2923 = ~n11258 | ~n11257;
  assign n11330 = ~n11405 & ~n11902;
  assign n11407 = ~n11259;
  assign n11260 = ~EAX_REG_16__SCAN_IN;
  assign n11261 = ~n11407 & ~n11260;
  assign n11265 = ~n11330 & ~n11261;
  assign n11262 = ~n13741 & ~n13431;
  assign n11264 = ~UWORD_REG_0__SCAN_IN | ~n11401;
  assign U2924 = ~n11265 | ~n11264;
  assign n11335 = ~n11405 & ~n11911;
  assign n11266 = ~EAX_REG_17__SCAN_IN;
  assign n11267 = ~n11407 & ~n11266;
  assign n11269 = ~n11335 & ~n11267;
  assign n11268 = ~UWORD_REG_1__SCAN_IN | ~n11401;
  assign U2925 = ~n11269 | ~n11268;
  assign n11340 = ~n11405 & ~n11921;
  assign n11270 = ~EAX_REG_18__SCAN_IN;
  assign n11271 = ~n11407 & ~n11270;
  assign n11273 = ~n11340 & ~n11271;
  assign n11272 = ~UWORD_REG_2__SCAN_IN | ~n11401;
  assign U2926 = ~n11273 | ~n11272;
  assign n11345 = ~n11405 & ~n11931;
  assign n11274 = ~EAX_REG_19__SCAN_IN;
  assign n11275 = ~n11407 & ~n11274;
  assign n11277 = ~n11345 & ~n11275;
  assign n11276 = ~UWORD_REG_3__SCAN_IN | ~n11401;
  assign U2927 = ~n11277 | ~n11276;
  assign n11350 = ~n11405 & ~n11941;
  assign n11278 = ~EAX_REG_20__SCAN_IN;
  assign n11279 = ~n11407 & ~n11278;
  assign n11281 = ~n11350 & ~n11279;
  assign n11280 = ~UWORD_REG_4__SCAN_IN | ~n11401;
  assign U2928 = ~n11281 | ~n11280;
  assign n11355 = ~n11405 & ~n11951;
  assign n11282 = ~EAX_REG_21__SCAN_IN;
  assign n11283 = ~n11407 & ~n11282;
  assign n11285 = ~n11355 & ~n11283;
  assign n11284 = ~UWORD_REG_5__SCAN_IN | ~n11401;
  assign U2929 = ~n11285 | ~n11284;
  assign n11960 = ~DATAI_6_;
  assign n11360 = ~n11405 & ~n11960;
  assign n11286 = ~EAX_REG_22__SCAN_IN;
  assign n11287 = ~n11407 & ~n11286;
  assign n11289 = ~n11360 & ~n11287;
  assign n11288 = ~UWORD_REG_6__SCAN_IN | ~n11401;
  assign U2930 = ~n11289 | ~n11288;
  assign n11972 = ~DATAI_7_;
  assign n11365 = ~n11405 & ~n11972;
  assign n11290 = ~EAX_REG_23__SCAN_IN;
  assign n11291 = ~n11407 & ~n11290;
  assign n11293 = ~n11365 & ~n11291;
  assign n11292 = ~UWORD_REG_7__SCAN_IN | ~n11401;
  assign U2931 = ~n11293 | ~n11292;
  assign n11294 = ~DATAI_8_;
  assign n11370 = ~n11405 & ~n11294;
  assign n11295 = ~EAX_REG_24__SCAN_IN;
  assign n11296 = ~n11407 & ~n11295;
  assign n11298 = ~n11370 & ~n11296;
  assign n11297 = ~UWORD_REG_8__SCAN_IN | ~n11401;
  assign U2932 = ~n11298 | ~n11297;
  assign n11299 = ~DATAI_9_;
  assign n11375 = ~n11405 & ~n11299;
  assign n11300 = ~EAX_REG_25__SCAN_IN;
  assign n11301 = ~n11407 & ~n11300;
  assign n11303 = ~n11375 & ~n11301;
  assign n11302 = ~UWORD_REG_9__SCAN_IN | ~n11401;
  assign U2933 = ~n11303 | ~n11302;
  assign n11304 = ~DATAI_10_;
  assign n11380 = ~n11405 & ~n11304;
  assign n11305 = ~EAX_REG_26__SCAN_IN;
  assign n11306 = ~n11407 & ~n11305;
  assign n11308 = ~n11380 & ~n11306;
  assign n11307 = ~UWORD_REG_10__SCAN_IN | ~n11401;
  assign U2934 = ~n11308 | ~n11307;
  assign n11309 = ~DATAI_11_;
  assign n11385 = ~n11405 & ~n11309;
  assign n11310 = ~EAX_REG_27__SCAN_IN;
  assign n11311 = ~n11407 & ~n11310;
  assign n11313 = ~n11385 & ~n11311;
  assign n11312 = ~UWORD_REG_11__SCAN_IN | ~n11401;
  assign U2935 = ~n11313 | ~n11312;
  assign n11314 = ~DATAI_12_;
  assign n11390 = ~n11405 & ~n11314;
  assign n11315 = ~EAX_REG_28__SCAN_IN;
  assign n11316 = ~n11407 & ~n11315;
  assign n11318 = ~n11390 & ~n11316;
  assign n11317 = ~UWORD_REG_12__SCAN_IN | ~n11401;
  assign U2936 = ~n11318 | ~n11317;
  assign n11319 = ~DATAI_13_;
  assign n11395 = ~n11405 & ~n11319;
  assign n11320 = ~EAX_REG_29__SCAN_IN;
  assign n11321 = ~n11407 & ~n11320;
  assign n11323 = ~n11395 & ~n11321;
  assign n11322 = ~UWORD_REG_13__SCAN_IN | ~n11401;
  assign U2937 = ~n11323 | ~n11322;
  assign n11324 = ~DATAI_14_;
  assign n11400 = ~n11405 & ~n11324;
  assign n11325 = ~n11407 & ~n9437;
  assign n11327 = ~n11400 & ~n11325;
  assign n11326 = ~UWORD_REG_14__SCAN_IN | ~n11401;
  assign U2938 = ~n11327 | ~n11326;
  assign n11328 = ~EAX_REG_0__SCAN_IN;
  assign n11329 = ~n11407 & ~n11328;
  assign n11332 = ~n11330 & ~n11329;
  assign n11331 = ~LWORD_REG_0__SCAN_IN | ~n11401;
  assign U2939 = ~n11332 | ~n11331;
  assign n11333 = ~EAX_REG_1__SCAN_IN;
  assign n11334 = ~n11407 & ~n11333;
  assign n11337 = ~n11335 & ~n11334;
  assign n11336 = ~LWORD_REG_1__SCAN_IN | ~n11401;
  assign U2940 = ~n11337 | ~n11336;
  assign n11338 = ~EAX_REG_2__SCAN_IN;
  assign n11339 = ~n11407 & ~n11338;
  assign n11342 = ~n11340 & ~n11339;
  assign n11341 = ~LWORD_REG_2__SCAN_IN | ~n11401;
  assign U2941 = ~n11342 | ~n11341;
  assign n11343 = ~EAX_REG_3__SCAN_IN;
  assign n11344 = ~n11407 & ~n11343;
  assign n11347 = ~n11345 & ~n11344;
  assign n11346 = ~LWORD_REG_3__SCAN_IN | ~n11401;
  assign U2942 = ~n11347 | ~n11346;
  assign n11348 = ~EAX_REG_4__SCAN_IN;
  assign n11349 = ~n11407 & ~n11348;
  assign n11352 = ~n11350 & ~n11349;
  assign n11351 = ~LWORD_REG_4__SCAN_IN | ~n11401;
  assign U2943 = ~n11352 | ~n11351;
  assign n11353 = ~EAX_REG_5__SCAN_IN;
  assign n11354 = ~n11407 & ~n11353;
  assign n11357 = ~n11355 & ~n11354;
  assign n11356 = ~LWORD_REG_5__SCAN_IN | ~n11401;
  assign U2944 = ~n11357 | ~n11356;
  assign n11359 = ~n11407 & ~n11358;
  assign n11362 = ~n11360 & ~n11359;
  assign n11361 = ~LWORD_REG_6__SCAN_IN | ~n11401;
  assign U2945 = ~n11362 | ~n11361;
  assign n11364 = ~n11407 & ~n11363;
  assign n11367 = ~n11365 & ~n11364;
  assign n11366 = ~LWORD_REG_7__SCAN_IN | ~n11401;
  assign U2946 = ~n11367 | ~n11366;
  assign n11369 = ~n11407 & ~n11368;
  assign n11372 = ~n11370 & ~n11369;
  assign n11371 = ~LWORD_REG_8__SCAN_IN | ~n11401;
  assign U2947 = ~n11372 | ~n11371;
  assign n11374 = ~n11407 & ~n11373;
  assign n11377 = ~n11375 & ~n11374;
  assign n11376 = ~LWORD_REG_9__SCAN_IN | ~n11401;
  assign U2948 = ~n11377 | ~n11376;
  assign n11379 = ~n11407 & ~n11378;
  assign n11382 = ~n11380 & ~n11379;
  assign n11381 = ~LWORD_REG_10__SCAN_IN | ~n11401;
  assign U2949 = ~n11382 | ~n11381;
  assign n11384 = ~n11407 & ~n11383;
  assign n11387 = ~n11385 & ~n11384;
  assign n11386 = ~LWORD_REG_11__SCAN_IN | ~n11401;
  assign U2950 = ~n11387 | ~n11386;
  assign n11389 = ~n11407 & ~n11388;
  assign n11392 = ~n11390 & ~n11389;
  assign n11391 = ~LWORD_REG_12__SCAN_IN | ~n11401;
  assign U2951 = ~n11392 | ~n11391;
  assign n11394 = ~n11407 & ~n11393;
  assign n11397 = ~n11395 & ~n11394;
  assign n11396 = ~LWORD_REG_13__SCAN_IN | ~n11401;
  assign U2952 = ~n11397 | ~n11396;
  assign n11399 = ~n11407 & ~n11398;
  assign n11403 = ~n11400 & ~n11399;
  assign n11402 = ~LWORD_REG_14__SCAN_IN | ~n11401;
  assign U2953 = ~n11403 | ~n11402;
  assign n11404 = ~DATAI_15_;
  assign n11409 = ~n11405 & ~n11404;
  assign n11408 = ~n11407 & ~n11406;
  assign n11411 = ~n11409 & ~n11408;
  assign n11410 = ~LWORD_REG_15__SCAN_IN | ~n11401;
  assign U2954 = ~n11411 | ~n11410;
  assign n11414 = ~n11412 & ~n11570;
  assign n11413 = n11581 & PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n11427 = ~n11414 & ~n11413;
  assign n11591 = ~n11559 & ~n13504;
  assign n11417 = ~n11591;
  assign n11416 = ~n11415 | ~n6996;
  assign n11425 = ~n11417 | ~n11416;
  assign n11453 = ~n11419;
  assign n11436 = ~n11418 | ~n11453;
  assign n11432 = ~n11436 & ~n7088;
  assign n11423 = ~n11432 & ~n11431;
  assign n11422 = ~n11421 & ~n11420;
  assign n11595 = n11423 ^ ~n11422;
  assign n11424 = ~n11595 & ~n11567;
  assign n11426 = ~n11425 & ~n11424;
  assign U2974 = ~n11427 | ~n11426;
  assign n11610 = ~n13499 & ~n11559;
  assign n11429 = ~n11610;
  assign n11428 = ~n11581 | ~PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n11442 = ~n11429 | ~n11428;
  assign n11440 = ~n11430 | ~n11548;
  assign n11434 = ~n11431;
  assign n11438 = ~n11432 | ~n11434;
  assign n11435 = ~n11434 | ~n11433;
  assign n11437 = ~n11436 | ~n11435;
  assign n11613 = ~n11438 | ~n11437;
  assign n11439 = ~n11613 | ~n11578;
  assign n11441 = ~n11440 | ~n11439;
  assign n11445 = ~n11442 & ~n11441;
  assign n11444 = ~n11443 | ~n6996;
  assign U2975 = ~n11445 | ~n11444;
  assign n11448 = ~n11446 & ~n11570;
  assign n11447 = n11581 & PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n11459 = ~n11448 & ~n11447;
  assign n13494 = ~REIP_REG_10__SCAN_IN;
  assign n11624 = ~n11559 & ~n13494;
  assign n11451 = ~n11624;
  assign n11450 = ~n11449 | ~n6996;
  assign n11457 = ~n11451 | ~n11450;
  assign n11455 = ~n11453 | ~n11452;
  assign n11635 = n11455 ^ n11454;
  assign n11456 = ~n11635 & ~n11567;
  assign n11458 = ~n11457 & ~n11456;
  assign U2976 = ~n11459 | ~n11458;
  assign n11641 = ~n11576 | ~REIP_REG_9__SCAN_IN;
  assign n11460 = ~n11581 | ~PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n11467 = ~n11641 | ~n11460;
  assign n11643 = n11461 ^ n11462;
  assign n11465 = ~n11643 | ~n11578;
  assign n11464 = ~n11548 | ~n11463;
  assign n11466 = ~n11465 | ~n11464;
  assign n11470 = ~n11467 & ~n11466;
  assign n11469 = ~n11468 | ~n6996;
  assign U2977 = ~n11470 | ~n11469;
  assign n11473 = ~n11471 & ~n11570;
  assign n11472 = n11581 & PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n11481 = ~n11473 & ~n11472;
  assign n11654 = ~n11576 | ~REIP_REG_8__SCAN_IN;
  assign n11475 = ~n11474 | ~n6996;
  assign n11479 = ~n11654 | ~n11475;
  assign n11656 = n11477 ^ ~n11476;
  assign n11478 = ~n11656 & ~n11567;
  assign n11480 = ~n11479 & ~n11478;
  assign U2978 = ~n11481 | ~n11480;
  assign n11674 = ~n11576 | ~REIP_REG_7__SCAN_IN;
  assign n11482 = ~n11581 | ~PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n11486 = ~n11674 | ~n11482;
  assign n11675 = n11483 ^ ~n11484;
  assign n11485 = ~n11675 & ~n11567;
  assign n11492 = ~n11486 & ~n11485;
  assign n11490 = ~n11487 & ~n11570;
  assign n11489 = ~n11488 & ~n11881;
  assign n11491 = ~n11490 & ~n11489;
  assign U2979 = ~n11492 | ~n11491;
  assign n11495 = ~n11548 | ~n11493;
  assign n11494 = ~n11581 | ~PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n11502 = ~n11495 | ~n11494;
  assign n11686 = ~n11576 | ~REIP_REG_6__SCAN_IN;
  assign n11498 = ~n11496 | ~n11497;
  assign n11696 = n11499 ^ n11498;
  assign n11500 = ~n11696 | ~n11578;
  assign n11501 = ~n11686 | ~n11500;
  assign n11505 = ~n11502 & ~n11501;
  assign n11504 = ~n11503 | ~n6996;
  assign U2980 = ~n11505 | ~n11504;
  assign n11708 = ~n13469 & ~n11559;
  assign n11507 = ~n11708;
  assign n11506 = ~n11581 | ~PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n11513 = ~n11507 | ~n11506;
  assign n11511 = ~n11719 | ~n11578;
  assign n11510 = ~n11548 | ~n11509;
  assign n11512 = ~n11511 | ~n11510;
  assign n11516 = ~n11513 & ~n11512;
  assign n11515 = ~n11514 | ~n6996;
  assign U2981 = ~n11516 | ~n11515;
  assign n11723 = ~n11576 | ~REIP_REG_4__SCAN_IN;
  assign n11517 = ~n11581 | ~PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n11521 = ~n11723 | ~n11517;
  assign n11725 = n11518 ^ ~n11519;
  assign n11520 = ~n11725 & ~n11567;
  assign n11527 = ~n11521 & ~n11520;
  assign n11525 = ~n11522 & ~n11570;
  assign n11524 = ~n11523 & ~n11881;
  assign n11526 = ~n11525 & ~n11524;
  assign U2982 = ~n11527 | ~n11526;
  assign n11532 = ~n11528 & ~n11570;
  assign n11531 = ~n11530 & ~n11529;
  assign n11546 = ~n11532 & ~n11531;
  assign n11740 = ~n11576 | ~REIP_REG_3__SCAN_IN;
  assign n11534 = ~n11533 | ~n6996;
  assign n11544 = ~n11740 | ~n11534;
  assign n11556 = n11537 ^ ~n11535;
  assign n11539 = ~n11556 | ~n11536;
  assign n11538 = ~n11537 | ~INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n11542 = ~n11539 | ~n11538;
  assign n11541 = n11540 ^ ~n11747;
  assign n11742 = n11542 ^ ~n11541;
  assign n11543 = ~n11742 & ~n11567;
  assign n11545 = ~n11544 & ~n11543;
  assign U2983 = ~n11546 | ~n11545;
  assign n11550 = ~n11548 | ~n11547;
  assign n11549 = ~n11581 | ~PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n11554 = ~n11550 | ~n11549;
  assign n11756 = ~n11576 | ~REIP_REG_2__SCAN_IN;
  assign n11552 = ~n11551 | ~n6996;
  assign n11553 = ~n11756 | ~n11552;
  assign n11558 = ~n11554 & ~n11553;
  assign n11761 = n11556 ^ ~n11555;
  assign n11557 = ~n11761 | ~n11578;
  assign U2984 = ~n11558 | ~n11557;
  assign n11776 = ~n13722 & ~n11559;
  assign n11561 = ~n11776;
  assign n11560 = ~n11581 | ~PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n11569 = ~n11561 | ~n11560;
  assign n11566 = ~n11563 | ~n11562;
  assign n11565 = n11564 ^ ~INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n11783 = n11566 ^ ~n11565;
  assign n11568 = ~n11783 & ~n11567;
  assign n11575 = ~n11569 & ~n11568;
  assign n11573 = ~PHYADDRPOINTER_REG_1__SCAN_IN & ~n11570;
  assign n11572 = ~n11571 & ~n11881;
  assign n11574 = ~n11573 & ~n11572;
  assign U2985 = ~n11575 | ~n11574;
  assign n11789 = ~n11576 | ~REIP_REG_0__SCAN_IN;
  assign n11802 = n11577 ^ INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n11579 = ~n11578 | ~n11802;
  assign n11585 = ~n11789 | ~n11579;
  assign n11583 = ~PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n11582 = ~n11581 & ~n11580;
  assign n11584 = ~n11583 & ~n11582;
  assign n11588 = ~n11585 & ~n11584;
  assign n11587 = ~n11586 | ~n6996;
  assign U2986 = ~n11588 | ~n11587;
  assign n11590 = ~n11792 & ~n11589;
  assign n11594 = ~n11591 & ~n11590;
  assign n11592 = ~INSTADDRPOINTER_REG_12__SCAN_IN & ~n11612;
  assign n11593 = ~INSTADDRPOINTER_REG_11__SCAN_IN | ~n11592;
  assign n11597 = ~n11594 | ~n11593;
  assign n11596 = ~n11595 & ~n11784;
  assign n11608 = ~n11597 & ~n11596;
  assign n11605 = ~n11616 | ~n11598;
  assign n11600 = ~n11599 | ~INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n11601 = ~n11600 | ~n11772;
  assign n11604 = ~n11601 | ~n11773;
  assign n11603 = ~n11663 & ~n11602;
  assign n11617 = ~n11604 & ~n11603;
  assign n11606 = ~n11605 | ~n11617;
  assign n11607 = ~n11606 | ~INSTADDRPOINTER_REG_12__SCAN_IN;
  assign U3006 = ~n11608 | ~n11607;
  assign n11611 = ~n11792 & ~n11609;
  assign n11621 = ~n11611 & ~n11610;
  assign n11615 = n11612 | INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n11614 = ~n11613 | ~n11803;
  assign n11619 = ~n11615 | ~n11614;
  assign n11618 = ~n11617 & ~n11616;
  assign n11620 = ~n11619 & ~n11618;
  assign U3007 = ~n11621 | ~n11620;
  assign n11623 = ~n11792 & ~n11622;
  assign n11639 = ~n11624 & ~n11623;
  assign n11649 = ~INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n11626 = INSTADDRPOINTER_REG_10__SCAN_IN ^ ~n11649;
  assign n11694 = ~n11625 & ~n11752;
  assign n11702 = ~n11772 & ~n11694;
  assign n11650 = ~n11702 & ~n11630;
  assign n11634 = ~n11626 | ~n11650;
  assign n11628 = n11689 & n11627;
  assign n11632 = ~n11629 & ~n11628;
  assign n11631 = ~n11772 | ~n11630;
  assign n11644 = ~n11632 | ~n11631;
  assign n11633 = ~INSTADDRPOINTER_REG_10__SCAN_IN | ~n11644;
  assign n11637 = ~n11634 | ~n11633;
  assign n11636 = ~n11635 & ~n11784;
  assign n11638 = ~n11637 & ~n11636;
  assign U3008 = ~n11639 | ~n11638;
  assign n11642 = n11792 | n11640;
  assign n11648 = ~n11642 | ~n11641;
  assign n11646 = ~n11643 | ~n11803;
  assign n11645 = ~INSTADDRPOINTER_REG_9__SCAN_IN | ~n11644;
  assign n11647 = ~n11646 | ~n11645;
  assign n11652 = ~n11648 & ~n11647;
  assign n11651 = ~n11650 | ~n11649;
  assign U3009 = ~n11652 | ~n11651;
  assign n11655 = ~n11739 | ~n11653;
  assign n11658 = ~n11655 | ~n11654;
  assign n11657 = ~n11656 & ~n11784;
  assign n11671 = ~n11658 & ~n11657;
  assign n11660 = ~n11659;
  assign n11746 = ~n11731 & ~n11702;
  assign n11680 = ~n11660 | ~n11746;
  assign n11661 = INSTADDRPOINTER_REG_7__SCAN_IN ^ ~INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n11669 = ~n11680 & ~n11661;
  assign n11664 = n11663 | n11662;
  assign n11667 = ~n11773 | ~n11664;
  assign n11666 = ~n11665 & ~n11732;
  assign n11679 = ~n11667 & ~n11666;
  assign n11668 = ~n11679 & ~n9021;
  assign n11670 = ~n11669 & ~n11668;
  assign U3010 = ~n11671 | ~n11670;
  assign n11673 = ~n11739 | ~n11672;
  assign n11677 = ~n11674 | ~n11673;
  assign n11676 = ~n11675 & ~n11784;
  assign n11684 = ~n11677 & ~n11676;
  assign n11682 = ~n11679 & ~n11678;
  assign n11681 = ~INSTADDRPOINTER_REG_7__SCAN_IN & ~n11680;
  assign n11683 = ~n11682 & ~n11681;
  assign U3011 = ~n11684 | ~n11683;
  assign n11687 = ~n11739 | ~n11685;
  assign n11700 = ~n11687 | ~n11686;
  assign n11688 = ~n11689 | ~n11752;
  assign n11762 = ~n11773 | ~n11688;
  assign n11712 = ~n11731 & ~n11728;
  assign n11701 = ~INSTADDRPOINTER_REG_5__SCAN_IN | ~n11712;
  assign n11691 = ~n11772 | ~n11701;
  assign n11690 = ~n11689 | ~n11728;
  assign n11692 = ~n11691 | ~n11690;
  assign n11716 = ~n11762 & ~n11692;
  assign n11693 = ~INSTADDRPOINTER_REG_5__SCAN_IN & ~n11728;
  assign n11710 = ~n11694 | ~n11693;
  assign n11695 = ~n11716 | ~n11710;
  assign n11698 = ~n11695 | ~INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n11697 = ~n11696 | ~n11803;
  assign n11699 = ~n11698 | ~n11697;
  assign n11706 = ~n11700 & ~n11699;
  assign n11704 = ~n11701;
  assign n11703 = ~INSTADDRPOINTER_REG_6__SCAN_IN & ~n11702;
  assign n11705 = ~n11704 | ~n11703;
  assign U3012 = ~n11706 | ~n11705;
  assign n11709 = ~n11792 & ~n11707;
  assign n11711 = ~n11709 & ~n11708;
  assign n11718 = ~n11711 | ~n11710;
  assign n11714 = ~n11712 | ~n11772;
  assign n11715 = n11714 & n11713;
  assign n11717 = ~n11716 & ~n11715;
  assign n11721 = ~n11718 & ~n11717;
  assign n11720 = ~n11719 | ~n11803;
  assign U3013 = ~n11721 | ~n11720;
  assign n11724 = ~n11739 | ~n11722;
  assign n11727 = ~n11724 | ~n11723;
  assign n11726 = ~n11725 & ~n11784;
  assign n11737 = ~n11727 & ~n11726;
  assign n11730 = ~n11746 | ~n11728;
  assign n11729 = ~INSTADDRPOINTER_REG_4__SCAN_IN & ~INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n11735 = ~n11730 & ~n11729;
  assign n11753 = ~n11731;
  assign n11733 = ~n11732 & ~n11753;
  assign n11745 = ~n11733 & ~n11762;
  assign n11734 = ~n11745 & ~n7066;
  assign n11736 = ~n11735 & ~n11734;
  assign U3014 = ~n11737 | ~n11736;
  assign n11741 = ~n11739 | ~n11738;
  assign n11744 = ~n11741 | ~n11740;
  assign n11743 = ~n11742 & ~n11784;
  assign n11751 = ~n11744 & ~n11743;
  assign n11749 = ~n11745 & ~n11747;
  assign n11748 = n11747 & n11746;
  assign n11750 = ~n11749 & ~n11748;
  assign U3015 = ~n11751 | ~n11750;
  assign n11754 = n11771 | n11752;
  assign n11755 = ~n11754 | ~n11753;
  assign n11757 = ~n11755 | ~n11772;
  assign n11760 = ~n11757 | ~n11756;
  assign n11759 = ~n11792 & ~n11758;
  assign n11770 = ~n11760 & ~n11759;
  assign n11764 = ~n11803 | ~n11761;
  assign n11763 = ~INSTADDRPOINTER_REG_2__SCAN_IN | ~n11762;
  assign n11768 = ~n11764 | ~n11763;
  assign n11766 = ~n11765 | ~INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n11767 = ~INSTADDRPOINTER_REG_2__SCAN_IN & ~n11766;
  assign n11769 = ~n11768 & ~n11767;
  assign U3016 = ~n11770 | ~n11769;
  assign n11790 = ~n11772 | ~n11771;
  assign n11774 = ~n11790 | ~n11773;
  assign n11788 = ~n11774 | ~INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n11777 = ~n11775 & ~n11792;
  assign n11782 = ~n11777 & ~n11776;
  assign n11779 = ~n11778 & ~INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n11781 = ~n11780 | ~n11779;
  assign n11786 = ~n11782 | ~n11781;
  assign n11785 = ~n11784 & ~n11783;
  assign n11787 = ~n11786 & ~n11785;
  assign U3017 = ~n11788 | ~n11787;
  assign n11801 = ~n11790 | ~n11789;
  assign n11793 = ~n11792 & ~n11791;
  assign n11799 = ~n11794 & ~n11793;
  assign n11797 = n11796 | n11795;
  assign n11798 = ~INSTADDRPOINTER_REG_0__SCAN_IN | ~n11797;
  assign n11800 = ~n11799 | ~n11798;
  assign n11805 = ~n11801 & ~n11800;
  assign n11804 = ~n11803 | ~n11802;
  assign U3018 = ~n11805 | ~n11804;
  assign n13749 = ~n13655 | ~n11983;
  assign n11807 = n13749 & n13304;
  assign n11872 = ~n11810 | ~STATE2_REG_1__SCAN_IN;
  assign n11859 = ~INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n11811 = ~n11872 & ~n11859;
  assign n11864 = ~INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~n11811;
  assign n11845 = n13350 & INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n11848 = ~n13342;
  assign n11822 = ~n11812;
  assign n11815 = ~n11826 | ~INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n11814 = ~n11813 | ~INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n11816 = ~n11815 | ~n11814;
  assign n11817 = ~n11822 | ~n11816;
  assign n11843 = ~n11848 & ~n11817;
  assign n11850 = ~n11819 & ~n11818;
  assign n11824 = ~n11820 | ~n11809;
  assign n11823 = ~n11822 | ~n13634;
  assign n11825 = ~n11824 | ~n11823;
  assign n11827 = ~n11826 | ~n11825;
  assign n11836 = ~n11850 & ~n11827;
  assign n11832 = ~n11867;
  assign n11830 = ~n9302 | ~n11828;
  assign n11831 = ~n11830 & ~n11829;
  assign n11833 = ~n11832 | ~n11831;
  assign n13341 = ~n11834 & ~n11833;
  assign n11835 = ~n12757 & ~n13341;
  assign n11841 = ~n11836 & ~n11835;
  assign n11837 = ~n11820 | ~INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n11838 = ~n11837 | ~n11809;
  assign n13620 = ~n8537 | ~n11838;
  assign n11839 = ~n13620;
  assign n11840 = ~n11847 | ~n11839;
  assign n11842 = ~n11841 | ~n11840;
  assign n13622 = ~n11843 & ~n11842;
  assign n11844 = ~n13622 & ~n13350;
  assign n11846 = ~n13367;
  assign n11858 = ~n13350;
  assign n11857 = ~n12248 & ~n13341;
  assign n11851 = n11820 ^ ~n11859;
  assign n11855 = ~n11847 | ~n11851;
  assign n11849 = INSTQUEUERD_ADDR_REG_1__SCAN_IN ^ ~INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n11853 = ~n11849 & ~n11848;
  assign n11852 = ~n11851 & ~n11850;
  assign n11854 = ~n11853 & ~n11852;
  assign n11856 = ~n11855 | ~n11854;
  assign n13630 = ~n11857 & ~n11856;
  assign n11861 = ~n11858 | ~n13630;
  assign n11860 = ~n13350 | ~n11859;
  assign n13362 = ~n11861 | ~n11860;
  assign n11862 = ~n13362;
  assign n11863 = ~n7226 | ~n11862;
  assign n13372 = ~n11864 | ~n11863;
  assign n11866 = ~n11865;
  assign n11877 = ~n13372 | ~n11866;
  assign n11870 = ~n11868 | ~n11867;
  assign n11869 = ~INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~n13350;
  assign n11871 = ~n11870 | ~n11869;
  assign n11875 = ~n11871 | ~n13655;
  assign n11874 = n11873 | n11872;
  assign n13334 = ~n11875 | ~n11874;
  assign n11876 = ~n13334;
  assign n13305 = ~n11877 | ~n11876;
  assign n11878 = ~FLUSH_REG_SCAN_IN & ~n13305;
  assign n11879 = ~n13618 & ~n11878;
  assign U3019 = INSTQUEUEWR_ADDR_REG_4__SCAN_IN & n13710;
  assign n13188 = ~n11967 & ~n13310;
  assign n12063 = ~n12841 | ~n12240;
  assign n11984 = ~n12063 & ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n11968 = ~n11984 | ~n13354;
  assign n11883 = ~n13093 & ~n11968;
  assign n13210 = ~DATAI_24_ | ~n6996;
  assign n11882 = ~n13290 & ~n13210;
  assign n11897 = ~n11883 & ~n11882;
  assign n12259 = ~n11903 | ~STATE2_REG_2__SCAN_IN;
  assign n12764 = ~n11901 | ~n12259;
  assign n11891 = ~STATE2_REG_3__SCAN_IN | ~n11968;
  assign n13695 = ~n10880;
  assign n12596 = ~n13695 & ~n10856;
  assign n11889 = ~n12596 | ~n12757;
  assign n11885 = ~n13290;
  assign n11886 = ~n11885 & ~n11898;
  assign n11887 = ~n13100 & ~n11886;
  assign n11888 = ~n13102 & ~n11887;
  assign n11890 = ~n11889 | ~n11888;
  assign n11892 = ~n11891 | ~n11890;
  assign n11895 = ~n12764 & ~n11892;
  assign n11893 = ~n12589;
  assign n12588 = ~n12765;
  assign n12260 = ~n11893 & ~n12588;
  assign n11894 = ~n12260;
  assign n12257 = ~n11894 | ~STATE2_REG_2__SCAN_IN;
  assign n11971 = ~n11895 | ~n12257;
  assign n11896 = ~INSTQUEUE_REG_0__0__SCAN_IN | ~n11971;
  assign n11900 = ~n11897 | ~n11896;
  assign n13189 = ~DATAI_16_ | ~n6996;
  assign n11899 = ~n12052 & ~n13189;
  assign n11907 = ~n11900 & ~n11899;
  assign n13207 = ~n11902 & ~n12246;
  assign n13675 = ~n12757;
  assign n12429 = ~n13675 & ~n13102;
  assign n12675 = ~n12596;
  assign n11905 = ~n12429 | ~n12596;
  assign n12064 = n11903 | n11983;
  assign n12774 = ~n12064;
  assign n11904 = ~n12260 | ~n12774;
  assign n11973 = ~n11905 | ~n11904;
  assign n11906 = ~n13207 | ~n11973;
  assign U3020 = ~n11907 | ~n11906;
  assign n13215 = ~n11967 & ~n11908;
  assign n11910 = ~n13121 & ~n11968;
  assign n13216 = ~DATAI_25_ | ~n6996;
  assign n11909 = ~n13290 & ~n13216;
  assign n11917 = ~n11910 & ~n11909;
  assign n11913 = ~INSTQUEUE_REG_0__1__SCAN_IN | ~n11971;
  assign n13219 = ~n11911 & ~n12246;
  assign n11912 = ~n13219 | ~n11973;
  assign n11915 = ~n11913 | ~n11912;
  assign n13222 = ~DATAI_17_ | ~n6996;
  assign n11914 = ~n12052 & ~n13222;
  assign n11916 = ~n11915 & ~n11914;
  assign U3021 = ~n11917 | ~n11916;
  assign n11920 = ~n13130 & ~n11968;
  assign n13228 = ~DATAI_26_ | ~n6996;
  assign n11919 = ~n13290 & ~n13228;
  assign n11927 = ~n11920 & ~n11919;
  assign n11923 = ~INSTQUEUE_REG_0__2__SCAN_IN | ~n11971;
  assign n13231 = ~n11921 & ~n12246;
  assign n11922 = ~n13231 | ~n11973;
  assign n11925 = ~n11923 | ~n11922;
  assign n13234 = ~DATAI_18_ | ~n6996;
  assign n11924 = ~n12052 & ~n13234;
  assign n11926 = ~n11925 & ~n11924;
  assign U3022 = ~n11927 | ~n11926;
  assign n13239 = ~n11967 & ~n11928;
  assign n11930 = ~n13139 & ~n11968;
  assign n13246 = ~DATAI_27_ | ~n6996;
  assign n11929 = ~n13290 & ~n13246;
  assign n11937 = ~n11930 & ~n11929;
  assign n11933 = ~INSTQUEUE_REG_0__3__SCAN_IN | ~n11971;
  assign n13243 = ~n11931 & ~n12246;
  assign n11932 = ~n13243 | ~n11973;
  assign n11935 = ~n11933 | ~n11932;
  assign n13240 = ~DATAI_19_ | ~n6996;
  assign n11934 = ~n12052 & ~n13240;
  assign n11936 = ~n11935 & ~n11934;
  assign U3023 = ~n11937 | ~n11936;
  assign n13251 = ~n11967 & ~n11938;
  assign n11940 = ~n13148 & ~n11968;
  assign n13258 = ~DATAI_28_ | ~n6996;
  assign n11939 = ~n13290 & ~n13258;
  assign n11947 = ~n11940 & ~n11939;
  assign n11943 = ~INSTQUEUE_REG_0__4__SCAN_IN | ~n11971;
  assign n13255 = ~n11941 & ~n12246;
  assign n11942 = ~n13255 | ~n11973;
  assign n11945 = ~n11943 | ~n11942;
  assign n13252 = ~DATAI_20_ | ~n6996;
  assign n11944 = ~n12052 & ~n13252;
  assign n11946 = ~n11945 & ~n11944;
  assign U3024 = ~n11947 | ~n11946;
  assign n11950 = ~n13157 & ~n11968;
  assign n13264 = ~DATAI_29_ | ~n6996;
  assign n11949 = ~n13290 & ~n13264;
  assign n11957 = ~n11950 & ~n11949;
  assign n11953 = ~INSTQUEUE_REG_0__5__SCAN_IN | ~n11971;
  assign n13267 = ~n11951 & ~n12246;
  assign n11952 = ~n13267 | ~n11973;
  assign n11955 = ~n11953 | ~n11952;
  assign n13270 = ~DATAI_21_ | ~n6996;
  assign n11954 = ~n12052 & ~n13270;
  assign n11956 = ~n11955 & ~n11954;
  assign U3025 = ~n11957 | ~n11956;
  assign n13275 = ~n11967 & ~n7773;
  assign n11959 = ~n13166 & ~n11968;
  assign n13282 = ~DATAI_30_ | ~n6996;
  assign n11958 = ~n13290 & ~n13282;
  assign n11966 = ~n11959 & ~n11958;
  assign n11962 = ~INSTQUEUE_REG_0__6__SCAN_IN | ~n11971;
  assign n13279 = ~n11960 & ~n12246;
  assign n11961 = ~n13279 | ~n11973;
  assign n11964 = ~n11962 | ~n11961;
  assign n13276 = ~DATAI_22_ | ~n6996;
  assign n11963 = ~n12052 & ~n13276;
  assign n11965 = ~n11964 & ~n11963;
  assign U3026 = ~n11966 | ~n11965;
  assign n13288 = ~n11967 & ~n13328;
  assign n11970 = ~n13176 & ~n11968;
  assign n13298 = ~DATAI_31_ | ~n6996;
  assign n11969 = ~n13290 & ~n13298;
  assign n11979 = ~n11970 & ~n11969;
  assign n11975 = ~INSTQUEUE_REG_0__7__SCAN_IN | ~n11971;
  assign n13295 = ~n11972 & ~n12246;
  assign n11974 = ~n13295 | ~n11973;
  assign n11977 = ~n11975 | ~n11974;
  assign n13289 = ~DATAI_23_ | ~n6996;
  assign n11976 = ~n12052 & ~n13289;
  assign n11978 = ~n11977 & ~n11976;
  assign U3027 = ~n11979 | ~n11978;
  assign n12051 = ~n11984 | ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n11982 = ~n13093 & ~n12051;
  assign n11981 = ~n12150 & ~n13189;
  assign n11993 = ~n11982 & ~n11981;
  assign n11985 = ~n11984 & ~n11983;
  assign n11991 = ~n12246 & ~n11985;
  assign n12499 = n12757 & n13703;
  assign n11996 = ~n12499 | ~n12596;
  assign n12850 = ~n11884;
  assign n11986 = ~n12850 | ~STATEBS16_REG_SCAN_IN;
  assign n11987 = ~n12673 & ~n11986;
  assign n11998 = ~n13102 & ~n11987;
  assign n11988 = ~n11996 | ~n11998;
  assign n13674 = ~STATE2_REG_3__SCAN_IN;
  assign n11989 = ~n11988 | ~n13674;
  assign n11990 = ~n11989 | ~n12051;
  assign n12055 = ~n11991 | ~n11990;
  assign n11992 = ~INSTQUEUE_REG_1__0__SCAN_IN | ~n12055;
  assign n11995 = ~n11993 | ~n11992;
  assign n11994 = ~n12052 & ~n13210;
  assign n12002 = ~n11995 & ~n11994;
  assign n11997 = ~n12051 | ~n11996;
  assign n12000 = ~n11998 | ~n11997;
  assign n12162 = ~n12063 & ~n11983;
  assign n11999 = ~n12162 | ~n13355;
  assign n12056 = ~n12000 | ~n11999;
  assign n12001 = ~n13207 | ~n12056;
  assign U3028 = ~n12002 | ~n12001;
  assign n12004 = ~n13121 & ~n12051;
  assign n12003 = ~n12150 & ~n13222;
  assign n12010 = ~n12004 & ~n12003;
  assign n12006 = ~INSTQUEUE_REG_1__1__SCAN_IN | ~n12055;
  assign n12005 = ~n13219 | ~n12056;
  assign n12008 = ~n12006 | ~n12005;
  assign n12007 = ~n12052 & ~n13216;
  assign n12009 = ~n12008 & ~n12007;
  assign U3029 = ~n12010 | ~n12009;
  assign n12012 = ~n13130 & ~n12051;
  assign n12011 = ~n12052 & ~n13228;
  assign n12018 = ~n12012 & ~n12011;
  assign n12014 = ~INSTQUEUE_REG_1__2__SCAN_IN | ~n12055;
  assign n12013 = ~n13231 | ~n12056;
  assign n12016 = ~n12014 | ~n12013;
  assign n12015 = ~n12150 & ~n13234;
  assign n12017 = ~n12016 & ~n12015;
  assign U3030 = ~n12018 | ~n12017;
  assign n12020 = ~n13139 & ~n12051;
  assign n12019 = ~n12150 & ~n13240;
  assign n12026 = ~n12020 & ~n12019;
  assign n12022 = ~INSTQUEUE_REG_1__3__SCAN_IN | ~n12055;
  assign n12021 = ~n13243 | ~n12056;
  assign n12024 = ~n12022 | ~n12021;
  assign n12023 = ~n12052 & ~n13246;
  assign n12025 = ~n12024 & ~n12023;
  assign U3031 = ~n12026 | ~n12025;
  assign n12028 = ~n13148 & ~n12051;
  assign n12027 = ~n12052 & ~n13258;
  assign n12034 = ~n12028 & ~n12027;
  assign n12030 = ~INSTQUEUE_REG_1__4__SCAN_IN | ~n12055;
  assign n12029 = ~n13255 | ~n12056;
  assign n12032 = ~n12030 | ~n12029;
  assign n12031 = ~n12150 & ~n13252;
  assign n12033 = ~n12032 & ~n12031;
  assign U3032 = ~n12034 | ~n12033;
  assign n12036 = ~n13157 & ~n12051;
  assign n12035 = ~n12052 & ~n13264;
  assign n12042 = ~n12036 & ~n12035;
  assign n12038 = ~INSTQUEUE_REG_1__5__SCAN_IN | ~n12055;
  assign n12037 = ~n13267 | ~n12056;
  assign n12040 = ~n12038 | ~n12037;
  assign n12039 = ~n12150 & ~n13270;
  assign n12041 = ~n12040 & ~n12039;
  assign U3033 = ~n12042 | ~n12041;
  assign n12044 = ~n13166 & ~n12051;
  assign n12043 = ~n12150 & ~n13276;
  assign n12050 = ~n12044 & ~n12043;
  assign n12046 = ~INSTQUEUE_REG_1__6__SCAN_IN | ~n12055;
  assign n12045 = ~n13279 | ~n12056;
  assign n12048 = ~n12046 | ~n12045;
  assign n12047 = ~n12052 & ~n13282;
  assign n12049 = ~n12048 & ~n12047;
  assign U3034 = ~n12050 | ~n12049;
  assign n12054 = ~n13176 & ~n12051;
  assign n12053 = ~n12052 & ~n13298;
  assign n12062 = ~n12054 & ~n12053;
  assign n12058 = ~INSTQUEUE_REG_1__7__SCAN_IN | ~n12055;
  assign n12057 = ~n13295 | ~n12056;
  assign n12060 = ~n12058 | ~n12057;
  assign n12059 = ~n12150 & ~n13289;
  assign n12061 = ~n12060 & ~n12059;
  assign U3035 = ~n12062 | ~n12061;
  assign n12174 = ~n12063 & ~n13355;
  assign n12144 = ~n12174 | ~n13354;
  assign n12069 = ~n13093 & ~n12144;
  assign n12067 = ~n13207;
  assign n12427 = n12765 | INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n12066 = ~n12064 & ~n12427;
  assign n12756 = ~n10856 & ~n10880;
  assign n12071 = ~n12756 | ~n12757;
  assign n12065 = ~n12071 & ~n13102;
  assign n12143 = ~n12066 & ~n12065;
  assign n12068 = ~n12067 & ~n12143;
  assign n12078 = ~n12069 & ~n12068;
  assign n12167 = ~n12759 | ~n12850;
  assign n12070 = ~n12150 | ~n12235;
  assign n13193 = ~n8937 | ~n13100;
  assign n12072 = ~n12070 | ~n13193;
  assign n12073 = ~n12072 | ~n12071;
  assign n12074 = ~n12073 | ~n13674;
  assign n12076 = ~n12074 | ~n12144;
  assign n12421 = n12427 & STATE2_REG_2__SCAN_IN;
  assign n12075 = ~n12421 & ~n12764;
  assign n12147 = ~n12076 | ~n12075;
  assign n12077 = ~INSTQUEUE_REG_2__0__SCAN_IN | ~n12147;
  assign n12080 = ~n12078 | ~n12077;
  assign n12079 = ~n12150 & ~n13210;
  assign n12083 = ~n12080 & ~n12079;
  assign n12081 = ~n13189;
  assign n12082 = ~n12154 | ~n12081;
  assign U3036 = ~n12083 | ~n12082;
  assign n12084 = ~n13219;
  assign n12086 = ~n12143 & ~n12084;
  assign n12085 = ~n13121 & ~n12144;
  assign n12088 = ~n12086 & ~n12085;
  assign n12087 = ~INSTQUEUE_REG_2__1__SCAN_IN | ~n12147;
  assign n12090 = ~n12088 | ~n12087;
  assign n12089 = ~n12150 & ~n13216;
  assign n12093 = ~n12090 & ~n12089;
  assign n12091 = ~n13222;
  assign n12092 = ~n12154 | ~n12091;
  assign U3037 = ~n12093 | ~n12092;
  assign n12094 = ~n13231;
  assign n12096 = ~n12143 & ~n12094;
  assign n12095 = ~n13130 & ~n12144;
  assign n12098 = ~n12096 & ~n12095;
  assign n12097 = ~INSTQUEUE_REG_2__2__SCAN_IN | ~n12147;
  assign n12100 = ~n12098 | ~n12097;
  assign n12099 = ~n12150 & ~n13228;
  assign n12103 = ~n12100 & ~n12099;
  assign n12101 = ~n13234;
  assign n12102 = ~n12154 | ~n12101;
  assign U3038 = ~n12103 | ~n12102;
  assign n12104 = ~n13243;
  assign n12106 = ~n12143 & ~n12104;
  assign n12105 = ~n13139 & ~n12144;
  assign n12108 = ~n12106 & ~n12105;
  assign n12107 = ~INSTQUEUE_REG_2__3__SCAN_IN | ~n12147;
  assign n12110 = ~n12108 | ~n12107;
  assign n12109 = ~n12150 & ~n13246;
  assign n12112 = ~n12110 & ~n12109;
  assign n12536 = ~n13240;
  assign n12111 = ~n12154 | ~n12536;
  assign U3039 = ~n12112 | ~n12111;
  assign n12113 = ~n13255;
  assign n12115 = ~n12143 & ~n12113;
  assign n12114 = ~n13148 & ~n12144;
  assign n12117 = ~n12115 & ~n12114;
  assign n12116 = ~INSTQUEUE_REG_2__4__SCAN_IN | ~n12147;
  assign n12119 = ~n12117 | ~n12116;
  assign n12118 = ~n12150 & ~n13258;
  assign n12121 = ~n12119 & ~n12118;
  assign n12545 = ~n13252;
  assign n12120 = ~n12154 | ~n12545;
  assign U3040 = ~n12121 | ~n12120;
  assign n12122 = ~n13267;
  assign n12124 = ~n12143 & ~n12122;
  assign n12123 = ~n13157 & ~n12144;
  assign n12126 = ~n12124 & ~n12123;
  assign n12125 = ~INSTQUEUE_REG_2__5__SCAN_IN | ~n12147;
  assign n12128 = ~n12126 | ~n12125;
  assign n12127 = ~n12150 & ~n13264;
  assign n12131 = ~n12128 & ~n12127;
  assign n12129 = ~n13270;
  assign n12130 = ~n12154 | ~n12129;
  assign U3041 = ~n12131 | ~n12130;
  assign n12132 = ~n13279;
  assign n12134 = ~n12143 & ~n12132;
  assign n12133 = ~n13166 & ~n12144;
  assign n12136 = ~n12134 & ~n12133;
  assign n12135 = ~INSTQUEUE_REG_2__6__SCAN_IN | ~n12147;
  assign n12138 = ~n12136 | ~n12135;
  assign n12137 = ~n12150 & ~n13282;
  assign n12141 = ~n12138 & ~n12137;
  assign n12139 = ~n13276;
  assign n12140 = ~n12154 | ~n12139;
  assign U3042 = ~n12141 | ~n12140;
  assign n12142 = ~n13295;
  assign n12146 = ~n12143 & ~n12142;
  assign n12145 = ~n13176 & ~n12144;
  assign n12149 = ~n12146 & ~n12145;
  assign n12148 = ~INSTQUEUE_REG_2__7__SCAN_IN | ~n12147;
  assign n12152 = ~n12149 | ~n12148;
  assign n12151 = ~n12150 & ~n13298;
  assign n12156 = ~n12152 & ~n12151;
  assign n12153 = ~n13289;
  assign n12155 = ~n12154 | ~n12153;
  assign U3043 = ~n12156 | ~n12155;
  assign n12228 = ~n12174 | ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n12158 = ~n13093 & ~n12228;
  assign n12157 = ~n12235 & ~n13210;
  assign n12166 = ~n12158 & ~n12157;
  assign n13684 = n13693 | n13100;
  assign n12159 = ~n13684;
  assign n13685 = ~n13683 | ~n12159;
  assign n12160 = ~n13685 & ~n11884;
  assign n12171 = ~n13102 & ~n12160;
  assign n12161 = ~n12499 | ~n12756;
  assign n12173 = ~n12228 | ~n12161;
  assign n12164 = ~n12171 | ~n12173;
  assign n12163 = ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~n12162;
  assign n12232 = ~n12164 | ~n12163;
  assign n12165 = ~n13207 | ~n12232;
  assign n12169 = ~n12166 | ~n12165;
  assign n12168 = ~n12324 & ~n13189;
  assign n12179 = ~n12169 & ~n12168;
  assign n12170 = ~n13674 & ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n12172 = ~n12171;
  assign n12176 = ~n12173 & ~n12172;
  assign n12175 = ~n12174 & ~n8937;
  assign n12177 = ~n12176 & ~n12175;
  assign n12231 = ~n13203 | ~n12177;
  assign n12178 = ~INSTQUEUE_REG_3__0__SCAN_IN | ~n12231;
  assign U3044 = ~n12179 | ~n12178;
  assign n12181 = ~n13121 & ~n12228;
  assign n12180 = ~n12324 & ~n13222;
  assign n12187 = ~n12181 & ~n12180;
  assign n12183 = ~INSTQUEUE_REG_3__1__SCAN_IN | ~n12231;
  assign n12182 = ~n13219 | ~n12232;
  assign n12185 = ~n12183 | ~n12182;
  assign n12184 = ~n12235 & ~n13216;
  assign n12186 = ~n12185 & ~n12184;
  assign U3045 = ~n12187 | ~n12186;
  assign n12189 = ~n13130 & ~n12228;
  assign n12188 = ~n12324 & ~n13234;
  assign n12195 = ~n12189 & ~n12188;
  assign n12191 = ~INSTQUEUE_REG_3__2__SCAN_IN | ~n12231;
  assign n12190 = ~n13231 | ~n12232;
  assign n12193 = ~n12191 | ~n12190;
  assign n12192 = ~n12235 & ~n13228;
  assign n12194 = ~n12193 & ~n12192;
  assign U3046 = ~n12195 | ~n12194;
  assign n12197 = ~n13139 & ~n12228;
  assign n12196 = ~n12324 & ~n13240;
  assign n12203 = ~n12197 & ~n12196;
  assign n12199 = ~INSTQUEUE_REG_3__3__SCAN_IN | ~n12231;
  assign n12198 = ~n13243 | ~n12232;
  assign n12201 = ~n12199 | ~n12198;
  assign n12200 = ~n12235 & ~n13246;
  assign n12202 = ~n12201 & ~n12200;
  assign U3047 = ~n12203 | ~n12202;
  assign n12205 = ~n13148 & ~n12228;
  assign n12204 = ~n12235 & ~n13258;
  assign n12211 = ~n12205 & ~n12204;
  assign n12207 = ~INSTQUEUE_REG_3__4__SCAN_IN | ~n12231;
  assign n12206 = ~n13255 | ~n12232;
  assign n12209 = ~n12207 | ~n12206;
  assign n12208 = ~n12324 & ~n13252;
  assign n12210 = ~n12209 & ~n12208;
  assign U3048 = ~n12211 | ~n12210;
  assign n12213 = ~n13157 & ~n12228;
  assign n12212 = ~n12324 & ~n13270;
  assign n12219 = ~n12213 & ~n12212;
  assign n12215 = ~INSTQUEUE_REG_3__5__SCAN_IN | ~n12231;
  assign n12214 = ~n13267 | ~n12232;
  assign n12217 = ~n12215 | ~n12214;
  assign n12216 = ~n12235 & ~n13264;
  assign n12218 = ~n12217 & ~n12216;
  assign U3049 = ~n12219 | ~n12218;
  assign n12221 = ~n13166 & ~n12228;
  assign n12220 = ~n12324 & ~n13276;
  assign n12227 = ~n12221 & ~n12220;
  assign n12223 = ~INSTQUEUE_REG_3__6__SCAN_IN | ~n12231;
  assign n12222 = ~n13279 | ~n12232;
  assign n12225 = ~n12223 | ~n12222;
  assign n12224 = ~n12235 & ~n13282;
  assign n12226 = ~n12225 & ~n12224;
  assign U3050 = ~n12227 | ~n12226;
  assign n12230 = ~n13176 & ~n12228;
  assign n12229 = ~n12324 & ~n13289;
  assign n12239 = ~n12230 & ~n12229;
  assign n12234 = ~INSTQUEUE_REG_3__7__SCAN_IN | ~n12231;
  assign n12233 = ~n13295 | ~n12232;
  assign n12237 = ~n12234 | ~n12233;
  assign n12236 = ~n12235 & ~n13298;
  assign n12238 = ~n12237 & ~n12236;
  assign U3051 = ~n12239 | ~n12238;
  assign n12241 = ~n12841 | ~n13355;
  assign n12344 = ~n12241 & ~n12240;
  assign n12317 = ~n12344 | ~n13354;
  assign n12245 = ~n13093 & ~n12317;
  assign n12243 = ~n12242;
  assign n12244 = ~n12399 & ~n13189;
  assign n12268 = ~n12245 & ~n12244;
  assign n12247 = ~STATE2_REG_3__SCAN_IN | ~n12317;
  assign n12256 = ~n13110 | ~n12247;
  assign n12932 = ~n12248 & ~n13695;
  assign n12254 = ~n12932 | ~n12757;
  assign n12250 = ~n12399;
  assign n12251 = ~n12250 & ~n12249;
  assign n12252 = ~n13100 & ~n12251;
  assign n12253 = ~n13102 & ~n12252;
  assign n12255 = n12254 & n12253;
  assign n12258 = ~n12256 & ~n12255;
  assign n12320 = ~n12258 | ~n12257;
  assign n12264 = ~INSTQUEUE_REG_4__0__SCAN_IN | ~n12320;
  assign n13112 = ~n12259;
  assign n12262 = ~n12260 | ~n13112;
  assign n12261 = ~n12932 | ~n12429;
  assign n12321 = ~n12262 | ~n12261;
  assign n12263 = ~n13207 | ~n12321;
  assign n12266 = ~n12264 | ~n12263;
  assign n12265 = ~n12324 & ~n13210;
  assign n12267 = ~n12266 & ~n12265;
  assign U3052 = ~n12268 | ~n12267;
  assign n12270 = ~n13121 & ~n12317;
  assign n12269 = ~n12399 & ~n13222;
  assign n12276 = ~n12270 & ~n12269;
  assign n12272 = ~INSTQUEUE_REG_4__1__SCAN_IN | ~n12320;
  assign n12271 = ~n13219 | ~n12321;
  assign n12274 = ~n12272 | ~n12271;
  assign n12273 = ~n12324 & ~n13216;
  assign n12275 = ~n12274 & ~n12273;
  assign U3053 = ~n12276 | ~n12275;
  assign n12278 = ~n13130 & ~n12317;
  assign n12277 = ~n12399 & ~n13234;
  assign n12284 = ~n12278 & ~n12277;
  assign n12280 = ~INSTQUEUE_REG_4__2__SCAN_IN | ~n12320;
  assign n12279 = ~n13231 | ~n12321;
  assign n12282 = ~n12280 | ~n12279;
  assign n12281 = ~n12324 & ~n13228;
  assign n12283 = ~n12282 & ~n12281;
  assign U3054 = ~n12284 | ~n12283;
  assign n12286 = ~n13139 & ~n12317;
  assign n12285 = ~n12399 & ~n13240;
  assign n12292 = ~n12286 & ~n12285;
  assign n12288 = ~INSTQUEUE_REG_4__3__SCAN_IN | ~n12320;
  assign n12287 = ~n13243 | ~n12321;
  assign n12290 = ~n12288 | ~n12287;
  assign n12289 = ~n12324 & ~n13246;
  assign n12291 = ~n12290 & ~n12289;
  assign U3055 = ~n12292 | ~n12291;
  assign n12294 = ~n13148 & ~n12317;
  assign n12293 = ~n12399 & ~n13252;
  assign n12300 = ~n12294 & ~n12293;
  assign n12296 = ~INSTQUEUE_REG_4__4__SCAN_IN | ~n12320;
  assign n12295 = ~n13255 | ~n12321;
  assign n12298 = ~n12296 | ~n12295;
  assign n12297 = ~n12324 & ~n13258;
  assign n12299 = ~n12298 & ~n12297;
  assign U3056 = ~n12300 | ~n12299;
  assign n12302 = ~n13157 & ~n12317;
  assign n12301 = ~n12399 & ~n13270;
  assign n12308 = ~n12302 & ~n12301;
  assign n12304 = ~INSTQUEUE_REG_4__5__SCAN_IN | ~n12320;
  assign n12303 = ~n13267 | ~n12321;
  assign n12306 = ~n12304 | ~n12303;
  assign n12305 = ~n12324 & ~n13264;
  assign n12307 = ~n12306 & ~n12305;
  assign U3057 = ~n12308 | ~n12307;
  assign n12310 = ~n13166 & ~n12317;
  assign n12309 = ~n12399 & ~n13276;
  assign n12316 = ~n12310 & ~n12309;
  assign n12312 = ~INSTQUEUE_REG_4__6__SCAN_IN | ~n12320;
  assign n12311 = ~n13279 | ~n12321;
  assign n12314 = ~n12312 | ~n12311;
  assign n12313 = ~n12324 & ~n13282;
  assign n12315 = ~n12314 & ~n12313;
  assign U3058 = ~n12316 | ~n12315;
  assign n12319 = ~n13176 & ~n12317;
  assign n12318 = ~n12399 & ~n13289;
  assign n12328 = ~n12319 & ~n12318;
  assign n12323 = ~INSTQUEUE_REG_4__7__SCAN_IN | ~n12320;
  assign n12322 = ~n13295 | ~n12321;
  assign n12326 = ~n12323 | ~n12322;
  assign n12325 = ~n12324 & ~n13298;
  assign n12327 = ~n12326 & ~n12325;
  assign U3059 = ~n12328 | ~n12327;
  assign n12398 = ~n12344 | ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n12331 = ~n13093 & ~n12398;
  assign n12330 = ~n12483 & ~n13189;
  assign n12338 = ~n12331 & ~n12330;
  assign n12332 = ~n12499 | ~n12932;
  assign n12342 = ~n12398 | ~n12332;
  assign n12333 = ~n13693 | ~STATEBS16_REG_SCAN_IN;
  assign n12334 = ~n13665 & ~n12333;
  assign n12341 = ~n13102 & ~n12334;
  assign n12336 = ~n12342 | ~n12341;
  assign n12335 = ~n12344 | ~STATE2_REG_2__SCAN_IN;
  assign n12403 = ~n12336 | ~n12335;
  assign n12337 = ~n13207 | ~n12403;
  assign n12340 = ~n12338 | ~n12337;
  assign n12339 = ~n12399 & ~n13210;
  assign n12349 = ~n12340 & ~n12339;
  assign n12343 = ~n12341;
  assign n12346 = ~n12343 & ~n12342;
  assign n12345 = ~n12344 & ~n8937;
  assign n12347 = ~n12346 & ~n12345;
  assign n12402 = ~n13203 | ~n12347;
  assign n12348 = ~INSTQUEUE_REG_5__0__SCAN_IN | ~n12402;
  assign U3060 = ~n12349 | ~n12348;
  assign n12351 = ~n13121 & ~n12398;
  assign n12350 = ~n12483 & ~n13222;
  assign n12357 = ~n12351 & ~n12350;
  assign n12353 = ~INSTQUEUE_REG_5__1__SCAN_IN | ~n12402;
  assign n12352 = ~n13219 | ~n12403;
  assign n12355 = ~n12353 | ~n12352;
  assign n12354 = ~n12399 & ~n13216;
  assign n12356 = ~n12355 & ~n12354;
  assign U3061 = ~n12357 | ~n12356;
  assign n12359 = ~n13130 & ~n12398;
  assign n12358 = ~n12399 & ~n13228;
  assign n12365 = ~n12359 & ~n12358;
  assign n12361 = ~INSTQUEUE_REG_5__2__SCAN_IN | ~n12402;
  assign n12360 = ~n13231 | ~n12403;
  assign n12363 = ~n12361 | ~n12360;
  assign n12362 = ~n12483 & ~n13234;
  assign n12364 = ~n12363 & ~n12362;
  assign U3062 = ~n12365 | ~n12364;
  assign n12367 = ~n13139 & ~n12398;
  assign n12366 = ~n12399 & ~n13246;
  assign n12373 = ~n12367 & ~n12366;
  assign n12369 = ~INSTQUEUE_REG_5__3__SCAN_IN | ~n12402;
  assign n12368 = ~n13243 | ~n12403;
  assign n12371 = ~n12369 | ~n12368;
  assign n12370 = ~n12483 & ~n13240;
  assign n12372 = ~n12371 & ~n12370;
  assign U3063 = ~n12373 | ~n12372;
  assign n12375 = ~n13148 & ~n12398;
  assign n12374 = ~n12483 & ~n13252;
  assign n12381 = ~n12375 & ~n12374;
  assign n12377 = ~INSTQUEUE_REG_5__4__SCAN_IN | ~n12402;
  assign n12376 = ~n13255 | ~n12403;
  assign n12379 = ~n12377 | ~n12376;
  assign n12378 = ~n12399 & ~n13258;
  assign n12380 = ~n12379 & ~n12378;
  assign U3064 = ~n12381 | ~n12380;
  assign n12383 = ~n13157 & ~n12398;
  assign n12382 = ~n12399 & ~n13264;
  assign n12389 = ~n12383 & ~n12382;
  assign n12385 = ~INSTQUEUE_REG_5__5__SCAN_IN | ~n12402;
  assign n12384 = ~n13267 | ~n12403;
  assign n12387 = ~n12385 | ~n12384;
  assign n12386 = ~n12483 & ~n13270;
  assign n12388 = ~n12387 & ~n12386;
  assign U3065 = ~n12389 | ~n12388;
  assign n12391 = ~n13166 & ~n12398;
  assign n12390 = ~n12483 & ~n13276;
  assign n12397 = ~n12391 & ~n12390;
  assign n12393 = ~INSTQUEUE_REG_5__6__SCAN_IN | ~n12402;
  assign n12392 = ~n13279 | ~n12403;
  assign n12395 = ~n12393 | ~n12392;
  assign n12394 = ~n12399 & ~n13282;
  assign n12396 = ~n12395 & ~n12394;
  assign U3066 = ~n12397 | ~n12396;
  assign n12401 = ~n13176 & ~n12398;
  assign n12400 = ~n12399 & ~n13298;
  assign n12409 = ~n12401 & ~n12400;
  assign n12405 = ~INSTQUEUE_REG_5__7__SCAN_IN | ~n12402;
  assign n12404 = ~n13295 | ~n12403;
  assign n12407 = ~n12405 | ~n12404;
  assign n12406 = ~n12483 & ~n13289;
  assign n12408 = ~n12407 & ~n12406;
  assign U3067 = ~n12409 | ~n12408;
  assign n12482 = ~n12508 | ~n13354;
  assign n12412 = ~n13093 & ~n12482;
  assign n12410 = n13693 | n13701;
  assign n12411 = ~n12550 & ~n13189;
  assign n12424 = ~n12412 & ~n12411;
  assign n13096 = n13695 & n10856;
  assign n12417 = ~n12757 | ~n13096;
  assign n12413 = ~n12483;
  assign n12414 = ~n12575 & ~n12413;
  assign n12415 = ~n13100 & ~n12414;
  assign n12416 = ~n13102 & ~n12415;
  assign n12419 = ~n12417 | ~n12416;
  assign n12418 = ~n12482 | ~STATE2_REG_3__SCAN_IN;
  assign n12420 = ~n12419 | ~n12418;
  assign n12422 = ~n12421 & ~n12420;
  assign n12486 = ~n13110 | ~n12422;
  assign n12423 = ~INSTQUEUE_REG_6__0__SCAN_IN | ~n12486;
  assign n12426 = ~n12424 | ~n12423;
  assign n12425 = ~n12483 & ~n13210;
  assign n12433 = ~n12426 & ~n12425;
  assign n12428 = ~n12427;
  assign n12431 = ~n13112 | ~n12428;
  assign n13195 = ~n13096;
  assign n12430 = ~n12429 | ~n13096;
  assign n12487 = ~n12431 | ~n12430;
  assign n12432 = ~n13207 | ~n12487;
  assign U3068 = ~n12433 | ~n12432;
  assign n12435 = ~n13121 & ~n12482;
  assign n12434 = ~n12550 & ~n13222;
  assign n12441 = ~n12435 & ~n12434;
  assign n12437 = ~INSTQUEUE_REG_6__1__SCAN_IN | ~n12486;
  assign n12436 = ~n13219 | ~n12487;
  assign n12439 = ~n12437 | ~n12436;
  assign n12438 = ~n12483 & ~n13216;
  assign n12440 = ~n12439 & ~n12438;
  assign U3069 = ~n12441 | ~n12440;
  assign n12443 = ~n13130 & ~n12482;
  assign n12442 = ~n12483 & ~n13228;
  assign n12449 = ~n12443 & ~n12442;
  assign n12445 = ~INSTQUEUE_REG_6__2__SCAN_IN | ~n12486;
  assign n12444 = ~n13231 | ~n12487;
  assign n12447 = ~n12445 | ~n12444;
  assign n12446 = ~n12550 & ~n13234;
  assign n12448 = ~n12447 & ~n12446;
  assign U3070 = ~n12449 | ~n12448;
  assign n12451 = ~n13139 & ~n12482;
  assign n12450 = ~n12550 & ~n13240;
  assign n12457 = ~n12451 & ~n12450;
  assign n12453 = ~INSTQUEUE_REG_6__3__SCAN_IN | ~n12486;
  assign n12452 = ~n13243 | ~n12487;
  assign n12455 = ~n12453 | ~n12452;
  assign n12454 = ~n12483 & ~n13246;
  assign n12456 = ~n12455 & ~n12454;
  assign U3071 = ~n12457 | ~n12456;
  assign n12459 = ~n13148 & ~n12482;
  assign n12458 = ~n12483 & ~n13258;
  assign n12465 = ~n12459 & ~n12458;
  assign n12461 = ~INSTQUEUE_REG_6__4__SCAN_IN | ~n12486;
  assign n12460 = ~n13255 | ~n12487;
  assign n12463 = ~n12461 | ~n12460;
  assign n12462 = ~n12550 & ~n13252;
  assign n12464 = ~n12463 & ~n12462;
  assign U3072 = ~n12465 | ~n12464;
  assign n12467 = ~n13157 & ~n12482;
  assign n12466 = ~n12550 & ~n13270;
  assign n12473 = ~n12467 & ~n12466;
  assign n12469 = ~INSTQUEUE_REG_6__5__SCAN_IN | ~n12486;
  assign n12468 = ~n13267 | ~n12487;
  assign n12471 = ~n12469 | ~n12468;
  assign n12470 = ~n12483 & ~n13264;
  assign n12472 = ~n12471 & ~n12470;
  assign U3073 = ~n12473 | ~n12472;
  assign n12475 = ~n13166 & ~n12482;
  assign n12474 = ~n12483 & ~n13282;
  assign n12481 = ~n12475 & ~n12474;
  assign n12477 = ~INSTQUEUE_REG_6__6__SCAN_IN | ~n12486;
  assign n12476 = ~n13279 | ~n12487;
  assign n12479 = ~n12477 | ~n12476;
  assign n12478 = ~n12550 & ~n13276;
  assign n12480 = ~n12479 & ~n12478;
  assign U3074 = ~n12481 | ~n12480;
  assign n12485 = ~n13176 & ~n12482;
  assign n12484 = ~n12483 & ~n13298;
  assign n12493 = ~n12485 & ~n12484;
  assign n12489 = ~INSTQUEUE_REG_6__7__SCAN_IN | ~n12486;
  assign n12488 = ~n13295 | ~n12487;
  assign n12491 = ~n12489 | ~n12488;
  assign n12490 = ~n12550 & ~n13289;
  assign n12492 = ~n12491 & ~n12490;
  assign U3075 = ~n12493 | ~n12492;
  assign n12573 = ~n12500;
  assign n12496 = ~n13188 | ~n12573;
  assign n12494 = ~n13210;
  assign n12495 = ~n12575 | ~n12494;
  assign n12517 = n12496 & n12495;
  assign n12497 = n13684 | n13683;
  assign n12498 = ~n12497 & ~n11884;
  assign n12505 = n12498 | n13102;
  assign n12501 = ~n12499 | ~n13096;
  assign n12506 = ~n12501 | ~n12500;
  assign n12503 = ~n12505 & ~n12506;
  assign n12502 = ~n12508 & ~n8937;
  assign n12504 = ~n12503 & ~n12502;
  assign n12578 = ~n13203 | ~n12504;
  assign n12512 = ~INSTQUEUE_REG_7__0__SCAN_IN | ~n12578;
  assign n12507 = ~n12505;
  assign n12510 = ~n12507 | ~n12506;
  assign n12509 = ~n12508 | ~STATE2_REG_2__SCAN_IN;
  assign n12579 = ~n12510 | ~n12509;
  assign n12511 = ~n13207 | ~n12579;
  assign n12515 = ~n12512 | ~n12511;
  assign n12513 = n13693 | n8939;
  assign n12514 = ~n12659 & ~n13189;
  assign n12516 = ~n12515 & ~n12514;
  assign U3076 = ~n12517 | ~n12516;
  assign n12520 = ~n13215 | ~n12573;
  assign n12518 = ~n13216;
  assign n12519 = ~n12575 | ~n12518;
  assign n12526 = n12520 & n12519;
  assign n12522 = ~INSTQUEUE_REG_7__1__SCAN_IN | ~n12578;
  assign n12521 = ~n13219 | ~n12579;
  assign n12524 = ~n12522 | ~n12521;
  assign n12523 = ~n12659 & ~n13222;
  assign n12525 = ~n12524 & ~n12523;
  assign U3077 = ~n12526 | ~n12525;
  assign n12529 = ~n13227 | ~n12573;
  assign n12527 = ~n13228;
  assign n12528 = ~n12575 | ~n12527;
  assign n12535 = n12529 & n12528;
  assign n12531 = ~INSTQUEUE_REG_7__2__SCAN_IN | ~n12578;
  assign n12530 = ~n13231 | ~n12579;
  assign n12533 = ~n12531 | ~n12530;
  assign n12532 = ~n12659 & ~n13234;
  assign n12534 = ~n12533 & ~n12532;
  assign U3078 = ~n12535 | ~n12534;
  assign n12538 = ~n13239 | ~n12573;
  assign n12537 = ~n12598 | ~n12536;
  assign n12544 = n12538 & n12537;
  assign n12540 = ~INSTQUEUE_REG_7__3__SCAN_IN | ~n12578;
  assign n12539 = ~n13243 | ~n12579;
  assign n12542 = ~n12540 | ~n12539;
  assign n12541 = ~n12550 & ~n13246;
  assign n12543 = ~n12542 & ~n12541;
  assign U3079 = ~n12544 | ~n12543;
  assign n12547 = ~n13251 | ~n12573;
  assign n12546 = ~n12598 | ~n12545;
  assign n12554 = n12547 & n12546;
  assign n12549 = ~INSTQUEUE_REG_7__4__SCAN_IN | ~n12578;
  assign n12548 = ~n13255 | ~n12579;
  assign n12552 = ~n12549 | ~n12548;
  assign n12551 = ~n12550 & ~n13258;
  assign n12553 = ~n12552 & ~n12551;
  assign U3080 = ~n12554 | ~n12553;
  assign n12557 = ~n13263 | ~n12573;
  assign n12555 = ~n13264;
  assign n12556 = ~n12575 | ~n12555;
  assign n12563 = n12557 & n12556;
  assign n12559 = ~INSTQUEUE_REG_7__5__SCAN_IN | ~n12578;
  assign n12558 = ~n13267 | ~n12579;
  assign n12561 = ~n12559 | ~n12558;
  assign n12560 = ~n12659 & ~n13270;
  assign n12562 = ~n12561 & ~n12560;
  assign U3081 = ~n12563 | ~n12562;
  assign n12566 = ~n13275 | ~n12573;
  assign n12564 = ~n13282;
  assign n12565 = ~n12575 | ~n12564;
  assign n12572 = n12566 & n12565;
  assign n12568 = ~INSTQUEUE_REG_7__6__SCAN_IN | ~n12578;
  assign n12567 = ~n13279 | ~n12579;
  assign n12570 = ~n12568 | ~n12567;
  assign n12569 = ~n12659 & ~n13276;
  assign n12571 = ~n12570 & ~n12569;
  assign U3082 = ~n12572 | ~n12571;
  assign n12577 = ~n13288 | ~n12573;
  assign n12574 = ~n13298;
  assign n12576 = ~n12575 | ~n12574;
  assign n12585 = n12577 & n12576;
  assign n12581 = ~INSTQUEUE_REG_7__7__SCAN_IN | ~n12578;
  assign n12580 = ~n13295 | ~n12579;
  assign n12583 = ~n12581 | ~n12580;
  assign n12582 = ~n12659 & ~n13289;
  assign n12584 = ~n12583 & ~n12582;
  assign U3083 = ~n12585 | ~n12584;
  assign n12587 = ~n12659 & ~n13210;
  assign n12753 = ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~n12240;
  assign n12687 = ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~n12753;
  assign n12658 = ~n12687 | ~n13354;
  assign n12586 = ~n13093 & ~n12658;
  assign n12593 = ~n12587 & ~n12586;
  assign n12943 = ~n12589 & ~n12588;
  assign n12591 = ~n12943 | ~n12774;
  assign n12590 = ~n12596 | ~n7228;
  assign n12663 = ~n12591 | ~n12590;
  assign n12592 = ~n13207 | ~n12663;
  assign n12595 = ~n12593 | ~n12592;
  assign n12760 = ~n11884 | ~n8939;
  assign n12594 = ~n12748 & ~n13189;
  assign n12609 = ~n12595 & ~n12594;
  assign n12604 = ~STATE2_REG_3__SCAN_IN | ~n12658;
  assign n12602 = ~n13675 | ~n12596;
  assign n12597 = ~n12748;
  assign n12599 = ~n12598 & ~n12597;
  assign n12600 = ~n13100 & ~n12599;
  assign n12601 = ~n13102 & ~n12600;
  assign n12603 = ~n12602 | ~n12601;
  assign n12605 = ~n12604 | ~n12603;
  assign n12607 = ~n12764 & ~n12605;
  assign n12606 = ~n12943;
  assign n12939 = ~n12606 | ~STATE2_REG_2__SCAN_IN;
  assign n12608 = ~INSTQUEUE_REG_8__0__SCAN_IN | ~n12662;
  assign U3084 = ~n12609 | ~n12608;
  assign n12611 = ~n13121 & ~n12658;
  assign n12610 = ~n12659 & ~n13216;
  assign n12617 = ~n12611 & ~n12610;
  assign n12613 = ~INSTQUEUE_REG_8__1__SCAN_IN | ~n12662;
  assign n12612 = ~n13219 | ~n12663;
  assign n12615 = ~n12613 | ~n12612;
  assign n12614 = ~n12748 & ~n13222;
  assign n12616 = ~n12615 & ~n12614;
  assign U3085 = ~n12617 | ~n12616;
  assign n12619 = ~n13130 & ~n12658;
  assign n12618 = ~n12659 & ~n13228;
  assign n12625 = ~n12619 & ~n12618;
  assign n12621 = ~INSTQUEUE_REG_8__2__SCAN_IN | ~n12662;
  assign n12620 = ~n13231 | ~n12663;
  assign n12623 = ~n12621 | ~n12620;
  assign n12622 = ~n12748 & ~n13234;
  assign n12624 = ~n12623 & ~n12622;
  assign U3086 = ~n12625 | ~n12624;
  assign n12627 = ~n13139 & ~n12658;
  assign n12626 = ~n12659 & ~n13246;
  assign n12633 = ~n12627 & ~n12626;
  assign n12629 = ~INSTQUEUE_REG_8__3__SCAN_IN | ~n12662;
  assign n12628 = ~n13243 | ~n12663;
  assign n12631 = ~n12629 | ~n12628;
  assign n12630 = ~n12748 & ~n13240;
  assign n12632 = ~n12631 & ~n12630;
  assign U3087 = ~n12633 | ~n12632;
  assign n12635 = ~n13148 & ~n12658;
  assign n12634 = ~n12659 & ~n13258;
  assign n12641 = ~n12635 & ~n12634;
  assign n12637 = ~INSTQUEUE_REG_8__4__SCAN_IN | ~n12662;
  assign n12636 = ~n13255 | ~n12663;
  assign n12639 = ~n12637 | ~n12636;
  assign n12638 = ~n12748 & ~n13252;
  assign n12640 = ~n12639 & ~n12638;
  assign U3088 = ~n12641 | ~n12640;
  assign n12643 = ~n13157 & ~n12658;
  assign n12642 = ~n12659 & ~n13264;
  assign n12649 = ~n12643 & ~n12642;
  assign n12645 = ~INSTQUEUE_REG_8__5__SCAN_IN | ~n12662;
  assign n12644 = ~n13267 | ~n12663;
  assign n12647 = ~n12645 | ~n12644;
  assign n12646 = ~n12748 & ~n13270;
  assign n12648 = ~n12647 & ~n12646;
  assign U3089 = ~n12649 | ~n12648;
  assign n12651 = ~n13166 & ~n12658;
  assign n12650 = ~n12659 & ~n13282;
  assign n12657 = ~n12651 & ~n12650;
  assign n12653 = ~INSTQUEUE_REG_8__6__SCAN_IN | ~n12662;
  assign n12652 = ~n13279 | ~n12663;
  assign n12655 = ~n12653 | ~n12652;
  assign n12654 = ~n12748 & ~n13276;
  assign n12656 = ~n12655 & ~n12654;
  assign U3090 = ~n12657 | ~n12656;
  assign n12661 = ~n13176 & ~n12658;
  assign n12660 = ~n12659 & ~n13298;
  assign n12669 = ~n12661 & ~n12660;
  assign n12665 = ~INSTQUEUE_REG_8__7__SCAN_IN | ~n12662;
  assign n12664 = ~n13295 | ~n12663;
  assign n12667 = ~n12665 | ~n12664;
  assign n12666 = ~n12748 & ~n13289;
  assign n12668 = ~n12667 & ~n12666;
  assign U3091 = ~n12669 | ~n12668;
  assign n12741 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~n12687;
  assign n12671 = ~n13093 & ~n12741;
  assign n12844 = ~n11884 | ~n13701;
  assign n12670 = ~n12830 & ~n13189;
  assign n12681 = ~n12671 & ~n12670;
  assign n12672 = ~n11884 | ~STATEBS16_REG_SCAN_IN;
  assign n12674 = ~n12673 & ~n12672;
  assign n12684 = ~n13102 & ~n12674;
  assign n13335 = ~n13703;
  assign n12676 = ~n12675 & ~n13335;
  assign n12677 = ~n12676 | ~n13675;
  assign n12685 = ~n12741 | ~n12677;
  assign n12679 = ~n12684 | ~n12685;
  assign n12859 = ~n11983 & ~n12753;
  assign n12678 = ~n13355 | ~n12859;
  assign n12745 = ~n12679 | ~n12678;
  assign n12680 = ~n13207 | ~n12745;
  assign n12683 = ~n12681 | ~n12680;
  assign n12682 = ~n12748 & ~n13210;
  assign n12692 = ~n12683 & ~n12682;
  assign n12686 = ~n12684;
  assign n12689 = ~n12686 & ~n12685;
  assign n12688 = ~n8937 & ~n12687;
  assign n12690 = ~n12689 & ~n12688;
  assign n12744 = ~n13203 | ~n12690;
  assign n12691 = ~INSTQUEUE_REG_9__0__SCAN_IN | ~n12744;
  assign U3092 = ~n12692 | ~n12691;
  assign n12694 = ~n13121 & ~n12741;
  assign n12693 = ~n12748 & ~n13216;
  assign n12700 = ~n12694 & ~n12693;
  assign n12696 = ~INSTQUEUE_REG_9__1__SCAN_IN | ~n12744;
  assign n12695 = ~n13219 | ~n12745;
  assign n12698 = ~n12696 | ~n12695;
  assign n12697 = ~n12830 & ~n13222;
  assign n12699 = ~n12698 & ~n12697;
  assign U3093 = ~n12700 | ~n12699;
  assign n12702 = ~n13130 & ~n12741;
  assign n12701 = ~n12748 & ~n13228;
  assign n12708 = ~n12702 & ~n12701;
  assign n12704 = ~INSTQUEUE_REG_9__2__SCAN_IN | ~n12744;
  assign n12703 = ~n13231 | ~n12745;
  assign n12706 = ~n12704 | ~n12703;
  assign n12705 = ~n12830 & ~n13234;
  assign n12707 = ~n12706 & ~n12705;
  assign U3094 = ~n12708 | ~n12707;
  assign n12710 = ~n13139 & ~n12741;
  assign n12709 = ~n12830 & ~n13240;
  assign n12716 = ~n12710 & ~n12709;
  assign n12712 = ~INSTQUEUE_REG_9__3__SCAN_IN | ~n12744;
  assign n12711 = ~n13243 | ~n12745;
  assign n12714 = ~n12712 | ~n12711;
  assign n12713 = ~n12748 & ~n13246;
  assign n12715 = ~n12714 & ~n12713;
  assign U3095 = ~n12716 | ~n12715;
  assign n12718 = ~n13148 & ~n12741;
  assign n12717 = ~n12830 & ~n13252;
  assign n12724 = ~n12718 & ~n12717;
  assign n12720 = ~INSTQUEUE_REG_9__4__SCAN_IN | ~n12744;
  assign n12719 = ~n13255 | ~n12745;
  assign n12722 = ~n12720 | ~n12719;
  assign n12721 = ~n12748 & ~n13258;
  assign n12723 = ~n12722 & ~n12721;
  assign U3096 = ~n12724 | ~n12723;
  assign n12726 = ~n13157 & ~n12741;
  assign n12725 = ~n12748 & ~n13264;
  assign n12732 = ~n12726 & ~n12725;
  assign n12728 = ~INSTQUEUE_REG_9__5__SCAN_IN | ~n12744;
  assign n12727 = ~n13267 | ~n12745;
  assign n12730 = ~n12728 | ~n12727;
  assign n12729 = ~n12830 & ~n13270;
  assign n12731 = ~n12730 & ~n12729;
  assign U3097 = ~n12732 | ~n12731;
  assign n12734 = ~n13166 & ~n12741;
  assign n12733 = ~n12830 & ~n13276;
  assign n12740 = ~n12734 & ~n12733;
  assign n12736 = ~INSTQUEUE_REG_9__6__SCAN_IN | ~n12744;
  assign n12735 = ~n13279 | ~n12745;
  assign n12738 = ~n12736 | ~n12735;
  assign n12737 = ~n12748 & ~n13282;
  assign n12739 = ~n12738 & ~n12737;
  assign U3098 = ~n12740 | ~n12739;
  assign n12743 = ~n13176 & ~n12741;
  assign n12742 = ~n12830 & ~n13289;
  assign n12752 = ~n12743 & ~n12742;
  assign n12747 = ~INSTQUEUE_REG_9__7__SCAN_IN | ~n12744;
  assign n12746 = ~n13295 | ~n12745;
  assign n12750 = ~n12747 | ~n12746;
  assign n12749 = ~n12748 & ~n13298;
  assign n12751 = ~n12750 & ~n12749;
  assign U3099 = ~n12752 | ~n12751;
  assign n12853 = ~n13355 & ~n12753;
  assign n12829 = ~n12853 | ~n13354;
  assign n12755 = ~n13093 & ~n12829;
  assign n12754 = ~n12830 & ~n13210;
  assign n12770 = ~n12755 & ~n12754;
  assign n12758 = ~n12756;
  assign n12848 = ~n12758 & ~n12757;
  assign n12761 = ~n12830 | ~n12923;
  assign n12762 = ~n12761 | ~STATEBS16_REG_SCAN_IN;
  assign n12775 = ~n8937 | ~n12762;
  assign n12763 = ~n12848 & ~n12775;
  assign n12768 = ~n12764 & ~n12763;
  assign n12773 = n12765 | n12841;
  assign n13108 = n12773 & STATE2_REG_2__SCAN_IN;
  assign n12766 = n12829 & STATE2_REG_3__SCAN_IN;
  assign n12767 = ~n13108 & ~n12766;
  assign n12833 = ~n12768 | ~n12767;
  assign n12769 = ~INSTQUEUE_REG_10__0__SCAN_IN | ~n12833;
  assign n12772 = ~n12770 | ~n12769;
  assign n12771 = ~n12923 & ~n13189;
  assign n12780 = ~n12772 & ~n12771;
  assign n13111 = ~n12773;
  assign n12778 = ~n12774 | ~n13111;
  assign n12776 = ~n12775;
  assign n12777 = ~n12848 | ~n12776;
  assign n12834 = ~n12778 | ~n12777;
  assign n12779 = ~n13207 | ~n12834;
  assign U3100 = ~n12780 | ~n12779;
  assign n12782 = ~n13121 & ~n12829;
  assign n12781 = ~n12830 & ~n13216;
  assign n12788 = ~n12782 & ~n12781;
  assign n12784 = ~INSTQUEUE_REG_10__1__SCAN_IN | ~n12833;
  assign n12783 = ~n13219 | ~n12834;
  assign n12786 = ~n12784 | ~n12783;
  assign n12785 = ~n12923 & ~n13222;
  assign n12787 = ~n12786 & ~n12785;
  assign U3101 = ~n12788 | ~n12787;
  assign n12790 = ~n13130 & ~n12829;
  assign n12789 = ~n12830 & ~n13228;
  assign n12796 = ~n12790 & ~n12789;
  assign n12792 = ~INSTQUEUE_REG_10__2__SCAN_IN | ~n12833;
  assign n12791 = ~n13231 | ~n12834;
  assign n12794 = ~n12792 | ~n12791;
  assign n12793 = ~n12923 & ~n13234;
  assign n12795 = ~n12794 & ~n12793;
  assign U3102 = ~n12796 | ~n12795;
  assign n12798 = ~n13139 & ~n12829;
  assign n12797 = ~n12830 & ~n13246;
  assign n12804 = ~n12798 & ~n12797;
  assign n12800 = ~INSTQUEUE_REG_10__3__SCAN_IN | ~n12833;
  assign n12799 = ~n13243 | ~n12834;
  assign n12802 = ~n12800 | ~n12799;
  assign n12801 = ~n12923 & ~n13240;
  assign n12803 = ~n12802 & ~n12801;
  assign U3103 = ~n12804 | ~n12803;
  assign n12806 = ~n13148 & ~n12829;
  assign n12805 = ~n12830 & ~n13258;
  assign n12812 = ~n12806 & ~n12805;
  assign n12808 = ~INSTQUEUE_REG_10__4__SCAN_IN | ~n12833;
  assign n12807 = ~n13255 | ~n12834;
  assign n12810 = ~n12808 | ~n12807;
  assign n12809 = ~n12923 & ~n13252;
  assign n12811 = ~n12810 & ~n12809;
  assign U3104 = ~n12812 | ~n12811;
  assign n12814 = ~n13157 & ~n12829;
  assign n12813 = ~n12830 & ~n13264;
  assign n12820 = ~n12814 & ~n12813;
  assign n12816 = ~INSTQUEUE_REG_10__5__SCAN_IN | ~n12833;
  assign n12815 = ~n13267 | ~n12834;
  assign n12818 = ~n12816 | ~n12815;
  assign n12817 = ~n12923 & ~n13270;
  assign n12819 = ~n12818 & ~n12817;
  assign U3105 = ~n12820 | ~n12819;
  assign n12822 = ~n13166 & ~n12829;
  assign n12821 = ~n12830 & ~n13282;
  assign n12828 = ~n12822 & ~n12821;
  assign n12824 = ~INSTQUEUE_REG_10__6__SCAN_IN | ~n12833;
  assign n12823 = ~n13279 | ~n12834;
  assign n12826 = ~n12824 | ~n12823;
  assign n12825 = ~n12923 & ~n13276;
  assign n12827 = ~n12826 & ~n12825;
  assign U3106 = ~n12828 | ~n12827;
  assign n12832 = ~n13176 & ~n12829;
  assign n12831 = ~n12830 & ~n13298;
  assign n12840 = ~n12832 & ~n12831;
  assign n12836 = ~INSTQUEUE_REG_10__7__SCAN_IN | ~n12833;
  assign n12835 = ~n13295 | ~n12834;
  assign n12838 = ~n12836 | ~n12835;
  assign n12837 = ~n12923 & ~n13289;
  assign n12839 = ~n12838 & ~n12837;
  assign U3107 = ~n12840 | ~n12839;
  assign n12843 = ~n12841 & ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n12842 = ~n13353;
  assign n12916 = ~n12843 | ~n12842;
  assign n12847 = ~n13093 & ~n12916;
  assign n12846 = ~n13007 & ~n13189;
  assign n12867 = ~n12847 & ~n12846;
  assign n12849 = ~n12848 | ~n13703;
  assign n12857 = ~n12916 | ~n12849;
  assign n12851 = ~n13685 & ~n12850;
  assign n12858 = ~n13102 & ~n12851;
  assign n12852 = ~n12858;
  assign n12855 = ~n12857 & ~n12852;
  assign n12854 = ~n12853 & ~n8937;
  assign n12856 = ~n12855 & ~n12854;
  assign n12919 = ~n13203 | ~n12856;
  assign n12863 = ~INSTQUEUE_REG_11__0__SCAN_IN | ~n12919;
  assign n12861 = ~n12858 | ~n12857;
  assign n12860 = ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~n12859;
  assign n12920 = ~n12861 | ~n12860;
  assign n12862 = ~n13207 | ~n12920;
  assign n12865 = ~n12863 | ~n12862;
  assign n12864 = ~n12923 & ~n13210;
  assign n12866 = ~n12865 & ~n12864;
  assign U3108 = ~n12867 | ~n12866;
  assign n12869 = ~n13121 & ~n12916;
  assign n12868 = ~n12923 & ~n13216;
  assign n12875 = ~n12869 & ~n12868;
  assign n12871 = ~INSTQUEUE_REG_11__1__SCAN_IN | ~n12919;
  assign n12870 = ~n13219 | ~n12920;
  assign n12873 = ~n12871 | ~n12870;
  assign n12872 = ~n13007 & ~n13222;
  assign n12874 = ~n12873 & ~n12872;
  assign U3109 = ~n12875 | ~n12874;
  assign n12877 = ~n13130 & ~n12916;
  assign n12876 = ~n12923 & ~n13228;
  assign n12883 = ~n12877 & ~n12876;
  assign n12879 = ~INSTQUEUE_REG_11__2__SCAN_IN | ~n12919;
  assign n12878 = ~n13231 | ~n12920;
  assign n12881 = ~n12879 | ~n12878;
  assign n12880 = ~n13007 & ~n13234;
  assign n12882 = ~n12881 & ~n12880;
  assign U3110 = ~n12883 | ~n12882;
  assign n12885 = ~n13139 & ~n12916;
  assign n12884 = ~n12923 & ~n13246;
  assign n12891 = ~n12885 & ~n12884;
  assign n12887 = ~INSTQUEUE_REG_11__3__SCAN_IN | ~n12919;
  assign n12886 = ~n13243 | ~n12920;
  assign n12889 = ~n12887 | ~n12886;
  assign n12888 = ~n13007 & ~n13240;
  assign n12890 = ~n12889 & ~n12888;
  assign U3111 = ~n12891 | ~n12890;
  assign n12893 = ~n13148 & ~n12916;
  assign n12892 = ~n12923 & ~n13258;
  assign n12899 = ~n12893 & ~n12892;
  assign n12895 = ~INSTQUEUE_REG_11__4__SCAN_IN | ~n12919;
  assign n12894 = ~n13255 | ~n12920;
  assign n12897 = ~n12895 | ~n12894;
  assign n12896 = ~n13007 & ~n13252;
  assign n12898 = ~n12897 & ~n12896;
  assign U3112 = ~n12899 | ~n12898;
  assign n12901 = ~n13157 & ~n12916;
  assign n12900 = ~n13007 & ~n13270;
  assign n12907 = ~n12901 & ~n12900;
  assign n12903 = ~INSTQUEUE_REG_11__5__SCAN_IN | ~n12919;
  assign n12902 = ~n13267 | ~n12920;
  assign n12905 = ~n12903 | ~n12902;
  assign n12904 = ~n12923 & ~n13264;
  assign n12906 = ~n12905 & ~n12904;
  assign U3113 = ~n12907 | ~n12906;
  assign n12909 = ~n13166 & ~n12916;
  assign n12908 = ~n12923 & ~n13282;
  assign n12915 = ~n12909 & ~n12908;
  assign n12911 = ~INSTQUEUE_REG_11__6__SCAN_IN | ~n12919;
  assign n12910 = ~n13279 | ~n12920;
  assign n12913 = ~n12911 | ~n12910;
  assign n12912 = ~n13007 & ~n13276;
  assign n12914 = ~n12913 & ~n12912;
  assign U3114 = ~n12915 | ~n12914;
  assign n12918 = ~n13176 & ~n12916;
  assign n12917 = ~n13007 & ~n13289;
  assign n12927 = ~n12918 & ~n12917;
  assign n12922 = ~INSTQUEUE_REG_11__7__SCAN_IN | ~n12919;
  assign n12921 = ~n13295 | ~n12920;
  assign n12925 = ~n12922 | ~n12921;
  assign n12924 = ~n12923 & ~n13298;
  assign n12926 = ~n12925 & ~n12924;
  assign U3115 = ~n12927 | ~n12926;
  assign n13024 = ~n12928 & ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n13000 = ~n13024 | ~n13354;
  assign n12931 = ~n13093 & ~n13000;
  assign n12930 = ~n13082 & ~n13189;
  assign n12951 = ~n12931 & ~n12930;
  assign n13014 = ~n12932 | ~n13675;
  assign n12934 = ~n13082;
  assign n12935 = ~n12934 & ~n12933;
  assign n12936 = ~n13100 & ~n12935;
  assign n12937 = ~n13102 & ~n12936;
  assign n12941 = n13014 & n12937;
  assign n12938 = ~STATE2_REG_3__SCAN_IN | ~n13000;
  assign n12940 = ~n12939 | ~n12938;
  assign n12942 = ~n12941 & ~n12940;
  assign n13003 = ~n13110 | ~n12942;
  assign n12947 = ~INSTQUEUE_REG_12__0__SCAN_IN | ~n13003;
  assign n12945 = ~n12932 | ~n7228;
  assign n12944 = ~n12943 | ~n13112;
  assign n13004 = ~n12945 | ~n12944;
  assign n12946 = ~n13207 | ~n13004;
  assign n12949 = ~n12947 | ~n12946;
  assign n12948 = ~n13007 & ~n13210;
  assign n12950 = ~n12949 & ~n12948;
  assign U3116 = ~n12951 | ~n12950;
  assign n12953 = ~n13121 & ~n13000;
  assign n12952 = ~n13082 & ~n13222;
  assign n12959 = ~n12953 & ~n12952;
  assign n12955 = ~INSTQUEUE_REG_12__1__SCAN_IN | ~n13003;
  assign n12954 = ~n13219 | ~n13004;
  assign n12957 = ~n12955 | ~n12954;
  assign n12956 = ~n13007 & ~n13216;
  assign n12958 = ~n12957 & ~n12956;
  assign U3117 = ~n12959 | ~n12958;
  assign n12961 = ~n13130 & ~n13000;
  assign n12960 = ~n13082 & ~n13234;
  assign n12967 = ~n12961 & ~n12960;
  assign n12963 = ~INSTQUEUE_REG_12__2__SCAN_IN | ~n13003;
  assign n12962 = ~n13231 | ~n13004;
  assign n12965 = ~n12963 | ~n12962;
  assign n12964 = ~n13007 & ~n13228;
  assign n12966 = ~n12965 & ~n12964;
  assign U3118 = ~n12967 | ~n12966;
  assign n12969 = ~n13139 & ~n13000;
  assign n12968 = ~n13082 & ~n13240;
  assign n12975 = ~n12969 & ~n12968;
  assign n12971 = ~INSTQUEUE_REG_12__3__SCAN_IN | ~n13003;
  assign n12970 = ~n13243 | ~n13004;
  assign n12973 = ~n12971 | ~n12970;
  assign n12972 = ~n13007 & ~n13246;
  assign n12974 = ~n12973 & ~n12972;
  assign U3119 = ~n12975 | ~n12974;
  assign n12977 = ~n13148 & ~n13000;
  assign n12976 = ~n13082 & ~n13252;
  assign n12983 = ~n12977 & ~n12976;
  assign n12979 = ~INSTQUEUE_REG_12__4__SCAN_IN | ~n13003;
  assign n12978 = ~n13255 | ~n13004;
  assign n12981 = ~n12979 | ~n12978;
  assign n12980 = ~n13007 & ~n13258;
  assign n12982 = ~n12981 & ~n12980;
  assign U3120 = ~n12983 | ~n12982;
  assign n12985 = ~n13157 & ~n13000;
  assign n12984 = ~n13082 & ~n13270;
  assign n12991 = ~n12985 & ~n12984;
  assign n12987 = ~INSTQUEUE_REG_12__5__SCAN_IN | ~n13003;
  assign n12986 = ~n13267 | ~n13004;
  assign n12989 = ~n12987 | ~n12986;
  assign n12988 = ~n13007 & ~n13264;
  assign n12990 = ~n12989 & ~n12988;
  assign U3121 = ~n12991 | ~n12990;
  assign n12993 = ~n13166 & ~n13000;
  assign n12992 = ~n13082 & ~n13276;
  assign n12999 = ~n12993 & ~n12992;
  assign n12995 = ~INSTQUEUE_REG_12__6__SCAN_IN | ~n13003;
  assign n12994 = ~n13279 | ~n13004;
  assign n12997 = ~n12995 | ~n12994;
  assign n12996 = ~n13007 & ~n13282;
  assign n12998 = ~n12997 & ~n12996;
  assign U3122 = ~n12999 | ~n12998;
  assign n13002 = ~n13176 & ~n13000;
  assign n13001 = ~n13082 & ~n13289;
  assign n13011 = ~n13002 & ~n13001;
  assign n13006 = ~INSTQUEUE_REG_12__7__SCAN_IN | ~n13003;
  assign n13005 = ~n13295 | ~n13004;
  assign n13009 = ~n13006 | ~n13005;
  assign n13008 = ~n13007 & ~n13298;
  assign n13010 = ~n13009 & ~n13008;
  assign U3123 = ~n13011 | ~n13010;
  assign n13081 = ~n13024 | ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n13013 = ~n13093 & ~n13081;
  assign n13012 = ~n13082 & ~n13210;
  assign n13032 = ~n13013 & ~n13012;
  assign n13015 = n13014 | n13335;
  assign n13022 = ~n13081 | ~n13015;
  assign n13016 = ~n13669;
  assign n13017 = ~n13016 & ~n13100;
  assign n13023 = ~n13102 & ~n13017;
  assign n13018 = ~n13023;
  assign n13020 = ~n13022 & ~n13018;
  assign n13019 = ~n13024 & ~n8937;
  assign n13021 = ~n13020 & ~n13019;
  assign n13085 = ~n13203 | ~n13021;
  assign n13028 = ~INSTQUEUE_REG_13__0__SCAN_IN | ~n13085;
  assign n13026 = ~n13023 | ~n13022;
  assign n13025 = ~n13024 | ~STATE2_REG_2__SCAN_IN;
  assign n13086 = ~n13026 | ~n13025;
  assign n13027 = ~n13207 | ~n13086;
  assign n13030 = ~n13028 | ~n13027;
  assign n13029 = ~n13177 & ~n13189;
  assign n13031 = ~n13030 & ~n13029;
  assign U3124 = ~n13032 | ~n13031;
  assign n13034 = ~n13121 & ~n13081;
  assign n13033 = ~n13082 & ~n13216;
  assign n13040 = ~n13034 & ~n13033;
  assign n13036 = ~INSTQUEUE_REG_13__1__SCAN_IN | ~n13085;
  assign n13035 = ~n13219 | ~n13086;
  assign n13038 = ~n13036 | ~n13035;
  assign n13037 = ~n13177 & ~n13222;
  assign n13039 = ~n13038 & ~n13037;
  assign U3125 = ~n13040 | ~n13039;
  assign n13042 = ~n13130 & ~n13081;
  assign n13041 = ~n13082 & ~n13228;
  assign n13048 = ~n13042 & ~n13041;
  assign n13044 = ~INSTQUEUE_REG_13__2__SCAN_IN | ~n13085;
  assign n13043 = ~n13231 | ~n13086;
  assign n13046 = ~n13044 | ~n13043;
  assign n13045 = ~n13177 & ~n13234;
  assign n13047 = ~n13046 & ~n13045;
  assign U3126 = ~n13048 | ~n13047;
  assign n13050 = ~n13139 & ~n13081;
  assign n13049 = ~n13177 & ~n13240;
  assign n13056 = ~n13050 & ~n13049;
  assign n13052 = ~INSTQUEUE_REG_13__3__SCAN_IN | ~n13085;
  assign n13051 = ~n13243 | ~n13086;
  assign n13054 = ~n13052 | ~n13051;
  assign n13053 = ~n13082 & ~n13246;
  assign n13055 = ~n13054 & ~n13053;
  assign U3127 = ~n13056 | ~n13055;
  assign n13058 = ~n13148 & ~n13081;
  assign n13057 = ~n13082 & ~n13258;
  assign n13064 = ~n13058 & ~n13057;
  assign n13060 = ~INSTQUEUE_REG_13__4__SCAN_IN | ~n13085;
  assign n13059 = ~n13255 | ~n13086;
  assign n13062 = ~n13060 | ~n13059;
  assign n13061 = ~n13177 & ~n13252;
  assign n13063 = ~n13062 & ~n13061;
  assign U3128 = ~n13064 | ~n13063;
  assign n13066 = ~n13157 & ~n13081;
  assign n13065 = ~n13082 & ~n13264;
  assign n13072 = ~n13066 & ~n13065;
  assign n13068 = ~INSTQUEUE_REG_13__5__SCAN_IN | ~n13085;
  assign n13067 = ~n13267 | ~n13086;
  assign n13070 = ~n13068 | ~n13067;
  assign n13069 = ~n13177 & ~n13270;
  assign n13071 = ~n13070 & ~n13069;
  assign U3129 = ~n13072 | ~n13071;
  assign n13074 = ~n13166 & ~n13081;
  assign n13073 = ~n13082 & ~n13282;
  assign n13080 = ~n13074 & ~n13073;
  assign n13076 = ~INSTQUEUE_REG_13__6__SCAN_IN | ~n13085;
  assign n13075 = ~n13279 | ~n13086;
  assign n13078 = ~n13076 | ~n13075;
  assign n13077 = ~n13177 & ~n13276;
  assign n13079 = ~n13078 & ~n13077;
  assign U3130 = ~n13080 | ~n13079;
  assign n13084 = ~n13176 & ~n13081;
  assign n13083 = ~n13082 & ~n13298;
  assign n13092 = ~n13084 & ~n13083;
  assign n13088 = ~INSTQUEUE_REG_13__7__SCAN_IN | ~n13085;
  assign n13087 = ~n13295 | ~n13086;
  assign n13090 = ~n13088 | ~n13087;
  assign n13089 = ~n13177 & ~n13289;
  assign n13091 = ~n13090 & ~n13089;
  assign U3131 = ~n13092 | ~n13091;
  assign n13175 = ~n13205 | ~n13354;
  assign n13095 = ~n13093 & ~n13175;
  assign n13094 = ~n13177 & ~n13210;
  assign n13120 = ~n13095 & ~n13094;
  assign n13118 = ~n13299 & ~n13189;
  assign n13106 = ~n13175 | ~STATE2_REG_3__SCAN_IN;
  assign n13104 = ~n13675 | ~n13096;
  assign n13098 = ~n13299;
  assign n13097 = ~n13177;
  assign n13099 = ~n13098 & ~n13097;
  assign n13101 = ~n13100 & ~n13099;
  assign n13103 = ~n13102 & ~n13101;
  assign n13105 = ~n13104 | ~n13103;
  assign n13107 = ~n13106 | ~n13105;
  assign n13109 = ~n13108 & ~n13107;
  assign n13180 = ~n13110 | ~n13109;
  assign n13116 = ~INSTQUEUE_REG_14__0__SCAN_IN | ~n13180;
  assign n13114 = ~n13096 | ~n7228;
  assign n13113 = ~n13112 | ~n13111;
  assign n13181 = ~n13114 | ~n13113;
  assign n13115 = ~n13207 | ~n13181;
  assign n13117 = ~n13116 | ~n13115;
  assign n13119 = ~n13118 & ~n13117;
  assign U3132 = ~n13120 | ~n13119;
  assign n13123 = ~n13121 & ~n13175;
  assign n13122 = ~n13177 & ~n13216;
  assign n13129 = ~n13123 & ~n13122;
  assign n13125 = ~INSTQUEUE_REG_14__1__SCAN_IN | ~n13180;
  assign n13124 = ~n13219 | ~n13181;
  assign n13127 = ~n13125 | ~n13124;
  assign n13126 = ~n13299 & ~n13222;
  assign n13128 = ~n13127 & ~n13126;
  assign U3133 = ~n13129 | ~n13128;
  assign n13132 = ~n13130 & ~n13175;
  assign n13131 = ~n13177 & ~n13228;
  assign n13138 = ~n13132 & ~n13131;
  assign n13134 = ~INSTQUEUE_REG_14__2__SCAN_IN | ~n13180;
  assign n13133 = ~n13231 | ~n13181;
  assign n13136 = ~n13134 | ~n13133;
  assign n13135 = ~n13299 & ~n13234;
  assign n13137 = ~n13136 & ~n13135;
  assign U3134 = ~n13138 | ~n13137;
  assign n13141 = ~n13139 & ~n13175;
  assign n13140 = ~n13177 & ~n13246;
  assign n13147 = ~n13141 & ~n13140;
  assign n13143 = ~INSTQUEUE_REG_14__3__SCAN_IN | ~n13180;
  assign n13142 = ~n13243 | ~n13181;
  assign n13145 = ~n13143 | ~n13142;
  assign n13144 = ~n13299 & ~n13240;
  assign n13146 = ~n13145 & ~n13144;
  assign U3135 = ~n13147 | ~n13146;
  assign n13150 = ~n13148 & ~n13175;
  assign n13149 = ~n13177 & ~n13258;
  assign n13156 = ~n13150 & ~n13149;
  assign n13152 = ~INSTQUEUE_REG_14__4__SCAN_IN | ~n13180;
  assign n13151 = ~n13255 | ~n13181;
  assign n13154 = ~n13152 | ~n13151;
  assign n13153 = ~n13299 & ~n13252;
  assign n13155 = ~n13154 & ~n13153;
  assign U3136 = ~n13156 | ~n13155;
  assign n13159 = ~n13157 & ~n13175;
  assign n13158 = ~n13177 & ~n13264;
  assign n13165 = ~n13159 & ~n13158;
  assign n13161 = ~INSTQUEUE_REG_14__5__SCAN_IN | ~n13180;
  assign n13160 = ~n13267 | ~n13181;
  assign n13163 = ~n13161 | ~n13160;
  assign n13162 = ~n13299 & ~n13270;
  assign n13164 = ~n13163 & ~n13162;
  assign U3137 = ~n13165 | ~n13164;
  assign n13168 = ~n13166 & ~n13175;
  assign n13167 = ~n13177 & ~n13282;
  assign n13174 = ~n13168 & ~n13167;
  assign n13170 = ~INSTQUEUE_REG_14__6__SCAN_IN | ~n13180;
  assign n13169 = ~n13279 | ~n13181;
  assign n13172 = ~n13170 | ~n13169;
  assign n13171 = ~n13299 & ~n13276;
  assign n13173 = ~n13172 & ~n13171;
  assign U3138 = ~n13174 | ~n13173;
  assign n13179 = ~n13176 & ~n13175;
  assign n13178 = ~n13177 & ~n13298;
  assign n13187 = ~n13179 & ~n13178;
  assign n13183 = ~INSTQUEUE_REG_14__7__SCAN_IN | ~n13180;
  assign n13182 = ~n13295 | ~n13181;
  assign n13185 = ~n13183 | ~n13182;
  assign n13184 = ~n13299 & ~n13289;
  assign n13186 = ~n13185 & ~n13184;
  assign U3139 = ~n13187 | ~n13186;
  assign n13287 = ~n13197;
  assign n13191 = ~n13188 | ~n13287;
  assign n13190 = n13290 | n13189;
  assign n13214 = n13191 & n13190;
  assign n13194 = ~n13192 & ~n11881;
  assign n13673 = ~n13193;
  assign n13199 = ~n13194 & ~n13673;
  assign n13196 = ~n13195 & ~n13335;
  assign n13198 = ~n13196 | ~n13675;
  assign n13204 = ~n13198 | ~n13197;
  assign n13201 = ~n13199 & ~n13204;
  assign n13200 = ~n13205 & ~n8937;
  assign n13202 = ~n13201 & ~n13200;
  assign n13293 = ~n13203 | ~n13202;
  assign n13209 = ~INSTQUEUE_REG_15__0__SCAN_IN | ~n13293;
  assign n13206 = ~n13205 | ~STATE2_REG_2__SCAN_IN;
  assign n13294 = ~n7227 | ~n13206;
  assign n13208 = ~n13207 | ~n13294;
  assign n13212 = ~n13209 | ~n13208;
  assign n13211 = ~n13299 & ~n13210;
  assign n13213 = ~n13212 & ~n13211;
  assign U3140 = ~n13214 | ~n13213;
  assign n13218 = ~n13215 | ~n13287;
  assign n13217 = n13299 | n13216;
  assign n13226 = n13218 & n13217;
  assign n13221 = ~INSTQUEUE_REG_15__1__SCAN_IN | ~n13293;
  assign n13220 = ~n13219 | ~n13294;
  assign n13224 = ~n13221 | ~n13220;
  assign n13223 = ~n13290 & ~n13222;
  assign n13225 = ~n13224 & ~n13223;
  assign U3141 = ~n13226 | ~n13225;
  assign n13230 = ~n13227 | ~n13287;
  assign n13229 = n13299 | n13228;
  assign n13238 = n13230 & n13229;
  assign n13233 = ~INSTQUEUE_REG_15__2__SCAN_IN | ~n13293;
  assign n13232 = ~n13231 | ~n13294;
  assign n13236 = ~n13233 | ~n13232;
  assign n13235 = ~n13290 & ~n13234;
  assign n13237 = ~n13236 & ~n13235;
  assign U3142 = ~n13238 | ~n13237;
  assign n13242 = ~n13239 | ~n13287;
  assign n13241 = n13290 | n13240;
  assign n13250 = n13242 & n13241;
  assign n13245 = ~INSTQUEUE_REG_15__3__SCAN_IN | ~n13293;
  assign n13244 = ~n13243 | ~n13294;
  assign n13248 = ~n13245 | ~n13244;
  assign n13247 = ~n13299 & ~n13246;
  assign n13249 = ~n13248 & ~n13247;
  assign U3143 = ~n13250 | ~n13249;
  assign n13254 = ~n13251 | ~n13287;
  assign n13253 = n13290 | n13252;
  assign n13262 = n13254 & n13253;
  assign n13257 = ~INSTQUEUE_REG_15__4__SCAN_IN | ~n13293;
  assign n13256 = ~n13255 | ~n13294;
  assign n13260 = ~n13257 | ~n13256;
  assign n13259 = ~n13299 & ~n13258;
  assign n13261 = ~n13260 & ~n13259;
  assign U3144 = ~n13262 | ~n13261;
  assign n13266 = ~n13263 | ~n13287;
  assign n13265 = n13299 | n13264;
  assign n13274 = n13266 & n13265;
  assign n13269 = ~INSTQUEUE_REG_15__5__SCAN_IN | ~n13293;
  assign n13268 = ~n13267 | ~n13294;
  assign n13272 = ~n13269 | ~n13268;
  assign n13271 = ~n13290 & ~n13270;
  assign n13273 = ~n13272 & ~n13271;
  assign U3145 = ~n13274 | ~n13273;
  assign n13278 = ~n13275 | ~n13287;
  assign n13277 = n13290 | n13276;
  assign n13286 = n13278 & n13277;
  assign n13281 = ~INSTQUEUE_REG_15__6__SCAN_IN | ~n13293;
  assign n13280 = ~n13279 | ~n13294;
  assign n13284 = ~n13281 | ~n13280;
  assign n13283 = ~n13299 & ~n13282;
  assign n13285 = ~n13284 & ~n13283;
  assign U3146 = ~n13286 | ~n13285;
  assign n13292 = ~n13288 | ~n13287;
  assign n13291 = n13290 | n13289;
  assign n13303 = n13292 & n13291;
  assign n13297 = ~INSTQUEUE_REG_15__7__SCAN_IN | ~n13293;
  assign n13296 = ~n13295 | ~n13294;
  assign n13301 = ~n13297 | ~n13296;
  assign n13300 = ~n13299 & ~n13298;
  assign n13302 = ~n13301 & ~n13300;
  assign U3147 = ~n13303 | ~n13302;
  assign n13707 = ~n13305 & ~n13304;
  assign n13306 = ~FLUSH_REG_SCAN_IN & ~MORE_REG_SCAN_IN;
  assign n13330 = ~n13307 & ~n13306;
  assign n13309 = ~n7773;
  assign n13313 = ~n13309 & ~n13308;
  assign n13312 = ~n13311 & ~n13310;
  assign n13314 = ~n13313 | ~n13312;
  assign n13316 = ~n13314 & ~n8946;
  assign n13317 = ~n13316 & ~n13315;
  assign n13319 = ~n13318 | ~n13317;
  assign n13323 = ~n13319 | ~n13325;
  assign n13322 = n13321 | n13320;
  assign n13327 = ~n13323 | ~n13322;
  assign n13326 = ~n13325 & ~n13324;
  assign n13329 = ~n13327 & ~n13326;
  assign n13332 = ~n13330 & ~n7023;
  assign n13333 = ~n13332 | ~n13331;
  assign n13374 = ~n13334 & ~n13333;
  assign n13361 = ~n13362 | ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n13340 = ~n13335 & ~n13341;
  assign n13338 = ~n13342 & ~n13336;
  assign n13337 = ~n13345 & ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n13339 = ~n13338 & ~n13337;
  assign n13654 = ~n13340 & ~n13339;
  assign n13349 = ~n10880 & ~n13341;
  assign n13347 = ~n13342 | ~n11813;
  assign n13646 = ~n13343 | ~n13344;
  assign n13346 = ~n13345 | ~n13646;
  assign n13348 = ~n13347 | ~n13346;
  assign n13641 = ~n13349 & ~n13348;
  assign n13352 = ~n13350 & ~n13641;
  assign n13351 = ~n13355 & ~n13352;
  assign n13359 = ~n13654 & ~n13351;
  assign n13357 = ~n13353 | ~n13352;
  assign n13356 = ~n13355 | ~n13354;
  assign n13358 = ~n13357 | ~n13356;
  assign n13360 = n13359 | n13358;
  assign n13366 = ~n13361 | ~n13360;
  assign n13364 = ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~n13362;
  assign n13363 = ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~n13367;
  assign n13365 = ~n13364 & ~n13363;
  assign n13369 = ~n13366 | ~n13365;
  assign n13368 = ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~n13367;
  assign n13370 = ~n13369 | ~n13368;
  assign n13371 = ~INSTQUEUEWR_ADDR_REG_4__SCAN_IN & ~n13370;
  assign n13373 = ~n13372 & ~n13371;
  assign n13391 = ~n13374 | ~n13373;
  assign n13378 = ~n13375 | ~STATE2_REG_0__SCAN_IN;
  assign n13376 = ~STATE2_REG_1__SCAN_IN | ~READY_N;
  assign n13377 = ~n13400 | ~n13376;
  assign n13382 = ~n13378 | ~n13377;
  assign n13381 = ~n13380 & ~n13379;
  assign n13383 = ~n13382 & ~n13381;
  assign n13616 = ~STATE2_REG_2__SCAN_IN | ~n13383;
  assign n13408 = ~READY_N | ~n11983;
  assign n13397 = ~n13616 | ~n13408;
  assign n13384 = ~n13707 & ~n13397;
  assign n13389 = ~STATE2_REG_0__SCAN_IN | ~n13384;
  assign n13385 = ~n13749;
  assign n13386 = ~n13652 | ~n13385;
  assign n13387 = ~n13616 | ~n13386;
  assign n13388 = ~n13387 | ~n13400;
  assign n13395 = ~n13389 | ~n13388;
  assign n13393 = ~n13391 | ~n13390;
  assign n13394 = n13393 & n13392;
  assign U3148 = ~n13395 | ~n13394;
  assign n13396 = ~n13409 & ~n13655;
  assign n13399 = ~n13397 | ~n13396;
  assign n13407 = n13399 & n13398;
  assign n13401 = ~n13400 & ~READY_N;
  assign n13403 = ~n13402 | ~n13401;
  assign n13405 = ~n13404 | ~n13403;
  assign n13406 = ~n13405 | ~n13616;
  assign U3149 = ~n13407 | ~n13406;
  assign n13412 = ~n13408 | ~n13618;
  assign n13410 = ~n13409;
  assign n13411 = ~n13410 | ~n13749;
  assign n13413 = ~n13412 & ~n13411;
  assign U3150 = n13414 | n13413;
  assign U3151 = DATAWIDTH_REG_31__SCAN_IN & n13613;
  assign U3152 = DATAWIDTH_REG_30__SCAN_IN & n13415;
  assign U3153 = DATAWIDTH_REG_29__SCAN_IN & n13613;
  assign U3154 = DATAWIDTH_REG_28__SCAN_IN & n13613;
  assign U3155 = DATAWIDTH_REG_27__SCAN_IN & n13613;
  assign U3156 = DATAWIDTH_REG_26__SCAN_IN & n13415;
  assign U3157 = DATAWIDTH_REG_25__SCAN_IN & n13415;
  assign U3158 = DATAWIDTH_REG_24__SCAN_IN & n13415;
  assign U3159 = DATAWIDTH_REG_23__SCAN_IN & n13415;
  assign U3160 = DATAWIDTH_REG_22__SCAN_IN & n13415;
  assign U3161 = DATAWIDTH_REG_21__SCAN_IN & n13415;
  assign U3162 = DATAWIDTH_REG_20__SCAN_IN & n13415;
  assign U3163 = DATAWIDTH_REG_19__SCAN_IN & n13415;
  assign U3164 = DATAWIDTH_REG_18__SCAN_IN & n13415;
  assign U3165 = DATAWIDTH_REG_17__SCAN_IN & n13415;
  assign U3166 = DATAWIDTH_REG_16__SCAN_IN & n13415;
  assign U3167 = DATAWIDTH_REG_15__SCAN_IN & n13415;
  assign U3168 = DATAWIDTH_REG_14__SCAN_IN & n13613;
  assign U3169 = DATAWIDTH_REG_13__SCAN_IN & n13613;
  assign U3170 = DATAWIDTH_REG_12__SCAN_IN & n13613;
  assign U3171 = DATAWIDTH_REG_11__SCAN_IN & n13613;
  assign U3172 = DATAWIDTH_REG_10__SCAN_IN & n13613;
  assign U3173 = DATAWIDTH_REG_9__SCAN_IN & n13415;
  assign U3174 = DATAWIDTH_REG_8__SCAN_IN & n13613;
  assign U3175 = DATAWIDTH_REG_7__SCAN_IN & n13613;
  assign U3176 = DATAWIDTH_REG_6__SCAN_IN & n13613;
  assign U3177 = DATAWIDTH_REG_5__SCAN_IN & n13613;
  assign U3178 = DATAWIDTH_REG_4__SCAN_IN & n13613;
  assign U3179 = DATAWIDTH_REG_3__SCAN_IN & n13613;
  assign U3180 = DATAWIDTH_REG_2__SCAN_IN & n13613;
  assign n13449 = ~STATE_REG_2__SCAN_IN;
  assign n13416 = NA_N & n13433;
  assign n13417 = ~n13449 & ~n13416;
  assign n13441 = ~STATE_REG_0__SCAN_IN & ~n13417;
  assign n13429 = ~STATE_REG_1__SCAN_IN | ~STATE_REG_2__SCAN_IN;
  assign n13418 = ~n13429;
  assign n13437 = ~HOLD;
  assign n13424 = ~n13449 & ~n13437;
  assign n13446 = ~n13433 & ~n13431;
  assign n13430 = ~n13424 & ~n13446;
  assign n13419 = ~n13418 & ~n13430;
  assign n13422 = ~n13441 & ~n13419;
  assign n13423 = ~STATE_REG_1__SCAN_IN | ~HOLD;
  assign n13420 = ~REQUESTPENDING_REG_SCAN_IN | ~n13423;
  assign n13421 = ~n13756 | ~n13420;
  assign U3181 = ~n13422 | ~n13421;
  assign n13444 = ~STATE_REG_0__SCAN_IN | ~REQUESTPENDING_REG_SCAN_IN;
  assign n13426 = ~n13423 | ~n13444;
  assign n13425 = ~n13424;
  assign n13428 = ~n13426 | ~n13425;
  assign n13427 = ~n13446 & ~n13739;
  assign U3182 = ~n13428 | ~n13427;
  assign n13443 = ~n13430 & ~n13429;
  assign n13432 = ~NA_N & ~n13431;
  assign n13434 = ~n13433 & ~n13432;
  assign n13435 = ~REQUESTPENDING_REG_SCAN_IN & ~n13434;
  assign n13436 = ~n13435 & ~STATE_REG_2__SCAN_IN;
  assign n13438 = ~n13437 & ~n13436;
  assign n13440 = ~n13439 & ~n13438;
  assign n13442 = ~n13441 & ~n13440;
  assign n13448 = ~n13443 & ~n13442;
  assign n13445 = ~NA_N & ~n13444;
  assign n13447 = ~n13446 | ~n13445;
  assign U3183 = ~n13448 | ~n13447;
  assign n13451 = ~n13454 & ~n13597;
  assign n13594 = ~STATE_REG_2__SCAN_IN | ~n13757;
  assign n13569 = n13594;
  assign n13450 = ~n13569 & ~n13722;
  assign n13453 = ~n13451 & ~n13450;
  assign n13452 = ~ADDRESS_REG_0__SCAN_IN | ~n13756;
  assign U3184 = ~n13453 | ~n13452;
  assign n13459 = ~REIP_REG_3__SCAN_IN;
  assign n13456 = ~n13459 & ~n13597;
  assign n13455 = ~n13569 & ~n13454;
  assign n13458 = ~n13456 & ~n13455;
  assign n13457 = ~ADDRESS_REG_1__SCAN_IN | ~n13756;
  assign U3185 = ~n13458 | ~n13457;
  assign n13464 = ~REIP_REG_4__SCAN_IN;
  assign n13461 = ~n13464 & ~n13597;
  assign n13460 = ~n13569 & ~n13459;
  assign n13463 = ~n13461 & ~n13460;
  assign n13462 = ~ADDRESS_REG_2__SCAN_IN | ~n13756;
  assign U3186 = ~n13463 | ~n13462;
  assign n13466 = ~n13464 & ~n13594;
  assign n13465 = ~n13597 & ~n13469;
  assign n13468 = ~n13466 & ~n13465;
  assign n13467 = ~ADDRESS_REG_3__SCAN_IN | ~n13756;
  assign U3187 = ~n13468 | ~n13467;
  assign n13474 = ~REIP_REG_6__SCAN_IN;
  assign n13471 = ~n13474 & ~n13597;
  assign n13470 = ~n13569 & ~n13469;
  assign n13473 = ~n13471 & ~n13470;
  assign n13472 = ~ADDRESS_REG_4__SCAN_IN | ~n13756;
  assign U3188 = ~n13473 | ~n13472;
  assign n13476 = ~n13474 & ~n13594;
  assign n13475 = ~n13597 & ~n13479;
  assign n13478 = ~n13476 & ~n13475;
  assign n13477 = ~ADDRESS_REG_5__SCAN_IN | ~n13756;
  assign U3189 = ~n13478 | ~n13477;
  assign n13481 = ~n13479 & ~n13594;
  assign n13480 = ~n13597 & ~n13484;
  assign n13483 = ~n13481 & ~n13480;
  assign n13482 = ~ADDRESS_REG_6__SCAN_IN | ~n13756;
  assign U3190 = ~n13483 | ~n13482;
  assign n13486 = ~n13484 & ~n13594;
  assign n13485 = ~n13597 & ~n13489;
  assign n13488 = ~n13486 & ~n13485;
  assign n13487 = ~ADDRESS_REG_7__SCAN_IN | ~n13756;
  assign U3191 = ~n13488 | ~n13487;
  assign n13491 = ~n13489 & ~n13594;
  assign n13490 = ~n13597 & ~n13494;
  assign n13493 = ~n13491 & ~n13490;
  assign n13492 = ~ADDRESS_REG_8__SCAN_IN | ~n13756;
  assign U3192 = ~n13493 | ~n13492;
  assign n13496 = ~n13494 & ~n13594;
  assign n13495 = ~n13597 & ~n13499;
  assign n13498 = ~n13496 & ~n13495;
  assign n13497 = ~ADDRESS_REG_9__SCAN_IN | ~n13756;
  assign U3193 = ~n13498 | ~n13497;
  assign n13501 = ~n13499 & ~n13594;
  assign n13500 = ~n13597 & ~n13504;
  assign n13503 = ~n13501 & ~n13500;
  assign n13502 = ~ADDRESS_REG_10__SCAN_IN | ~n13756;
  assign U3194 = ~n13503 | ~n13502;
  assign n13506 = ~n13504 & ~n13594;
  assign n13505 = ~n13597 & ~n13509;
  assign n13508 = ~n13506 & ~n13505;
  assign n13507 = ~ADDRESS_REG_11__SCAN_IN | ~n13756;
  assign U3195 = ~n13508 | ~n13507;
  assign n13514 = ~REIP_REG_14__SCAN_IN;
  assign n13511 = ~n13514 & ~n13597;
  assign n13510 = ~n13569 & ~n13509;
  assign n13513 = ~n13511 & ~n13510;
  assign n13512 = ~ADDRESS_REG_12__SCAN_IN | ~n13756;
  assign U3196 = ~n13513 | ~n13512;
  assign n13516 = ~n13514 & ~n13594;
  assign n13515 = ~n13597 & ~n13519;
  assign n13518 = ~n13516 & ~n13515;
  assign n13517 = ~ADDRESS_REG_13__SCAN_IN | ~n13756;
  assign U3197 = ~n13518 | ~n13517;
  assign n13524 = ~REIP_REG_16__SCAN_IN;
  assign n13521 = ~n13524 & ~n13597;
  assign n13520 = ~n13594 & ~n13519;
  assign n13523 = ~n13521 & ~n13520;
  assign n13522 = ~ADDRESS_REG_14__SCAN_IN | ~n13756;
  assign U3198 = ~n13523 | ~n13522;
  assign n13526 = ~n13524 & ~n13594;
  assign n13525 = ~n13597 & ~n13529;
  assign n13528 = ~n13526 & ~n13525;
  assign n13527 = ~ADDRESS_REG_15__SCAN_IN | ~n13756;
  assign U3199 = ~n13528 | ~n13527;
  assign n13531 = ~n13529 & ~n13594;
  assign n13530 = ~n13597 & ~n13534;
  assign n13533 = ~n13531 & ~n13530;
  assign n13532 = ~ADDRESS_REG_16__SCAN_IN | ~n13756;
  assign U3200 = ~n13533 | ~n13532;
  assign n13536 = ~n13539 & ~n13597;
  assign n13535 = ~n13569 & ~n13534;
  assign n13538 = ~n13536 & ~n13535;
  assign n13537 = ~ADDRESS_REG_17__SCAN_IN | ~n13756;
  assign U3201 = ~n13538 | ~n13537;
  assign n13541 = ~n10045 & ~n13597;
  assign n13540 = ~n13594 & ~n13539;
  assign n13543 = ~n13541 & ~n13540;
  assign n13542 = ~ADDRESS_REG_18__SCAN_IN | ~n13756;
  assign U3202 = ~n13543 | ~n13542;
  assign n13545 = ~n10045 & ~n13594;
  assign n13544 = ~n13597 & ~n13548;
  assign n13547 = ~n13545 & ~n13544;
  assign n13546 = ~ADDRESS_REG_19__SCAN_IN | ~n13756;
  assign U3203 = ~n13547 | ~n13546;
  assign n13550 = ~n13548 & ~n13594;
  assign n13549 = ~n13597 & ~n13553;
  assign n13552 = ~n13550 & ~n13549;
  assign n13551 = ~ADDRESS_REG_20__SCAN_IN | ~n13756;
  assign U3204 = ~n13552 | ~n13551;
  assign n13555 = ~n13553 & ~n13594;
  assign n13554 = ~n13597 & ~n13558;
  assign n13557 = ~n13555 & ~n13554;
  assign n13556 = ~ADDRESS_REG_21__SCAN_IN | ~n13756;
  assign U3205 = ~n13557 | ~n13556;
  assign n13560 = ~n13558 & ~n13594;
  assign n13559 = ~n13597 & ~n13563;
  assign n13562 = ~n13560 & ~n13559;
  assign n13561 = ~ADDRESS_REG_22__SCAN_IN | ~n13756;
  assign U3206 = ~n13562 | ~n13561;
  assign n13565 = ~n13563 & ~n13594;
  assign n13564 = ~n13597 & ~n13568;
  assign n13567 = ~n13565 & ~n13564;
  assign n13566 = ~ADDRESS_REG_23__SCAN_IN | ~n13756;
  assign U3207 = ~n13567 | ~n13566;
  assign n13574 = ~REIP_REG_26__SCAN_IN;
  assign n13571 = ~n13574 & ~n13597;
  assign n13570 = ~n13569 & ~n13568;
  assign n13573 = ~n13571 & ~n13570;
  assign n13572 = ~ADDRESS_REG_24__SCAN_IN | ~n13756;
  assign U3208 = ~n13573 | ~n13572;
  assign n13576 = ~n13574 & ~n13594;
  assign n13579 = ~REIP_REG_27__SCAN_IN;
  assign n13575 = ~n13597 & ~n13579;
  assign n13578 = ~n13576 & ~n13575;
  assign n13577 = ~ADDRESS_REG_25__SCAN_IN | ~n13756;
  assign U3209 = ~n13578 | ~n13577;
  assign n13581 = ~n13579 & ~n13594;
  assign n13580 = ~n13597 & ~n13584;
  assign n13583 = ~n13581 & ~n13580;
  assign n13582 = ~ADDRESS_REG_26__SCAN_IN | ~n13756;
  assign U3210 = ~n13583 | ~n13582;
  assign n13586 = ~n13584 & ~n13594;
  assign n13585 = ~n13597 & ~n13589;
  assign n13588 = ~n13586 & ~n13585;
  assign n13587 = ~ADDRESS_REG_27__SCAN_IN | ~n13756;
  assign U3211 = ~n13588 | ~n13587;
  assign n13591 = ~n13589 & ~n13594;
  assign n13595 = ~REIP_REG_30__SCAN_IN;
  assign n13590 = ~n13597 & ~n13595;
  assign n13593 = ~n13591 & ~n13590;
  assign n13592 = ~ADDRESS_REG_28__SCAN_IN | ~n13756;
  assign U3212 = ~n13593 | ~n13592;
  assign n13599 = ~n13595 & ~n13594;
  assign n13596 = ~REIP_REG_31__SCAN_IN;
  assign n13598 = ~n13597 & ~n13596;
  assign n13601 = ~n13599 & ~n13598;
  assign n13600 = ~ADDRESS_REG_29__SCAN_IN | ~n13756;
  assign U3213 = ~n13601 | ~n13600;
  assign n13603 = ~BE_N_REG_3__SCAN_IN | ~n13756;
  assign n13602 = ~BYTEENABLE_REG_3__SCAN_IN | ~n13757;
  assign U3445 = ~n13603 | ~n13602;
  assign n13605 = ~BE_N_REG_2__SCAN_IN | ~n13756;
  assign n13604 = ~BYTEENABLE_REG_2__SCAN_IN | ~n13757;
  assign U3446 = ~n13605 | ~n13604;
  assign n13607 = ~BE_N_REG_1__SCAN_IN | ~n13756;
  assign n13606 = ~BYTEENABLE_REG_1__SCAN_IN | ~n13757;
  assign U3447 = ~n13607 | ~n13606;
  assign n13609 = ~BE_N_REG_0__SCAN_IN | ~n13756;
  assign n13608 = ~BYTEENABLE_REG_0__SCAN_IN | ~n13757;
  assign U3448 = ~n13609 | ~n13608;
  assign n13612 = ~n13615;
  assign n13611 = ~DATAWIDTH_REG_0__SCAN_IN & ~n13610;
  assign U3451 = ~n13612 & ~n13611;
  assign n13614 = ~DATAWIDTH_REG_1__SCAN_IN | ~n13613;
  assign U3452 = ~n13615 | ~n13614;
  assign n13617 = ~n13616 | ~STATE2_REG_0__SCAN_IN;
  assign n13619 = ~n13617 | ~STATE2_REG_3__SCAN_IN;
  assign U3453 = ~n13619 | ~n13618;
  assign n13621 = ~n13652;
  assign n13624 = ~n13621 & ~n13620;
  assign n13623 = ~n13622 & ~n13653;
  assign n13625 = n13624 | n13623;
  assign n13627 = ~n13625 | ~n13661;
  assign n13626 = ~INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~n13662;
  assign U3456 = ~n13627 | ~n13626;
  assign n13628 = ~n13652 | ~n13634;
  assign n13629 = ~n13661 | ~n13628;
  assign n13640 = ~n13629 | ~INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n13633 = ~n13630 & ~n13653;
  assign n13643 = INSTADDRPOINTER_REG_31__SCAN_IN ^ INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n13631 = ~n13643;
  assign n13642 = ~STATE2_REG_1__SCAN_IN | ~INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n13632 = ~n13631 & ~n13642;
  assign n13637 = ~n13633 & ~n13632;
  assign n13635 = ~n13634 & ~INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n13636 = ~n13652 | ~n13635;
  assign n13638 = ~n13637 | ~n13636;
  assign n13639 = ~n13638 | ~n13661;
  assign U3459 = ~n13640 | ~n13639;
  assign n13645 = ~n13641 & ~n13653;
  assign n13644 = ~n13643 & ~n13642;
  assign n13648 = ~n13645 & ~n13644;
  assign n13647 = ~n13652 | ~n13646;
  assign n13649 = ~n13648 | ~n13647;
  assign n13651 = ~n13661 | ~n13649;
  assign n13650 = ~INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~n13662;
  assign U3460 = ~n13651 | ~n13650;
  assign n13659 = ~n13652 | ~n13336;
  assign n13657 = ~n13654 & ~n13653;
  assign n13656 = ~n13655 & ~INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n13658 = ~n13657 & ~n13656;
  assign n13660 = ~n13659 | ~n13658;
  assign n13664 = ~n13661 | ~n13660;
  assign n13663 = ~INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~n13662;
  assign U3461 = ~n13664 | ~n13663;
  assign n13709 = ~n13710;
  assign n13666 = ~n13665;
  assign n13668 = ~n13666 | ~n7848;
  assign n13667 = ~n13683 | ~n11884;
  assign n13670 = ~n13668 | ~n13667;
  assign n13672 = ~n13670 & ~n13669;
  assign n13671 = ~n8937 | ~STATEBS16_REG_SCAN_IN;
  assign n13679 = ~n13672 & ~n13671;
  assign n13677 = ~n11884 | ~n13673;
  assign n13702 = ~n13674 | ~STATE2_REG_1__SCAN_IN;
  assign n13676 = ~n13675 | ~n13702;
  assign n13678 = ~n13677 | ~n13676;
  assign n13680 = n13679 | n13678;
  assign n13682 = ~n13709 | ~n13680;
  assign n13681 = ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~n13710;
  assign U3462 = ~n13682 | ~n13681;
  assign n13686 = ~n7833 | ~n13684;
  assign n13687 = ~n13686 | ~n13685;
  assign n13689 = ~n13687 | ~n8937;
  assign n13688 = ~n10856 | ~n13702;
  assign n13690 = ~n13689 | ~n13688;
  assign n13692 = ~n13709 | ~n13690;
  assign n13691 = ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~n13710;
  assign U3463 = ~n13692 | ~n13691;
  assign n13694 = n13693 ^ ~STATEBS16_REG_SCAN_IN;
  assign n13697 = ~n13694 | ~n8937;
  assign n13696 = ~n13695 | ~n13702;
  assign n13698 = ~n13697 | ~n13696;
  assign n13700 = ~n13709 | ~n13698;
  assign n13699 = ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~n13710;
  assign U3464 = ~n13700 | ~n13699;
  assign n13705 = ~n13701 | ~n8937;
  assign n13704 = ~n13703 | ~n13702;
  assign n13706 = ~n13705 | ~n13704;
  assign n13708 = n13707 | n13706;
  assign n13712 = ~n13709 | ~n13708;
  assign n13711 = ~n13710 | ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign U3465 = ~n13712 | ~n13711;
  assign n13721 = ~BYTEENABLE_REG_2__SCAN_IN | ~n13726;
  assign n13715 = ~n13713;
  assign n13714 = ~DATAWIDTH_REG_0__SCAN_IN | ~n13723;
  assign n13716 = ~n13715 | ~n13714;
  assign n13718 = ~n13722 | ~n13716;
  assign n13717 = ~REIP_REG_1__SCAN_IN | ~REIP_REG_0__SCAN_IN;
  assign n13719 = ~n13718 | ~n13717;
  assign n13720 = ~n13724 | ~n13719;
  assign U3468 = ~n13721 | ~n13720;
  assign n13725 = ~n13723 | ~n13722;
  assign n13728 = ~n13725 | ~n13724;
  assign n13727 = ~BYTEENABLE_REG_0__SCAN_IN | ~n13726;
  assign U3469 = ~n13728 | ~n13727;
  assign n13730 = ~W_R_N_REG_SCAN_IN | ~n13756;
  assign n13729 = READREQUEST_REG_SCAN_IN | n13756;
  assign U3470 = ~n13730 | ~n13729;
  assign n13734 = ~MORE_REG_SCAN_IN | ~n13731;
  assign n13732 = ~n13731;
  assign n13733 = ~n13732 | ~n7023;
  assign U3471 = ~n13734 | ~n13733;
  assign n13738 = ~n13735 & ~READY_N;
  assign n13761 = ~n13764;
  assign n13737 = n13761 | n13736;
  assign n13753 = ~n13738 & ~n13737;
  assign n13752 = ~n13753;
  assign n13740 = ~n13739 | ~STATEBS16_REG_SCAN_IN;
  assign n13745 = ~n13741 | ~n13740;
  assign n13744 = ~n13743 | ~n13742;
  assign n13746 = ~n13745 | ~n13744;
  assign n13747 = ~READY_N & ~n13746;
  assign n13748 = ~STATE2_REG_2__SCAN_IN | ~n13747;
  assign n13750 = ~STATE2_REG_0__SCAN_IN | ~n13748;
  assign n13751 = ~n13750 | ~n13749;
  assign n13755 = ~n13752 | ~n13751;
  assign n13754 = ~n13753 | ~REQUESTPENDING_REG_SCAN_IN;
  assign U3472 = ~n13755 | ~n13754;
  assign n13759 = ~M_IO_N_REG_SCAN_IN | ~n13756;
  assign n13758 = ~MEMORYFETCH_REG_SCAN_IN | ~n13757;
  assign U3473 = ~n13759 | ~n13758;
  assign n13766 = ~n13761 | ~n13760;
  assign n13763 = n13762 | READREQUEST_REG_SCAN_IN;
  assign n13765 = ~n13764 | ~n13763;
  assign U3474 = ~n13766 | ~n13765;
  assign n11918 = n7325 & n7324;
  assign n7512 = n7460 | n7459;
  assign n13336 = ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
endmodule


