

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125;

  NOR3_X1 U11161 ( .A1(n16077), .A2(n13826), .A3(n18792), .ZN(n17334) );
  NAND2_X1 U11162 ( .A1(n11681), .A2(n19106), .ZN(n11705) );
  INV_X2 U11163 ( .A(n11763), .ZN(n12139) );
  OAI21_X1 U11164 ( .B1(n13485), .B2(n11075), .A(n10984), .ZN(n13566) );
  CLKBUF_X2 U11165 ( .A(n12107), .Z(n9719) );
  OR2_X1 U11166 ( .A1(n11487), .A2(n11483), .ZN(n19462) );
  OR2_X1 U11167 ( .A1(n11487), .A2(n11486), .ZN(n13709) );
  NAND2_X1 U11168 ( .A1(n9844), .A2(n11470), .ZN(n19537) );
  OAI21_X1 U11169 ( .B1(n20207), .B2(n11075), .A(n10987), .ZN(n13043) );
  AND2_X1 U11170 ( .A1(n14140), .A2(n20841), .ZN(n11588) );
  NAND2_X1 U11171 ( .A1(n13272), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14153) );
  AND2_X1 U11172 ( .A1(n14129), .A2(n11510), .ZN(n14163) );
  CLKBUF_X2 U11173 ( .A(n12598), .Z(n17291) );
  CLKBUF_X1 U11174 ( .A(n12479), .Z(n13891) );
  INV_X1 U11175 ( .A(n13871), .ZN(n17063) );
  CLKBUF_X1 U11176 ( .A(n12598), .Z(n17190) );
  CLKBUF_X2 U11177 ( .A(n10353), .Z(n10875) );
  CLKBUF_X2 U11178 ( .A(n10320), .Z(n10900) );
  NOR2_X1 U11179 ( .A1(n10447), .A2(n20135), .ZN(n13055) );
  CLKBUF_X2 U11180 ( .A(n10315), .Z(n10870) );
  CLKBUF_X2 U11181 ( .A(n11379), .Z(n12957) );
  AND4_X1 U11182 ( .A1(n10306), .A2(n10305), .A3(n10304), .A4(n10303), .ZN(
        n10312) );
  INV_X1 U11183 ( .A(n12954), .ZN(n11381) );
  CLKBUF_X1 U11184 ( .A(n19096), .Z(n9717) );
  NOR2_X1 U11185 ( .A1(n19060), .A2(n19757), .ZN(n19096) );
  AND2_X1 U11186 ( .A1(n9849), .A2(n9848), .ZN(n9847) );
  CLKBUF_X2 U11187 ( .A(n10868), .Z(n10890) );
  AND4_X1 U11188 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        n10298) );
  AOI22_X1 U11190 ( .A1(n20875), .A2(keyinput108), .B1(n20874), .B2(keyinput24), .ZN(n20873) );
  OR2_X1 U11191 ( .A1(n11478), .A2(n11483), .ZN(n19349) );
  NAND2_X1 U11192 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18900), .ZN(
        n12397) );
  OAI221_X1 U11193 ( .B1(n20875), .B2(keyinput108), .C1(n20874), .C2(
        keyinput24), .A(n20873), .ZN(n20879) );
  NAND2_X1 U11194 ( .A1(n11306), .A2(n11370), .ZN(n12367) );
  AND2_X1 U11195 ( .A1(n11500), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11571) );
  AND2_X1 U11196 ( .A1(n11353), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11575) );
  NAND2_X1 U11197 ( .A1(n9844), .A2(n11484), .ZN(n19572) );
  NOR2_X1 U11198 ( .A1(n12397), .A2(n12406), .ZN(n12439) );
  AND3_X1 U11199 ( .A1(n10184), .A2(n10183), .A3(n10182), .ZN(n10185) );
  AND2_X1 U11200 ( .A1(n10629), .A2(n10628), .ZN(n13412) );
  AND2_X1 U11201 ( .A1(n14714), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14715) );
  AND2_X1 U11202 ( .A1(n11069), .A2(n14912), .ZN(n14724) );
  OAI21_X1 U11203 ( .B1(n14795), .B2(n9721), .A(n11066), .ZN(n14765) );
  NAND2_X1 U11204 ( .A1(n11366), .A2(n12954), .ZN(n11386) );
  CLKBUF_X3 U11205 ( .A(n11457), .Z(n11464) );
  INV_X1 U11206 ( .A(n9740), .ZN(n19098) );
  INV_X1 U11207 ( .A(n12359), .ZN(n19943) );
  INV_X1 U11208 ( .A(n9771), .ZN(n17269) );
  NOR2_X1 U11209 ( .A1(n18104), .A2(n12680), .ZN(n18008) );
  XNOR2_X1 U11210 ( .A(n11705), .B(n20980), .ZN(n13686) );
  INV_X1 U11211 ( .A(n13961), .ZN(n13962) );
  INV_X1 U11212 ( .A(n20039), .ZN(n20030) );
  AOI211_X1 U11213 ( .C1(n16151), .C2(n14760), .A(n14759), .B(n14758), .ZN(
        n14761) );
  INV_X1 U11214 ( .A(n17730), .ZN(n17817) );
  INV_X1 U11215 ( .A(n11366), .ZN(n11689) );
  INV_X2 U11216 ( .A(n18280), .ZN(n18198) );
  NAND2_X2 U11217 ( .A1(n15601), .A2(n15571), .ZN(n15595) );
  NOR2_X4 U11218 ( .A1(n13997), .A2(n16296), .ZN(n14016) );
  XNOR2_X2 U11219 ( .A(n11758), .B(n16471), .ZN(n13767) );
  INV_X1 U11220 ( .A(n10163), .ZN(n9718) );
  BUF_X2 U11221 ( .A(n10977), .Z(n13485) );
  AND2_X1 U11222 ( .A1(n12088), .A2(n19757), .ZN(n12107) );
  INV_X8 U11223 ( .A(n9772), .ZN(n17220) );
  AND2_X4 U11224 ( .A1(n10181), .A2(n13188), .ZN(n10356) );
  BUF_X4 U11225 ( .A(n12439), .Z(n17256) );
  INV_X1 U11226 ( .A(n11689), .ZN(n9720) );
  NAND2_X2 U11227 ( .A1(n11277), .A2(n11276), .ZN(n11366) );
  INV_X2 U11228 ( .A(n9720), .ZN(n19325) );
  XNOR2_X2 U11229 ( .A(n11985), .B(n11986), .ZN(n11983) );
  NAND2_X2 U11230 ( .A1(n11382), .A2(n12742), .ZN(n15928) );
  AOI21_X2 U11231 ( .B1(n15816), .B2(n15814), .A(n15569), .ZN(n15614) );
  NAND2_X2 U11232 ( .A1(n15568), .A2(n15838), .ZN(n15816) );
  XNOR2_X2 U11233 ( .A(n9920), .B(n10551), .ZN(n20207) );
  NAND2_X1 U11234 ( .A1(n9838), .A2(n14261), .ZN(n14264) );
  OR2_X1 U11235 ( .A1(n12515), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12518) );
  NAND2_X1 U11236 ( .A1(n9901), .A2(n11023), .ZN(n13655) );
  AND2_X1 U11237 ( .A1(n15259), .A2(n9826), .ZN(n15195) );
  INV_X4 U11238 ( .A(n14734), .ZN(n9721) );
  OR2_X1 U11239 ( .A1(n11489), .A2(n11488), .ZN(n11603) );
  AND2_X2 U11240 ( .A1(n13049), .A2(n11463), .ZN(n9844) );
  AND2_X1 U11241 ( .A1(n10574), .A2(n10573), .ZN(n15065) );
  INV_X2 U11242 ( .A(n18029), .ZN(n18767) );
  AND2_X1 U11243 ( .A1(n11778), .A2(n11776), .ZN(n11782) );
  OAI21_X1 U11244 ( .B1(n16662), .B2(n12627), .A(n18784), .ZN(n15966) );
  BUF_X4 U11245 ( .A(n12012), .Z(n12076) );
  INV_X2 U11246 ( .A(n17491), .ZN(n12477) );
  AND3_X1 U11247 ( .A1(n9785), .A2(n12448), .A3(n10061), .ZN(n17491) );
  CLKBUF_X2 U11248 ( .A(n11308), .Z(n12358) );
  CLKBUF_X2 U11250 ( .A(n10391), .Z(n20161) );
  CLKBUF_X2 U11251 ( .A(n12479), .Z(n17288) );
  CLKBUF_X3 U11252 ( .A(n12556), .Z(n9726) );
  INV_X1 U11253 ( .A(n12418), .ZN(n17006) );
  INV_X4 U11254 ( .A(n12446), .ZN(n9722) );
  BUF_X2 U11255 ( .A(n12450), .Z(n17157) );
  BUF_X1 U11256 ( .A(n12450), .Z(n17292) );
  BUF_X2 U11257 ( .A(n10313), .Z(n10856) );
  BUF_X2 U11258 ( .A(n10673), .Z(n10892) );
  CLKBUF_X2 U11259 ( .A(n10352), .Z(n10851) );
  OR2_X1 U11260 ( .A1(n12407), .A2(n17039), .ZN(n9772) );
  OR2_X1 U11261 ( .A1(n17039), .A2(n12402), .ZN(n10163) );
  INV_X1 U11262 ( .A(n9771), .ZN(n15952) );
  CLKBUF_X2 U11263 ( .A(n10397), .Z(n9723) );
  CLKBUF_X2 U11264 ( .A(n10398), .Z(n10877) );
  BUF_X2 U11265 ( .A(n10321), .Z(n10898) );
  AND2_X2 U11266 ( .A1(n10575), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13457) );
  NAND2_X2 U11267 ( .A1(n18908), .A2(n18914), .ZN(n17039) );
  NAND2_X1 U11268 ( .A1(n10051), .A2(n10052), .ZN(n11126) );
  AOI211_X1 U11269 ( .C1(n15651), .C2(n16460), .A(n15650), .B(n15649), .ZN(
        n15652) );
  AOI211_X1 U11270 ( .C1(n15638), .C2(n16460), .A(n15637), .B(n15636), .ZN(
        n15639) );
  XNOR2_X1 U11271 ( .A(n14741), .B(n14740), .ZN(n14942) );
  NAND2_X1 U11272 ( .A1(n14264), .A2(n9837), .ZN(n15400) );
  AND3_X1 U11273 ( .A1(n14745), .A2(n11068), .A3(n9836), .ZN(n14723) );
  NOR2_X1 U11274 ( .A1(n15789), .A2(n15790), .ZN(n16339) );
  AND2_X1 U11275 ( .A1(n10139), .A2(n10140), .ZN(n15515) );
  XNOR2_X1 U11276 ( .A(n10113), .B(n14070), .ZN(n14721) );
  NAND2_X1 U11277 ( .A1(n15408), .A2(n9748), .ZN(n9838) );
  AND2_X2 U11278 ( .A1(n14393), .A2(n10111), .ZN(n14066) );
  AND2_X1 U11279 ( .A1(n14784), .A2(n14753), .ZN(n11068) );
  OR2_X1 U11280 ( .A1(n15708), .A2(n11982), .ZN(n15551) );
  OR2_X1 U11281 ( .A1(n15706), .A2(n15705), .ZN(n15708) );
  NAND2_X1 U11282 ( .A1(n15598), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16381) );
  OR2_X1 U11283 ( .A1(n14217), .A2(n14216), .ZN(n14218) );
  NAND2_X1 U11284 ( .A1(n9915), .A2(n9721), .ZN(n14794) );
  AND2_X1 U11285 ( .A1(n10085), .A2(n10081), .ZN(n16060) );
  AND2_X1 U11286 ( .A1(n16287), .A2(n14195), .ZN(n14172) );
  AOI22_X1 U11287 ( .A1(n18265), .A2(n17985), .B1(n18181), .B2(n17984), .ZN(
        n17987) );
  AOI21_X1 U11288 ( .B1(n15148), .B2(n16493), .A(n15494), .ZN(n12382) );
  NAND2_X1 U11289 ( .A1(n9971), .A2(n13688), .ZN(n13692) );
  NAND2_X1 U11290 ( .A1(n13721), .A2(n13720), .ZN(n13719) );
  NAND2_X1 U11291 ( .A1(n13953), .A2(n10723), .ZN(n14629) );
  NAND2_X1 U11292 ( .A1(n10087), .A2(n10088), .ZN(n9971) );
  AOI211_X1 U11293 ( .C1(n15647), .C2(n16493), .A(n15646), .B(n15645), .ZN(
        n15648) );
  OAI21_X1 U11294 ( .B1(n13655), .B2(n13656), .A(n11030), .ZN(n13721) );
  NAND2_X1 U11295 ( .A1(n15138), .A2(n12341), .ZN(n14337) );
  NOR2_X1 U11296 ( .A1(n9919), .A2(n9918), .ZN(n9917) );
  CLKBUF_X1 U11297 ( .A(n11961), .Z(n11966) );
  AND2_X1 U11298 ( .A1(n9778), .A2(n15161), .ZN(n15656) );
  NAND2_X1 U11299 ( .A1(n17641), .A2(n17995), .ZN(n17640) );
  OAI21_X1 U11300 ( .B1(n14347), .B2(n12335), .A(n9775), .ZN(n16280) );
  MUX2_X1 U11301 ( .A(n17983), .B(n17982), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n17985) );
  AND2_X1 U11302 ( .A1(n12512), .A2(n12511), .ZN(n17641) );
  NAND2_X1 U11303 ( .A1(n9902), .A2(n11013), .ZN(n13537) );
  OR3_X2 U11304 ( .A1(n15171), .A2(n10025), .A3(n14346), .ZN(n9775) );
  NOR2_X1 U11305 ( .A1(n11839), .A2(n15839), .ZN(n10138) );
  INV_X1 U11306 ( .A(n17098), .ZN(n17103) );
  NAND2_X1 U11307 ( .A1(n10648), .A2(n10647), .ZN(n10974) );
  AND2_X1 U11308 ( .A1(n11587), .A2(n11586), .ZN(n11682) );
  OR2_X1 U11309 ( .A1(n15249), .A2(n12139), .ZN(n11848) );
  NAND2_X1 U11310 ( .A1(n15153), .A2(n9882), .ZN(n16270) );
  AND2_X1 U11311 ( .A1(n9884), .A2(n9883), .ZN(n15153) );
  OR2_X1 U11312 ( .A1(n15218), .A2(n11847), .ZN(n15249) );
  NAND2_X1 U11313 ( .A1(n12679), .A2(n17865), .ZN(n17777) );
  AND2_X1 U11314 ( .A1(n12508), .A2(n12507), .ZN(n17757) );
  CLKBUF_X1 U11315 ( .A(n13017), .Z(n13048) );
  AND2_X1 U11316 ( .A1(n15279), .A2(n11763), .ZN(n11827) );
  INV_X1 U11317 ( .A(n17881), .ZN(n17808) );
  OAI21_X2 U11318 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18929), .A(n16669), 
        .ZN(n17968) );
  AOI21_X1 U11319 ( .B1(n11851), .B2(n10164), .A(n11841), .ZN(n11846) );
  INV_X2 U11320 ( .A(n9739), .ZN(n9740) );
  OR2_X1 U11321 ( .A1(n11840), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10164) );
  NAND2_X1 U11322 ( .A1(n9844), .A2(n11466), .ZN(n19605) );
  OR2_X1 U11323 ( .A1(n11487), .A2(n11482), .ZN(n11612) );
  OR2_X1 U11324 ( .A1(n11487), .A2(n11488), .ZN(n19425) );
  NAND2_X1 U11325 ( .A1(n9844), .A2(n10133), .ZN(n19627) );
  OR2_X1 U11326 ( .A1(n11489), .A2(n11482), .ZN(n11615) );
  OR2_X1 U11327 ( .A1(n11478), .A2(n11486), .ZN(n19399) );
  NAND2_X1 U11328 ( .A1(n11456), .A2(n19295), .ZN(n11487) );
  NAND2_X1 U11329 ( .A1(n9839), .A2(n12987), .ZN(n12991) );
  OR2_X1 U11330 ( .A1(n11478), .A2(n11482), .ZN(n13931) );
  OR2_X1 U11331 ( .A1(n11489), .A2(n11486), .ZN(n11608) );
  OR2_X1 U11332 ( .A1(n11478), .A2(n11488), .ZN(n19300) );
  BUF_X1 U11333 ( .A(n12982), .Z(n13049) );
  NAND2_X1 U11334 ( .A1(n11851), .A2(n11817), .ZN(n11812) );
  OR2_X1 U11335 ( .A1(n12982), .A2(n19295), .ZN(n11478) );
  OR2_X1 U11336 ( .A1(n12937), .A2(n12936), .ZN(n12938) );
  INV_X2 U11337 ( .A(n16074), .ZN(n13387) );
  NAND2_X2 U11338 ( .A1(n14661), .A2(n13065), .ZN(n14712) );
  OR2_X1 U11339 ( .A1(n11800), .A2(n10022), .ZN(n11817) );
  BUF_X2 U11340 ( .A(n12930), .Z(n19295) );
  INV_X2 U11341 ( .A(n13179), .ZN(n13252) );
  NAND2_X1 U11342 ( .A1(n20245), .A2(n9734), .ZN(n20180) );
  NOR2_X2 U11343 ( .A1(n19943), .A2(n19340), .ZN(n19759) );
  NOR2_X1 U11344 ( .A1(n19259), .A2(n19269), .ZN(n12970) );
  NOR2_X1 U11345 ( .A1(n20906), .A2(n17250), .ZN(n17237) );
  INV_X2 U11346 ( .A(n19164), .ZN(n19161) );
  NAND2_X1 U11347 ( .A1(n10041), .A2(n10505), .ZN(n9920) );
  INV_X1 U11348 ( .A(n9745), .ZN(n9746) );
  AND2_X1 U11349 ( .A1(n11438), .A2(n11437), .ZN(n11448) );
  NAND2_X1 U11350 ( .A1(n11453), .A2(n11452), .ZN(n11458) );
  AND2_X1 U11351 ( .A1(n10482), .A2(n10480), .ZN(n10531) );
  OR2_X1 U11352 ( .A1(n11435), .A2(n11436), .ZN(n11438) );
  AND2_X1 U11353 ( .A1(n11775), .A2(n21042), .ZN(n11778) );
  NAND2_X1 U11354 ( .A1(n11442), .A2(n11441), .ZN(n11986) );
  NAND2_X1 U11355 ( .A1(n10437), .A2(n10436), .ZN(n10439) );
  CLKBUF_X1 U11356 ( .A(n17581), .Z(n17599) );
  NAND2_X1 U11357 ( .A1(n17919), .A2(n12494), .ZN(n12497) );
  AND2_X1 U11358 ( .A1(n11756), .A2(n10005), .ZN(n11771) );
  NAND2_X1 U11359 ( .A1(n11756), .A2(n10006), .ZN(n11851) );
  INV_X1 U11360 ( .A(n10032), .ZN(n12121) );
  AOI21_X1 U11361 ( .B1(n11400), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n11399), .ZN(n11423) );
  NOR2_X1 U11362 ( .A1(n11430), .A2(n11429), .ZN(n11431) );
  AND2_X1 U11363 ( .A1(n11687), .A2(n11688), .ZN(n11701) );
  OAI211_X1 U11364 ( .C1(n11401), .C2(n19839), .A(n11398), .B(n11397), .ZN(
        n11399) );
  NOR2_X1 U11365 ( .A1(n11695), .A2(n11694), .ZN(n11687) );
  AND2_X1 U11366 ( .A1(n10525), .A2(n10524), .ZN(n10526) );
  AND2_X1 U11367 ( .A1(n11395), .A2(n11937), .ZN(n13349) );
  NOR2_X1 U11368 ( .A1(n11139), .A2(n10446), .ZN(n10427) );
  CLKBUF_X1 U11369 ( .A(n10365), .Z(n9729) );
  INV_X1 U11370 ( .A(n14049), .ZN(n13062) );
  CLKBUF_X1 U11371 ( .A(n10364), .Z(n10331) );
  AND2_X1 U11372 ( .A1(n11167), .A2(n10420), .ZN(n11139) );
  AND2_X1 U11373 ( .A1(n11392), .A2(n12365), .ZN(n9973) );
  AOI21_X1 U11374 ( .B1(n10505), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10043), 
        .ZN(n10042) );
  AND2_X1 U11376 ( .A1(n13579), .A2(n11233), .ZN(n12873) );
  AND2_X2 U11377 ( .A1(n11381), .A2(n11305), .ZN(n11370) );
  AND2_X1 U11378 ( .A1(n11278), .A2(n11689), .ZN(n11306) );
  AND2_X1 U11379 ( .A1(n19319), .A2(n11380), .ZN(n12365) );
  AND2_X1 U11380 ( .A1(n12553), .A2(n9932), .ZN(n18932) );
  OR2_X1 U11381 ( .A1(n11585), .A2(n11584), .ZN(n11674) );
  OR2_X1 U11382 ( .A1(n11601), .A2(n11600), .ZN(n11955) );
  OR2_X1 U11384 ( .A1(n10000), .A2(n11548), .ZN(n9999) );
  OR2_X1 U11385 ( .A1(n10518), .A2(n10517), .ZN(n10989) );
  NOR2_X1 U11386 ( .A1(n9934), .A2(n9933), .ZN(n9932) );
  NAND2_X2 U11387 ( .A1(n10447), .A2(n20157), .ZN(n11246) );
  AOI211_X1 U11388 ( .C1(n17288), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n12552), .B(n12551), .ZN(n12553) );
  OR2_X1 U11389 ( .A1(n12544), .A2(n12545), .ZN(n17554) );
  NAND2_X1 U11390 ( .A1(n11292), .A2(n11291), .ZN(n12954) );
  AND2_X2 U11391 ( .A1(n20135), .A2(n10447), .ZN(n13587) );
  NAND2_X2 U11392 ( .A1(n11321), .A2(n11320), .ZN(n12350) );
  NAND2_X1 U11393 ( .A1(n11362), .A2(n11361), .ZN(n11380) );
  NAND2_X1 U11394 ( .A1(n11304), .A2(n11303), .ZN(n11308) );
  OR2_X1 U11395 ( .A1(n10492), .A2(n10491), .ZN(n11044) );
  OR2_X1 U11396 ( .A1(n10502), .A2(n10501), .ZN(n10990) );
  NAND2_X1 U11397 ( .A1(n11265), .A2(n9865), .ZN(n11379) );
  AND4_X1 U11398 ( .A1(n11653), .A2(n11652), .A3(n11651), .A4(n11650), .ZN(
        n11654) );
  NAND2_X1 U11399 ( .A1(n11284), .A2(n11283), .ZN(n11292) );
  NAND2_X1 U11400 ( .A1(n11319), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11320) );
  INV_X1 U11401 ( .A(n12555), .ZN(n9933) );
  NAND2_X1 U11402 ( .A1(n11360), .A2(n20841), .ZN(n11361) );
  NAND2_X1 U11403 ( .A1(n11314), .A2(n20841), .ZN(n11321) );
  OAI21_X1 U11404 ( .B1(n9864), .B2(n9863), .A(n20841), .ZN(n9865) );
  BUF_X2 U11405 ( .A(n10322), .Z(n10806) );
  INV_X2 U11406 ( .A(n20820), .ZN(n13442) );
  NOR2_X2 U11407 ( .A1(n20130), .A2(n20129), .ZN(n20131) );
  AND2_X1 U11408 ( .A1(n10324), .A2(n10323), .ZN(n10325) );
  AND4_X1 U11409 ( .A1(n10319), .A2(n10318), .A3(n10317), .A4(n10316), .ZN(
        n10165) );
  AND4_X1 U11410 ( .A1(n10177), .A2(n10176), .A3(n10175), .A4(n10174), .ZN(
        n10187) );
  AND4_X1 U11411 ( .A1(n10410), .A2(n10409), .A3(n10408), .A4(n10407), .ZN(
        n10411) );
  AND4_X1 U11412 ( .A1(n10406), .A2(n10405), .A3(n10404), .A4(n10403), .ZN(
        n10412) );
  AND4_X1 U11413 ( .A1(n10402), .A2(n10401), .A3(n10400), .A4(n10399), .ZN(
        n10413) );
  AND4_X1 U11414 ( .A1(n10396), .A2(n10395), .A3(n10394), .A4(n10393), .ZN(
        n10414) );
  AND4_X1 U11415 ( .A1(n10382), .A2(n10381), .A3(n10380), .A4(n10379), .ZN(
        n10383) );
  AND4_X1 U11416 ( .A1(n10378), .A2(n10377), .A3(n10376), .A4(n10375), .ZN(
        n10384) );
  AND4_X1 U11417 ( .A1(n10374), .A2(n10373), .A3(n10372), .A4(n10371), .ZN(
        n10385) );
  AND4_X1 U11418 ( .A1(n10293), .A2(n10292), .A3(n10291), .A4(n10290), .ZN(
        n10299) );
  AND4_X1 U11419 ( .A1(n10289), .A2(n10288), .A3(n10287), .A4(n10286), .ZN(
        n10300) );
  AND4_X1 U11420 ( .A1(n10285), .A2(n10284), .A3(n10283), .A4(n10282), .ZN(
        n10301) );
  INV_X2 U11421 ( .A(n16656), .ZN(U215) );
  AND2_X1 U11422 ( .A1(n11282), .A2(n11281), .ZN(n11283) );
  AND3_X1 U11423 ( .A1(n11280), .A2(n20841), .A3(n11279), .ZN(n11284) );
  AND4_X1 U11424 ( .A1(n11359), .A2(n11358), .A3(n11357), .A4(n11356), .ZN(
        n11360) );
  NAND2_X2 U11425 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19960), .ZN(n19875) );
  NAND2_X2 U11426 ( .A1(n19960), .A2(n19838), .ZN(n19876) );
  INV_X2 U11427 ( .A(n19276), .ZN(n9725) );
  NOR2_X1 U11428 ( .A1(n18893), .A2(n18804), .ZN(n20824) );
  BUF_X2 U11429 ( .A(n10302), .Z(n10811) );
  BUF_X2 U11430 ( .A(n10314), .Z(n10891) );
  BUF_X2 U11431 ( .A(n10199), .Z(n10876) );
  OR2_X2 U11432 ( .A1(n11129), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16200) );
  INV_X2 U11433 ( .A(n16658), .ZN(n16660) );
  NOR2_X2 U11434 ( .A1(n18298), .A2(n18356), .ZN(n18664) );
  NOR2_X2 U11435 ( .A1(n18356), .A2(n18377), .ZN(n18434) );
  NOR2_X2 U11436 ( .A1(n18755), .A2(n18377), .ZN(n18396) );
  BUF_X2 U11437 ( .A(n10356), .Z(n10899) );
  OR2_X1 U11438 ( .A1(n12402), .A2(n12406), .ZN(n14035) );
  OR2_X1 U11439 ( .A1(n12407), .A2(n12406), .ZN(n13859) );
  CLKBUF_X2 U11440 ( .A(n11334), .Z(n11354) );
  CLKBUF_X1 U11441 ( .A(n10869), .Z(n10893) );
  CLKBUF_X1 U11442 ( .A(n13384), .Z(n19117) );
  NAND2_X1 U11443 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18908), .ZN(
        n12403) );
  AND2_X2 U11444 ( .A1(n11257), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11509) );
  NAND2_X1 U11445 ( .A1(n18900), .A2(n20949), .ZN(n12407) );
  NAND2_X1 U11446 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20949), .ZN(
        n12402) );
  AND2_X1 U11447 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9845) );
  INV_X1 U11448 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11257) );
  NOR2_X2 U11449 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10181) );
  NOR2_X1 U11450 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11258) );
  NOR2_X1 U11451 ( .A1(n13411), .A2(n13412), .ZN(n9727) );
  INV_X1 U11452 ( .A(n10537), .ZN(n9728) );
  OR2_X1 U11453 ( .A1(n14419), .A2(n14421), .ZN(n9730) );
  NAND2_X1 U11454 ( .A1(n9730), .A2(n14420), .ZN(n14757) );
  NOR2_X1 U11455 ( .A1(n13411), .A2(n13412), .ZN(n13413) );
  XNOR2_X1 U11456 ( .A(n13819), .B(n10721), .ZN(n13952) );
  NAND2_X1 U11457 ( .A1(n10534), .A2(n10533), .ZN(n9731) );
  NAND2_X1 U11458 ( .A1(n10534), .A2(n10533), .ZN(n10546) );
  AOI22_X2 U11459 ( .A1(n16332), .A2(n19285), .B1(n19288), .B2(n16331), .ZN(
        n16333) );
  AOI21_X2 U11460 ( .B1(n15614), .B2(n15611), .A(n15570), .ZN(n15603) );
  NAND2_X1 U11461 ( .A1(n12095), .A2(n9720), .ZN(n12304) );
  AND2_X1 U11463 ( .A1(n10165), .A2(n10328), .ZN(n9733) );
  AND2_X1 U11464 ( .A1(n10165), .A2(n10328), .ZN(n10449) );
  XNOR2_X1 U11465 ( .A(n13476), .B(n20285), .ZN(n20406) );
  NOR2_X2 U11466 ( .A1(n13619), .A2(n19143), .ZN(n13620) );
  NAND2_X1 U11467 ( .A1(n10482), .A2(n10480), .ZN(n9734) );
  AND2_X1 U11468 ( .A1(n11426), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11400) );
  AND2_X2 U11469 ( .A1(n13256), .A2(n13258), .ZN(n9735) );
  NAND2_X1 U11470 ( .A1(n10442), .A2(n10441), .ZN(n9736) );
  NAND2_X1 U11471 ( .A1(n10442), .A2(n10441), .ZN(n10482) );
  AND2_X4 U11472 ( .A1(n11464), .A2(n11458), .ZN(n12816) );
  NAND2_X1 U11473 ( .A1(n10050), .A2(n10049), .ZN(n14716) );
  INV_X1 U11474 ( .A(n14508), .ZN(n9737) );
  INV_X1 U11476 ( .A(n14508), .ZN(n10096) );
  INV_X1 U11478 ( .A(n19113), .ZN(n9739) );
  OAI22_X1 U11479 ( .A1(n16510), .A2(n13629), .B1(n15488), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n19113) );
  OAI21_X2 U11480 ( .B1(n15401), .B2(n14283), .A(n15396), .ZN(n14344) );
  NOR2_X2 U11481 ( .A1(n15400), .A2(n15402), .ZN(n15401) );
  OAI22_X1 U11482 ( .A1(n13181), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n10979), 
        .B2(n10561), .ZN(n10479) );
  NAND2_X1 U11483 ( .A1(n10048), .A2(n13476), .ZN(n13181) );
  INV_X4 U11484 ( .A(n10423), .ZN(n10387) );
  NAND3_X4 U11485 ( .A1(n10187), .A2(n10186), .A3(n10185), .ZN(n10389) );
  NAND2_X1 U11487 ( .A1(n9734), .A2(n10459), .ZN(n10045) );
  NAND2_X2 U11488 ( .A1(n10434), .A2(n10433), .ZN(n10463) );
  OAI21_X2 U11489 ( .B1(n10438), .B2(n10428), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10434) );
  AND2_X2 U11490 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10179) );
  OAI21_X2 U11491 ( .B1(n10977), .B2(n10104), .A(n10544), .ZN(n10545) );
  AOI21_X1 U11492 ( .B1(n11136), .B2(n11135), .A(n14066), .ZN(n14729) );
  AND2_X2 U11493 ( .A1(n10545), .A2(n10556), .ZN(n9822) );
  NOR2_X2 U11494 ( .A1(n14344), .A2(n14345), .ZN(n14343) );
  NAND2_X2 U11495 ( .A1(n13133), .A2(n10556), .ZN(n13256) );
  AND2_X1 U11496 ( .A1(n14265), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9741) );
  INV_X2 U11497 ( .A(n10388), .ZN(n11149) );
  AND2_X2 U11498 ( .A1(n13457), .A2(n13188), .ZN(n10397) );
  NAND2_X1 U11499 ( .A1(n20180), .A2(n10529), .ZN(n13582) );
  OR2_X1 U11501 ( .A1(n10422), .A2(n11246), .ZN(n13160) );
  NAND2_X2 U11502 ( .A1(n11162), .A2(n11246), .ZN(n11167) );
  AND2_X4 U11503 ( .A1(n10178), .A2(n13457), .ZN(n10353) );
  AND2_X2 U11504 ( .A1(n10180), .A2(n13457), .ZN(n10868) );
  AND2_X2 U11505 ( .A1(n13457), .A2(n13473), .ZN(n10314) );
  AND2_X1 U11506 ( .A1(n13188), .A2(n10179), .ZN(n9743) );
  AND2_X1 U11507 ( .A1(n13188), .A2(n10179), .ZN(n9744) );
  AND2_X1 U11508 ( .A1(n13188), .A2(n10179), .ZN(n10321) );
  AND2_X4 U11509 ( .A1(n13458), .A2(n13188), .ZN(n10352) );
  AND2_X4 U11510 ( .A1(n10094), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13458) );
  XNOR2_X2 U11511 ( .A(n10584), .B(n15066), .ZN(n10999) );
  NAND2_X2 U11512 ( .A1(n10537), .A2(n10536), .ZN(n10584) );
  NAND2_X2 U11513 ( .A1(n14629), .A2(n10752), .ZN(n14557) );
  NAND2_X2 U11514 ( .A1(n14524), .A2(n14525), .ZN(n14508) );
  NOR2_X4 U11515 ( .A1(n14557), .A2(n10105), .ZN(n14524) );
  INV_X1 U11516 ( .A(n18737), .ZN(n9745) );
  NOR2_X4 U11517 ( .A1(n14409), .A2(n14410), .ZN(n14393) );
  XNOR2_X2 U11518 ( .A(n14065), .B(n14066), .ZN(n10972) );
  NAND2_X1 U11519 ( .A1(n12472), .A2(n12653), .ZN(n12500) );
  NAND2_X1 U11520 ( .A1(n9740), .A2(n15155), .ZN(n9882) );
  AND2_X1 U11521 ( .A1(n13272), .A2(n11515), .ZN(n14155) );
  NAND2_X1 U11522 ( .A1(n10597), .A2(n9873), .ZN(n10645) );
  NOR2_X1 U11523 ( .A1(n10619), .A2(n9874), .ZN(n9873) );
  AND2_X1 U11524 ( .A1(n11396), .A2(n12365), .ZN(n11415) );
  NAND2_X1 U11525 ( .A1(n11665), .A2(n11664), .ZN(n11673) );
  INV_X1 U11526 ( .A(n11662), .ZN(n11665) );
  NAND2_X1 U11527 ( .A1(n12632), .A2(n12631), .ZN(n9938) );
  INV_X1 U11528 ( .A(n14068), .ZN(n10886) );
  OR3_X1 U11529 ( .A1(n9947), .A2(n9814), .A3(n9946), .ZN(n9945) );
  INV_X1 U11530 ( .A(n14395), .ZN(n9946) );
  OR2_X1 U11531 ( .A1(n11799), .A2(n11821), .ZN(n10024) );
  NOR2_X1 U11532 ( .A1(n10011), .A2(n11761), .ZN(n10010) );
  INV_X1 U11533 ( .A(n11755), .ZN(n10011) );
  NAND2_X1 U11534 ( .A1(n11264), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11265) );
  NAND2_X1 U11535 ( .A1(n11857), .A2(n11851), .ZN(n15093) );
  NAND2_X1 U11536 ( .A1(n15704), .A2(n9823), .ZN(n10140) );
  NAND2_X1 U11537 ( .A1(n9985), .A2(n15754), .ZN(n9984) );
  NAND2_X1 U11538 ( .A1(n9986), .A2(n15574), .ZN(n9985) );
  INV_X1 U11539 ( .A(n9987), .ZN(n9986) );
  INV_X1 U11540 ( .A(n13692), .ZN(n11962) );
  NOR2_X1 U11541 ( .A1(n17040), .A2(n12407), .ZN(n14030) );
  AND2_X1 U11542 ( .A1(n10074), .A2(n10071), .ZN(n10070) );
  AND2_X1 U11543 ( .A1(n10073), .A2(n10072), .ZN(n10071) );
  NAND2_X1 U11544 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10074) );
  AOI22_X1 U11545 ( .A1(n12479), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12418), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10073) );
  NAND2_X1 U11546 ( .A1(n17756), .A2(n17868), .ZN(n12510) );
  NAND2_X1 U11547 ( .A1(n17883), .A2(n12503), .ZN(n12506) );
  NOR2_X1 U11548 ( .A1(n10389), .A2(n20811), .ZN(n14068) );
  AND2_X1 U11549 ( .A1(n20811), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14067) );
  NAND2_X1 U11550 ( .A1(n11812), .A2(n10020), .ZN(n11811) );
  OR2_X1 U11551 ( .A1(n10024), .A2(n9818), .ZN(n10023) );
  NAND2_X1 U11552 ( .A1(n11851), .A2(n11792), .ZN(n11791) );
  BUF_X1 U11553 ( .A(n11443), .Z(n15101) );
  AND4_X1 U11554 ( .A1(n11649), .A2(n11648), .A3(n11647), .A4(n11646), .ZN(
        n11655) );
  OR2_X1 U11555 ( .A1(n15208), .A2(n15192), .ZN(n10160) );
  OAI21_X1 U11556 ( .B1(n15595), .B2(n15572), .A(n15594), .ZN(n16338) );
  NAND2_X1 U11557 ( .A1(n11897), .A2(n11896), .ZN(n13330) );
  OR2_X1 U11558 ( .A1(n19567), .A2(n19925), .ZN(n19683) );
  OAI21_X1 U11559 ( .B1(n16722), .B2(n9970), .A(n9968), .ZN(n16711) );
  NAND2_X1 U11560 ( .A1(n16933), .A2(n9969), .ZN(n9968) );
  OR2_X1 U11561 ( .A1(n17610), .A2(n16713), .ZN(n9970) );
  INV_X1 U11562 ( .A(n16713), .ZN(n9969) );
  BUF_X1 U11563 ( .A(n14030), .Z(n15950) );
  OAI21_X1 U11564 ( .B1(n16281), .B2(n19085), .A(n9879), .ZN(n9878) );
  AOI21_X1 U11565 ( .B1(n15483), .B2(n19125), .A(n9880), .ZN(n9879) );
  AND2_X1 U11566 ( .A1(n9717), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9880) );
  NAND2_X1 U11567 ( .A1(n9740), .A2(n15532), .ZN(n9883) );
  NAND2_X1 U11568 ( .A1(n9846), .A2(n11376), .ZN(n11405) );
  INV_X1 U11569 ( .A(n12343), .ZN(n9846) );
  NAND2_X1 U11570 ( .A1(n9850), .A2(n12356), .ZN(n11410) );
  NOR2_X1 U11571 ( .A1(n11895), .A2(n14263), .ZN(n11396) );
  INV_X1 U11572 ( .A(n11427), .ZN(n11430) );
  NAND2_X1 U11573 ( .A1(n9853), .A2(n9851), .ZN(n11409) );
  NAND2_X1 U11574 ( .A1(n12367), .A2(n9852), .ZN(n9851) );
  NAND2_X1 U11575 ( .A1(n12348), .A2(n12350), .ZN(n9853) );
  OR2_X1 U11576 ( .A1(n11881), .A2(n11880), .ZN(n11882) );
  NAND2_X1 U11577 ( .A1(n10597), .A2(n10598), .ZN(n10620) );
  INV_X1 U11578 ( .A(n10505), .ZN(n10044) );
  INV_X1 U11579 ( .A(n10551), .ZN(n10043) );
  AND2_X2 U11580 ( .A1(n10173), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10178) );
  OR2_X1 U11581 ( .A1(n11639), .A2(n11638), .ZN(n11680) );
  NOR2_X1 U11582 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14129) );
  AND2_X1 U11583 ( .A1(n11882), .A2(n11660), .ZN(n11662) );
  INV_X1 U11584 ( .A(n12584), .ZN(n9931) );
  NAND2_X1 U11585 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n9930) );
  NAND2_X1 U11586 ( .A1(n13143), .A2(n10331), .ZN(n10454) );
  NOR2_X1 U11587 ( .A1(n11136), .A2(n10112), .ZN(n10111) );
  INV_X1 U11588 ( .A(n14394), .ZN(n10112) );
  INV_X1 U11589 ( .A(n14488), .ZN(n10099) );
  INV_X1 U11590 ( .A(n10968), .ZN(n10956) );
  NAND2_X1 U11591 ( .A1(n15076), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10968) );
  NAND2_X1 U11592 ( .A1(n9809), .A2(n10770), .ZN(n10108) );
  INV_X1 U11593 ( .A(n13787), .ZN(n10095) );
  INV_X1 U11594 ( .A(n10886), .ZN(n10965) );
  XNOR2_X1 U11595 ( .A(n10974), .B(n10651), .ZN(n11032) );
  OR2_X1 U11596 ( .A1(n14517), .A2(n9943), .ZN(n9942) );
  OR2_X1 U11597 ( .A1(n13587), .A2(n11194), .ZN(n11196) );
  NAND2_X1 U11598 ( .A1(n14058), .A2(n13587), .ZN(n11243) );
  OAI21_X2 U11599 ( .B1(n13582), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10532), 
        .ZN(n10988) );
  OAI211_X1 U11600 ( .C1(n20144), .C2(n11129), .A(n10465), .B(n10464), .ZN(
        n10466) );
  NAND2_X1 U11601 ( .A1(n10313), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10370) );
  NAND2_X1 U11602 ( .A1(n10302), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10368) );
  NAND4_X2 U11603 ( .A1(n10301), .A2(n10300), .A3(n10299), .A4(n10298), .ZN(
        n10391) );
  NAND3_X1 U11604 ( .A1(n20161), .A2(n20135), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11109) );
  NAND2_X1 U11605 ( .A1(n10430), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10562) );
  CLKBUF_X1 U11606 ( .A(n11144), .Z(n11145) );
  NOR2_X1 U11607 ( .A1(n11808), .A2(n10021), .ZN(n10020) );
  INV_X1 U11608 ( .A(n11756), .ZN(n10009) );
  NAND2_X1 U11609 ( .A1(n13635), .A2(n11667), .ZN(n9998) );
  AND3_X1 U11610 ( .A1(n11689), .A2(n14263), .A3(n12957), .ZN(n12088) );
  INV_X1 U11611 ( .A(n11499), .ZN(n14128) );
  NAND2_X1 U11612 ( .A1(n9842), .A2(n10151), .ZN(n14217) );
  NAND2_X1 U11613 ( .A1(n9820), .A2(n15419), .ZN(n10151) );
  INV_X1 U11614 ( .A(n15241), .ZN(n10034) );
  OR2_X1 U11615 ( .A1(n11371), .A2(n12359), .ZN(n12352) );
  INV_X1 U11616 ( .A(n12367), .ZN(n12355) );
  NOR2_X1 U11617 ( .A1(n13726), .A2(n15289), .ZN(n15288) );
  NAND2_X1 U11618 ( .A1(n10119), .A2(n13223), .ZN(n10118) );
  INV_X1 U11619 ( .A(n10120), .ZN(n10119) );
  INV_X1 U11620 ( .A(n13630), .ZN(n9898) );
  NAND2_X1 U11621 ( .A1(n15158), .A2(n15388), .ZN(n10127) );
  NOR2_X1 U11622 ( .A1(n10013), .A2(n10016), .ZN(n10012) );
  INV_X1 U11623 ( .A(n11871), .ZN(n10016) );
  INV_X1 U11624 ( .A(n10014), .ZN(n10013) );
  AND2_X1 U11625 ( .A1(n10132), .A2(n10131), .ZN(n10130) );
  AND2_X1 U11626 ( .A1(n15762), .A2(n15270), .ZN(n10132) );
  INV_X1 U11627 ( .A(n15336), .ZN(n10028) );
  AOI21_X1 U11628 ( .B1(n12140), .B2(n12141), .A(n10031), .ZN(n10030) );
  INV_X1 U11629 ( .A(n16477), .ZN(n10031) );
  NAND2_X1 U11630 ( .A1(n11972), .A2(n11971), .ZN(n11976) );
  INV_X1 U11631 ( .A(n11970), .ZN(n11972) );
  NOR2_X1 U11632 ( .A1(n11752), .A2(n11751), .ZN(n12135) );
  NAND2_X1 U11633 ( .A1(n13517), .A2(n13516), .ZN(n10090) );
  NAND2_X1 U11634 ( .A1(n11454), .A2(n11425), .ZN(n11449) );
  NAND2_X1 U11635 ( .A1(n14161), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11508) );
  NOR2_X1 U11636 ( .A1(n17040), .A2(n12402), .ZN(n12479) );
  NOR2_X1 U11637 ( .A1(n17039), .A2(n12404), .ZN(n12405) );
  NOR2_X1 U11638 ( .A1(n17040), .A2(n12397), .ZN(n12556) );
  OAI21_X1 U11639 ( .B1(n15974), .B2(n18733), .A(n17552), .ZN(n15965) );
  INV_X1 U11640 ( .A(n12515), .ZN(n10079) );
  NOR2_X1 U11641 ( .A1(n10084), .A2(n17613), .ZN(n10081) );
  AND2_X1 U11642 ( .A1(n18101), .A2(n12505), .ZN(n10077) );
  NAND2_X1 U11643 ( .A1(n17898), .A2(n12499), .ZN(n12501) );
  NOR2_X1 U11644 ( .A1(n18322), .A2(n12647), .ZN(n15987) );
  XNOR2_X1 U11645 ( .A(n17479), .B(n12477), .ZN(n12478) );
  INV_X1 U11646 ( .A(n9938), .ZN(n12645) );
  NOR3_X1 U11647 ( .A1(n18326), .A2(n17347), .A3(n12637), .ZN(n13825) );
  NAND2_X1 U11648 ( .A1(n18322), .A2(n12646), .ZN(n12622) );
  INV_X1 U11649 ( .A(n11144), .ZN(n9871) );
  AND2_X1 U11650 ( .A1(n14585), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13597) );
  AND4_X1 U11651 ( .A1(n13071), .A2(n13210), .A3(n13072), .A4(n16055), .ZN(
        n13073) );
  INV_X1 U11652 ( .A(n10945), .ZN(n10952) );
  OR2_X1 U11653 ( .A1(n10943), .A2(n10942), .ZN(n10945) );
  NAND2_X1 U11654 ( .A1(n10925), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10935) );
  OR2_X1 U11655 ( .A1(n10910), .A2(n10909), .ZN(n10918) );
  OAI211_X1 U11656 ( .C1(n10886), .C2(n10644), .A(n10643), .B(n10642), .ZN(
        n13506) );
  NAND2_X1 U11657 ( .A1(n10605), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10623) );
  AND3_X1 U11658 ( .A1(n13144), .A2(n11074), .A3(n16055), .ZN(n16037) );
  NAND2_X1 U11660 ( .A1(n9944), .A2(n14057), .ZN(n14356) );
  INV_X1 U11661 ( .A(n14714), .ZN(n10054) );
  NAND2_X1 U11662 ( .A1(n14714), .A2(n10055), .ZN(n10050) );
  NOR3_X1 U11663 ( .A1(n14463), .A2(n9947), .A3(n9814), .ZN(n14408) );
  OR2_X1 U11664 ( .A1(n9770), .A2(n14465), .ZN(n14463) );
  NAND2_X1 U11665 ( .A1(n14616), .A2(n11212), .ZN(n14619) );
  NAND2_X1 U11666 ( .A1(n13719), .A2(n9917), .ZN(n11048) );
  INV_X1 U11667 ( .A(n11042), .ZN(n9918) );
  INV_X1 U11668 ( .A(n10162), .ZN(n9919) );
  INV_X1 U11669 ( .A(n13587), .ZN(n14358) );
  AND2_X1 U11670 ( .A1(n13154), .A2(n13210), .ZN(n13169) );
  NOR2_X1 U11671 ( .A1(n20286), .A2(n20291), .ZN(n20469) );
  NOR2_X1 U11672 ( .A1(n20292), .A2(n20291), .ZN(n20611) );
  NAND2_X1 U11673 ( .A1(n20815), .A2(n20134), .ZN(n20291) );
  INV_X1 U11674 ( .A(n12947), .ZN(n13321) );
  OR2_X1 U11675 ( .A1(n10023), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10022) );
  NOR2_X1 U11676 ( .A1(n11800), .A2(n10024), .ZN(n11819) );
  NAND2_X1 U11677 ( .A1(n11782), .A2(n11781), .ZN(n11792) );
  NOR2_X1 U11678 ( .A1(n10008), .A2(n19325), .ZN(n10006) );
  INV_X1 U11679 ( .A(n10008), .ZN(n10005) );
  INV_X1 U11680 ( .A(n14153), .ZN(n12292) );
  NAND2_X1 U11681 ( .A1(n13026), .A2(n9805), .ZN(n10148) );
  OR2_X1 U11682 ( .A1(n12158), .A2(n12157), .ZN(n13023) );
  AND2_X1 U11683 ( .A1(n12992), .A2(n15351), .ZN(n13015) );
  INV_X1 U11684 ( .A(n11451), .ZN(n11452) );
  NAND2_X1 U11685 ( .A1(n15413), .A2(n15415), .ZN(n15414) );
  AND2_X1 U11686 ( .A1(n14258), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n15351) );
  OR2_X1 U11687 ( .A1(n12949), .A2(n16516), .ZN(n12752) );
  NOR2_X1 U11688 ( .A1(n15866), .A2(n13376), .ZN(n15826) );
  AOI21_X1 U11689 ( .B1(n15557), .B2(n15558), .A(n11850), .ZN(n15704) );
  INV_X1 U11690 ( .A(n9984), .ZN(n9979) );
  NOR2_X1 U11691 ( .A1(n9984), .A2(n9982), .ZN(n9981) );
  INV_X1 U11692 ( .A(n15571), .ZN(n9982) );
  NAND2_X1 U11693 ( .A1(n15595), .A2(n15594), .ZN(n9983) );
  AOI21_X1 U11694 ( .B1(n15572), .B2(n15594), .A(n9988), .ZN(n9987) );
  INV_X1 U11695 ( .A(n15573), .ZN(n9988) );
  OR2_X1 U11696 ( .A1(n15844), .A2(n15834), .ZN(n15789) );
  OAI21_X1 U11697 ( .B1(n15880), .B2(n15883), .A(n11789), .ZN(n15870) );
  NAND2_X1 U11698 ( .A1(n9993), .A2(n9990), .ZN(n15880) );
  AND2_X1 U11699 ( .A1(n9991), .A2(n16374), .ZN(n9990) );
  AND2_X1 U11700 ( .A1(n11773), .A2(n9992), .ZN(n9991) );
  INV_X1 U11701 ( .A(n15898), .ZN(n9992) );
  OAI211_X1 U11702 ( .C1(n11967), .C2(n11965), .A(n11964), .B(n11963), .ZN(
        n13765) );
  NAND2_X1 U11703 ( .A1(n11962), .A2(n11965), .ZN(n11963) );
  NOR2_X2 U11704 ( .A1(n13527), .A2(n13528), .ZN(n13694) );
  NAND2_X1 U11705 ( .A1(n12817), .A2(n19757), .ZN(n12986) );
  AND2_X1 U11706 ( .A1(n14130), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13272) );
  INV_X1 U11707 ( .A(n11482), .ZN(n11466) );
  NAND2_X1 U11708 ( .A1(n19210), .A2(n19917), .ZN(n19888) );
  OR2_X1 U11709 ( .A1(n19567), .A2(n13708), .ZN(n19713) );
  NAND2_X1 U11710 ( .A1(n19907), .A2(n19917), .ZN(n19712) );
  NAND2_X1 U11711 ( .A1(n12876), .A2(n12875), .ZN(n19765) );
  NAND2_X1 U11712 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19765), .ZN(n19340) );
  NAND2_X1 U11713 ( .A1(n18932), .A2(n17554), .ZN(n12627) );
  AOI21_X1 U11714 ( .B1(n12642), .B2(n12644), .A(n12641), .ZN(n18772) );
  OAI21_X1 U11715 ( .B1(n16767), .B2(n9967), .A(n9965), .ZN(n16755) );
  OR2_X1 U11716 ( .A1(n17660), .A2(n17677), .ZN(n9967) );
  NAND2_X1 U11717 ( .A1(n16933), .A2(n9966), .ZN(n9965) );
  INV_X1 U11718 ( .A(n17660), .ZN(n9966) );
  NOR2_X1 U11719 ( .A1(n16767), .A2(n17677), .ZN(n16766) );
  INV_X1 U11720 ( .A(n17721), .ZN(n9963) );
  NAND2_X1 U11721 ( .A1(n17190), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10068) );
  NAND2_X1 U11722 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10069) );
  NAND2_X1 U11723 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10067) );
  NAND2_X1 U11724 ( .A1(n15950), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10064) );
  NAND2_X1 U11725 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10065) );
  NAND2_X1 U11726 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10063) );
  AND3_X1 U11727 ( .A1(n18772), .A2(n18927), .A3(n15965), .ZN(n16079) );
  INV_X1 U11728 ( .A(n18932), .ZN(n17494) );
  NOR2_X1 U11729 ( .A1(n17762), .A2(n12680), .ZN(n17666) );
  INV_X1 U11730 ( .A(n16560), .ZN(n10082) );
  NOR2_X1 U11731 ( .A1(n17761), .A2(n10153), .ZN(n12508) );
  XNOR2_X1 U11732 ( .A(n12501), .B(n10058), .ZN(n17884) );
  INV_X1 U11733 ( .A(n12502), .ZN(n10058) );
  XNOR2_X1 U11734 ( .A(n17491), .B(n10060), .ZN(n17958) );
  AND2_X1 U11735 ( .A1(n11152), .A2(n13210), .ZN(n16118) );
  NOR2_X1 U11737 ( .A1(n12752), .A2(n13321), .ZN(n19953) );
  NAND2_X1 U11738 ( .A1(n15185), .A2(n15543), .ZN(n9885) );
  INV_X1 U11739 ( .A(n19165), .ZN(n19151) );
  AND2_X1 U11740 ( .A1(n19205), .A2(n12958), .ZN(n19172) );
  OAI21_X1 U11741 ( .B1(n12084), .B2(n12083), .A(n9768), .ZN(n15497) );
  OR2_X1 U11742 ( .A1(n15156), .A2(n15388), .ZN(n15389) );
  OAI21_X1 U11743 ( .B1(n19291), .B2(n16343), .A(n16342), .ZN(n9859) );
  INV_X1 U11744 ( .A(n16417), .ZN(n19291) );
  INV_X1 U11745 ( .A(n16421), .ZN(n19285) );
  XNOR2_X1 U11746 ( .A(n9768), .B(n15102), .ZN(n16281) );
  NAND2_X1 U11747 ( .A1(n9752), .A2(n10091), .ZN(n15499) );
  OAI21_X1 U11748 ( .B1(n15551), .B2(n10092), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10091) );
  XNOR2_X1 U11749 ( .A(n16338), .B(n9801), .ZN(n16438) );
  NAND2_X1 U11750 ( .A1(n9855), .A2(n9854), .ZN(n16437) );
  NAND2_X1 U11751 ( .A1(n15590), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9854) );
  NAND2_X1 U11752 ( .A1(n16339), .A2(n9856), .ZN(n9855) );
  NOR2_X1 U11753 ( .A1(n16340), .A2(n21013), .ZN(n9856) );
  AND2_X1 U11754 ( .A1(n12372), .A2(n19937), .ZN(n16485) );
  INV_X1 U11755 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19931) );
  OR2_X1 U11756 ( .A1(n12829), .A2(n12821), .ZN(n19925) );
  OAI21_X1 U11757 ( .B1(n12990), .B2(n13048), .A(n15350), .ZN(n19567) );
  INV_X1 U11758 ( .A(n19818), .ZN(n19792) );
  NOR2_X1 U11759 ( .A1(n16721), .A2(n16933), .ZN(n16712) );
  NAND2_X1 U11760 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17053), .ZN(n17035) );
  INV_X1 U11761 ( .A(n17045), .ZN(n17053) );
  INV_X1 U11762 ( .A(n17392), .ZN(n18332) );
  AOI21_X1 U11763 ( .B1(n17351), .B2(n9925), .A(n9924), .ZN(n9923) );
  INV_X1 U11764 ( .A(P3_EAX_REG_31__SCAN_IN), .ZN(n9924) );
  OR2_X1 U11765 ( .A1(n17427), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n9925) );
  NOR2_X1 U11766 ( .A1(n17383), .A2(n19337), .ZN(n9922) );
  NAND2_X1 U11767 ( .A1(n17352), .A2(n17471), .ZN(n17351) );
  INV_X1 U11768 ( .A(n17358), .ZN(n17353) );
  NAND2_X1 U11769 ( .A1(n17393), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n17388) );
  INV_X1 U11770 ( .A(n17453), .ZN(n17344) );
  NOR2_X1 U11771 ( .A1(n18332), .A2(n17486), .ZN(n17478) );
  AND2_X1 U11772 ( .A1(n18265), .A2(n18044), .ZN(n18092) );
  NOR2_X1 U11773 ( .A1(n9779), .A2(n10003), .ZN(n10002) );
  NAND2_X1 U11774 ( .A1(n11538), .A2(n10004), .ZN(n10003) );
  NAND2_X1 U11775 ( .A1(n11571), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10004) );
  NAND2_X1 U11776 ( .A1(n12262), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10001) );
  AND2_X1 U11777 ( .A1(n11386), .A2(n14263), .ZN(n11347) );
  AOI22_X1 U11778 ( .A1(n11353), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14127), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11301) );
  NAND2_X1 U11779 ( .A1(n11673), .A2(n11672), .ZN(n11675) );
  XNOR2_X1 U11780 ( .A(n20841), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11676) );
  OR2_X1 U11781 ( .A1(n12529), .A2(n12530), .ZN(n12525) );
  INV_X1 U11782 ( .A(n11090), .ZN(n11087) );
  AND2_X1 U11783 ( .A1(n10425), .A2(n10389), .ZN(n10443) );
  OR2_X1 U11784 ( .A1(n10618), .A2(n10617), .ZN(n11018) );
  OR2_X1 U11785 ( .A1(n10594), .A2(n10593), .ZN(n11015) );
  OR2_X1 U11786 ( .A1(n10476), .A2(n10475), .ZN(n10980) );
  NAND2_X1 U11787 ( .A1(n10527), .A2(n10526), .ZN(n10535) );
  OR2_X1 U11788 ( .A1(n10422), .A2(n10387), .ZN(n10346) );
  NAND2_X1 U11789 ( .A1(n10438), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10458) );
  INV_X1 U11790 ( .A(n14172), .ZN(n10150) );
  AOI22_X1 U11791 ( .A1(n11498), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n11514), .ZN(n9868) );
  NAND2_X1 U11792 ( .A1(n14127), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n9867) );
  NAND2_X1 U11793 ( .A1(n13775), .A2(n12140), .ZN(n10029) );
  NAND2_X1 U11794 ( .A1(n11432), .A2(n11431), .ZN(n11435) );
  NAND2_X1 U11795 ( .A1(n12012), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n11397) );
  INV_X1 U11796 ( .A(n9999), .ZN(n12117) );
  AOI21_X1 U11797 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19903), .A(
        n11678), .ZN(n11878) );
  NOR2_X1 U11798 ( .A1(n11677), .A2(n11676), .ZN(n11678) );
  INV_X1 U11799 ( .A(n11675), .ZN(n11677) );
  AND2_X1 U11800 ( .A1(n11911), .A2(n11379), .ZN(n11309) );
  NAND2_X1 U11801 ( .A1(n11484), .A2(n11474), .ZN(n11616) );
  AOI22_X1 U11802 ( .A1(n11514), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11334), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11285) );
  NAND2_X1 U11803 ( .A1(n12439), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10072) );
  NOR2_X1 U11804 ( .A1(n17464), .A2(n12474), .ZN(n12472) );
  AOI21_X1 U11805 ( .B1(n18754), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12524), .ZN(n12530) );
  AND2_X1 U11806 ( .A1(n12640), .A2(n12639), .ZN(n12524) );
  OAI22_X1 U11807 ( .A1(n18900), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n21008), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12529) );
  NAND2_X1 U11808 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12404) );
  NOR2_X1 U11809 ( .A1(n12634), .A2(n12618), .ZN(n12646) );
  NOR2_X1 U11810 ( .A1(n21125), .A2(n20161), .ZN(n10392) );
  NOR2_X1 U11811 ( .A1(n9796), .A2(n10098), .ZN(n10097) );
  INV_X1 U11812 ( .A(n14476), .ZN(n10098) );
  OR2_X1 U11813 ( .A1(n9948), .A2(n14451), .ZN(n9947) );
  INV_X1 U11814 ( .A(n10646), .ZN(n10647) );
  INV_X1 U11815 ( .A(n10645), .ZN(n10648) );
  NAND2_X1 U11816 ( .A1(n10040), .A2(n10998), .ZN(n11004) );
  NAND2_X1 U11817 ( .A1(n13567), .A2(n13566), .ZN(n10040) );
  NOR2_X1 U11818 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11153), .ZN(
        n9911) );
  NAND2_X1 U11819 ( .A1(n13140), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9914) );
  NAND2_X1 U11820 ( .A1(n10995), .A2(n9907), .ZN(n9913) );
  NAND2_X1 U11821 ( .A1(n11157), .A2(n11156), .ZN(n11160) );
  AOI22_X1 U11822 ( .A1(n10322), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9744), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10357) );
  NAND2_X1 U11823 ( .A1(n10353), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10354) );
  AOI22_X1 U11824 ( .A1(n10352), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10322), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10309) );
  AOI22_X1 U11825 ( .A1(n10353), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10352), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U11826 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10673), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10175) );
  INV_X1 U11827 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20541) );
  NAND2_X1 U11828 ( .A1(n20406), .A2(n20815), .ZN(n10574) );
  INV_X1 U11829 ( .A(n13483), .ZN(n20134) );
  AOI21_X1 U11830 ( .B1(n20814), .B2(n13490), .A(n13482), .ZN(n13483) );
  OR2_X1 U11831 ( .A1(n20161), .A2(n20815), .ZN(n10561) );
  INV_X1 U11832 ( .A(n11109), .ZN(n11115) );
  OR2_X1 U11833 ( .A1(n13472), .A2(n13471), .ZN(n16034) );
  NOR2_X1 U11834 ( .A1(n11860), .A2(n10015), .ZN(n10014) );
  NOR2_X1 U11835 ( .A1(n10019), .A2(n11805), .ZN(n10018) );
  INV_X1 U11836 ( .A(n10020), .ZN(n10019) );
  AND2_X1 U11837 ( .A1(n11812), .A2(n10018), .ZN(n11807) );
  NAND2_X1 U11838 ( .A1(n10010), .A2(n11768), .ZN(n10008) );
  NAND2_X1 U11839 ( .A1(n10121), .A2(n16377), .ZN(n10120) );
  INV_X1 U11840 ( .A(n13028), .ZN(n10121) );
  INV_X1 U11841 ( .A(n14155), .ZN(n14099) );
  INV_X1 U11842 ( .A(n14161), .ZN(n14095) );
  NAND2_X1 U11843 ( .A1(n11400), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10146) );
  CLKBUF_X1 U11844 ( .A(n11500), .Z(n14307) );
  CLKBUF_X1 U11845 ( .A(n11353), .Z(n14326) );
  NAND2_X1 U11846 ( .A1(n10026), .A2(n15160), .ZN(n10025) );
  INV_X1 U11847 ( .A(n15172), .ZN(n10026) );
  INV_X1 U11848 ( .A(n15229), .ZN(n10033) );
  NAND2_X1 U11849 ( .A1(n15463), .A2(n15464), .ZN(n9843) );
  INV_X1 U11850 ( .A(n13743), .ZN(n10147) );
  AND2_X1 U11851 ( .A1(n12827), .A2(n19944), .ZN(n14258) );
  NAND2_X1 U11852 ( .A1(n12982), .A2(n12981), .ZN(n9839) );
  NAND2_X1 U11853 ( .A1(n12359), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11895) );
  NAND2_X1 U11854 ( .A1(n15129), .A2(n9886), .ZN(n9889) );
  NOR2_X1 U11855 ( .A1(n15559), .A2(n9887), .ZN(n9886) );
  INV_X1 U11856 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n9887) );
  NAND2_X1 U11857 ( .A1(n15123), .A2(n9894), .ZN(n9897) );
  NOR2_X1 U11858 ( .A1(n15109), .A2(n9895), .ZN(n9894) );
  INV_X1 U11859 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n9895) );
  NAND2_X1 U11860 ( .A1(n15117), .A2(n9890), .ZN(n9893) );
  NOR2_X1 U11861 ( .A1(n16370), .A2(n9891), .ZN(n9890) );
  INV_X1 U11862 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n9891) );
  NOR2_X1 U11863 ( .A1(n15537), .A2(n10141), .ZN(n10139) );
  NAND2_X1 U11864 ( .A1(n10143), .A2(n10142), .ZN(n10141) );
  NAND2_X1 U11865 ( .A1(n10144), .A2(n15705), .ZN(n10142) );
  AND2_X1 U11866 ( .A1(n10036), .A2(n13959), .ZN(n10035) );
  INV_X1 U11867 ( .A(n15304), .ZN(n10122) );
  AND2_X1 U11868 ( .A1(n10038), .A2(n10037), .ZN(n10036) );
  INV_X1 U11869 ( .A(n15299), .ZN(n10037) );
  AND2_X1 U11870 ( .A1(n9829), .A2(n15823), .ZN(n10038) );
  INV_X1 U11871 ( .A(n9862), .ZN(n9861) );
  OAI21_X1 U11872 ( .B1(n11968), .B2(n9774), .A(n11974), .ZN(n9862) );
  OR2_X1 U11873 ( .A1(n11976), .A2(n12139), .ZN(n11975) );
  AND2_X1 U11874 ( .A1(n11754), .A2(n11753), .ZN(n11971) );
  AOI21_X1 U11875 ( .B1(n11443), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n11447), .ZN(n11985) );
  NOR2_X1 U11876 ( .A1(n12359), .A2(n12350), .ZN(n11387) );
  NOR2_X1 U11877 ( .A1(n11535), .A2(n11534), .ZN(n12112) );
  OR2_X1 U11878 ( .A1(n14236), .A2(n12828), .ZN(n12926) );
  NAND2_X1 U11879 ( .A1(n12935), .A2(n12934), .ZN(n12937) );
  INV_X1 U11880 ( .A(n14156), .ZN(n14101) );
  NAND2_X1 U11881 ( .A1(n9972), .A2(n11912), .ZN(n11385) );
  NAND2_X1 U11882 ( .A1(n9975), .A2(n12088), .ZN(n9972) );
  AND2_X1 U11883 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14130) );
  AND4_X1 U11884 ( .A1(n19319), .A2(n11367), .A3(n11366), .A4(n11379), .ZN(
        n11368) );
  INV_X1 U11885 ( .A(n11486), .ZN(n10133) );
  OR2_X1 U11886 ( .A1(n15917), .A2(n12816), .ZN(n11488) );
  AND2_X1 U11887 ( .A1(n11891), .A2(n11890), .ZN(n11899) );
  AND2_X1 U11888 ( .A1(n11666), .A2(n11673), .ZN(n11900) );
  AND2_X1 U11889 ( .A1(n13285), .A2(n13284), .ZN(n13319) );
  NOR2_X1 U11890 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18914), .ZN(
        n12639) );
  INV_X1 U11891 ( .A(n17039), .ZN(n10057) );
  INV_X1 U11892 ( .A(n12397), .ZN(n10056) );
  NAND2_X1 U11893 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18914), .ZN(
        n12406) );
  NAND2_X1 U11894 ( .A1(n12721), .A2(n9760), .ZN(n16536) );
  OR2_X1 U11895 ( .A1(n12404), .A2(n12403), .ZN(n9769) );
  NOR2_X1 U11896 ( .A1(n17040), .A2(n12404), .ZN(n12418) );
  NOR2_X1 U11897 ( .A1(n9938), .A2(n9936), .ZN(n12638) );
  INV_X1 U11898 ( .A(n9937), .ZN(n9936) );
  AOI21_X1 U11899 ( .B1(n12634), .B2(n12635), .A(n15967), .ZN(n9937) );
  INV_X1 U11900 ( .A(n12554), .ZN(n9934) );
  NAND2_X1 U11901 ( .A1(n9777), .A2(n9753), .ZN(n12647) );
  NOR2_X1 U11902 ( .A1(n13183), .A2(n13141), .ZN(n13190) );
  NAND2_X1 U11903 ( .A1(n10788), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10785) );
  INV_X1 U11904 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14538) );
  OR2_X1 U11905 ( .A1(n20817), .A2(n13574), .ZN(n14585) );
  AND4_X1 U11906 ( .A1(n10452), .A2(n10451), .A3(n10450), .A4(n13159), .ZN(
        n10453) );
  OAI21_X1 U11907 ( .B1(n9731), .B2(n10104), .A(n10103), .ZN(n13064) );
  AOI21_X1 U11908 ( .B1(n10102), .B2(n10797), .A(n10550), .ZN(n10103) );
  INV_X1 U11909 ( .A(n10547), .ZN(n10102) );
  OAI21_X1 U11910 ( .B1(n13074), .B2(n13583), .A(n13409), .ZN(n13096) );
  INV_X2 U11911 ( .A(n10447), .ZN(n13165) );
  NOR2_X1 U11912 ( .A1(n10110), .A2(n10114), .ZN(n10109) );
  INV_X1 U11913 ( .A(n10111), .ZN(n10110) );
  INV_X1 U11914 ( .A(n14065), .ZN(n10114) );
  AOI22_X1 U11915 ( .A1(n14733), .A2(n10960), .B1(n10959), .B2(n10958), .ZN(
        n14394) );
  OR2_X1 U11916 ( .A1(n10935), .A2(n14756), .ZN(n10943) );
  OAI21_X1 U11917 ( .B1(n14748), .B2(n10971), .A(n10951), .ZN(n14410) );
  AOI22_X1 U11918 ( .A1(n14760), .A2(n10960), .B1(n10941), .B2(n10940), .ZN(
        n14421) );
  NOR2_X1 U11919 ( .A1(n10918), .A2(n14773), .ZN(n10925) );
  OAI21_X1 U11920 ( .B1(n14769), .B2(n10971), .A(n10934), .ZN(n14437) );
  CLKBUF_X1 U11921 ( .A(n14435), .Z(n14436) );
  OAI21_X1 U11922 ( .B1(n14787), .B2(n10971), .A(n10917), .ZN(n14462) );
  CLKBUF_X1 U11923 ( .A(n14460), .Z(n14461) );
  OAI21_X1 U11924 ( .B1(n14805), .B2(n10971), .A(n10887), .ZN(n14488) );
  AND2_X1 U11925 ( .A1(n14497), .A2(n10101), .ZN(n10100) );
  INV_X1 U11926 ( .A(n14509), .ZN(n10101) );
  NOR2_X1 U11927 ( .A1(n10820), .A2(n10167), .ZN(n10834) );
  NAND2_X1 U11928 ( .A1(n10834), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10848) );
  NAND2_X1 U11929 ( .A1(n10805), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10820) );
  NOR2_X1 U11930 ( .A1(n10785), .A2(n14538), .ZN(n10805) );
  NAND2_X1 U11931 ( .A1(n10106), .A2(n14611), .ZN(n10105) );
  INV_X1 U11932 ( .A(n10108), .ZN(n10106) );
  OR2_X1 U11933 ( .A1(n10724), .A2(n16091), .ZN(n10753) );
  NOR2_X1 U11934 ( .A1(n20875), .A2(n10753), .ZN(n10788) );
  INV_X1 U11935 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n20875) );
  NOR2_X1 U11936 ( .A1(n10684), .A2(n13795), .ZN(n10689) );
  NAND2_X1 U11937 ( .A1(n10668), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10684) );
  AND3_X1 U11938 ( .A1(n10688), .A2(n10687), .A3(n10686), .ZN(n13787) );
  CLKBUF_X1 U11939 ( .A(n13605), .Z(n13606) );
  AND2_X1 U11940 ( .A1(n10640), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10652) );
  NOR2_X1 U11941 ( .A1(n10623), .A2(n10626), .ZN(n10640) );
  INV_X1 U11942 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10626) );
  AOI21_X1 U11943 ( .B1(n11007), .B2(n10797), .A(n10607), .ZN(n13449) );
  NAND2_X1 U11944 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10576) );
  AND2_X1 U11945 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n10166), .ZN(
        n10605) );
  INV_X1 U11946 ( .A(n10576), .ZN(n10166) );
  NOR2_X1 U11947 ( .A1(n14463), .A2(n9947), .ZN(n14434) );
  INV_X1 U11948 ( .A(n14765), .ZN(n14784) );
  OR3_X1 U11949 ( .A1(n9942), .A2(n14489), .A3(n14477), .ZN(n9941) );
  NAND2_X1 U11950 ( .A1(n11064), .A2(n9916), .ZN(n9915) );
  AND2_X1 U11951 ( .A1(n14821), .A2(n9834), .ZN(n9916) );
  NOR2_X1 U11952 ( .A1(n14528), .A2(n14517), .ZN(n14519) );
  OR2_X1 U11953 ( .A1(n14619), .A2(n14526), .ZN(n14528) );
  AND2_X1 U11954 ( .A1(n11209), .A2(n11208), .ZN(n14614) );
  AND2_X1 U11955 ( .A1(n14563), .A2(n11204), .ZN(n14616) );
  NAND2_X1 U11956 ( .A1(n9951), .A2(n9804), .ZN(n14633) );
  NOR2_X1 U11957 ( .A1(n14633), .A2(n14562), .ZN(n14563) );
  INV_X1 U11958 ( .A(n9776), .ZN(n16148) );
  NOR2_X1 U11959 ( .A1(n13811), .A2(n13790), .ZN(n13927) );
  NAND2_X1 U11960 ( .A1(n13610), .A2(n13609), .ZN(n13813) );
  AND3_X1 U11961 ( .A1(n11183), .A2(n11196), .A3(n11182), .ZN(n13814) );
  NAND2_X1 U11962 ( .A1(n9940), .A2(n9939), .ZN(n13811) );
  INV_X1 U11963 ( .A(n13814), .ZN(n9939) );
  INV_X1 U11964 ( .A(n13813), .ZN(n9940) );
  NOR2_X1 U11965 ( .A1(n10996), .A2(n20113), .ZN(n16209) );
  AND2_X1 U11966 ( .A1(n13511), .A2(n13510), .ZN(n13610) );
  NOR2_X1 U11967 ( .A1(n13453), .A2(n13415), .ZN(n13511) );
  NAND2_X1 U11968 ( .A1(n13260), .A2(n9949), .ZN(n13453) );
  NOR2_X1 U11969 ( .A1(n9950), .A2(n13450), .ZN(n9949) );
  INV_X1 U11970 ( .A(n13259), .ZN(n9950) );
  AND2_X1 U11971 ( .A1(n13135), .A2(n13134), .ZN(n13260) );
  NAND2_X1 U11972 ( .A1(n13260), .A2(n13259), .ZN(n13451) );
  AND2_X1 U11973 ( .A1(n13169), .A2(n13164), .ZN(n15035) );
  NAND2_X1 U11974 ( .A1(n10529), .A2(n10046), .ZN(n10048) );
  NOR2_X1 U11975 ( .A1(n10466), .A2(n10047), .ZN(n10046) );
  CLKBUF_X1 U11976 ( .A(n13473), .Z(n13474) );
  CLKBUF_X1 U11977 ( .A(n12858), .Z(n12859) );
  INV_X1 U11978 ( .A(n19964), .ZN(n13210) );
  AND4_X1 U11979 ( .A1(n10370), .A2(n10369), .A3(n10368), .A4(n10367), .ZN(
        n10386) );
  AND3_X1 U11980 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20815), .A3(n20134), 
        .ZN(n20172) );
  INV_X1 U11981 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21022) );
  NOR2_X1 U11982 ( .A1(n11109), .A2(n11075), .ZN(n11111) );
  NAND2_X1 U11983 ( .A1(n10562), .A2(n10561), .ZN(n11089) );
  OR2_X1 U11984 ( .A1(n11113), .A2(n11082), .ZN(n11083) );
  XNOR2_X1 U11985 ( .A(n15094), .B(n11873), .ZN(n11874) );
  NAND2_X1 U11986 ( .A1(n15107), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15105) );
  AND2_X1 U11987 ( .A1(n15134), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15107) );
  OR2_X1 U11988 ( .A1(n11800), .A2(n11799), .ZN(n11823) );
  NOR2_X1 U11989 ( .A1(n10009), .A2(n10007), .ZN(n11769) );
  INV_X1 U11990 ( .A(n10010), .ZN(n10007) );
  OR2_X1 U11991 ( .A1(n9900), .A2(n9899), .ZN(n13912) );
  NAND2_X1 U11992 ( .A1(n11756), .A2(n11755), .ZN(n11762) );
  NAND2_X1 U11993 ( .A1(n11929), .A2(n9720), .ZN(n11669) );
  NAND2_X1 U11994 ( .A1(n13374), .A2(n13373), .ZN(n13619) );
  NOR2_X1 U11995 ( .A1(n15331), .A2(n10120), .ZN(n16379) );
  NOR2_X1 U11996 ( .A1(n15171), .A2(n15172), .ZN(n15174) );
  NAND2_X1 U11997 ( .A1(n15259), .A2(n9817), .ZN(n15243) );
  CLKBUF_X1 U11998 ( .A(n15425), .Z(n15426) );
  CLKBUF_X1 U11999 ( .A(n13997), .Z(n13760) );
  CLKBUF_X1 U12000 ( .A(n15824), .Z(n15852) );
  AND2_X1 U12001 ( .A1(n12236), .A2(n12235), .ZN(n15868) );
  CLKBUF_X1 U12002 ( .A(n15902), .Z(n16454) );
  INV_X1 U12003 ( .A(n12365), .ZN(n12353) );
  INV_X1 U12004 ( .A(n12711), .ZN(n13961) );
  NOR2_X1 U12005 ( .A1(n15105), .A2(n16272), .ZN(n15103) );
  AND2_X1 U12006 ( .A1(n15132), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15134) );
  NOR2_X1 U12007 ( .A1(n15130), .A2(n15210), .ZN(n15132) );
  OR2_X1 U12008 ( .A1(n9889), .A2(n9888), .ZN(n15130) );
  NAND2_X1 U12009 ( .A1(n9751), .A2(n9806), .ZN(n15239) );
  INV_X1 U12010 ( .A(n15237), .ZN(n10129) );
  NOR2_X1 U12011 ( .A1(n15239), .A2(n15226), .ZN(n15228) );
  NAND2_X1 U12012 ( .A1(n15129), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15128) );
  NOR2_X1 U12013 ( .A1(n15577), .A2(n15126), .ZN(n15129) );
  NAND2_X1 U12014 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n15127), .ZN(
        n15126) );
  AND2_X1 U12015 ( .A1(n9751), .A2(n15762), .ZN(n15764) );
  OR2_X1 U12016 ( .A1(n9897), .A2(n9896), .ZN(n15124) );
  INV_X1 U12017 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9896) );
  NOR2_X1 U12018 ( .A1(n15124), .A2(n18993), .ZN(n15127) );
  NOR2_X1 U12019 ( .A1(n15616), .A2(n15120), .ZN(n15123) );
  NAND2_X1 U12020 ( .A1(n15123), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15122) );
  NAND2_X1 U12021 ( .A1(n15826), .A2(n15827), .ZN(n15829) );
  NAND2_X1 U12022 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n15121), .ZN(
        n15120) );
  NOR2_X1 U12023 ( .A1(n15118), .A2(n16354), .ZN(n15121) );
  OR2_X1 U12024 ( .A1(n9893), .A2(n9892), .ZN(n15118) );
  NOR2_X1 U12025 ( .A1(n10118), .A2(n10117), .ZN(n10116) );
  INV_X1 U12026 ( .A(n15864), .ZN(n10117) );
  NOR2_X1 U12027 ( .A1(n15331), .A2(n10118), .ZN(n15865) );
  NAND2_X1 U12028 ( .A1(n15117), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15116) );
  NOR2_X1 U12029 ( .A1(n16392), .A2(n15114), .ZN(n15117) );
  NOR2_X1 U12030 ( .A1(n13913), .A2(n13912), .ZN(n15115) );
  NAND2_X1 U12031 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n15115), .ZN(
        n15114) );
  NOR2_X1 U12032 ( .A1(n13630), .A2(n16429), .ZN(n15113) );
  NAND2_X1 U12033 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13630) );
  NAND2_X1 U12034 ( .A1(n10126), .A2(n10125), .ZN(n10124) );
  INV_X1 U12035 ( .A(n15170), .ZN(n10126) );
  NOR2_X1 U12036 ( .A1(n10127), .A2(n12082), .ZN(n10125) );
  NOR2_X1 U12037 ( .A1(n9803), .A2(n15479), .ZN(n15480) );
  OR2_X1 U12038 ( .A1(n10093), .A2(n12380), .ZN(n10092) );
  NOR2_X1 U12039 ( .A1(n15515), .A2(n15514), .ZN(n15516) );
  NAND2_X1 U12040 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10093) );
  NOR2_X1 U12041 ( .A1(n15551), .A2(n15538), .ZN(n15540) );
  NAND2_X1 U12042 ( .A1(n10137), .A2(n15729), .ZN(n10134) );
  INV_X1 U12043 ( .A(n11838), .ZN(n10137) );
  NAND2_X1 U12044 ( .A1(n9751), .A2(n10130), .ZN(n15257) );
  NAND2_X1 U12046 ( .A1(n15826), .A2(n9759), .ZN(n15305) );
  AND2_X1 U12047 ( .A1(n15826), .A2(n9800), .ZN(n15303) );
  NAND2_X1 U12048 ( .A1(n12284), .A2(n10038), .ZN(n16443) );
  OR3_X1 U12049 ( .A1(n11830), .A2(n12139), .A3(n16446), .ZN(n15611) );
  NAND2_X1 U12050 ( .A1(n9977), .A2(n9765), .ZN(n15844) );
  INV_X1 U12051 ( .A(n15886), .ZN(n9976) );
  NAND2_X1 U12052 ( .A1(n9977), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15886) );
  AND2_X1 U12053 ( .A1(n12388), .A2(n12387), .ZN(n15818) );
  AND2_X1 U12054 ( .A1(n12163), .A2(n12162), .ZN(n15336) );
  NAND2_X1 U12055 ( .A1(n10089), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10088) );
  INV_X1 U12056 ( .A(n13517), .ZN(n10089) );
  NOR2_X1 U12057 ( .A1(n11522), .A2(n11521), .ZN(n12880) );
  AOI21_X1 U12058 ( .B1(n15917), .B2(n12981), .A(n12826), .ZN(n12830) );
  XNOR2_X1 U12059 ( .A(n12121), .B(n12120), .ZN(n12891) );
  CLKBUF_X1 U12060 ( .A(n13016), .Z(n12990) );
  NAND2_X1 U12061 ( .A1(n13048), .A2(n12990), .ZN(n15350) );
  AND3_X1 U12062 ( .A1(n19425), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19428), 
        .ZN(n19433) );
  AND2_X1 U12063 ( .A1(n19532), .A2(n19890), .ZN(n19541) );
  INV_X1 U12064 ( .A(n12358), .ZN(n13939) );
  CLKBUF_X1 U12065 ( .A(n12954), .Z(n12955) );
  INV_X1 U12066 ( .A(n19334), .ZN(n19336) );
  INV_X1 U12067 ( .A(n19335), .ZN(n19338) );
  INV_X1 U12068 ( .A(n19765), .ZN(n19343) );
  NOR2_X1 U12069 ( .A1(n13962), .A2(n13674), .ZN(n19335) );
  NOR2_X1 U12070 ( .A1(n16755), .A2(n16933), .ZN(n16745) );
  NOR2_X1 U12071 ( .A1(n16781), .A2(n17693), .ZN(n16780) );
  NAND2_X1 U12072 ( .A1(n9960), .A2(n9959), .ZN(n9962) );
  NOR2_X1 U12073 ( .A1(n17873), .A2(n9954), .ZN(n9953) );
  NOR2_X1 U12074 ( .A1(n17501), .A2(n17503), .ZN(n9927) );
  AOI221_X1 U12075 ( .B1(n18933), .B2(n18784), .C1(n17552), .C2(n18784), .A(
        n17551), .ZN(n17553) );
  AND2_X1 U12076 ( .A1(n12721), .A2(n9825), .ZN(n16535) );
  NOR2_X1 U12077 ( .A1(n17655), .A2(n17656), .ZN(n12721) );
  NAND2_X1 U12078 ( .A1(n17751), .A2(n9797), .ZN(n17694) );
  NOR2_X1 U12079 ( .A1(n17731), .A2(n9958), .ZN(n9957) );
  NOR2_X1 U12080 ( .A1(n12724), .A2(n17765), .ZN(n17751) );
  NOR2_X1 U12081 ( .A1(n17801), .A2(n17803), .ZN(n17789) );
  NOR2_X1 U12082 ( .A1(n16906), .A2(n16917), .ZN(n17829) );
  NAND2_X1 U12083 ( .A1(n9833), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17827) );
  NOR2_X1 U12084 ( .A1(n17873), .A2(n17886), .ZN(n17869) );
  NOR2_X1 U12085 ( .A1(n17901), .A2(n17905), .ZN(n17871) );
  NOR2_X1 U12086 ( .A1(n18778), .A2(n18792), .ZN(n12682) );
  OAI211_X1 U12087 ( .C1(n16565), .C2(n10080), .A(n17795), .B(n10078), .ZN(
        n10086) );
  INV_X1 U12088 ( .A(n10081), .ZN(n10080) );
  NAND2_X1 U12089 ( .A1(n10079), .A2(n10081), .ZN(n10078) );
  NAND2_X1 U12090 ( .A1(n17640), .A2(n10059), .ZN(n12514) );
  AND2_X1 U12091 ( .A1(n17651), .A2(n9802), .ZN(n10059) );
  NAND2_X1 U12092 ( .A1(n18305), .A2(n18229), .ZN(n18029) );
  AND2_X1 U12093 ( .A1(n12510), .A2(n9787), .ZN(n17668) );
  NAND2_X1 U12094 ( .A1(n17668), .A2(n18018), .ZN(n17667) );
  NOR2_X1 U12095 ( .A1(n20842), .A2(n17686), .ZN(n17673) );
  INV_X1 U12096 ( .A(n12510), .ZN(n17715) );
  NAND2_X1 U12097 ( .A1(n17757), .A2(n20847), .ZN(n17756) );
  AOI21_X1 U12098 ( .B1(n17867), .B2(n10075), .A(n17795), .ZN(n17761) );
  AND2_X1 U12099 ( .A1(n12504), .A2(n10076), .ZN(n10075) );
  AND2_X1 U12100 ( .A1(n10159), .A2(n10077), .ZN(n10076) );
  NOR2_X1 U12101 ( .A1(n12506), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17867) );
  INV_X1 U12102 ( .A(n17777), .ZN(n18156) );
  NAND2_X1 U12103 ( .A1(n17884), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17883) );
  NAND2_X1 U12104 ( .A1(n17912), .A2(n12498), .ZN(n17899) );
  NAND2_X1 U12105 ( .A1(n17899), .A2(n17900), .ZN(n17898) );
  XNOR2_X1 U12106 ( .A(n12497), .B(n12496), .ZN(n17913) );
  INV_X1 U12107 ( .A(n12495), .ZN(n12496) );
  NOR2_X1 U12108 ( .A1(n15966), .A2(n12625), .ZN(n12715) );
  INV_X1 U12109 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18754) );
  NAND2_X1 U12110 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17040) );
  NOR2_X2 U12111 ( .A1(n18947), .A2(n13823), .ZN(n18768) );
  NAND2_X1 U12112 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18736) );
  INV_X1 U12113 ( .A(n17554), .ZN(n18305) );
  INV_X1 U12114 ( .A(n12647), .ZN(n18309) );
  NOR2_X1 U12115 ( .A1(n12576), .A2(n12575), .ZN(n18322) );
  NOR2_X1 U12116 ( .A1(n12566), .A2(n12565), .ZN(n18326) );
  OR2_X1 U12117 ( .A1(n12633), .A2(n12622), .ZN(n18784) );
  NAND2_X1 U12118 ( .A1(n14353), .A2(n14354), .ZN(n20817) );
  INV_X1 U12119 ( .A(n20041), .ZN(n20000) );
  INV_X1 U12120 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n13972) );
  INV_X1 U12121 ( .A(n19987), .ZN(n20043) );
  NOR2_X1 U12122 ( .A1(n14479), .A2(n19967), .ZN(n19987) );
  OR2_X1 U12123 ( .A1(n14590), .A2(n14362), .ZN(n20028) );
  AND2_X1 U12124 ( .A1(n14585), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20042) );
  OR2_X1 U12125 ( .A1(n14053), .A2(n20128), .ZN(n14683) );
  OR2_X1 U12126 ( .A1(n14679), .A2(n13065), .ZN(n14711) );
  NOR2_X1 U12127 ( .A1(n13096), .A2(n20820), .ZN(n16074) );
  INV_X1 U12128 ( .A(n13096), .ZN(n13445) );
  XNOR2_X1 U12129 ( .A(n13577), .B(n14369), .ZN(n14719) );
  INV_X1 U12130 ( .A(n16127), .ZN(n16151) );
  AND2_X1 U12131 ( .A1(n19970), .A2(n11127), .ZN(n16135) );
  INV_X1 U12132 ( .A(n16135), .ZN(n14818) );
  XNOR2_X1 U12133 ( .A(n14360), .B(n14359), .ZN(n14883) );
  NAND2_X1 U12134 ( .A1(n14723), .A2(n11070), .ZN(n10053) );
  AND2_X1 U12135 ( .A1(n14397), .A2(n14396), .ZN(n14941) );
  NAND2_X1 U12136 ( .A1(n9904), .A2(n9903), .ZN(n14746) );
  OR2_X1 U12137 ( .A1(n14778), .A2(n14777), .ZN(n14779) );
  NAND2_X1 U12138 ( .A1(n11048), .A2(n13802), .ZN(n13946) );
  NOR2_X1 U12139 ( .A1(n13657), .A2(n16228), .ZN(n16231) );
  INV_X1 U12140 ( .A(n15051), .ZN(n20122) );
  AND2_X1 U12141 ( .A1(n13169), .A2(n13168), .ZN(n20116) );
  NAND2_X1 U12142 ( .A1(n9731), .A2(n10547), .ZN(n20208) );
  INV_X1 U12143 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20459) );
  CLKBUF_X1 U12144 ( .A(n13181), .Z(n13182) );
  INV_X1 U12145 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20127) );
  NAND2_X1 U12146 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n16055), .ZN(n15089) );
  OAI22_X1 U12147 ( .A1(n20148), .A2(n20147), .B1(n20472), .B2(n20287), .ZN(
        n20175) );
  INV_X1 U12148 ( .A(n20374), .ZN(n20334) );
  OAI211_X1 U12149 ( .C1(n20427), .C2(n20547), .A(n20469), .B(n20411), .ZN(
        n20429) );
  INV_X1 U12150 ( .A(n20399), .ZN(n20428) );
  AND2_X1 U12151 ( .A1(n20602), .A2(n20540), .ZN(n20597) );
  OAI211_X1 U12152 ( .C1(n20642), .C2(n20612), .A(n20611), .B(n20610), .ZN(
        n20645) );
  INV_X1 U12153 ( .A(n20477), .ZN(n20668) );
  INV_X1 U12154 ( .A(n20481), .ZN(n20674) );
  INV_X1 U12155 ( .A(n20489), .ZN(n20686) );
  INV_X1 U12156 ( .A(n20493), .ZN(n20692) );
  AND2_X1 U12157 ( .A1(n20602), .A2(n20382), .ZN(n20708) );
  INV_X1 U12158 ( .A(n20501), .ZN(n20706) );
  INV_X1 U12159 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20714) );
  INV_X2 U12160 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20811) );
  NAND2_X1 U12161 ( .A1(n15218), .A2(n15223), .ZN(n15201) );
  NAND2_X1 U12162 ( .A1(n11812), .A2(n11813), .ZN(n11809) );
  OR2_X1 U12163 ( .A1(n11800), .A2(n10023), .ZN(n11815) );
  AND2_X1 U12164 ( .A1(n19272), .A2(n13642), .ZN(n19123) );
  NAND2_X1 U12165 ( .A1(n15140), .A2(n13647), .ZN(n19126) );
  AND2_X1 U12166 ( .A1(n11784), .A2(n11783), .ZN(n15323) );
  AND2_X1 U12167 ( .A1(n19953), .A2(n13636), .ZN(n19125) );
  OR2_X1 U12168 ( .A1(n19953), .A2(n13640), .ZN(n19129) );
  INV_X1 U12169 ( .A(n19123), .ZN(n19121) );
  INV_X1 U12170 ( .A(n19085), .ZN(n19133) );
  CLKBUF_X1 U12171 ( .A(n13743), .Z(n13621) );
  AND2_X1 U12172 ( .A1(n12278), .A2(n12277), .ZN(n19143) );
  CLKBUF_X1 U12173 ( .A(n13619), .Z(n13375) );
  OR2_X1 U12174 ( .A1(n12195), .A2(n12194), .ZN(n19150) );
  AND2_X1 U12175 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n13015), .ZN(
        n13020) );
  INV_X1 U12176 ( .A(n19925), .ZN(n13708) );
  AND2_X1 U12177 ( .A1(n12815), .A2(n15925), .ZN(n19164) );
  CLKBUF_X1 U12178 ( .A(n15406), .Z(n15407) );
  INV_X1 U12179 ( .A(n19180), .ZN(n19232) );
  OR2_X1 U12180 ( .A1(n12959), .A2(n19172), .ZN(n19207) );
  AND2_X1 U12181 ( .A1(n12837), .A2(n19825), .ZN(n19259) );
  INV_X1 U12182 ( .A(n19951), .ZN(n19269) );
  INV_X1 U12183 ( .A(n19261), .ZN(n19268) );
  XNOR2_X1 U12184 ( .A(n16339), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9997) );
  INV_X1 U12185 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16370) );
  INV_X1 U12186 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13913) );
  AND2_X1 U12187 ( .A1(n16428), .A2(n13779), .ZN(n16417) );
  INV_X1 U12188 ( .A(n19288), .ZN(n16418) );
  INV_X1 U12189 ( .A(n16428), .ZN(n19284) );
  NAND2_X1 U12190 ( .A1(n19168), .A2(n16493), .ZN(n15635) );
  OR2_X1 U12191 ( .A1(n16275), .A2(n16466), .ZN(n10152) );
  OR2_X1 U12192 ( .A1(n15156), .A2(n15159), .ZN(n15659) );
  NAND2_X1 U12193 ( .A1(n11798), .A2(n10138), .ZN(n10136) );
  NAND2_X1 U12194 ( .A1(n9980), .A2(n9978), .ZN(n15575) );
  NAND2_X1 U12195 ( .A1(n9979), .A2(n9807), .ZN(n9978) );
  NAND2_X1 U12196 ( .A1(n9983), .A2(n9987), .ZN(n15756) );
  CLKBUF_X1 U12197 ( .A(n15841), .Z(n15842) );
  CLKBUF_X1 U12198 ( .A(n15870), .Z(n15875) );
  AND2_X1 U12199 ( .A1(n9989), .A2(n9991), .ZN(n16372) );
  NAND2_X1 U12200 ( .A1(n9989), .A2(n11773), .ZN(n15900) );
  OAI21_X1 U12201 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15598), .A(
        n16381), .ZN(n16388) );
  INV_X1 U12202 ( .A(n15818), .ZN(n15907) );
  OAI21_X1 U12203 ( .B1(n13775), .B2(n12141), .A(n12140), .ZN(n16478) );
  NAND2_X1 U12204 ( .A1(n11969), .A2(n11968), .ZN(n13908) );
  AND2_X1 U12205 ( .A1(n12372), .A2(n12345), .ZN(n16493) );
  INV_X1 U12206 ( .A(n16493), .ZN(n16479) );
  INV_X1 U12207 ( .A(n16466), .ZN(n16494) );
  AND2_X1 U12208 ( .A1(n15793), .A2(n15798), .ZN(n16491) );
  INV_X1 U12209 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19922) );
  INV_X1 U12210 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19912) );
  INV_X1 U12211 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19903) );
  NAND2_X1 U12212 ( .A1(n12816), .A2(n12981), .ZN(n12819) );
  AND2_X1 U12213 ( .A1(n13330), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15935) );
  INV_X1 U12214 ( .A(n19915), .ZN(n19917) );
  CLKBUF_X1 U12215 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n21077) );
  INV_X1 U12216 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n20966) );
  CLKBUF_X1 U12217 ( .A(n11912), .Z(n11913) );
  NOR2_X1 U12218 ( .A1(n19458), .A2(n19888), .ZN(n19447) );
  INV_X1 U12219 ( .A(n19481), .ZN(n19482) );
  NOR2_X2 U12220 ( .A1(n19712), .A2(n19458), .ZN(n19560) );
  OAI21_X1 U12221 ( .B1(n19606), .B2(n19621), .A(n19765), .ZN(n19624) );
  INV_X1 U12222 ( .A(n19813), .ZN(n19754) );
  INV_X1 U12223 ( .A(n19731), .ZN(n19773) );
  AND2_X1 U12224 ( .A1(n19944), .A2(n19312), .ZN(n19771) );
  INV_X1 U12225 ( .A(n19653), .ZN(n19799) );
  NAND2_X1 U12226 ( .A1(n19298), .A2(n19895), .ZN(n19818) );
  AND2_X1 U12227 ( .A1(n12983), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19810) );
  NOR2_X1 U12228 ( .A1(n19713), .A2(n19712), .ZN(n19814) );
  INV_X1 U12229 ( .A(n19117), .ZN(n19090) );
  AND2_X1 U12230 ( .A1(n13351), .A2(n13350), .ZN(n16509) );
  NOR2_X1 U12231 ( .A1(n18771), .A2(n17551), .ZN(n18948) );
  NAND2_X1 U12232 ( .A1(n18930), .A2(n18772), .ZN(n17551) );
  INV_X1 U12233 ( .A(n12682), .ZN(n16669) );
  OR2_X1 U12234 ( .A1(n16711), .A2(n16933), .ZN(n16699) );
  NOR2_X1 U12235 ( .A1(n16722), .A2(n17610), .ZN(n16721) );
  NOR2_X1 U12236 ( .A1(n12733), .A2(n17639), .ZN(n16683) );
  NOR2_X1 U12237 ( .A1(n16766), .A2(n16933), .ZN(n16756) );
  AND2_X1 U12238 ( .A1(n9962), .A2(n9961), .ZN(n16790) );
  INV_X1 U12239 ( .A(n17712), .ZN(n9961) );
  INV_X1 U12240 ( .A(n9962), .ZN(n16791) );
  INV_X1 U12241 ( .A(n9964), .ZN(n16803) );
  AND2_X1 U12242 ( .A1(n9964), .A2(n9963), .ZN(n16802) );
  NOR2_X1 U12243 ( .A1(n16933), .A2(n12726), .ZN(n16814) );
  NOR2_X1 U12244 ( .A1(n16814), .A2(n17729), .ZN(n16813) );
  NOR2_X1 U12245 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16861), .ZN(n16848) );
  NOR2_X1 U12246 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16929), .ZN(n16922) );
  INV_X1 U12247 ( .A(n17031), .ZN(n17041) );
  AND2_X1 U12248 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17112), .ZN(n17107) );
  AND2_X1 U12249 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17113), .ZN(n17118) );
  NAND2_X1 U12250 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17169), .ZN(n17154) );
  NOR2_X1 U12251 ( .A1(n16823), .A2(n17170), .ZN(n17169) );
  NOR2_X1 U12252 ( .A1(n16930), .A2(n17281), .ZN(n17253) );
  INV_X1 U12253 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17307) );
  INV_X1 U12254 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17329) );
  INV_X1 U12255 ( .A(n17334), .ZN(n17337) );
  NAND2_X1 U12256 ( .A1(n17371), .A2(n9767), .ZN(n17358) );
  NAND2_X1 U12257 ( .A1(n17371), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n17367) );
  NOR2_X1 U12258 ( .A1(n17505), .A2(n17378), .ZN(n17371) );
  NOR2_X1 U12259 ( .A1(n17388), .A2(n17509), .ZN(n17345) );
  OR2_X1 U12260 ( .A1(n17507), .A2(n17377), .ZN(n17378) );
  NOR2_X1 U12261 ( .A1(n17419), .A2(n9935), .ZN(n17393) );
  NAND2_X1 U12262 ( .A1(n17423), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17419) );
  INV_X1 U12263 ( .A(n17383), .ZN(n17417) );
  NAND2_X1 U12264 ( .A1(n9929), .A2(n9747), .ZN(n17453) );
  INV_X1 U12265 ( .A(n17428), .ZN(n9928) );
  NOR2_X1 U12266 ( .A1(n12413), .A2(n12412), .ZN(n17458) );
  NOR2_X1 U12267 ( .A1(n17428), .A2(n17467), .ZN(n17463) );
  NOR2_X1 U12268 ( .A1(n12434), .A2(n12433), .ZN(n17472) );
  INV_X1 U12269 ( .A(n17478), .ZN(n17471) );
  INV_X1 U12270 ( .A(n17490), .ZN(n17480) );
  NOR2_X1 U12271 ( .A1(n10066), .A2(n10062), .ZN(n10061) );
  NOR2_X1 U12272 ( .A1(n12489), .A2(n12488), .ZN(n17967) );
  NOR3_X1 U12273 ( .A1(n16077), .A2(n17494), .A3(n17554), .ZN(n16078) );
  NOR2_X1 U12274 ( .A1(n20824), .A2(n20825), .ZN(n17512) );
  NOR2_X1 U12275 ( .A1(n17551), .A2(n17492), .ZN(n20825) );
  AOI21_X1 U12276 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17692), .A(
        n18678), .ZN(n17802) );
  AND2_X1 U12277 ( .A1(n17751), .A2(n9955), .ZN(n17676) );
  AND2_X1 U12278 ( .A1(n9797), .A2(n9956), .ZN(n9955) );
  INV_X1 U12279 ( .A(n17695), .ZN(n9956) );
  AND2_X1 U12280 ( .A1(n17751), .A2(n9957), .ZN(n17720) );
  NOR2_X1 U12281 ( .A1(n18080), .A2(n17864), .ZN(n17769) );
  INV_X1 U12282 ( .A(n17847), .ZN(n17864) );
  INV_X1 U12283 ( .A(n17861), .ZN(n17879) );
  NAND2_X1 U12284 ( .A1(n17911), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17901) );
  INV_X1 U12285 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17905) );
  NOR2_X1 U12286 ( .A1(n17926), .A2(n17928), .ZN(n17911) );
  INV_X1 U12287 ( .A(n17962), .ZN(n17952) );
  NAND2_X1 U12288 ( .A1(n17968), .A2(n17872), .ZN(n17963) );
  NAND2_X1 U12289 ( .A1(n18305), .A2(n12682), .ZN(n17972) );
  INV_X1 U12290 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18893) );
  NAND2_X1 U12291 ( .A1(n10085), .A2(n10083), .ZN(n15995) );
  AOI21_X1 U12292 ( .B1(n12715), .B2(n16010), .A(n16011), .ZN(n18737) );
  NOR2_X1 U12293 ( .A1(n18768), .A2(n18282), .ZN(n18162) );
  INV_X1 U12294 ( .A(n18162), .ZN(n18167) );
  INV_X1 U12295 ( .A(n18170), .ZN(n18184) );
  NOR2_X2 U12296 ( .A1(n18167), .A2(n9745), .ZN(n18229) );
  AOI21_X2 U12297 ( .B1(n15994), .B2(n15993), .A(n18792), .ZN(n18265) );
  INV_X1 U12298 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21008) );
  INV_X2 U12299 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18914) );
  INV_X1 U12300 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18908) );
  INV_X2 U12301 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20949) );
  NOR2_X1 U12302 ( .A1(n18301), .A2(n15973), .ZN(n18915) );
  INV_X1 U12303 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18887) );
  AOI21_X1 U12305 ( .B1(n11254), .B2(n16115), .A(n11253), .ZN(n11255) );
  NAND2_X1 U12306 ( .A1(n9881), .A2(n9876), .ZN(P2_U2824) );
  AND2_X1 U12307 ( .A1(n15142), .A2(n9877), .ZN(n9876) );
  INV_X1 U12308 ( .A(n9878), .ZN(n9877) );
  NAND2_X1 U12309 ( .A1(n15394), .A2(n9840), .ZN(P2_U2858) );
  INV_X1 U12310 ( .A(n9841), .ZN(n9840) );
  OAI21_X1 U12311 ( .B1(n16275), .B2(n19161), .A(n15393), .ZN(n9841) );
  AOI21_X1 U12312 ( .B1(n16436), .B2(n19294), .A(n9859), .ZN(n9858) );
  NAND2_X1 U12313 ( .A1(n16437), .A2(n19288), .ZN(n9860) );
  NAND2_X1 U12314 ( .A1(n16438), .A2(n19285), .ZN(n9857) );
  OAI211_X1 U12315 ( .C1(n15805), .C2(n16421), .A(n9996), .B(n9994), .ZN(
        P2_U2997) );
  NOR2_X1 U12316 ( .A1(n15600), .A2(n9995), .ZN(n9994) );
  OR2_X1 U12317 ( .A1(n9997), .A2(n16418), .ZN(n9996) );
  AND2_X1 U12318 ( .A1(n16417), .A2(n19005), .ZN(n9995) );
  NOR2_X1 U12319 ( .A1(n12393), .A2(n12392), .ZN(n12394) );
  AOI211_X1 U12320 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n16716), .A(n16715), 
        .B(n16714), .ZN(n16717) );
  NAND2_X1 U12321 ( .A1(n9926), .A2(n9921), .ZN(P3_U2704) );
  NAND2_X1 U12322 ( .A1(n17346), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n9926) );
  NOR2_X1 U12323 ( .A1(n9923), .A2(n9922), .ZN(n9921) );
  AND4_X1 U12324 ( .A1(n9928), .A2(n9831), .A3(P3_EAX_REG_2__SCAN_IN), .A4(
        P3_EAX_REG_1__SCAN_IN), .ZN(n9747) );
  NOR2_X1 U12325 ( .A1(n12403), .A2(n12397), .ZN(n12598) );
  NAND2_X1 U12326 ( .A1(n14241), .A2(n9815), .ZN(n9748) );
  AND3_X1 U12327 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9749) );
  AND2_X1 U12328 ( .A1(n9762), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9750) );
  INV_X2 U12329 ( .A(n10163), .ZN(n17274) );
  AND2_X1 U12330 ( .A1(n15288), .A2(n12049), .ZN(n9751) );
  NAND2_X1 U12331 ( .A1(n10057), .A2(n10056), .ZN(n12446) );
  NOR2_X1 U12332 ( .A1(n14508), .A2(n9796), .ZN(n14475) );
  NAND2_X1 U12333 ( .A1(n10974), .A2(n10976), .ZN(n11054) );
  AND2_X1 U12334 ( .A1(n10027), .A2(n9798), .ZN(n15335) );
  OR3_X1 U12335 ( .A1(n15551), .A2(n10092), .A3(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n9752) );
  AND4_X1 U12336 ( .A1(n12583), .A2(n12582), .A3(n12581), .A4(n12580), .ZN(
        n9753) );
  NAND2_X1 U12337 ( .A1(n15598), .A2(n9750), .ZN(n15556) );
  NAND2_X1 U12338 ( .A1(n15414), .A2(n14218), .ZN(n14241) );
  NAND2_X1 U12339 ( .A1(n11812), .A2(n9821), .ZN(n11840) );
  OR2_X1 U12340 ( .A1(n10148), .A2(n9816), .ZN(n9754) );
  AND2_X1 U12341 ( .A1(n13802), .A2(n9782), .ZN(n9755) );
  AND2_X1 U12342 ( .A1(n9748), .A2(n14260), .ZN(n9756) );
  INV_X1 U12343 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16429) );
  NAND2_X1 U12344 ( .A1(n15259), .A2(n15260), .ZN(n15240) );
  NOR2_X1 U12345 ( .A1(n15418), .A2(n15419), .ZN(n9757) );
  NOR3_X1 U12346 ( .A1(n14528), .A2(n9942), .A3(n14489), .ZN(n9758) );
  AND2_X1 U12347 ( .A1(n13605), .A2(n9799), .ZN(n13788) );
  INV_X1 U12348 ( .A(n10797), .ZN(n10104) );
  INV_X1 U12349 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17886) );
  AND2_X1 U12350 ( .A1(n10123), .A2(n15827), .ZN(n9759) );
  INV_X1 U12351 ( .A(n10598), .ZN(n9874) );
  AND2_X1 U12352 ( .A1(n14016), .A2(n9819), .ZN(n15424) );
  NAND2_X1 U12353 ( .A1(n19156), .A2(n13026), .ZN(n13219) );
  INV_X2 U12354 ( .A(n13266), .ZN(n14325) );
  AND2_X1 U12355 ( .A1(n9749), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9760) );
  AND2_X1 U12356 ( .A1(n9817), .A2(n10033), .ZN(n9761) );
  AND2_X1 U12357 ( .A1(n15767), .A2(n15769), .ZN(n9762) );
  AND2_X1 U12358 ( .A1(n9750), .A2(n15721), .ZN(n9763) );
  AND2_X1 U12359 ( .A1(n15223), .A2(n10017), .ZN(n9764) );
  AND2_X1 U12360 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15599), .ZN(
        n9765) );
  AND2_X1 U12361 ( .A1(n9764), .A2(n15189), .ZN(n9766) );
  AND2_X1 U12362 ( .A1(n9927), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n9767) );
  OR2_X1 U12363 ( .A1(n10160), .A2(n10124), .ZN(n9768) );
  OR2_X1 U12364 ( .A1(n14528), .A2(n9941), .ZN(n9770) );
  NAND2_X1 U12365 ( .A1(n10107), .A2(n10770), .ZN(n14534) );
  OR3_X1 U12366 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20949), .A3(
        n18736), .ZN(n9771) );
  NOR2_X1 U12367 ( .A1(n14508), .A2(n14509), .ZN(n14496) );
  AND2_X1 U12368 ( .A1(n14265), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13998) );
  NAND2_X1 U12369 ( .A1(n10140), .A2(n10142), .ZN(n15535) );
  AND2_X1 U12370 ( .A1(n15259), .A2(n9761), .ZN(n9773) );
  NAND2_X1 U12371 ( .A1(n11064), .A2(n14821), .ZN(n14800) );
  NAND2_X1 U12372 ( .A1(n11851), .A2(n11765), .ZN(n11775) );
  NOR2_X1 U12373 ( .A1(n14557), .A2(n10108), .ZN(n14535) );
  NAND2_X1 U12374 ( .A1(n11066), .A2(n9721), .ZN(n14752) );
  AND2_X1 U12375 ( .A1(n13906), .A2(n16482), .ZN(n9774) );
  OR2_X1 U12376 ( .A1(n15551), .A2(n10093), .ZN(n15506) );
  INV_X1 U12377 ( .A(n9944), .ZN(n14396) );
  NOR2_X1 U12378 ( .A1(n14463), .A2(n9945), .ZN(n9944) );
  NAND2_X1 U12379 ( .A1(n10136), .A2(n11838), .ZN(n15730) );
  AND2_X1 U12380 ( .A1(n14873), .A2(n11049), .ZN(n9776) );
  INV_X1 U12381 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n16510) );
  NAND2_X1 U12382 ( .A1(n12819), .A2(n12818), .ZN(n12829) );
  AND4_X1 U12383 ( .A1(n12586), .A2(n12585), .A3(n9931), .A4(n9930), .ZN(n9777) );
  AND2_X1 U12384 ( .A1(n15598), .A2(n9762), .ZN(n15565) );
  NAND2_X1 U12385 ( .A1(n10096), .A2(n10100), .ZN(n14487) );
  INV_X1 U12386 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11658) );
  INV_X1 U12387 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11256) );
  INV_X1 U12388 ( .A(n12405), .ZN(n17075) );
  INV_X1 U12389 ( .A(n17075), .ZN(n17268) );
  OR2_X1 U12390 ( .A1(n15171), .A2(n10025), .ZN(n9778) );
  AND2_X1 U12391 ( .A1(n11523), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n9779) );
  INV_X1 U12392 ( .A(n14557), .ZN(n10107) );
  NOR2_X1 U12393 ( .A1(n16399), .A2(n13910), .ZN(n9780) );
  NAND2_X1 U12394 ( .A1(n9729), .A2(n10366), .ZN(n9781) );
  NOR3_X1 U12395 ( .A1(n10160), .A2(n15170), .A3(n10128), .ZN(n15156) );
  NAND2_X1 U12396 ( .A1(n15598), .A2(n15767), .ZN(n15590) );
  OR2_X1 U12397 ( .A1(n9721), .A2(n16233), .ZN(n9782) );
  INV_X1 U12398 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11515) );
  INV_X2 U12399 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20841) );
  INV_X1 U12400 ( .A(n9977), .ZN(n16383) );
  OR2_X1 U12401 ( .A1(n10458), .A2(n10457), .ZN(n10459) );
  INV_X1 U12402 ( .A(n10459), .ZN(n10047) );
  AND2_X1 U12403 ( .A1(n11363), .A2(n11380), .ZN(n9783) );
  OR2_X2 U12404 ( .A1(n10362), .A2(n10361), .ZN(n20157) );
  INV_X1 U12405 ( .A(n20157), .ZN(n10415) );
  AND3_X1 U12406 ( .A1(n11171), .A2(n11196), .A3(n11170), .ZN(n13450) );
  NOR2_X1 U12407 ( .A1(n10160), .A2(n15170), .ZN(n15157) );
  NAND2_X1 U12408 ( .A1(n15195), .A2(n15194), .ZN(n15171) );
  OR2_X1 U12409 ( .A1(n12113), .A2(n12114), .ZN(n9784) );
  AND2_X1 U12410 ( .A1(n12447), .A2(n12449), .ZN(n9785) );
  AND2_X1 U12411 ( .A1(n9907), .A2(n10996), .ZN(n9786) );
  OR2_X1 U12412 ( .A1(n17666), .A2(n10156), .ZN(n9787) );
  AND2_X1 U12413 ( .A1(n10085), .A2(n10082), .ZN(n9788) );
  AND2_X1 U12414 ( .A1(n11759), .A2(n9780), .ZN(n9789) );
  AND2_X1 U12415 ( .A1(n11679), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9790) );
  INV_X1 U12416 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16415) );
  INV_X1 U12417 ( .A(n11401), .ZN(n12003) );
  NAND4_X2 U12418 ( .A1(n11657), .A2(n11656), .A3(n11655), .A4(n11654), .ZN(
        n11763) );
  NOR2_X1 U12419 ( .A1(n15108), .A2(n15132), .ZN(n9791) );
  INV_X1 U12420 ( .A(n11513), .ZN(n11738) );
  NAND2_X1 U12421 ( .A1(n11760), .A2(n11759), .ZN(n13909) );
  AND2_X1 U12422 ( .A1(n14016), .A2(n14018), .ZN(n14089) );
  NAND2_X1 U12423 ( .A1(n10147), .A2(n13757), .ZN(n13758) );
  OAI21_X1 U12424 ( .B1(n16079), .B2(n16078), .A(n18930), .ZN(n17486) );
  INV_X1 U12425 ( .A(n17486), .ZN(n9929) );
  OR2_X1 U12426 ( .A1(n14528), .A2(n9942), .ZN(n9792) );
  AND2_X1 U12427 ( .A1(n12284), .A2(n15823), .ZN(n9793) );
  INV_X1 U12428 ( .A(n9951), .ZN(n16101) );
  NOR2_X1 U12429 ( .A1(n13955), .A2(n13956), .ZN(n9951) );
  XOR2_X1 U12430 ( .A(n12905), .B(n11951), .Z(n9794) );
  AND2_X1 U12431 ( .A1(n17371), .A2(n9927), .ZN(n9795) );
  NAND2_X1 U12432 ( .A1(n10100), .A2(n10099), .ZN(n9796) );
  NAND2_X1 U12433 ( .A1(n13605), .A2(n10672), .ZN(n13786) );
  AND2_X1 U12434 ( .A1(n10426), .A2(n10443), .ZN(n11071) );
  AND2_X1 U12435 ( .A1(n9957), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9797) );
  NAND2_X1 U12436 ( .A1(n13719), .A2(n11042), .ZN(n13801) );
  NAND2_X1 U12437 ( .A1(n17690), .A2(n17968), .ZN(n17750) );
  AND2_X1 U12438 ( .A1(n10030), .A2(n10028), .ZN(n9798) );
  AND2_X1 U12439 ( .A1(n10672), .A2(n10095), .ZN(n9799) );
  AND2_X1 U12440 ( .A1(n9759), .A2(n10122), .ZN(n9800) );
  AND2_X1 U12441 ( .A1(n16337), .A2(n16336), .ZN(n9801) );
  INV_X1 U12442 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20815) );
  XNOR2_X1 U12443 ( .A(n14171), .B(n14195), .ZN(n15463) );
  OR2_X1 U12444 ( .A1(n17868), .A2(n17974), .ZN(n9802) );
  AND2_X1 U12445 ( .A1(n15765), .A2(n15272), .ZN(n15259) );
  NOR3_X1 U12446 ( .A1(n15152), .A2(n12139), .A3(n20856), .ZN(n9803) );
  NAND2_X1 U12447 ( .A1(n9751), .A2(n10132), .ZN(n15255) );
  NOR2_X1 U12448 ( .A1(n15465), .A2(n14172), .ZN(n15418) );
  INV_X1 U12449 ( .A(n9843), .ZN(n15465) );
  NAND2_X1 U12450 ( .A1(n11309), .A2(n11922), .ZN(n12348) );
  INV_X1 U12451 ( .A(n9884), .ZN(n15180) );
  NAND2_X1 U12452 ( .A1(n9740), .A2(n9885), .ZN(n9884) );
  AND2_X1 U12453 ( .A1(n14632), .A2(n16100), .ZN(n9804) );
  AND2_X1 U12454 ( .A1(n11701), .A2(n11700), .ZN(n11756) );
  AND2_X1 U12455 ( .A1(n19150), .A2(n13218), .ZN(n9805) );
  NAND2_X1 U12456 ( .A1(n11386), .A2(n11308), .ZN(n11911) );
  NOR2_X1 U12457 ( .A1(n13958), .A2(n15283), .ZN(n14019) );
  AND2_X1 U12458 ( .A1(n10130), .A2(n10129), .ZN(n9806) );
  NAND2_X1 U12459 ( .A1(n15574), .A2(n15594), .ZN(n9807) );
  AND2_X1 U12460 ( .A1(n12284), .A2(n10036), .ZN(n9808) );
  AOI21_X1 U12461 ( .B1(n11032), .B2(n10797), .A(n10657), .ZN(n13604) );
  OR3_X1 U12462 ( .A1(n11828), .A2(n12139), .A3(n21013), .ZN(n15593) );
  NOR2_X1 U12463 ( .A1(n14536), .A2(n14546), .ZN(n9809) );
  AND2_X1 U12464 ( .A1(n11070), .A2(n10055), .ZN(n9810) );
  XNOR2_X1 U12465 ( .A(n14217), .B(n14214), .ZN(n15413) );
  AND2_X1 U12466 ( .A1(n9799), .A2(n13820), .ZN(n9811) );
  AND2_X1 U12467 ( .A1(n9800), .A2(n13727), .ZN(n9812) );
  AND2_X1 U12468 ( .A1(n9798), .A2(n15901), .ZN(n9813) );
  NAND2_X1 U12471 ( .A1(n14406), .A2(n14422), .ZN(n9814) );
  INV_X1 U12472 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9958) );
  INV_X1 U12473 ( .A(n17795), .ZN(n17868) );
  NOR2_X2 U12474 ( .A1(n17458), .A2(n12500), .ZN(n17795) );
  AND2_X1 U12475 ( .A1(n14242), .A2(n14239), .ZN(n9815) );
  NOR2_X1 U12476 ( .A1(n12231), .A2(n12230), .ZN(n9816) );
  NAND2_X1 U12477 ( .A1(n10027), .A2(n10030), .ZN(n15334) );
  NOR2_X1 U12478 ( .A1(n15331), .A2(n13028), .ZN(n13027) );
  AND2_X1 U12479 ( .A1(n10034), .A2(n15260), .ZN(n9817) );
  NOR2_X1 U12480 ( .A1(n13523), .A2(n13007), .ZN(n12999) );
  AND3_X1 U12481 ( .A1(n11393), .A2(n11392), .A3(n12357), .ZN(n12342) );
  NOR2_X1 U12482 ( .A1(n12993), .A2(n12995), .ZN(n12994) );
  NOR2_X1 U12483 ( .A1(n12892), .A2(n12122), .ZN(n13358) );
  AND2_X1 U12484 ( .A1(n19325), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n9818) );
  AND2_X1 U12485 ( .A1(n16291), .A2(n14018), .ZN(n9819) );
  NAND2_X1 U12486 ( .A1(n14195), .A2(n14194), .ZN(n9820) );
  INV_X1 U12487 ( .A(n11813), .ZN(n10021) );
  AND2_X1 U12488 ( .A1(n10018), .A2(n16293), .ZN(n9821) );
  OR2_X1 U12489 ( .A1(n10144), .A2(n15705), .ZN(n9823) );
  INV_X1 U12490 ( .A(n10084), .ZN(n10083) );
  OR2_X1 U12491 ( .A1(n16560), .A2(n16015), .ZN(n10084) );
  INV_X1 U12492 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10173) );
  OR2_X1 U12493 ( .A1(n13024), .A2(n10148), .ZN(n10149) );
  AND2_X1 U12494 ( .A1(n9819), .A2(n15427), .ZN(n9824) );
  AND2_X1 U12495 ( .A1(n9760), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9825) );
  AND2_X1 U12496 ( .A1(n9761), .A2(n15209), .ZN(n9826) );
  AND2_X1 U12497 ( .A1(n13759), .A2(n13757), .ZN(n9827) );
  INV_X1 U12498 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10060) );
  NAND2_X1 U12499 ( .A1(n17751), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16826) );
  NAND2_X1 U12500 ( .A1(n12721), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17604) );
  AND2_X1 U12501 ( .A1(n12721), .A2(n9749), .ZN(n9828) );
  INV_X1 U12502 ( .A(n15546), .ZN(n10143) );
  INV_X1 U12503 ( .A(n13623), .ZN(n10123) );
  INV_X1 U12504 ( .A(n15256), .ZN(n10131) );
  INV_X1 U12505 ( .A(n11856), .ZN(n10015) );
  NAND2_X1 U12506 ( .A1(n12307), .A2(n12306), .ZN(n9829) );
  AND2_X1 U12507 ( .A1(n11845), .A2(n9766), .ZN(n9830) );
  AND3_X1 U12508 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .ZN(n9831) );
  AND2_X1 U12509 ( .A1(n11845), .A2(n9764), .ZN(n9832) );
  INV_X1 U12510 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9888) );
  INV_X1 U12511 ( .A(n12350), .ZN(n19319) );
  INV_X1 U12512 ( .A(n12350), .ZN(n9852) );
  INV_X1 U12513 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n9892) );
  AND3_X1 U12514 ( .A1(n12255), .A2(n12254), .A3(n12253), .ZN(n13372) );
  INV_X1 U12515 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17873) );
  AND2_X1 U12516 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n9833) );
  AND2_X1 U12517 ( .A1(n14904), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9834) );
  INV_X1 U12518 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n10017) );
  AND3_X1 U12519 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .ZN(n9835) );
  AND2_X1 U12520 ( .A1(n14740), .A2(n14958), .ZN(n9836) );
  INV_X1 U12521 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10055) );
  NAND3_X2 U12522 ( .A1(n18946), .A2(n18945), .A3(n18935), .ZN(n18280) );
  AOI22_X2 U12523 ( .A1(DATAI_17_), .A2(n20131), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20171), .ZN(n20620) );
  NAND2_X1 U12524 ( .A1(n9756), .A2(n15408), .ZN(n9837) );
  OR2_X2 U12525 ( .A1(n15406), .A2(n15410), .ZN(n15408) );
  XNOR2_X2 U12526 ( .A(n11984), .B(n11983), .ZN(n12982) );
  NAND2_X2 U12527 ( .A1(n11439), .A2(n11438), .ZN(n11984) );
  NAND2_X1 U12528 ( .A1(n13620), .A2(n13622), .ZN(n13743) );
  NOR2_X2 U12529 ( .A1(n13024), .A2(n9754), .ZN(n13374) );
  AND2_X2 U12530 ( .A1(n11415), .A2(n12355), .ZN(n12012) );
  NAND3_X1 U12531 ( .A1(n9843), .A2(n9820), .A3(n10150), .ZN(n9842) );
  AND2_X4 U12532 ( .A1(n11511), .A2(n13290), .ZN(n11353) );
  INV_X2 U12533 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13290) );
  AND2_X2 U12534 ( .A1(n11658), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11511) );
  AND2_X2 U12535 ( .A1(n9845), .A2(n11256), .ZN(n14140) );
  NAND2_X2 U12536 ( .A1(n9847), .A2(n11405), .ZN(n11440) );
  NAND2_X1 U12537 ( .A1(n11409), .A2(n9790), .ZN(n9848) );
  NAND2_X1 U12538 ( .A1(n11410), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9849) );
  NAND3_X1 U12539 ( .A1(n11369), .A2(n19943), .A3(n11377), .ZN(n12356) );
  NAND2_X1 U12540 ( .A1(n11408), .A2(n19943), .ZN(n9850) );
  NAND2_X1 U12541 ( .A1(n11374), .A2(n11375), .ZN(n12343) );
  NAND3_X1 U12542 ( .A1(n9860), .A2(n9858), .A3(n9857), .ZN(P2_U2996) );
  XNOR2_X2 U12543 ( .A(n11958), .B(n11708), .ZN(n11960) );
  NAND3_X1 U12544 ( .A1(n10145), .A2(n11955), .A3(n11682), .ZN(n11958) );
  OAI21_X2 U12545 ( .B1(n11969), .B2(n9774), .A(n9861), .ZN(n16395) );
  NAND2_X1 U12546 ( .A1(n16395), .A2(n16393), .ZN(n11979) );
  NOR2_X2 U12547 ( .A1(n16381), .A2(n16380), .ZN(n9977) );
  NAND3_X1 U12548 ( .A1(n9870), .A2(n9869), .A3(n9866), .ZN(n9863) );
  NAND3_X1 U12549 ( .A1(n11259), .A2(n9867), .A3(n9868), .ZN(n9864) );
  NAND2_X1 U12550 ( .A1(n11355), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n9866) );
  NAND2_X1 U12551 ( .A1(n14292), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n9869) );
  NAND2_X1 U12552 ( .A1(n14140), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n9870) );
  NAND2_X1 U12553 ( .A1(n12858), .A2(n12868), .ZN(n13071) );
  NAND2_X2 U12554 ( .A1(n9871), .A2(n20135), .ZN(n12868) );
  NAND3_X1 U12555 ( .A1(n10365), .A2(n10366), .A3(n9872), .ZN(n12858) );
  NOR2_X1 U12556 ( .A1(n10422), .A2(n20135), .ZN(n9872) );
  NAND2_X1 U12557 ( .A1(n13071), .A2(n12918), .ZN(n13155) );
  INV_X1 U12558 ( .A(n10988), .ZN(n10533) );
  NAND2_X2 U12559 ( .A1(n9875), .A2(n11063), .ZN(n11064) );
  NAND3_X1 U12560 ( .A1(n11059), .A2(n14873), .A3(n11049), .ZN(n9875) );
  NAND3_X1 U12561 ( .A1(n10974), .A2(n11031), .A3(n11024), .ZN(n11027) );
  NAND2_X1 U12562 ( .A1(n14765), .A2(n14734), .ZN(n14762) );
  NAND2_X1 U12563 ( .A1(n15143), .A2(n19034), .ZN(n9881) );
  INV_X1 U12564 ( .A(n9889), .ZN(n15131) );
  INV_X1 U12565 ( .A(n9893), .ZN(n15119) );
  INV_X1 U12566 ( .A(n9897), .ZN(n15125) );
  NAND3_X1 U12567 ( .A1(n9898), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n15112) );
  NAND4_X1 U12568 ( .A1(n9898), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9900) );
  INV_X1 U12569 ( .A(n9900), .ZN(n15110) );
  INV_X1 U12570 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9899) );
  NAND2_X1 U12571 ( .A1(n13537), .A2(n13536), .ZN(n9901) );
  NAND2_X1 U12572 ( .A1(n13543), .A2(n13544), .ZN(n9902) );
  NAND2_X1 U12573 ( .A1(n14745), .A2(n11068), .ZN(n9905) );
  NAND2_X1 U12574 ( .A1(n14745), .A2(n9721), .ZN(n9903) );
  NAND2_X1 U12575 ( .A1(n9905), .A2(n14734), .ZN(n9904) );
  NAND2_X1 U12576 ( .A1(n9786), .A2(n10995), .ZN(n9912) );
  NAND2_X1 U12577 ( .A1(n9914), .A2(n9906), .ZN(n9908) );
  AND2_X1 U12578 ( .A1(n9913), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n9906) );
  INV_X1 U12579 ( .A(n13045), .ZN(n9907) );
  NAND2_X1 U12580 ( .A1(n13140), .A2(n9911), .ZN(n9910) );
  NAND2_X1 U12581 ( .A1(n9909), .A2(n9908), .ZN(n13567) );
  AND2_X1 U12582 ( .A1(n9912), .A2(n9910), .ZN(n9909) );
  NAND2_X1 U12583 ( .A1(n9914), .A2(n9913), .ZN(n10997) );
  OAI211_X1 U12584 ( .C1(n18322), .C2(n13822), .A(n12627), .B(n18309), .ZN(
        n12628) );
  NAND3_X1 U12585 ( .A1(n9835), .A2(P3_EAX_REG_21__SCAN_IN), .A3(
        P3_EAX_REG_20__SCAN_IN), .ZN(n9935) );
  INV_X1 U12586 ( .A(n14498), .ZN(n9943) );
  NOR2_X1 U12587 ( .A1(n14463), .A2(n14451), .ZN(n14450) );
  INV_X1 U12588 ( .A(n14432), .ZN(n9948) );
  AOI21_X1 U12589 ( .B1(n10447), .B2(n16072), .A(n20724), .ZN(n13146) );
  NOR2_X1 U12590 ( .A1(n10388), .A2(n10447), .ZN(n11146) );
  NAND2_X1 U12591 ( .A1(n10388), .A2(n10447), .ZN(n11075) );
  NAND2_X1 U12592 ( .A1(n10430), .A2(n10447), .ZN(n13583) );
  OAI21_X1 U12593 ( .B1(n11141), .B2(n11140), .A(n10447), .ZN(n11142) );
  NOR2_X1 U12594 ( .A1(n12859), .A2(n10447), .ZN(n16256) );
  NAND2_X1 U12595 ( .A1(n11098), .A2(n10447), .ZN(n11117) );
  AOI21_X1 U12596 ( .B1(n11089), .B2(n10447), .A(n9952), .ZN(n11098) );
  AND2_X1 U12597 ( .A1(n11149), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U12598 ( .A1(n20172), .A2(n10447), .ZN(n20477) );
  NAND2_X1 U12599 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n9954) );
  NAND2_X1 U12600 ( .A1(n9953), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16906) );
  INV_X1 U12601 ( .A(n16933), .ZN(n9959) );
  NAND2_X1 U12602 ( .A1(n16813), .A2(n9963), .ZN(n9960) );
  OR2_X1 U12603 ( .A1(n16813), .A2(n16933), .ZN(n9964) );
  OAI22_X1 U12604 ( .A1(n13690), .A2(n9971), .B1(n13691), .B2(n13692), .ZN(
        n16410) );
  NAND2_X1 U12605 ( .A1(n12352), .A2(n13635), .ZN(n12357) );
  INV_X1 U12606 ( .A(n11385), .ZN(n9974) );
  NAND3_X1 U12607 ( .A1(n11393), .A2(n9973), .A3(n12357), .ZN(n11416) );
  NAND3_X1 U12608 ( .A1(n11394), .A2(n9974), .A3(n11416), .ZN(n11426) );
  AND3_X2 U12609 ( .A1(n15348), .A2(n12365), .A3(n19943), .ZN(n9975) );
  NAND2_X1 U12610 ( .A1(n9976), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16356) );
  NAND2_X1 U12611 ( .A1(n15886), .A2(n11794), .ZN(n16355) );
  NAND2_X1 U12612 ( .A1(n15601), .A2(n9981), .ZN(n9980) );
  NAND2_X1 U12613 ( .A1(n11760), .A2(n9789), .ZN(n9993) );
  CLKBUF_X1 U12614 ( .A(n9993), .Z(n9989) );
  OAI21_X1 U12615 ( .B1(n9999), .B2(n13635), .A(n9998), .ZN(n11929) );
  NAND3_X1 U12616 ( .A1(n10002), .A2(n11539), .A3(n10001), .ZN(n10000) );
  AND2_X1 U12617 ( .A1(n15093), .A2(n10014), .ZN(n11872) );
  NAND2_X1 U12618 ( .A1(n15093), .A2(n10012), .ZN(n15094) );
  NAND2_X1 U12619 ( .A1(n15093), .A2(n11856), .ZN(n11859) );
  AND2_X1 U12620 ( .A1(n11846), .A2(n9832), .ZN(n11852) );
  AND2_X1 U12621 ( .A1(n11846), .A2(n11845), .ZN(n15218) );
  NAND2_X1 U12622 ( .A1(n11846), .A2(n9830), .ZN(n11857) );
  NAND2_X1 U12623 ( .A1(n10029), .A2(n9813), .ZN(n15902) );
  CLKBUF_X1 U12624 ( .A(n10029), .Z(n10027) );
  XNOR2_X1 U12625 ( .A(n12113), .B(n12114), .ZN(n13032) );
  OAI21_X1 U12626 ( .B1(n13032), .B2(n13031), .A(n9784), .ZN(n10032) );
  NAND2_X1 U12627 ( .A1(n12284), .A2(n10035), .ZN(n13958) );
  INV_X1 U12628 ( .A(n10039), .ZN(n10534) );
  NAND2_X1 U12629 ( .A1(n10039), .A2(n10988), .ZN(n10547) );
  NAND2_X1 U12630 ( .A1(n10528), .A2(n10535), .ZN(n10039) );
  NAND2_X1 U12631 ( .A1(n10552), .A2(n20815), .ZN(n10041) );
  XNOR2_X2 U12632 ( .A(n9736), .B(n10481), .ZN(n10552) );
  OAI21_X2 U12633 ( .B1(n10552), .B2(n10044), .A(n10042), .ZN(n10527) );
  NAND2_X1 U12634 ( .A1(n10530), .A2(n10531), .ZN(n10529) );
  OAI211_X2 U12635 ( .C1(n10530), .C2(n10047), .A(n10045), .B(n10466), .ZN(
        n13476) );
  NAND2_X1 U12636 ( .A1(n14723), .A2(n9810), .ZN(n10049) );
  INV_X1 U12637 ( .A(n14716), .ZN(n10051) );
  INV_X1 U12638 ( .A(n11126), .ZN(n14931) );
  NAND3_X1 U12639 ( .A1(n10054), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n10053), .ZN(n10052) );
  NAND2_X2 U12640 ( .A1(n11048), .A2(n9755), .ZN(n14873) );
  INV_X2 U12641 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18900) );
  NOR2_X2 U12642 ( .A1(n12514), .A2(n17988), .ZN(n17625) );
  NAND3_X1 U12643 ( .A1(n10065), .A2(n10064), .A3(n10063), .ZN(n10062) );
  NAND4_X1 U12644 ( .A1(n10070), .A2(n10069), .A3(n10068), .A4(n10067), .ZN(
        n10066) );
  NAND2_X1 U12645 ( .A1(n16565), .A2(n12515), .ZN(n10085) );
  NAND2_X1 U12646 ( .A1(n10086), .A2(n12518), .ZN(n12516) );
  AND2_X4 U12647 ( .A1(n11512), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11355) );
  AND2_X2 U12648 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11512) );
  NAND2_X1 U12649 ( .A1(n13519), .A2(n10090), .ZN(n10087) );
  NAND2_X1 U12650 ( .A1(n15598), .A2(n9763), .ZN(n15706) );
  NOR2_X1 U12651 ( .A1(n15551), .A2(n10092), .ZN(n15508) );
  AND2_X2 U12652 ( .A1(n13473), .A2(n13458), .ZN(n10313) );
  NOR2_X4 U12653 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13473) );
  NAND2_X1 U12654 ( .A1(n13605), .A2(n9811), .ZN(n13819) );
  NAND2_X1 U12655 ( .A1(n9737), .A2(n10097), .ZN(n14460) );
  NAND2_X1 U12656 ( .A1(n13063), .A2(n13064), .ZN(n13132) );
  NAND2_X1 U12657 ( .A1(n14393), .A2(n14394), .ZN(n11135) );
  NAND2_X1 U12658 ( .A1(n14393), .A2(n10109), .ZN(n10113) );
  INV_X1 U12659 ( .A(n15331), .ZN(n10115) );
  NAND2_X1 U12660 ( .A1(n10115), .A2(n10116), .ZN(n15866) );
  NAND2_X1 U12661 ( .A1(n15826), .A2(n9812), .ZN(n13726) );
  OR3_X1 U12662 ( .A1(n10160), .A2(n10127), .A3(n15170), .ZN(n15390) );
  INV_X1 U12663 ( .A(n15158), .ZN(n10128) );
  NAND2_X2 U12664 ( .A1(n12359), .A2(n11371), .ZN(n13635) );
  NAND2_X2 U12665 ( .A1(n11332), .A2(n11333), .ZN(n12359) );
  NAND2_X1 U12666 ( .A1(n11798), .A2(n11797), .ZN(n15568) );
  NAND3_X1 U12667 ( .A1(n10135), .A2(n10134), .A3(n15728), .ZN(n15557) );
  NAND3_X1 U12668 ( .A1(n11798), .A2(n10138), .A3(n15729), .ZN(n10135) );
  NAND2_X1 U12669 ( .A1(n15515), .A2(n10157), .ZN(n11863) );
  INV_X1 U12670 ( .A(n10158), .ZN(n10144) );
  INV_X1 U12671 ( .A(n11683), .ZN(n10145) );
  NAND2_X1 U12672 ( .A1(n10145), .A2(n11682), .ZN(n11956) );
  AND2_X4 U12673 ( .A1(n11512), .A2(n13290), .ZN(n11498) );
  NAND3_X1 U12674 ( .A1(n11414), .A2(n11413), .A3(n10146), .ZN(n11450) );
  INV_X4 U12675 ( .A(n11371), .ZN(n14263) );
  NAND2_X2 U12676 ( .A1(n11345), .A2(n11346), .ZN(n11371) );
  NAND2_X1 U12677 ( .A1(n10147), .A2(n9827), .ZN(n13997) );
  INV_X1 U12678 ( .A(n10149), .ZN(n13371) );
  NAND2_X1 U12679 ( .A1(n14016), .A2(n9824), .ZN(n15425) );
  INV_X1 U12680 ( .A(n15425), .ZN(n14126) );
  NAND2_X1 U12681 ( .A1(n14419), .A2(n14421), .ZN(n14409) );
  NOR2_X2 U12682 ( .A1(n14435), .A2(n14437), .ZN(n14419) );
  NAND2_X1 U12683 ( .A1(n15499), .A2(n16460), .ZN(n12395) );
  AND2_X1 U12684 ( .A1(n20208), .A2(n20207), .ZN(n20601) );
  NOR2_X1 U12685 ( .A1(n20208), .A2(n20207), .ZN(n20572) );
  NOR2_X1 U12686 ( .A1(n20208), .A2(n20133), .ZN(n20540) );
  CLKBUF_X1 U12687 ( .A(n13049), .Z(n16425) );
  CLKBUF_X1 U12688 ( .A(n13766), .Z(n13768) );
  NAND2_X1 U12689 ( .A1(n14448), .A2(n14449), .ZN(n14435) );
  NAND2_X1 U12690 ( .A1(n11956), .A2(n11685), .ZN(n11947) );
  NAND2_X1 U12691 ( .A1(n12994), .A2(n15330), .ZN(n15331) );
  NOR2_X2 U12692 ( .A1(n14460), .A2(n14462), .ZN(n14448) );
  XNOR2_X1 U12693 ( .A(n14241), .B(n9815), .ZN(n15406) );
  OAI22_X1 U12694 ( .A1(n11440), .A2(n11415), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n12012), .ZN(n11421) );
  AOI21_X1 U12695 ( .B1(n14721), .B2(n16152), .A(n14720), .ZN(n14722) );
  AOI22_X1 U12696 ( .A1(n14140), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11330) );
  NAND2_X1 U12697 ( .A1(n10868), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10369) );
  AOI22_X1 U12698 ( .A1(n10868), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10302), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10305) );
  INV_X1 U12699 ( .A(n19970), .ZN(n11125) );
  AND2_X1 U12700 ( .A1(n17795), .A2(n18093), .ZN(n10153) );
  AND4_X1 U12701 ( .A1(n12438), .A2(n12437), .A3(n12436), .A4(n12435), .ZN(
        n10154) );
  AND3_X1 U12702 ( .A1(n12442), .A2(n12441), .A3(n12440), .ZN(n10155) );
  NAND2_X1 U12703 ( .A1(n11347), .A2(n12367), .ZN(n11408) );
  AND3_X1 U12704 ( .A1(n17685), .A2(n18012), .A3(n20842), .ZN(n10156) );
  INV_X1 U12705 ( .A(n13132), .ZN(n10555) );
  NAND2_X1 U12706 ( .A1(n16118), .A2(n14071), .ZN(n14636) );
  INV_X1 U12707 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10455) );
  OR2_X1 U12708 ( .A1(n15518), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10157) );
  AND2_X1 U12709 ( .A1(n11851), .A2(n11763), .ZN(n10158) );
  INV_X2 U12710 ( .A(n17338), .ZN(n17332) );
  OR2_X1 U12711 ( .A1(n17554), .A2(n17599), .ZN(n17602) );
  AND2_X1 U12712 ( .A1(n18143), .A2(n18117), .ZN(n10159) );
  INV_X1 U12713 ( .A(n11483), .ZN(n11484) );
  AND3_X1 U12714 ( .A1(n11350), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11349), .ZN(n10161) );
  AND2_X1 U12715 ( .A1(n12960), .A2(n12961), .ZN(n12113) );
  INV_X1 U12716 ( .A(n20207), .ZN(n20133) );
  NOR2_X2 U12717 ( .A1(n21125), .A2(n20811), .ZN(n10797) );
  INV_X1 U12718 ( .A(n14932), .ZN(n11254) );
  OR2_X1 U12719 ( .A1(n11047), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10162) );
  INV_X1 U12720 ( .A(n11443), .ZN(n12002) );
  NOR2_X1 U12721 ( .A1(n12407), .A2(n12403), .ZN(n12450) );
  INV_X1 U12722 ( .A(n12579), .ZN(n13871) );
  INV_X1 U12723 ( .A(n13674), .ZN(n19294) );
  NAND3_X1 U12724 ( .A1(n19894), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19765), 
        .ZN(n13674) );
  INV_X1 U12725 ( .A(n12087), .ZN(n12338) );
  INV_X1 U12726 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n12874) );
  OR2_X1 U12727 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n10971) );
  INV_X1 U12728 ( .A(n20135), .ZN(n10430) );
  INV_X1 U12729 ( .A(n11089), .ZN(n11106) );
  NAND2_X1 U12730 ( .A1(n11388), .A2(n11387), .ZN(n11389) );
  OR3_X1 U12731 ( .A1(n11106), .A2(n11105), .A3(n12862), .ZN(n11107) );
  OAI21_X1 U12732 ( .B1(n9781), .B2(n10432), .A(n10431), .ZN(n10433) );
  AND2_X2 U12733 ( .A1(n11515), .A2(n11258), .ZN(n11334) );
  NAND2_X1 U12734 ( .A1(n19912), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11672) );
  OAI22_X1 U12735 ( .A1(n11552), .A2(n19627), .B1(n11608), .B2(n11551), .ZN(
        n11553) );
  NOR2_X1 U12736 ( .A1(n11401), .A2(n11428), .ZN(n11429) );
  AOI22_X1 U12737 ( .A1(n11514), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14292), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11300) );
  NAND2_X1 U12738 ( .A1(n10388), .A2(n10449), .ZN(n10424) );
  NAND2_X1 U12739 ( .A1(n13020), .A2(n13019), .ZN(n13021) );
  OR2_X1 U12740 ( .A1(n14212), .A2(n14215), .ZN(n14238) );
  AOI22_X1 U12741 ( .A1(n14127), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14140), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11338) );
  AND2_X1 U12742 ( .A1(n11641), .A2(n11640), .ZN(n11708) );
  NAND2_X1 U12743 ( .A1(n11443), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11432) );
  AOI22_X1 U12744 ( .A1(n11353), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11498), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11325) );
  NOR2_X1 U12745 ( .A1(n11113), .A2(n11112), .ZN(n12863) );
  INV_X1 U12746 ( .A(n13449), .ZN(n10608) );
  OR2_X1 U12747 ( .A1(n13819), .A2(n10722), .ZN(n10723) );
  INV_X1 U12748 ( .A(n13806), .ZN(n10672) );
  OR2_X1 U12749 ( .A1(n10639), .A2(n10638), .ZN(n11034) );
  NAND2_X1 U12750 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10367) );
  AND2_X1 U12751 ( .A1(n10355), .A2(n10354), .ZN(n10360) );
  INV_X1 U12752 ( .A(n11911), .ZN(n11914) );
  NAND2_X1 U12753 ( .A1(n9741), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11501) );
  NOR2_X1 U12754 ( .A1(n12402), .A2(n12403), .ZN(n12579) );
  OR2_X1 U12755 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20127), .ZN(
        n11112) );
  AND2_X1 U12756 ( .A1(n13166), .A2(n13583), .ZN(n12918) );
  INV_X1 U12757 ( .A(n10888), .ZN(n10170) );
  NAND2_X1 U12758 ( .A1(n10748), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10724) );
  NAND2_X1 U12759 ( .A1(n10689), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10703) );
  INV_X1 U12760 ( .A(n10980), .ZN(n10979) );
  AND2_X1 U12761 ( .A1(n11202), .A2(n11201), .ZN(n14562) );
  INV_X1 U12762 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10575) );
  AND2_X1 U12763 ( .A1(n20511), .A2(n10462), .ZN(n20144) );
  AND2_X1 U12764 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n20966), .ZN(
        n11877) );
  NAND2_X1 U12765 ( .A1(n19325), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11668) );
  INV_X1 U12766 ( .A(n13372), .ZN(n13373) );
  AND2_X1 U12767 ( .A1(n14258), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12936) );
  INV_X1 U12768 ( .A(n14216), .ZN(n14214) );
  INV_X1 U12769 ( .A(n14162), .ZN(n14096) );
  INV_X1 U12770 ( .A(n15430), .ZN(n12049) );
  INV_X1 U12771 ( .A(n11450), .ZN(n11453) );
  INV_X1 U12772 ( .A(n15839), .ZN(n11797) );
  OR2_X1 U12773 ( .A1(n19049), .A2(n12139), .ZN(n11795) );
  AND4_X1 U12774 ( .A1(n11645), .A2(n11644), .A3(n11643), .A4(n11642), .ZN(
        n11657) );
  NAND2_X1 U12775 ( .A1(n12102), .A2(n12101), .ZN(n12960) );
  INV_X1 U12776 ( .A(n11488), .ZN(n11470) );
  AND3_X1 U12777 ( .A1(n11380), .A2(n12350), .A3(n11379), .ZN(n11372) );
  INV_X1 U12778 ( .A(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n20889) );
  NAND2_X1 U12779 ( .A1(n17256), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12440) );
  AND2_X1 U12780 ( .A1(n13825), .A2(n12623), .ZN(n12624) );
  AND2_X1 U12781 ( .A1(n11083), .A2(n11112), .ZN(n12865) );
  NAND2_X1 U12782 ( .A1(n10952), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10961) );
  INV_X1 U12783 ( .A(n10848), .ZN(n10168) );
  NAND2_X1 U12784 ( .A1(n10622), .A2(n10797), .ZN(n10629) );
  AOI22_X1 U12785 ( .A1(n14383), .A2(n10960), .B1(n10334), .B2(n10333), .ZN(
        n14065) );
  NAND2_X1 U12786 ( .A1(n10170), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10910) );
  NOR2_X1 U12787 ( .A1(n13972), .A2(n10703), .ZN(n10748) );
  INV_X1 U12788 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13795) );
  AND2_X1 U12789 ( .A1(n10652), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10668) );
  OR2_X1 U12790 ( .A1(n10572), .A2(n10571), .ZN(n11001) );
  OR2_X1 U12791 ( .A1(n13158), .A2(n11148), .ZN(n13183) );
  AND2_X1 U12792 ( .A1(n11181), .A2(n11180), .ZN(n13609) );
  NAND2_X1 U12793 ( .A1(n13587), .A2(n11224), .ZN(n11229) );
  INV_X1 U12794 ( .A(n20179), .ZN(n20248) );
  NAND2_X1 U12795 ( .A1(n10560), .A2(n10559), .ZN(n20285) );
  AND2_X1 U12796 ( .A1(n10557), .A2(n20649), .ZN(n20407) );
  AOI221_X1 U12797 ( .B1(n11878), .B2(n20966), .C1(n11878), .C2(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n11877), .ZN(n11903) );
  NAND2_X1 U12798 ( .A1(n11669), .A2(n11668), .ZN(n11695) );
  NAND2_X1 U12799 ( .A1(n12937), .A2(n12936), .ZN(n12979) );
  INV_X1 U12800 ( .A(n11514), .ZN(n14310) );
  INV_X1 U12801 ( .A(n9719), .ZN(n12333) );
  AND2_X1 U12802 ( .A1(n16510), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12981) );
  NOR2_X1 U12803 ( .A1(n15644), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15646) );
  AND2_X1 U12804 ( .A1(n12309), .A2(n12308), .ZN(n15299) );
  OR3_X1 U12805 ( .A1(n12896), .A2(n12895), .A3(n12373), .ZN(n13361) );
  INV_X1 U12806 ( .A(n13329), .ZN(n12951) );
  OR2_X1 U12807 ( .A1(n19592), .A2(n19531), .ZN(n19532) );
  INV_X1 U12808 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19757) );
  AND2_X1 U12809 ( .A1(n12531), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12533) );
  AND2_X1 U12810 ( .A1(n12727), .A2(n16857), .ZN(n12726) );
  AOI211_X1 U12811 ( .C1(n17220), .C2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n12604), .B(n12603), .ZN(n12605) );
  NOR2_X1 U12812 ( .A1(n12622), .A2(n13826), .ZN(n12716) );
  NAND2_X1 U12813 ( .A1(n16550), .A2(n17881), .ZN(n12684) );
  INV_X1 U12814 ( .A(n17750), .ZN(n17692) );
  NAND2_X1 U12815 ( .A1(n12513), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12511) );
  NAND2_X1 U12816 ( .A1(n17762), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12507) );
  NOR2_X1 U12817 ( .A1(n17888), .A2(n18203), .ZN(n12674) );
  OR2_X1 U12818 ( .A1(n12716), .A2(n12624), .ZN(n12625) );
  OR2_X1 U12819 ( .A1(n10961), .A2(n10171), .ZN(n13575) );
  INV_X1 U12820 ( .A(n10866), .ZN(n10169) );
  NAND2_X1 U12821 ( .A1(n10168), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10866) );
  INV_X1 U12822 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16091) );
  INV_X1 U12823 ( .A(n20042), .ZN(n19999) );
  NAND2_X1 U12824 ( .A1(n13597), .A2(n13586), .ZN(n14590) );
  INV_X1 U12825 ( .A(n14069), .ZN(n14070) );
  AND3_X1 U12826 ( .A1(n10671), .A2(n10670), .A3(n10669), .ZN(n13806) );
  AND3_X1 U12827 ( .A1(n11071), .A2(n11073), .A3(n11072), .ZN(n13144) );
  AND2_X1 U12828 ( .A1(n13550), .A2(n15037), .ZN(n20097) );
  INV_X1 U12829 ( .A(n20099), .ZN(n16201) );
  INV_X1 U12830 ( .A(n15089), .ZN(n13482) );
  OR2_X1 U12831 ( .A1(n10999), .A2(n20132), .ZN(n20242) );
  INV_X1 U12832 ( .A(n15065), .ZN(n15066) );
  AOI21_X1 U12833 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20573), .A(n20291), 
        .ZN(n20660) );
  OR2_X1 U12834 ( .A1(n12371), .A2(n12370), .ZN(n13329) );
  INV_X1 U12835 ( .A(n19126), .ZN(n19109) );
  INV_X2 U12836 ( .A(n12003), .ZN(n15099) );
  INV_X1 U12837 ( .A(n13520), .ZN(n11994) );
  OR2_X1 U12838 ( .A1(n12814), .A2(n12367), .ZN(n13265) );
  INV_X1 U12839 ( .A(n15408), .ZN(n15409) );
  AND2_X1 U12840 ( .A1(n12134), .A2(n12133), .ZN(n13528) );
  XOR2_X1 U12841 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n13628), .Z(
        n15488) );
  OR2_X1 U12842 ( .A1(n12389), .A2(n15907), .ZN(n15736) );
  NAND2_X1 U12843 ( .A1(n13368), .A2(n13367), .ZN(n13366) );
  AND2_X1 U12844 ( .A1(n11945), .A2(n15925), .ZN(n12372) );
  NAND2_X1 U12845 ( .A1(n15935), .A2(n16510), .ZN(n12876) );
  NAND2_X1 U12846 ( .A1(n19567), .A2(n13708), .ZN(n19458) );
  AND2_X1 U12847 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19714), .ZN(
        n12983) );
  AOI21_X1 U12848 ( .B1(n12530), .B2(n12529), .A(n12528), .ZN(n12644) );
  NOR2_X1 U12849 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16889), .ZN(n16871) );
  NOR2_X1 U12850 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16964), .ZN(n16942) );
  NAND2_X1 U12851 ( .A1(n18948), .A2(n17494), .ZN(n12734) );
  NOR2_X1 U12852 ( .A1(n15988), .A2(n13823), .ZN(n15972) );
  NAND3_X1 U12853 ( .A1(n12607), .A2(n12606), .A3(n12605), .ZN(n17392) );
  NOR2_X1 U12854 ( .A1(n17429), .A2(n17342), .ZN(n17343) );
  INV_X1 U12855 ( .A(n18322), .ZN(n17347) );
  OAI21_X1 U12856 ( .B1(n16558), .B2(n17972), .A(n12684), .ZN(n12685) );
  INV_X1 U12857 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17928) );
  NOR2_X1 U12858 ( .A1(n17890), .A2(n17889), .ZN(n17888) );
  NAND2_X1 U12859 ( .A1(n12673), .A2(n17896), .ZN(n17889) );
  OR2_X1 U12860 ( .A1(n18909), .A2(n18800), .ZN(n18300) );
  INV_X1 U12861 ( .A(n18445), .ZN(n18589) );
  NAND2_X1 U12862 ( .A1(n18589), .A2(n18641), .ZN(n18313) );
  AOI22_X1 U12863 ( .A1(n18769), .A2(n18767), .B1(n18773), .B2(n18766), .ZN(
        n18778) );
  NAND2_X1 U12864 ( .A1(n11124), .A2(n11123), .ZN(n16055) );
  NAND2_X1 U12865 ( .A1(n10169), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10888) );
  INV_X1 U12866 ( .A(n14571), .ZN(n20018) );
  AND2_X1 U12867 ( .A1(n13597), .A2(n13589), .ZN(n20024) );
  NOR2_X1 U12868 ( .A1(n16118), .A2(n11252), .ZN(n11253) );
  INV_X1 U12869 ( .A(n16118), .ZN(n14623) );
  INV_X1 U12870 ( .A(n14636), .ZN(n16115) );
  INV_X1 U12871 ( .A(n14638), .ZN(n16116) );
  BUF_X1 U12872 ( .A(n14409), .Z(n14420) );
  INV_X1 U12873 ( .A(n14683), .ZN(n14701) );
  NAND2_X1 U12874 ( .A1(n13060), .A2(n13210), .ZN(n14679) );
  INV_X1 U12875 ( .A(n13228), .ZN(n13253) );
  AND2_X1 U12876 ( .A1(n13179), .A2(n13165), .ZN(n20083) );
  NOR2_X1 U12877 ( .A1(n10107), .A2(n14631), .ZN(n16096) );
  INV_X1 U12878 ( .A(n20129), .ZN(n16152) );
  AND2_X1 U12879 ( .A1(n13169), .A2(n13190), .ZN(n16207) );
  OR2_X1 U12880 ( .A1(n15035), .A2(n20122), .ZN(n20099) );
  AND2_X1 U12881 ( .A1(n13169), .A2(n13157), .ZN(n20117) );
  NOR2_X1 U12882 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16255) );
  OAI22_X1 U12883 ( .A1(n20214), .A2(n20213), .B1(n20472), .B2(n20345), .ZN(
        n20238) );
  INV_X1 U12884 ( .A(n20242), .ZN(n20251) );
  AND2_X1 U12885 ( .A1(n20208), .A2(n20133), .ZN(n20382) );
  NOR2_X1 U12886 ( .A1(n13485), .A2(n15066), .ZN(n20383) );
  INV_X1 U12887 ( .A(n20508), .ZN(n20462) );
  INV_X1 U12888 ( .A(n20533), .ZN(n20536) );
  INV_X1 U12889 ( .A(n20382), .ZN(n20509) );
  NAND2_X1 U12890 ( .A1(n13485), .A2(n10999), .ZN(n20510) );
  INV_X1 U12891 ( .A(n20606), .ZN(n20644) );
  INV_X1 U12892 ( .A(n20460), .ZN(n20655) );
  INV_X1 U12893 ( .A(n20485), .ZN(n20680) );
  INV_X1 U12894 ( .A(n20497), .ZN(n20698) );
  OR2_X1 U12895 ( .A1(n16043), .A2(n16042), .ZN(n16049) );
  INV_X1 U12896 ( .A(n13334), .ZN(n19937) );
  INV_X1 U12897 ( .A(n19129), .ZN(n19060) );
  INV_X1 U12898 ( .A(n15288), .ZN(n15431) );
  AND2_X1 U12899 ( .A1(n12980), .A2(n12943), .ZN(n19907) );
  INV_X1 U12900 ( .A(n19205), .ZN(n19231) );
  AND2_X1 U12901 ( .A1(n13378), .A2(n13377), .ZN(n19045) );
  AND2_X1 U12902 ( .A1(n12878), .A2(n14263), .ZN(n19288) );
  OAI21_X1 U12903 ( .B1(n15482), .B2(n15481), .A(n15480), .ZN(n15486) );
  NAND2_X1 U12904 ( .A1(n19210), .A2(n19915), .ZN(n19568) );
  INV_X1 U12905 ( .A(n19424), .ZN(n19412) );
  INV_X1 U12906 ( .A(n19438), .ZN(n19454) );
  NAND2_X1 U12907 ( .A1(n19907), .A2(n19915), .ZN(n19687) );
  OAI21_X1 U12908 ( .B1(n19494), .B2(n19509), .A(n19765), .ZN(n19512) );
  NOR2_X1 U12909 ( .A1(n19427), .A2(n19712), .ZN(n19492) );
  NOR2_X1 U12910 ( .A1(n19713), .A2(n19888), .ZN(n19603) );
  INV_X1 U12911 ( .A(n19808), .ZN(n19673) );
  NOR2_X1 U12912 ( .A1(n19683), .A2(n19687), .ZN(n19744) );
  NOR2_X1 U12913 ( .A1(n13961), .A2(n13674), .ZN(n19334) );
  AND2_X1 U12914 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n11944), .ZN(n15925) );
  INV_X1 U12915 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19838) );
  INV_X1 U12916 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n18956) );
  NOR2_X1 U12917 ( .A1(n15966), .A2(n15965), .ZN(n18771) );
  INV_X1 U12918 ( .A(n17015), .ZN(n17049) );
  NOR2_X1 U12919 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16820), .ZN(n16804) );
  NOR2_X1 U12920 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16839), .ZN(n16824) );
  NOR2_X1 U12921 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16914), .ZN(n16895) );
  NOR2_X1 U12922 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16988), .ZN(n16969) );
  INV_X1 U12923 ( .A(n17035), .ZN(n16992) );
  NOR2_X1 U12924 ( .A1(n18785), .A2(n12734), .ZN(n17031) );
  NOR2_X1 U12925 ( .A1(n13827), .A2(n17130), .ZN(n17113) );
  NOR2_X1 U12926 ( .A1(n17337), .A2(n17284), .ZN(n17316) );
  AOI21_X1 U12927 ( .B1(n13825), .B2(n13824), .A(n15972), .ZN(n16077) );
  INV_X1 U12928 ( .A(n18326), .ZN(n17341) );
  NOR2_X1 U12929 ( .A1(n17603), .A2(n17431), .ZN(n17423) );
  NAND2_X1 U12930 ( .A1(n17344), .A2(n17343), .ZN(n17431) );
  NOR2_X1 U12931 ( .A1(n17545), .A2(n17477), .ZN(n17476) );
  INV_X1 U12932 ( .A(n17475), .ZN(n17485) );
  INV_X1 U12933 ( .A(n17526), .ZN(n20823) );
  INV_X1 U12934 ( .A(n17553), .ZN(n17581) );
  NOR2_X2 U12935 ( .A1(n18893), .A2(n17963), .ZN(n17730) );
  NOR2_X2 U12936 ( .A1(n17458), .A2(n17971), .ZN(n17861) );
  NAND2_X1 U12937 ( .A1(n17750), .A2(n17817), .ZN(n17962) );
  NOR2_X1 U12938 ( .A1(n17650), .A2(n15999), .ZN(n17978) );
  NAND2_X1 U12939 ( .A1(n18749), .A2(n18734), .ZN(n18735) );
  INV_X1 U12940 ( .A(n18280), .ZN(n18125) );
  NOR2_X1 U12941 ( .A1(n15968), .A2(n15982), .ZN(n18766) );
  NAND2_X1 U12942 ( .A1(n18935), .A2(n18300), .ZN(n18445) );
  INV_X1 U12943 ( .A(n18562), .ZN(n18553) );
  INV_X1 U12944 ( .A(n18671), .ZN(n18663) );
  NOR2_X1 U12945 ( .A1(n18945), .A2(n18796), .ZN(n18930) );
  INV_X1 U12946 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18809) );
  INV_X1 U12947 ( .A(U212), .ZN(n16621) );
  NAND3_X1 U12948 ( .A1(n12869), .A2(n13210), .A3(n16055), .ZN(n14354) );
  OR2_X1 U12949 ( .A1(n14719), .A2(n13580), .ZN(n14571) );
  INV_X1 U12950 ( .A(n20024), .ZN(n20053) );
  INV_X1 U12951 ( .A(n16116), .ZN(n14628) );
  NAND2_X1 U12952 ( .A1(n16118), .A2(n10389), .ZN(n14638) );
  NAND2_X1 U12953 ( .A1(n13073), .A2(n20813), .ZN(n13409) );
  NOR2_X1 U12954 ( .A1(n14354), .A2(n13110), .ZN(n13179) );
  OR2_X1 U12955 ( .A1(n16135), .A2(n13041), .ZN(n16127) );
  NAND2_X2 U12956 ( .A1(n16037), .A2(n13210), .ZN(n19970) );
  INV_X1 U12957 ( .A(n20116), .ZN(n20107) );
  AND2_X1 U12958 ( .A1(n14990), .A2(n14891), .ZN(n16199) );
  INV_X1 U12959 ( .A(n20117), .ZN(n20091) );
  INV_X1 U12960 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20573) );
  NAND2_X1 U12961 ( .A1(n20251), .A2(n20540), .ZN(n20206) );
  NAND2_X1 U12962 ( .A1(n20251), .A2(n20572), .ZN(n20236) );
  NAND2_X1 U12963 ( .A1(n20251), .A2(n20601), .ZN(n20284) );
  NAND2_X1 U12964 ( .A1(n20383), .A2(n20540), .ZN(n20338) );
  NAND2_X1 U12965 ( .A1(n20383), .A2(n20601), .ZN(n20405) );
  NAND2_X1 U12966 ( .A1(n20433), .A2(n20540), .ZN(n20457) );
  OR2_X1 U12967 ( .A1(n20510), .A2(n20437), .ZN(n20508) );
  OR2_X1 U12968 ( .A1(n20510), .A2(n20458), .ZN(n20533) );
  OR2_X1 U12969 ( .A1(n20510), .A2(n20509), .ZN(n20571) );
  NAND2_X1 U12970 ( .A1(n20602), .A2(n20601), .ZN(n20712) );
  INV_X1 U12971 ( .A(n20798), .ZN(n20718) );
  INV_X1 U12972 ( .A(n20787), .ZN(n20780) );
  INV_X1 U12973 ( .A(n19125), .ZN(n19107) );
  INV_X1 U12974 ( .A(n19907), .ZN(n19210) );
  AND2_X1 U12975 ( .A1(n12929), .A2(n12832), .ZN(n19915) );
  AND2_X1 U12976 ( .A1(n12953), .A2(n15925), .ZN(n19205) );
  AND2_X1 U12977 ( .A1(n19236), .A2(n19180), .ZN(n19215) );
  INV_X1 U12978 ( .A(n19207), .ZN(n19240) );
  INV_X1 U12979 ( .A(n12970), .ZN(n19261) );
  INV_X1 U12980 ( .A(n19272), .ZN(n12835) );
  INV_X1 U12981 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16354) );
  INV_X1 U12982 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16392) );
  NAND2_X1 U12983 ( .A1(n12884), .A2(n12883), .ZN(n16428) );
  AND2_X1 U12984 ( .A1(n12395), .A2(n12394), .ZN(n12396) );
  INV_X1 U12985 ( .A(n16485), .ZN(n16498) );
  INV_X1 U12986 ( .A(n16460), .ZN(n16503) );
  OR2_X1 U12987 ( .A1(n19568), .A2(n19427), .ZN(n19378) );
  NOR2_X1 U12988 ( .A1(n13934), .A2(n19343), .ZN(n19394) );
  OR2_X1 U12989 ( .A1(n19427), .A2(n19888), .ZN(n19424) );
  NOR2_X1 U12990 ( .A1(n19433), .A2(n19431), .ZN(n19438) );
  INV_X1 U12991 ( .A(n19447), .ZN(n19457) );
  OR2_X1 U12992 ( .A1(n19427), .A2(n19687), .ZN(n19481) );
  INV_X1 U12993 ( .A(n19492), .ZN(n19529) );
  AOI21_X1 U12994 ( .B1(n19536), .B2(n19539), .A(n19535), .ZN(n19565) );
  INV_X1 U12995 ( .A(n19603), .ZN(n19662) );
  AOI211_X2 U12996 ( .C1(n13673), .C2(n13677), .A(n19343), .B(n13672), .ZN(
        n19682) );
  INV_X1 U12997 ( .A(n19744), .ZN(n19753) );
  INV_X1 U12998 ( .A(n19814), .ZN(n19795) );
  AND2_X1 U12999 ( .A1(n13344), .A2(n13343), .ZN(n16517) );
  INV_X1 U13000 ( .A(n19887), .ZN(n19884) );
  INV_X1 U13001 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16666) );
  INV_X1 U13002 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16917) );
  INV_X1 U13003 ( .A(n17019), .ZN(n17050) );
  AND2_X1 U13004 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17118), .ZN(n17112) );
  NOR2_X2 U13005 ( .A1(n18332), .A2(n17337), .ZN(n17338) );
  NOR2_X1 U13006 ( .A1(n17429), .A2(n17457), .ZN(n17443) );
  NOR2_X1 U13007 ( .A1(n12424), .A2(n12423), .ZN(n17464) );
  NAND2_X1 U13008 ( .A1(n18748), .A2(n9929), .ZN(n17490) );
  INV_X1 U13009 ( .A(n17512), .ZN(n17526) );
  INV_X1 U13010 ( .A(n20825), .ZN(n17549) );
  INV_X1 U13011 ( .A(n17600), .ZN(n17592) );
  INV_X1 U13012 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18176) );
  NAND2_X1 U13013 ( .A1(n12682), .A2(n17554), .ZN(n17971) );
  INV_X1 U13014 ( .A(n18265), .ZN(n18281) );
  INV_X1 U13015 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18752) );
  INV_X1 U13016 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18762) );
  INV_X1 U13017 ( .A(n18915), .ZN(n18912) );
  INV_X1 U13018 ( .A(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n21100) );
  INV_X1 U13019 ( .A(n18930), .ZN(n18792) );
  INV_X1 U13020 ( .A(n17690), .ZN(n18804) );
  INV_X1 U13021 ( .A(n18884), .ZN(n18882) );
  OR2_X1 U13022 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18809), .ZN(n18943) );
  INV_X1 U13023 ( .A(n16619), .ZN(n16624) );
  OAI21_X1 U13024 ( .B1(n14644), .B2(n14638), .A(n11255), .ZN(P1_U2843) );
  NAND2_X1 U13025 ( .A1(n12689), .A2(n12688), .ZN(P3_U2799) );
  INV_X1 U13026 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10167) );
  INV_X1 U13027 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10909) );
  INV_X1 U13028 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14773) );
  INV_X1 U13029 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14756) );
  INV_X1 U13030 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10942) );
  INV_X1 U13031 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10171) );
  XNOR2_X1 U13032 ( .A(n13575), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14383) );
  INV_X1 U13033 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U13035 ( .A1(n10313), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10868), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10177) );
  AND2_X2 U13036 ( .A1(n13458), .A2(n10178), .ZN(n10199) );
  AOI22_X1 U13037 ( .A1(n10199), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10314), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10176) );
  AND2_X2 U13038 ( .A1(n13458), .A2(n10180), .ZN(n10315) );
  AND2_X2 U13039 ( .A1(n10180), .A2(n10181), .ZN(n10673) );
  AND2_X2 U13040 ( .A1(n10178), .A2(n10181), .ZN(n10302) );
  AND2_X4 U13041 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13188) );
  AOI22_X1 U13042 ( .A1(n10302), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10397), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10174) );
  AND2_X4 U13044 ( .A1(n13473), .A2(n10179), .ZN(n10869) );
  AOI22_X1 U13045 ( .A1(n10320), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10869), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10186) );
  AND2_X2 U13046 ( .A1(n10180), .A2(n10179), .ZN(n10322) );
  AOI22_X1 U13047 ( .A1(n9744), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n10322), .ZN(n10183) );
  AND2_X2 U13048 ( .A1(n13473), .A2(n10181), .ZN(n10398) );
  AOI22_X1 U13049 ( .A1(n10398), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10356), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10182) );
  INV_X1 U13050 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n20950) );
  NOR2_X1 U13051 ( .A1(n20950), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10188) );
  INV_X2 U13052 ( .A(n10971), .ZN(n10960) );
  AOI211_X1 U13053 ( .C1(n10965), .C2(P1_EAX_REG_30__SCAN_IN), .A(n10188), .B(
        n10960), .ZN(n10334) );
  AOI22_X1 U13054 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10806), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10192) );
  AOI22_X1 U13055 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10900), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10191) );
  AOI22_X1 U13056 ( .A1(n9723), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U13057 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10869), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10189) );
  NAND4_X1 U13058 ( .A1(n10192), .A2(n10191), .A3(n10190), .A4(n10189), .ZN(
        n10198) );
  AOI22_X1 U13059 ( .A1(n10891), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U13060 ( .A1(n10856), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10811), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10195) );
  AOI22_X1 U13061 ( .A1(n10899), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10194) );
  AOI22_X1 U13062 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10877), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10193) );
  NAND4_X1 U13063 ( .A1(n10196), .A2(n10195), .A3(n10194), .A4(n10193), .ZN(
        n10197) );
  NOR2_X1 U13064 ( .A1(n10198), .A2(n10197), .ZN(n10964) );
  AOI22_X1 U13065 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n10890), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U13066 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n9723), .B1(
        n10811), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10202) );
  AOI22_X1 U13067 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n10876), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10201) );
  AOI22_X1 U13068 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10356), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10200) );
  NAND4_X1 U13069 ( .A1(n10203), .A2(n10202), .A3(n10201), .A4(n10200), .ZN(
        n10209) );
  AOI22_X1 U13070 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10352), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10207) );
  AOI22_X1 U13071 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10869), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10206) );
  AOI22_X1 U13072 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10856), .B1(
        n10877), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10205) );
  AOI22_X1 U13073 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10204) );
  NAND4_X1 U13074 ( .A1(n10207), .A2(n10206), .A3(n10205), .A4(n10204), .ZN(
        n10208) );
  NOR2_X1 U13075 ( .A1(n10209), .A2(n10208), .ZN(n10947) );
  AOI22_X1 U13076 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10900), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10213) );
  AOI22_X1 U13077 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10212) );
  AOI22_X1 U13078 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10211) );
  AOI22_X1 U13079 ( .A1(n10892), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10877), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10210) );
  NAND4_X1 U13080 ( .A1(n10213), .A2(n10212), .A3(n10211), .A4(n10210), .ZN(
        n10219) );
  AOI22_X1 U13081 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10217) );
  AOI22_X1 U13082 ( .A1(n10313), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10216) );
  AOI22_X1 U13083 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10215) );
  AOI22_X1 U13084 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10214) );
  NAND4_X1 U13085 ( .A1(n10217), .A2(n10216), .A3(n10215), .A4(n10214), .ZN(
        n10218) );
  NOR2_X1 U13086 ( .A1(n10219), .A2(n10218), .ZN(n10930) );
  AOI22_X1 U13087 ( .A1(n10891), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10223) );
  AOI22_X1 U13088 ( .A1(n10313), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10222) );
  AOI22_X1 U13089 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10806), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10221) );
  AOI22_X1 U13090 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10220) );
  NAND4_X1 U13091 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        n10229) );
  AOI22_X1 U13092 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10811), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10227) );
  AOI22_X1 U13093 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10673), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10226) );
  AOI22_X1 U13094 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10225) );
  AOI22_X1 U13095 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10224) );
  NAND4_X1 U13096 ( .A1(n10227), .A2(n10226), .A3(n10225), .A4(n10224), .ZN(
        n10228) );
  NOR2_X1 U13097 ( .A1(n10229), .A2(n10228), .ZN(n10912) );
  AOI22_X1 U13098 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10851), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10233) );
  AOI22_X1 U13099 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10232) );
  AOI22_X1 U13100 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10231) );
  AOI22_X1 U13101 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10230) );
  NAND4_X1 U13102 ( .A1(n10233), .A2(n10232), .A3(n10231), .A4(n10230), .ZN(
        n10239) );
  AOI22_X1 U13103 ( .A1(n10891), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10856), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10237) );
  AOI22_X1 U13104 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10236) );
  AOI22_X1 U13105 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10235) );
  AOI22_X1 U13106 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10234) );
  NAND4_X1 U13107 ( .A1(n10237), .A2(n10236), .A3(n10235), .A4(n10234), .ZN(
        n10238) );
  NOR2_X1 U13108 ( .A1(n10239), .A2(n10238), .ZN(n10913) );
  NOR2_X1 U13109 ( .A1(n10912), .A2(n10913), .ZN(n10920) );
  AOI22_X1 U13110 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10243) );
  AOI22_X1 U13111 ( .A1(n10856), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10242) );
  AOI22_X1 U13112 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10241) );
  INV_X1 U13113 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n20874) );
  AOI22_X1 U13114 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10673), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10240) );
  NAND4_X1 U13115 ( .A1(n10243), .A2(n10242), .A3(n10241), .A4(n10240), .ZN(
        n10249) );
  AOI22_X1 U13116 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10352), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10247) );
  AOI22_X1 U13117 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10246) );
  AOI22_X1 U13118 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10245) );
  AOI22_X1 U13119 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10244) );
  NAND4_X1 U13120 ( .A1(n10247), .A2(n10246), .A3(n10245), .A4(n10244), .ZN(
        n10248) );
  OR2_X1 U13121 ( .A1(n10249), .A2(n10248), .ZN(n10921) );
  NAND2_X1 U13122 ( .A1(n10920), .A2(n10921), .ZN(n10929) );
  NOR2_X1 U13123 ( .A1(n10930), .A2(n10929), .ZN(n10937) );
  AOI22_X1 U13124 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10253) );
  AOI22_X1 U13125 ( .A1(n10313), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10252) );
  AOI22_X1 U13126 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10251) );
  AOI22_X1 U13127 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10673), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10250) );
  NAND4_X1 U13128 ( .A1(n10253), .A2(n10252), .A3(n10251), .A4(n10250), .ZN(
        n10259) );
  AOI22_X1 U13129 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10352), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10257) );
  AOI22_X1 U13130 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10869), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10256) );
  AOI22_X1 U13131 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10356), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U13132 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10254) );
  NAND4_X1 U13133 ( .A1(n10257), .A2(n10256), .A3(n10255), .A4(n10254), .ZN(
        n10258) );
  OR2_X1 U13134 ( .A1(n10259), .A2(n10258), .ZN(n10938) );
  NAND2_X1 U13135 ( .A1(n10937), .A2(n10938), .ZN(n10946) );
  NOR2_X1 U13136 ( .A1(n10947), .A2(n10946), .ZN(n10954) );
  INV_X1 U13137 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n20990) );
  AOI22_X1 U13138 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10263) );
  AOI22_X1 U13139 ( .A1(n10313), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10262) );
  AOI22_X1 U13140 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10261) );
  AOI22_X1 U13141 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10260) );
  NAND4_X1 U13142 ( .A1(n10263), .A2(n10262), .A3(n10261), .A4(n10260), .ZN(
        n10269) );
  AOI22_X1 U13143 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10851), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10267) );
  AOI22_X1 U13144 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10869), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10266) );
  AOI22_X1 U13145 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10356), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10265) );
  AOI22_X1 U13146 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10264) );
  NAND4_X1 U13147 ( .A1(n10267), .A2(n10266), .A3(n10265), .A4(n10264), .ZN(
        n10268) );
  OR2_X1 U13148 ( .A1(n10269), .A2(n10268), .ZN(n10955) );
  NAND2_X1 U13149 ( .A1(n10954), .A2(n10955), .ZN(n10963) );
  NOR2_X1 U13150 ( .A1(n10964), .A2(n10963), .ZN(n10281) );
  AOI22_X1 U13151 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10851), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10273) );
  AOI22_X1 U13152 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10272) );
  AOI22_X1 U13153 ( .A1(n10891), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10271) );
  AOI22_X1 U13154 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10356), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10270) );
  NAND4_X1 U13155 ( .A1(n10273), .A2(n10272), .A3(n10271), .A4(n10270), .ZN(
        n10279) );
  AOI22_X1 U13156 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10277) );
  AOI22_X1 U13157 ( .A1(n10313), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10811), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10276) );
  AOI22_X1 U13158 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10275) );
  AOI22_X1 U13159 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10869), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10274) );
  NAND4_X1 U13160 ( .A1(n10277), .A2(n10276), .A3(n10275), .A4(n10274), .ZN(
        n10278) );
  NOR2_X1 U13161 ( .A1(n10279), .A2(n10278), .ZN(n10280) );
  XNOR2_X1 U13162 ( .A(n10281), .B(n10280), .ZN(n10332) );
  NAND2_X1 U13163 ( .A1(n10313), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10285) );
  NAND2_X1 U13164 ( .A1(n10868), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10284) );
  NAND2_X1 U13165 ( .A1(n10302), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10283) );
  NAND2_X1 U13166 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10282) );
  NAND2_X1 U13167 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10289) );
  NAND2_X1 U13168 ( .A1(n10199), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10288) );
  NAND2_X1 U13169 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10287) );
  NAND2_X1 U13170 ( .A1(n10673), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10286) );
  NAND2_X1 U13171 ( .A1(n10353), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10293) );
  NAND2_X1 U13172 ( .A1(n10352), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10292) );
  NAND2_X1 U13173 ( .A1(n10322), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10291) );
  NAND2_X1 U13174 ( .A1(n10321), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10290) );
  NAND2_X1 U13175 ( .A1(n10320), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10297) );
  NAND2_X1 U13176 ( .A1(n10869), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10296) );
  NAND2_X1 U13177 ( .A1(n10398), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10295) );
  NAND2_X1 U13178 ( .A1(n10356), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10294) );
  NAND2_X1 U13179 ( .A1(n10391), .A2(n10389), .ZN(n10363) );
  INV_X1 U13180 ( .A(n10363), .ZN(n10330) );
  AOI22_X1 U13181 ( .A1(n10199), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10314), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U13182 ( .A1(n10353), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10321), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13183 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10356), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10303) );
  AOI22_X1 U13184 ( .A1(n10313), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10397), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10310) );
  AOI22_X1 U13185 ( .A1(n10673), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10398), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10308) );
  AOI22_X1 U13186 ( .A1(n10320), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10869), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10307) );
  AND4_X2 U13187 ( .A1(n10310), .A2(n10309), .A3(n10308), .A4(n10307), .ZN(
        n10311) );
  NAND2_X4 U13188 ( .A1(n10312), .A2(n10311), .ZN(n10388) );
  AOI22_X1 U13189 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10313), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U13190 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10673), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10318) );
  AOI22_X1 U13191 ( .A1(n10353), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10869), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U13192 ( .A1(n10398), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10356), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10316) );
  AOI22_X1 U13193 ( .A1(n10199), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10868), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U13194 ( .A1(n10302), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10397), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U13195 ( .A1(n10352), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10320), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U13196 ( .A1(n10322), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9743), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10323) );
  AND3_X2 U13197 ( .A1(n10327), .A2(n10326), .A3(n10325), .ZN(n10328) );
  INV_X1 U13198 ( .A(n10424), .ZN(n10329) );
  NAND2_X1 U13199 ( .A1(n10330), .A2(n10329), .ZN(n10364) );
  INV_X1 U13200 ( .A(n10331), .ZN(n15076) );
  NAND2_X1 U13201 ( .A1(n10332), .A2(n10956), .ZN(n10333) );
  NAND2_X1 U13202 ( .A1(n21125), .A2(n10388), .ZN(n10345) );
  AOI22_X1 U13203 ( .A1(n10199), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10314), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10338) );
  AOI22_X1 U13204 ( .A1(n10313), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10868), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10337) );
  AOI22_X1 U13205 ( .A1(n10302), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10397), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13206 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10673), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10335) );
  NAND4_X1 U13207 ( .A1(n10338), .A2(n10337), .A3(n10336), .A4(n10335), .ZN(
        n10344) );
  AOI22_X1 U13208 ( .A1(n10353), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10352), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10342) );
  AOI22_X1 U13209 ( .A1(n10320), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10869), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10341) );
  AOI22_X1 U13210 ( .A1(n10398), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10356), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10340) );
  AOI22_X1 U13211 ( .A1(n10322), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10321), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10339) );
  NAND4_X1 U13212 ( .A1(n10342), .A2(n10341), .A3(n10340), .A4(n10339), .ZN(
        n10343) );
  OR2_X2 U13213 ( .A1(n10344), .A2(n10343), .ZN(n10423) );
  NAND2_X1 U13214 ( .A1(n10345), .A2(n10387), .ZN(n10347) );
  INV_X2 U13215 ( .A(n10391), .ZN(n10421) );
  NAND2_X2 U13216 ( .A1(n10388), .A2(n10421), .ZN(n10422) );
  NAND2_X1 U13217 ( .A1(n10347), .A2(n10346), .ZN(n10366) );
  AOI22_X1 U13218 ( .A1(n10199), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10314), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10351) );
  AOI22_X1 U13219 ( .A1(n10313), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10868), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U13220 ( .A1(n10302), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10397), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U13221 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10673), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10348) );
  NAND4_X1 U13222 ( .A1(n10351), .A2(n10350), .A3(n10349), .A4(n10348), .ZN(
        n10362) );
  NAND2_X1 U13223 ( .A1(n10352), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10355) );
  AOI22_X1 U13224 ( .A1(n10320), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10869), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10359) );
  AOI22_X1 U13225 ( .A1(n10398), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10356), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10358) );
  NAND4_X1 U13226 ( .A1(n10360), .A2(n10359), .A3(n10358), .A4(n10357), .ZN(
        n10361) );
  NAND2_X1 U13227 ( .A1(n21125), .A2(n10389), .ZN(n10416) );
  AOI22_X1 U13228 ( .A1(n10364), .A2(n20157), .B1(n10416), .B2(n10363), .ZN(
        n10365) );
  INV_X1 U13229 ( .A(n10422), .ZN(n11074) );
  NAND2_X1 U13230 ( .A1(n10673), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10374) );
  NAND2_X1 U13231 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10373) );
  NAND2_X1 U13232 ( .A1(n10199), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10372) );
  NAND2_X1 U13233 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10371) );
  NAND2_X1 U13234 ( .A1(n10353), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10378) );
  NAND2_X1 U13235 ( .A1(n10352), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10377) );
  NAND2_X1 U13236 ( .A1(n10322), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10376) );
  NAND2_X1 U13237 ( .A1(n10321), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10375) );
  NAND2_X1 U13238 ( .A1(n10320), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10382) );
  NAND2_X1 U13239 ( .A1(n10869), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10381) );
  NAND2_X1 U13240 ( .A1(n10398), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10380) );
  NAND2_X1 U13241 ( .A1(n10356), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10379) );
  NAND4_X4 U13242 ( .A1(n10386), .A2(n10385), .A3(n10384), .A4(n10383), .ZN(
        n20135) );
  AND2_X2 U13243 ( .A1(n10387), .A2(n20157), .ZN(n10419) );
  AND2_X2 U13244 ( .A1(n11149), .A2(n10389), .ZN(n13061) );
  NAND3_X1 U13245 ( .A1(n10419), .A2(n13061), .A3(n10392), .ZN(n11144) );
  NAND2_X1 U13246 ( .A1(n10199), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10396) );
  NAND2_X1 U13247 ( .A1(n10868), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10395) );
  NAND2_X1 U13248 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10394) );
  NAND2_X1 U13249 ( .A1(n10673), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10393) );
  NAND2_X1 U13250 ( .A1(n10313), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10402) );
  NAND2_X1 U13251 ( .A1(n10302), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10401) );
  NAND2_X1 U13252 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10400) );
  NAND2_X1 U13253 ( .A1(n10398), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10399) );
  NAND2_X1 U13254 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10406) );
  NAND2_X1 U13255 ( .A1(n10320), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10405) );
  NAND2_X1 U13256 ( .A1(n10322), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10404) );
  NAND2_X1 U13257 ( .A1(n10321), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10403) );
  NAND2_X1 U13258 ( .A1(n10353), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10410) );
  NAND2_X1 U13259 ( .A1(n10352), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10409) );
  NAND2_X1 U13260 ( .A1(n10356), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10408) );
  NAND2_X1 U13261 ( .A1(n10869), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10407) );
  NAND4_X4 U13262 ( .A1(n10414), .A2(n10413), .A3(n10412), .A4(n10411), .ZN(
        n10447) );
  NAND2_X2 U13263 ( .A1(n13165), .A2(n20135), .ZN(n13166) );
  XNOR2_X1 U13264 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12915) );
  NOR2_X2 U13266 ( .A1(n10429), .A2(n20135), .ZN(n11141) );
  NAND3_X1 U13267 ( .A1(n11141), .A2(n13062), .A3(n11146), .ZN(n13167) );
  OAI21_X1 U13268 ( .B1(n12868), .B2(n12915), .A(n13167), .ZN(n10417) );
  INV_X1 U13269 ( .A(n10417), .ZN(n10418) );
  NAND2_X1 U13270 ( .A1(n13155), .A2(n10418), .ZN(n10438) );
  NAND2_X1 U13271 ( .A1(n10415), .A2(n20135), .ZN(n11162) );
  INV_X1 U13272 ( .A(n11073), .ZN(n10420) );
  NAND2_X1 U13273 ( .A1(n10423), .A2(n20135), .ZN(n11137) );
  OAI211_X1 U13274 ( .C1(n13166), .C2(n10421), .A(n13160), .B(n11137), .ZN(
        n10446) );
  OR2_X1 U13275 ( .A1(n10424), .A2(n20161), .ZN(n10426) );
  NAND2_X1 U13276 ( .A1(n21125), .A2(n11149), .ZN(n10425) );
  NAND2_X1 U13277 ( .A1(n11071), .A2(n10421), .ZN(n13143) );
  NAND2_X1 U13278 ( .A1(n10427), .A2(n10454), .ZN(n10428) );
  NAND2_X1 U13279 ( .A1(n10429), .A2(n13165), .ZN(n10432) );
  INV_X1 U13280 ( .A(n10562), .ZN(n10431) );
  NAND2_X1 U13281 ( .A1(n10463), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10437) );
  NAND2_X1 U13282 ( .A1(n16255), .A2(n20815), .ZN(n11129) );
  NAND2_X1 U13283 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10461) );
  OAI21_X1 U13284 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n10461), .ZN(n20466) );
  NAND2_X1 U13285 ( .A1(n20714), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16052) );
  NAND2_X1 U13286 ( .A1(n16052), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10456) );
  OAI21_X1 U13287 ( .B1(n11129), .B2(n20466), .A(n10456), .ZN(n10435) );
  INV_X1 U13288 ( .A(n10435), .ZN(n10436) );
  XNOR2_X2 U13289 ( .A(n10439), .B(n10458), .ZN(n10530) );
  NAND2_X1 U13290 ( .A1(n10463), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10442) );
  INV_X1 U13291 ( .A(n16052), .ZN(n10440) );
  MUX2_X1 U13292 ( .A(n10440), .B(n11129), .S(n20573), .Z(n10441) );
  INV_X1 U13293 ( .A(n13166), .ZN(n20813) );
  INV_X1 U13294 ( .A(n10443), .ZN(n10445) );
  NAND3_X1 U13295 ( .A1(n13583), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n16255), 
        .ZN(n10444) );
  AOI21_X1 U13296 ( .B1(n20813), .B2(n10445), .A(n10444), .ZN(n10452) );
  INV_X1 U13297 ( .A(n10446), .ZN(n10451) );
  INV_X1 U13298 ( .A(n13055), .ZN(n13579) );
  NAND2_X1 U13299 ( .A1(n10424), .A2(n20157), .ZN(n10448) );
  NAND2_X1 U13300 ( .A1(n12873), .A2(n10448), .ZN(n10450) );
  NAND2_X1 U13301 ( .A1(n11141), .A2(n9733), .ZN(n13159) );
  NAND2_X1 U13302 ( .A1(n9781), .A2(n13055), .ZN(n13185) );
  OAI211_X1 U13303 ( .C1(n10454), .C2(n13165), .A(n10453), .B(n13185), .ZN(
        n10480) );
  AND2_X1 U13304 ( .A1(n10456), .A2(n10455), .ZN(n10457) );
  INV_X1 U13305 ( .A(n10461), .ZN(n10460) );
  NAND2_X1 U13306 ( .A1(n10460), .A2(n20459), .ZN(n20511) );
  NAND2_X1 U13307 ( .A1(n10461), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10462) );
  NAND2_X1 U13308 ( .A1(n10463), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10465) );
  NAND2_X1 U13309 ( .A1(n16052), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10464) );
  AOI22_X1 U13310 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10470) );
  AOI22_X1 U13311 ( .A1(n10856), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10469) );
  AOI22_X1 U13312 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10468) );
  AOI22_X1 U13313 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10467) );
  NAND4_X1 U13314 ( .A1(n10470), .A2(n10469), .A3(n10468), .A4(n10467), .ZN(
        n10476) );
  AOI22_X1 U13315 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10851), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10474) );
  AOI22_X1 U13316 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10869), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10473) );
  AOI22_X1 U13317 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U13318 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10471) );
  NAND4_X1 U13319 ( .A1(n10474), .A2(n10473), .A3(n10472), .A4(n10471), .ZN(
        n10475) );
  INV_X1 U13320 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10477) );
  OAI22_X1 U13321 ( .A1(n10562), .A2(n10979), .B1(n11109), .B2(n10477), .ZN(
        n10478) );
  XNOR2_X1 U13322 ( .A(n10479), .B(n10478), .ZN(n10538) );
  INV_X1 U13323 ( .A(n10538), .ZN(n10537) );
  INV_X1 U13324 ( .A(n10480), .ZN(n10481) );
  AOI22_X1 U13325 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10900), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13326 ( .A1(n10891), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10811), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13327 ( .A1(n10353), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10322), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U13328 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10483) );
  NAND4_X1 U13329 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n10483), .ZN(
        n10492) );
  AOI22_X1 U13330 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13331 ( .A1(n10856), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U13332 ( .A1(n10869), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13333 ( .A1(n10398), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10356), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10487) );
  NAND4_X1 U13334 ( .A1(n10490), .A2(n10489), .A3(n10488), .A4(n10487), .ZN(
        n10491) );
  INV_X1 U13335 ( .A(n11044), .ZN(n10503) );
  AOI22_X1 U13336 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10496) );
  AOI22_X1 U13337 ( .A1(n10891), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10495) );
  AOI22_X1 U13338 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10494) );
  AOI22_X1 U13339 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10493) );
  NAND4_X1 U13340 ( .A1(n10496), .A2(n10495), .A3(n10494), .A4(n10493), .ZN(
        n10502) );
  AOI22_X1 U13341 ( .A1(n10353), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10322), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U13342 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10900), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U13343 ( .A1(n10856), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10498) );
  AOI22_X1 U13344 ( .A1(n10869), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10356), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10497) );
  NAND4_X1 U13345 ( .A1(n10500), .A2(n10499), .A3(n10498), .A4(n10497), .ZN(
        n10501) );
  XNOR2_X1 U13346 ( .A(n10503), .B(n10990), .ZN(n10504) );
  INV_X1 U13347 ( .A(n10561), .ZN(n10975) );
  NAND2_X1 U13348 ( .A1(n10504), .A2(n10975), .ZN(n10505) );
  INV_X1 U13349 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10508) );
  AOI21_X1 U13350 ( .B1(n10421), .B2(n11044), .A(n20815), .ZN(n10507) );
  NAND2_X1 U13351 ( .A1(n10430), .A2(n10990), .ZN(n10506) );
  OAI211_X1 U13352 ( .C1(n11109), .C2(n10508), .A(n10507), .B(n10506), .ZN(
        n10551) );
  NAND2_X1 U13353 ( .A1(n10975), .A2(n11044), .ZN(n10524) );
  NAND2_X1 U13354 ( .A1(n10527), .A2(n10524), .ZN(n10522) );
  AOI22_X1 U13355 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10512) );
  AOI22_X1 U13356 ( .A1(n10891), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10856), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10511) );
  AOI22_X1 U13357 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10322), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10510) );
  AOI22_X1 U13358 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10869), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10509) );
  NAND4_X1 U13359 ( .A1(n10512), .A2(n10511), .A3(n10510), .A4(n10509), .ZN(
        n10518) );
  AOI22_X1 U13360 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10516) );
  AOI22_X1 U13361 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U13362 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U13363 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10513) );
  NAND4_X1 U13364 ( .A1(n10516), .A2(n10515), .A3(n10514), .A4(n10513), .ZN(
        n10517) );
  INV_X1 U13365 ( .A(n10989), .ZN(n10519) );
  OR2_X1 U13366 ( .A1(n10562), .A2(n10519), .ZN(n10521) );
  NAND2_X1 U13367 ( .A1(n11115), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10520) );
  OAI211_X1 U13368 ( .C1(n10561), .C2(n11044), .A(n10521), .B(n10520), .ZN(
        n10523) );
  NAND2_X1 U13369 ( .A1(n10522), .A2(n10523), .ZN(n10528) );
  INV_X1 U13370 ( .A(n10523), .ZN(n10525) );
  INV_X1 U13371 ( .A(n10530), .ZN(n20245) );
  NAND2_X1 U13372 ( .A1(n10975), .A2(n10989), .ZN(n10532) );
  NAND2_X1 U13373 ( .A1(n10546), .A2(n10535), .ZN(n10539) );
  INV_X1 U13374 ( .A(n10539), .ZN(n10536) );
  NAND2_X1 U13375 ( .A1(n9728), .A2(n10539), .ZN(n10540) );
  NAND2_X1 U13376 ( .A1(n10584), .A2(n10540), .ZN(n10977) );
  NAND2_X1 U13377 ( .A1(n13062), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10604) );
  NAND2_X1 U13378 ( .A1(n14068), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n10542) );
  OAI21_X1 U13379 ( .B1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n10576), .ZN(n14584) );
  OAI21_X1 U13380 ( .B1(n14584), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20811), 
        .ZN(n10541) );
  OAI211_X1 U13381 ( .C1(n10604), .C2(n10094), .A(n10542), .B(n10541), .ZN(
        n10543) );
  INV_X1 U13382 ( .A(n10543), .ZN(n10544) );
  NAND2_X1 U13383 ( .A1(n14067), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10556) );
  NAND2_X1 U13384 ( .A1(n14068), .A2(P1_EAX_REG_1__SCAN_IN), .ZN(n10549) );
  NAND2_X1 U13385 ( .A1(n20811), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10548) );
  OAI211_X1 U13386 ( .C1(n10604), .C2(n10455), .A(n10549), .B(n10548), .ZN(
        n10550) );
  AOI21_X1 U13387 ( .B1(n20207), .B2(n9733), .A(n20811), .ZN(n13014) );
  NAND2_X1 U13388 ( .A1(n10552), .A2(n10797), .ZN(n10554) );
  AOI22_X1 U13389 ( .A1(n14068), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20811), .ZN(n10553) );
  OAI211_X1 U13390 ( .C1(n10604), .C2(n10173), .A(n10554), .B(n10553), .ZN(
        n13013) );
  MUX2_X1 U13391 ( .A(n10960), .B(n13014), .S(n13013), .Z(n13063) );
  NAND2_X1 U13392 ( .A1(n9822), .A2(n10555), .ZN(n13133) );
  NAND2_X1 U13393 ( .A1(n10463), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10560) );
  INV_X1 U13394 ( .A(n11129), .ZN(n10558) );
  NOR3_X1 U13395 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20459), .A3(
        n20541), .ZN(n20381) );
  NAND2_X1 U13396 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20381), .ZN(
        n20375) );
  NAND2_X1 U13397 ( .A1(n21022), .A2(n20375), .ZN(n10557) );
  NAND3_X1 U13398 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20652) );
  INV_X1 U13399 ( .A(n20652), .ZN(n20662) );
  NAND2_X1 U13400 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20662), .ZN(
        n20649) );
  AOI22_X1 U13401 ( .A1(n10558), .A2(n20407), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16052), .ZN(n10559) );
  AOI22_X1 U13402 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U13403 ( .A1(n10856), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10565) );
  AOI22_X1 U13404 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10564) );
  AOI22_X1 U13405 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10563) );
  NAND4_X1 U13406 ( .A1(n10566), .A2(n10565), .A3(n10564), .A4(n10563), .ZN(
        n10572) );
  AOI22_X1 U13407 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10851), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10570) );
  AOI22_X1 U13408 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U13409 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U13410 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10567) );
  NAND4_X1 U13411 ( .A1(n10570), .A2(n10569), .A3(n10568), .A4(n10567), .ZN(
        n10571) );
  AOI22_X1 U13412 ( .A1(n11089), .A2(n11001), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n11115), .ZN(n10573) );
  NAND2_X1 U13413 ( .A1(n10999), .A2(n10797), .ZN(n10583) );
  NAND2_X1 U13414 ( .A1(n10965), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n10580) );
  INV_X1 U13415 ( .A(n10605), .ZN(n10578) );
  INV_X1 U13416 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14573) );
  NAND2_X1 U13417 ( .A1(n14573), .A2(n10576), .ZN(n10577) );
  NAND2_X1 U13418 ( .A1(n10578), .A2(n10577), .ZN(n14572) );
  AOI22_X1 U13419 ( .A1(n14572), .A2(n10960), .B1(n14067), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10579) );
  OAI211_X1 U13420 ( .C1(n10604), .C2(n10575), .A(n10580), .B(n10579), .ZN(
        n10581) );
  INV_X1 U13421 ( .A(n10581), .ZN(n10582) );
  NAND2_X1 U13422 ( .A1(n10583), .A2(n10582), .ZN(n13258) );
  NAND2_X1 U13423 ( .A1(n13256), .A2(n13258), .ZN(n13257) );
  NOR2_X2 U13424 ( .A1(n10584), .A2(n15065), .ZN(n10597) );
  AOI22_X1 U13425 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10876), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10588) );
  AOI22_X1 U13426 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10890), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10587) );
  AOI22_X1 U13427 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10806), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10586) );
  AOI22_X1 U13428 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10585) );
  NAND4_X1 U13429 ( .A1(n10588), .A2(n10587), .A3(n10586), .A4(n10585), .ZN(
        n10594) );
  AOI22_X1 U13430 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10811), .B1(
        n10856), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10592) );
  AOI22_X1 U13431 ( .A1(n10891), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10591) );
  AOI22_X1 U13432 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10590) );
  AOI22_X1 U13433 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n10900), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10589) );
  NAND4_X1 U13434 ( .A1(n10592), .A2(n10591), .A3(n10590), .A4(n10589), .ZN(
        n10593) );
  NAND2_X1 U13435 ( .A1(n11089), .A2(n11015), .ZN(n10596) );
  NAND2_X1 U13436 ( .A1(n11115), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10595) );
  NAND2_X1 U13437 ( .A1(n10596), .A2(n10595), .ZN(n10598) );
  INV_X1 U13438 ( .A(n10597), .ZN(n10599) );
  NAND2_X1 U13439 ( .A1(n10599), .A2(n9874), .ZN(n10600) );
  AND2_X1 U13440 ( .A1(n10620), .A2(n10600), .ZN(n11007) );
  INV_X1 U13441 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n10603) );
  NAND2_X1 U13442 ( .A1(n10965), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n10602) );
  NAND2_X1 U13443 ( .A1(n20811), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10601) );
  OAI211_X1 U13444 ( .C1(n10604), .C2(n10603), .A(n10602), .B(n10601), .ZN(
        n10606) );
  OAI21_X1 U13445 ( .B1(n10605), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n10623), .ZN(n20035) );
  MUX2_X1 U13446 ( .A(n10606), .B(n20035), .S(n10960), .Z(n10607) );
  NAND2_X1 U13447 ( .A1(n9735), .A2(n10608), .ZN(n13411) );
  AOI22_X1 U13448 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10612) );
  AOI22_X1 U13449 ( .A1(n10856), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10611) );
  INV_X1 U13450 ( .A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n21039) );
  AOI22_X1 U13451 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10610) );
  AOI22_X1 U13452 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10609) );
  NAND4_X1 U13453 ( .A1(n10612), .A2(n10611), .A3(n10610), .A4(n10609), .ZN(
        n10618) );
  AOI22_X1 U13454 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10851), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10616) );
  AOI22_X1 U13455 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U13456 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10614) );
  AOI22_X1 U13457 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10613) );
  NAND4_X1 U13458 ( .A1(n10616), .A2(n10615), .A3(n10614), .A4(n10613), .ZN(
        n10617) );
  AOI22_X1 U13459 ( .A1(n11089), .A2(n11018), .B1(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .B2(n11115), .ZN(n10619) );
  NAND2_X1 U13460 ( .A1(n10620), .A2(n10619), .ZN(n10621) );
  NAND2_X1 U13461 ( .A1(n10645), .A2(n10621), .ZN(n11014) );
  INV_X1 U13462 ( .A(n11014), .ZN(n10622) );
  INV_X1 U13463 ( .A(n14067), .ZN(n10706) );
  AND2_X1 U13464 ( .A1(n10623), .A2(n10626), .ZN(n10624) );
  OR2_X1 U13465 ( .A1(n10624), .A2(n10640), .ZN(n20029) );
  NAND2_X1 U13466 ( .A1(n20029), .A2(n10960), .ZN(n10625) );
  OAI21_X1 U13467 ( .B1(n10626), .B2(n10706), .A(n10625), .ZN(n10627) );
  AOI21_X1 U13468 ( .B1(n10965), .B2(P1_EAX_REG_5__SCAN_IN), .A(n10627), .ZN(
        n10628) );
  INV_X1 U13469 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n10644) );
  AOI22_X1 U13470 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10633) );
  AOI22_X1 U13471 ( .A1(n10856), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10811), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10632) );
  AOI22_X1 U13472 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10631) );
  AOI22_X1 U13473 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10877), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10630) );
  NAND4_X1 U13474 ( .A1(n10633), .A2(n10632), .A3(n10631), .A4(n10630), .ZN(
        n10639) );
  AOI22_X1 U13475 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10900), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10637) );
  AOI22_X1 U13476 ( .A1(n10891), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10636) );
  AOI22_X1 U13477 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10635) );
  AOI22_X1 U13478 ( .A1(n10892), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10634) );
  NAND4_X1 U13479 ( .A1(n10637), .A2(n10636), .A3(n10635), .A4(n10634), .ZN(
        n10638) );
  AOI22_X1 U13480 ( .A1(n11089), .A2(n11034), .B1(n11115), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10646) );
  NAND2_X1 U13481 ( .A1(n10645), .A2(n10646), .ZN(n11024) );
  NAND2_X1 U13482 ( .A1(n11024), .A2(n10797), .ZN(n10643) );
  NOR2_X1 U13483 ( .A1(n10640), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10641) );
  OR2_X1 U13484 ( .A1(n10652), .A2(n10641), .ZN(n20012) );
  AOI22_X1 U13485 ( .A1(n20012), .A2(n10960), .B1(n14067), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10642) );
  NAND2_X1 U13486 ( .A1(n13413), .A2(n13506), .ZN(n13507) );
  INV_X1 U13487 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10650) );
  NAND2_X1 U13488 ( .A1(n11089), .A2(n11044), .ZN(n10649) );
  OAI21_X1 U13489 ( .B1(n10650), .B2(n11109), .A(n10649), .ZN(n10651) );
  INV_X1 U13490 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n10656) );
  NOR2_X1 U13491 ( .A1(n10652), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10653) );
  OR2_X1 U13492 ( .A1(n10668), .A2(n10653), .ZN(n20002) );
  INV_X1 U13493 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19998) );
  NOR2_X1 U13494 ( .A1(n10706), .A2(n19998), .ZN(n10654) );
  AOI21_X1 U13495 ( .B1(n20002), .B2(n10960), .A(n10654), .ZN(n10655) );
  OAI21_X1 U13496 ( .B1(n10886), .B2(n10656), .A(n10655), .ZN(n10657) );
  NOR2_X2 U13497 ( .A1(n13507), .A2(n13604), .ZN(n13605) );
  AOI22_X1 U13498 ( .A1(n10856), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10661) );
  AOI22_X1 U13499 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10806), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10660) );
  AOI22_X1 U13500 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10877), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10659) );
  AOI22_X1 U13501 ( .A1(n10869), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10658) );
  NAND4_X1 U13502 ( .A1(n10661), .A2(n10660), .A3(n10659), .A4(n10658), .ZN(
        n10667) );
  AOI22_X1 U13503 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10665) );
  AOI22_X1 U13504 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10664) );
  AOI22_X1 U13505 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10663) );
  AOI22_X1 U13506 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10662) );
  NAND4_X1 U13507 ( .A1(n10665), .A2(n10664), .A3(n10663), .A4(n10662), .ZN(
        n10666) );
  OAI21_X1 U13508 ( .B1(n10667), .B2(n10666), .A(n10797), .ZN(n10671) );
  XOR2_X1 U13509 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n10668), .Z(n19986) );
  INV_X1 U13510 ( .A(n19986), .ZN(n13808) );
  AOI22_X1 U13511 ( .A1(n14067), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n10960), .B2(n13808), .ZN(n10670) );
  NAND2_X1 U13512 ( .A1(n10965), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n10669) );
  AOI22_X1 U13513 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10900), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10677) );
  AOI22_X1 U13514 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10676) );
  AOI22_X1 U13515 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10675) );
  AOI22_X1 U13516 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10674) );
  NAND4_X1 U13517 ( .A1(n10677), .A2(n10676), .A3(n10675), .A4(n10674), .ZN(
        n10683) );
  AOI22_X1 U13518 ( .A1(n10891), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10856), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U13519 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U13520 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U13521 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10678) );
  NAND4_X1 U13522 ( .A1(n10681), .A2(n10680), .A3(n10679), .A4(n10678), .ZN(
        n10682) );
  OAI21_X1 U13523 ( .B1(n10683), .B2(n10682), .A(n10797), .ZN(n10688) );
  NAND2_X1 U13524 ( .A1(n10965), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n10687) );
  INV_X1 U13525 ( .A(n10684), .ZN(n10685) );
  XNOR2_X1 U13526 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n10685), .ZN(
        n13947) );
  AOI22_X1 U13527 ( .A1(n10960), .A2(n13947), .B1(n14067), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10686) );
  XOR2_X1 U13528 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B(n10689), .Z(
        n16150) );
  AOI22_X1 U13529 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10900), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U13530 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10811), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U13531 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10691) );
  AOI22_X1 U13532 ( .A1(n10869), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10690) );
  NAND4_X1 U13533 ( .A1(n10693), .A2(n10692), .A3(n10691), .A4(n10690), .ZN(
        n10699) );
  AOI22_X1 U13534 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10697) );
  AOI22_X1 U13535 ( .A1(n10856), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10696) );
  AOI22_X1 U13536 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10695) );
  AOI22_X1 U13537 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10877), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10694) );
  NAND4_X1 U13538 ( .A1(n10697), .A2(n10696), .A3(n10695), .A4(n10694), .ZN(
        n10698) );
  OR2_X1 U13539 ( .A1(n10699), .A2(n10698), .ZN(n10700) );
  AOI22_X1 U13540 ( .A1(n10797), .A2(n10700), .B1(n14067), .B2(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10702) );
  NAND2_X1 U13541 ( .A1(n10965), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n10701) );
  OAI211_X1 U13542 ( .C1(n16150), .C2(n10971), .A(n10702), .B(n10701), .ZN(
        n13820) );
  NAND2_X1 U13543 ( .A1(n10703), .A2(n13972), .ZN(n10705) );
  INV_X1 U13544 ( .A(n10748), .ZN(n10704) );
  NAND2_X1 U13545 ( .A1(n10705), .A2(n10704), .ZN(n14878) );
  NAND2_X1 U13546 ( .A1(n14878), .A2(n10960), .ZN(n10709) );
  NOR2_X1 U13547 ( .A1(n10706), .A2(n13972), .ZN(n10707) );
  AOI21_X1 U13548 ( .B1(n10965), .B2(P1_EAX_REG_11__SCAN_IN), .A(n10707), .ZN(
        n10708) );
  NAND2_X1 U13549 ( .A1(n10709), .A2(n10708), .ZN(n10721) );
  AOI22_X1 U13550 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10713) );
  AOI22_X1 U13551 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10856), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13552 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13553 ( .A1(n9723), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10710) );
  NAND4_X1 U13554 ( .A1(n10713), .A2(n10712), .A3(n10711), .A4(n10710), .ZN(
        n10719) );
  AOI22_X1 U13555 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10811), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U13556 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10806), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13557 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10715) );
  AOI22_X1 U13558 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10714) );
  NAND4_X1 U13559 ( .A1(n10717), .A2(n10716), .A3(n10715), .A4(n10714), .ZN(
        n10718) );
  OR2_X1 U13560 ( .A1(n10719), .A2(n10718), .ZN(n10720) );
  AND2_X1 U13561 ( .A1(n10797), .A2(n10720), .ZN(n13954) );
  NAND2_X1 U13562 ( .A1(n13952), .A2(n13954), .ZN(n13953) );
  INV_X1 U13563 ( .A(n10721), .ZN(n10722) );
  XNOR2_X1 U13564 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n10724), .ZN(
        n16089) );
  AOI22_X1 U13565 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10900), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10728) );
  AOI22_X1 U13566 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10727) );
  AOI22_X1 U13567 ( .A1(n10891), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U13568 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10725) );
  NAND4_X1 U13569 ( .A1(n10728), .A2(n10727), .A3(n10726), .A4(n10725), .ZN(
        n10734) );
  AOI22_X1 U13570 ( .A1(n10856), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10811), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10732) );
  AOI22_X1 U13571 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U13572 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10877), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10730) );
  AOI22_X1 U13573 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10729) );
  NAND4_X1 U13574 ( .A1(n10732), .A2(n10731), .A3(n10730), .A4(n10729), .ZN(
        n10733) );
  OR2_X1 U13575 ( .A1(n10734), .A2(n10733), .ZN(n10735) );
  AOI22_X1 U13576 ( .A1(n10797), .A2(n10735), .B1(n14067), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10737) );
  NAND2_X1 U13577 ( .A1(n10965), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n10736) );
  OAI211_X1 U13578 ( .C1(n16089), .C2(n10971), .A(n10737), .B(n10736), .ZN(
        n14630) );
  AOI22_X1 U13579 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10856), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10741) );
  AOI22_X1 U13580 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n9723), .B1(
        n10811), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10740) );
  AOI22_X1 U13581 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10806), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10739) );
  AOI22_X1 U13582 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10892), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10738) );
  NAND4_X1 U13583 ( .A1(n10741), .A2(n10740), .A3(n10739), .A4(n10738), .ZN(
        n10747) );
  AOI22_X1 U13584 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10876), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10745) );
  AOI22_X1 U13585 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U13586 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10870), .B1(
        n10877), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10743) );
  AOI22_X1 U13587 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10742) );
  NAND4_X1 U13588 ( .A1(n10745), .A2(n10744), .A3(n10743), .A4(n10742), .ZN(
        n10746) );
  NOR2_X1 U13589 ( .A1(n10747), .A2(n10746), .ZN(n10751) );
  XNOR2_X1 U13590 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n10748), .ZN(
        n16102) );
  AOI22_X1 U13591 ( .A1(n10960), .A2(n16102), .B1(n14067), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10750) );
  NAND2_X1 U13592 ( .A1(n10965), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n10749) );
  OAI211_X1 U13593 ( .C1(n10104), .C2(n10751), .A(n10750), .B(n10749), .ZN(
        n14710) );
  AND2_X1 U13594 ( .A1(n14630), .A2(n14710), .ZN(n10752) );
  NAND2_X1 U13595 ( .A1(n10753), .A2(n20875), .ZN(n10755) );
  INV_X1 U13596 ( .A(n10788), .ZN(n10754) );
  NAND2_X1 U13597 ( .A1(n10755), .A2(n10754), .ZN(n14857) );
  AOI22_X1 U13598 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10759) );
  AOI22_X1 U13599 ( .A1(n10856), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U13600 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10757) );
  AOI22_X1 U13601 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10756) );
  NAND4_X1 U13602 ( .A1(n10759), .A2(n10758), .A3(n10757), .A4(n10756), .ZN(
        n10765) );
  AOI22_X1 U13603 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10900), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10763) );
  AOI22_X1 U13604 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U13605 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10761) );
  AOI22_X1 U13606 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10760) );
  NAND4_X1 U13607 ( .A1(n10763), .A2(n10762), .A3(n10761), .A4(n10760), .ZN(
        n10764) );
  OAI21_X1 U13608 ( .B1(n10765), .B2(n10764), .A(n10797), .ZN(n10768) );
  NAND2_X1 U13609 ( .A1(n10965), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n10767) );
  NAND2_X1 U13610 ( .A1(n14067), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10766) );
  NAND3_X1 U13611 ( .A1(n10768), .A2(n10767), .A3(n10766), .ZN(n10769) );
  AOI21_X1 U13612 ( .B1(n14857), .B2(n10960), .A(n10769), .ZN(n14559) );
  INV_X1 U13613 ( .A(n14559), .ZN(n10770) );
  AOI22_X1 U13614 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13615 ( .A1(n10856), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U13616 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10806), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U13617 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10771) );
  NAND4_X1 U13618 ( .A1(n10774), .A2(n10773), .A3(n10772), .A4(n10771), .ZN(
        n10780) );
  AOI22_X1 U13619 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10778) );
  AOI22_X1 U13620 ( .A1(n10891), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10777) );
  AOI22_X1 U13621 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10776) );
  AOI22_X1 U13622 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10775) );
  NAND4_X1 U13623 ( .A1(n10778), .A2(n10777), .A3(n10776), .A4(n10775), .ZN(
        n10779) );
  NOR2_X1 U13624 ( .A1(n10780), .A2(n10779), .ZN(n10784) );
  NAND2_X1 U13625 ( .A1(n20811), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10781) );
  NAND2_X1 U13626 ( .A1(n10971), .A2(n10781), .ZN(n10782) );
  AOI21_X1 U13627 ( .B1(n10965), .B2(P1_EAX_REG_16__SCAN_IN), .A(n10782), .ZN(
        n10783) );
  OAI21_X1 U13628 ( .B1(n10968), .B2(n10784), .A(n10783), .ZN(n10787) );
  XNOR2_X1 U13629 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B(n10785), .ZN(
        n14828) );
  NAND2_X1 U13630 ( .A1(n10960), .A2(n14828), .ZN(n10786) );
  NAND2_X1 U13631 ( .A1(n10787), .A2(n10786), .ZN(n14536) );
  INV_X1 U13632 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14550) );
  XNOR2_X1 U13633 ( .A(n14550), .B(n10788), .ZN(n14846) );
  INV_X1 U13634 ( .A(n14846), .ZN(n10804) );
  AOI22_X1 U13635 ( .A1(n10856), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10792) );
  AOI22_X1 U13636 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10791) );
  AOI22_X1 U13637 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10790) );
  AOI22_X1 U13638 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10789) );
  NAND4_X1 U13639 ( .A1(n10792), .A2(n10791), .A3(n10790), .A4(n10789), .ZN(
        n10799) );
  AOI22_X1 U13640 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10851), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10796) );
  AOI22_X1 U13641 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10795) );
  AOI22_X1 U13642 ( .A1(n10891), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10794) );
  AOI22_X1 U13643 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10793) );
  NAND4_X1 U13644 ( .A1(n10796), .A2(n10795), .A3(n10794), .A4(n10793), .ZN(
        n10798) );
  OAI21_X1 U13645 ( .B1(n10799), .B2(n10798), .A(n10797), .ZN(n10802) );
  NAND2_X1 U13646 ( .A1(n10965), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n10801) );
  NAND2_X1 U13647 ( .A1(n14067), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10800) );
  NAND3_X1 U13648 ( .A1(n10802), .A2(n10801), .A3(n10800), .ZN(n10803) );
  AOI21_X1 U13649 ( .B1(n10804), .B2(n10960), .A(n10803), .ZN(n14546) );
  XOR2_X1 U13650 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n10805), .Z(
        n16136) );
  AOI22_X1 U13651 ( .A1(n10965), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n14067), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10819) );
  AOI22_X1 U13652 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10810) );
  AOI22_X1 U13653 ( .A1(n10352), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10806), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U13654 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10869), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U13655 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10807) );
  NAND4_X1 U13656 ( .A1(n10810), .A2(n10809), .A3(n10808), .A4(n10807), .ZN(
        n10817) );
  AOI22_X1 U13657 ( .A1(n10856), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10815) );
  AOI22_X1 U13658 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U13659 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10813) );
  AOI22_X1 U13660 ( .A1(n10892), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10877), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10812) );
  NAND4_X1 U13661 ( .A1(n10815), .A2(n10814), .A3(n10813), .A4(n10812), .ZN(
        n10816) );
  OAI21_X1 U13662 ( .B1(n10817), .B2(n10816), .A(n10956), .ZN(n10818) );
  OAI211_X1 U13663 ( .C1(n16136), .C2(n10971), .A(n10819), .B(n10818), .ZN(
        n14611) );
  XNOR2_X1 U13664 ( .A(n10820), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14820) );
  AOI21_X1 U13665 ( .B1(n10167), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10821) );
  AOI21_X1 U13666 ( .B1(n10965), .B2(P1_EAX_REG_18__SCAN_IN), .A(n10821), .ZN(
        n10833) );
  AOI22_X1 U13667 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10352), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10825) );
  AOI22_X1 U13668 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10869), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U13669 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U13670 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10822) );
  NAND4_X1 U13671 ( .A1(n10825), .A2(n10824), .A3(n10823), .A4(n10822), .ZN(
        n10831) );
  AOI22_X1 U13672 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10829) );
  AOI22_X1 U13673 ( .A1(n10856), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U13674 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U13675 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10826) );
  NAND4_X1 U13676 ( .A1(n10829), .A2(n10828), .A3(n10827), .A4(n10826), .ZN(
        n10830) );
  OAI21_X1 U13677 ( .B1(n10831), .B2(n10830), .A(n10956), .ZN(n10832) );
  AOI22_X1 U13678 ( .A1(n14820), .A2(n10960), .B1(n10833), .B2(n10832), .ZN(
        n14525) );
  OAI21_X1 U13679 ( .B1(n10834), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n10848), .ZN(n16126) );
  INV_X1 U13680 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14687) );
  AOI22_X1 U13681 ( .A1(n10856), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10811), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U13682 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10837) );
  AOI22_X1 U13683 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10877), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U13684 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10835) );
  NAND4_X1 U13685 ( .A1(n10838), .A2(n10837), .A3(n10836), .A4(n10835), .ZN(
        n10844) );
  AOI22_X1 U13686 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10842) );
  AOI22_X1 U13687 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10806), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U13688 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10869), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U13689 ( .A1(n10891), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10839) );
  NAND4_X1 U13690 ( .A1(n10842), .A2(n10841), .A3(n10840), .A4(n10839), .ZN(
        n10843) );
  OAI21_X1 U13691 ( .B1(n10844), .B2(n10843), .A(n10956), .ZN(n10846) );
  AOI21_X1 U13692 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20811), .A(
        n10960), .ZN(n10845) );
  OAI211_X1 U13693 ( .C1(n10886), .C2(n14687), .A(n10846), .B(n10845), .ZN(
        n10847) );
  OAI21_X1 U13694 ( .B1(n16126), .B2(n10971), .A(n10847), .ZN(n14509) );
  INV_X1 U13695 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n21040) );
  NAND2_X1 U13696 ( .A1(n10848), .A2(n21040), .ZN(n10849) );
  AND2_X1 U13697 ( .A1(n10866), .A2(n10849), .ZN(n14813) );
  AOI21_X1 U13698 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n21040), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10850) );
  AOI21_X1 U13699 ( .B1(n10965), .B2(P1_EAX_REG_20__SCAN_IN), .A(n10850), .ZN(
        n10864) );
  AOI22_X1 U13700 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10870), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U13701 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10890), .B1(
        n10811), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U13702 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U13703 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10852) );
  NAND4_X1 U13704 ( .A1(n10855), .A2(n10854), .A3(n10853), .A4(n10852), .ZN(
        n10862) );
  AOI22_X1 U13705 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10900), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10860) );
  AOI22_X1 U13706 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10856), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10859) );
  AOI22_X1 U13707 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10876), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U13708 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10869), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10857) );
  NAND4_X1 U13709 ( .A1(n10860), .A2(n10859), .A3(n10858), .A4(n10857), .ZN(
        n10861) );
  OAI21_X1 U13710 ( .B1(n10862), .B2(n10861), .A(n10956), .ZN(n10863) );
  AOI22_X1 U13711 ( .A1(n14813), .A2(n10960), .B1(n10864), .B2(n10863), .ZN(
        n14497) );
  INV_X1 U13712 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10865) );
  NAND2_X1 U13713 ( .A1(n10866), .A2(n10865), .ZN(n10867) );
  NAND2_X1 U13714 ( .A1(n10888), .A2(n10867), .ZN(n14805) );
  INV_X1 U13715 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14674) );
  AOI22_X1 U13716 ( .A1(n10891), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10874) );
  AOI22_X1 U13717 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10869), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10873) );
  AOI22_X1 U13718 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10872) );
  AOI22_X1 U13719 ( .A1(n10806), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10871) );
  NAND4_X1 U13720 ( .A1(n10874), .A2(n10873), .A3(n10872), .A4(n10871), .ZN(
        n10883) );
  AOI22_X1 U13721 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10352), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10881) );
  AOI22_X1 U13722 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10856), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U13723 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U13724 ( .A1(n10892), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10877), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10878) );
  NAND4_X1 U13725 ( .A1(n10881), .A2(n10880), .A3(n10879), .A4(n10878), .ZN(
        n10882) );
  OAI21_X1 U13726 ( .B1(n10883), .B2(n10882), .A(n10956), .ZN(n10885) );
  AOI21_X1 U13727 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20811), .A(
        n10960), .ZN(n10884) );
  OAI211_X1 U13728 ( .C1(n10886), .C2(n14674), .A(n10885), .B(n10884), .ZN(
        n10887) );
  XNOR2_X1 U13729 ( .A(n10888), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14793) );
  INV_X1 U13730 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14791) );
  NOR2_X1 U13731 ( .A1(n14791), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10889) );
  AOI211_X1 U13732 ( .C1(n10965), .C2(P1_EAX_REG_22__SCAN_IN), .A(n10960), .B(
        n10889), .ZN(n10908) );
  AOI22_X1 U13733 ( .A1(n10875), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10806), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10897) );
  AOI22_X1 U13734 ( .A1(n10891), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10896) );
  AOI22_X1 U13735 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U13736 ( .A1(n10877), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10894) );
  NAND4_X1 U13737 ( .A1(n10897), .A2(n10896), .A3(n10895), .A4(n10894), .ZN(
        n10906) );
  AOI22_X1 U13738 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10856), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10904) );
  AOI22_X1 U13739 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10903) );
  AOI22_X1 U13740 ( .A1(n10851), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10898), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10902) );
  AOI22_X1 U13741 ( .A1(n10900), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10899), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10901) );
  NAND4_X1 U13742 ( .A1(n10904), .A2(n10903), .A3(n10902), .A4(n10901), .ZN(
        n10905) );
  OAI21_X1 U13743 ( .B1(n10906), .B2(n10905), .A(n10956), .ZN(n10907) );
  AOI22_X1 U13744 ( .A1(n14793), .A2(n10960), .B1(n10908), .B2(n10907), .ZN(
        n14476) );
  NAND2_X1 U13745 ( .A1(n10910), .A2(n10909), .ZN(n10911) );
  NAND2_X1 U13746 ( .A1(n10918), .A2(n10911), .ZN(n14787) );
  XNOR2_X1 U13747 ( .A(n10913), .B(n10912), .ZN(n10916) );
  AOI21_X1 U13748 ( .B1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20811), .A(
        n10960), .ZN(n10915) );
  NAND2_X1 U13749 ( .A1(n10965), .A2(P1_EAX_REG_23__SCAN_IN), .ZN(n10914) );
  OAI211_X1 U13750 ( .C1(n10968), .C2(n10916), .A(n10915), .B(n10914), .ZN(
        n10917) );
  XNOR2_X1 U13751 ( .A(n10918), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14775) );
  NOR2_X1 U13752 ( .A1(n14773), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10919) );
  AOI211_X1 U13753 ( .C1(n10965), .C2(P1_EAX_REG_24__SCAN_IN), .A(n10960), .B(
        n10919), .ZN(n10924) );
  XOR2_X1 U13754 ( .A(n10921), .B(n10920), .Z(n10922) );
  NAND2_X1 U13755 ( .A1(n10922), .A2(n10956), .ZN(n10923) );
  AOI22_X1 U13756 ( .A1(n14775), .A2(n10960), .B1(n10924), .B2(n10923), .ZN(
        n14449) );
  INV_X1 U13757 ( .A(n10925), .ZN(n10927) );
  INV_X1 U13758 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10926) );
  NAND2_X1 U13759 ( .A1(n10927), .A2(n10926), .ZN(n10928) );
  NAND2_X1 U13760 ( .A1(n10935), .A2(n10928), .ZN(n14769) );
  XNOR2_X1 U13761 ( .A(n10930), .B(n10929), .ZN(n10933) );
  AOI21_X1 U13762 ( .B1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20811), .A(
        n10960), .ZN(n10932) );
  NAND2_X1 U13763 ( .A1(n10965), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n10931) );
  OAI211_X1 U13764 ( .C1(n10933), .C2(n10968), .A(n10932), .B(n10931), .ZN(
        n10934) );
  XNOR2_X1 U13765 ( .A(n10935), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14760) );
  AOI21_X1 U13766 ( .B1(n14756), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10936) );
  AOI21_X1 U13767 ( .B1(n10965), .B2(P1_EAX_REG_26__SCAN_IN), .A(n10936), .ZN(
        n10941) );
  XOR2_X1 U13768 ( .A(n10938), .B(n10937), .Z(n10939) );
  NAND2_X1 U13769 ( .A1(n10939), .A2(n10956), .ZN(n10940) );
  NAND2_X1 U13770 ( .A1(n10943), .A2(n10942), .ZN(n10944) );
  NAND2_X1 U13771 ( .A1(n10945), .A2(n10944), .ZN(n14748) );
  XNOR2_X1 U13772 ( .A(n10947), .B(n10946), .ZN(n10950) );
  AOI21_X1 U13773 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20811), .A(
        n10960), .ZN(n10949) );
  NAND2_X1 U13774 ( .A1(n10965), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n10948) );
  OAI211_X1 U13775 ( .C1(n10950), .C2(n10968), .A(n10949), .B(n10948), .ZN(
        n10951) );
  XOR2_X1 U13776 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B(n10952), .Z(
        n14733) );
  INV_X1 U13777 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14731) );
  AOI21_X1 U13778 ( .B1(n14731), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10953) );
  AOI21_X1 U13779 ( .B1(n10965), .B2(P1_EAX_REG_28__SCAN_IN), .A(n10953), .ZN(
        n10959) );
  XOR2_X1 U13780 ( .A(n10955), .B(n10954), .Z(n10957) );
  NAND2_X1 U13781 ( .A1(n10957), .A2(n10956), .ZN(n10958) );
  INV_X1 U13782 ( .A(n10961), .ZN(n10962) );
  OAI21_X1 U13783 ( .B1(n10962), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n13575), .ZN(n14727) );
  XNOR2_X1 U13784 ( .A(n10964), .B(n10963), .ZN(n10969) );
  AOI21_X1 U13785 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20811), .A(
        n10960), .ZN(n10967) );
  NAND2_X1 U13786 ( .A1(n10965), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n10966) );
  OAI211_X1 U13787 ( .C1(n10969), .C2(n10968), .A(n10967), .B(n10966), .ZN(
        n10970) );
  OAI21_X1 U13788 ( .B1(n14727), .B2(n10971), .A(n10970), .ZN(n11136) );
  INV_X1 U13789 ( .A(n10972), .ZN(n14376) );
  NAND3_X1 U13790 ( .A1(n20815), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16261) );
  INV_X1 U13791 ( .A(n16261), .ZN(n10973) );
  NOR2_X2 U13792 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20661) );
  NAND2_X1 U13793 ( .A1(n10973), .A2(n20661), .ZN(n20129) );
  NAND2_X1 U13794 ( .A1(n14376), .A2(n16152), .ZN(n11134) );
  INV_X1 U13795 ( .A(n11075), .ZN(n11031) );
  AND3_X1 U13796 ( .A1(n10975), .A2(n11031), .A3(n11044), .ZN(n10976) );
  NOR2_X1 U13797 ( .A1(n9721), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11070) );
  NAND2_X1 U13798 ( .A1(n10990), .A2(n10989), .ZN(n10978) );
  NAND2_X1 U13799 ( .A1(n10979), .A2(n10978), .ZN(n11000) );
  NAND3_X1 U13800 ( .A1(n10980), .A2(n10990), .A3(n10989), .ZN(n10981) );
  NAND2_X1 U13801 ( .A1(n11000), .A2(n10981), .ZN(n10983) );
  NAND2_X1 U13802 ( .A1(n10430), .A2(n20157), .ZN(n10985) );
  INV_X1 U13803 ( .A(n10985), .ZN(n10982) );
  AOI21_X1 U13804 ( .B1(n10983), .B2(n20813), .A(n10982), .ZN(n10984) );
  OAI21_X1 U13805 ( .B1(n13166), .B2(n10990), .A(n10985), .ZN(n10986) );
  INV_X1 U13806 ( .A(n10986), .ZN(n10987) );
  NAND2_X2 U13807 ( .A1(n13043), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13045) );
  OR2_X1 U13808 ( .A1(n10988), .A2(n13165), .ZN(n10994) );
  XNOR2_X1 U13809 ( .A(n10990), .B(n10989), .ZN(n10991) );
  OAI211_X1 U13810 ( .C1(n10991), .C2(n13166), .A(n11073), .B(n10388), .ZN(
        n10992) );
  INV_X1 U13811 ( .A(n10992), .ZN(n10993) );
  NAND2_X1 U13812 ( .A1(n10994), .A2(n10993), .ZN(n10995) );
  XNOR2_X2 U13813 ( .A(n13045), .B(n10995), .ZN(n13140) );
  INV_X1 U13814 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10996) );
  NAND2_X1 U13815 ( .A1(n10997), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10998) );
  XNOR2_X1 U13816 ( .A(n11004), .B(n20095), .ZN(n13500) );
  NAND2_X1 U13817 ( .A1(n10999), .A2(n11031), .ZN(n11003) );
  NAND2_X1 U13818 ( .A1(n11000), .A2(n11001), .ZN(n11017) );
  OAI211_X1 U13819 ( .C1(n11001), .C2(n11000), .A(n11017), .B(n20813), .ZN(
        n11002) );
  NAND2_X1 U13820 ( .A1(n11003), .A2(n11002), .ZN(n13501) );
  NAND2_X1 U13821 ( .A1(n13500), .A2(n13501), .ZN(n11006) );
  NAND2_X1 U13822 ( .A1(n11004), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11005) );
  NAND2_X1 U13823 ( .A1(n11006), .A2(n11005), .ZN(n13543) );
  INV_X1 U13824 ( .A(n11007), .ZN(n11008) );
  OR2_X1 U13825 ( .A1(n11008), .A2(n11075), .ZN(n11011) );
  XNOR2_X1 U13826 ( .A(n11017), .B(n11015), .ZN(n11009) );
  NAND2_X1 U13827 ( .A1(n11009), .A2(n20813), .ZN(n11010) );
  NAND2_X1 U13828 ( .A1(n11011), .A2(n11010), .ZN(n11012) );
  INV_X1 U13829 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21014) );
  XNOR2_X1 U13830 ( .A(n11012), .B(n21014), .ZN(n13544) );
  NAND2_X1 U13831 ( .A1(n11012), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11013) );
  OR2_X1 U13832 ( .A1(n11014), .A2(n11075), .ZN(n11021) );
  INV_X1 U13833 ( .A(n11015), .ZN(n11016) );
  NOR2_X1 U13834 ( .A1(n11017), .A2(n11016), .ZN(n11019) );
  NAND2_X1 U13835 ( .A1(n11019), .A2(n11018), .ZN(n11033) );
  OAI211_X1 U13836 ( .C1(n11019), .C2(n11018), .A(n11033), .B(n20813), .ZN(
        n11020) );
  NAND2_X1 U13837 ( .A1(n11021), .A2(n11020), .ZN(n11022) );
  INV_X1 U13838 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13558) );
  XNOR2_X1 U13839 ( .A(n11022), .B(n13558), .ZN(n13536) );
  NAND2_X1 U13840 ( .A1(n11022), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11023) );
  XNOR2_X1 U13841 ( .A(n11033), .B(n11034), .ZN(n11025) );
  NAND2_X1 U13842 ( .A1(n11025), .A2(n20813), .ZN(n11026) );
  NAND2_X1 U13843 ( .A1(n11027), .A2(n11026), .ZN(n11028) );
  XNOR2_X1 U13844 ( .A(n11028), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13656) );
  INV_X1 U13845 ( .A(n11028), .ZN(n11029) );
  INV_X1 U13846 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14886) );
  NAND2_X1 U13847 ( .A1(n11029), .A2(n14886), .ZN(n11030) );
  NAND2_X1 U13848 ( .A1(n11032), .A2(n11031), .ZN(n11038) );
  INV_X1 U13849 ( .A(n11033), .ZN(n11035) );
  NAND2_X1 U13850 ( .A1(n11035), .A2(n11034), .ZN(n11043) );
  XNOR2_X1 U13851 ( .A(n11043), .B(n11044), .ZN(n11036) );
  NAND2_X1 U13852 ( .A1(n11036), .A2(n20813), .ZN(n11037) );
  NAND2_X1 U13853 ( .A1(n11038), .A2(n11037), .ZN(n11039) );
  INV_X1 U13854 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11040) );
  XNOR2_X1 U13855 ( .A(n11039), .B(n11040), .ZN(n13720) );
  INV_X1 U13856 ( .A(n11039), .ZN(n11041) );
  NAND2_X1 U13857 ( .A1(n11041), .A2(n11040), .ZN(n11042) );
  INV_X1 U13858 ( .A(n11043), .ZN(n11045) );
  NAND3_X1 U13859 ( .A1(n11045), .A2(n20813), .A3(n11044), .ZN(n11046) );
  NAND2_X1 U13860 ( .A1(n9721), .A2(n11046), .ZN(n11047) );
  NAND2_X1 U13861 ( .A1(n11047), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13802) );
  INV_X1 U13862 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16233) );
  INV_X2 U13863 ( .A(n11054), .ZN(n14734) );
  NAND2_X1 U13864 ( .A1(n9721), .A2(n16233), .ZN(n11049) );
  NAND2_X1 U13865 ( .A1(n14734), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14852) );
  INV_X1 U13866 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15055) );
  NAND2_X1 U13867 ( .A1(n9721), .A2(n15055), .ZN(n11050) );
  NAND2_X1 U13868 ( .A1(n14852), .A2(n11050), .ZN(n14867) );
  INV_X1 U13869 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16214) );
  NAND2_X1 U13870 ( .A1(n9721), .A2(n16214), .ZN(n14866) );
  NAND2_X1 U13871 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11051) );
  NAND2_X1 U13872 ( .A1(n9721), .A2(n11051), .ZN(n14863) );
  NAND2_X1 U13873 ( .A1(n14866), .A2(n14863), .ZN(n11052) );
  NOR2_X1 U13874 ( .A1(n14867), .A2(n11052), .ZN(n14851) );
  INV_X1 U13875 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16198) );
  NAND2_X1 U13876 ( .A1(n9721), .A2(n16198), .ZN(n11053) );
  NAND2_X1 U13877 ( .A1(n14851), .A2(n11053), .ZN(n14825) );
  NAND2_X1 U13878 ( .A1(n14734), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14836) );
  OAI21_X1 U13879 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(n14734), .ZN(n11055) );
  AND2_X1 U13880 ( .A1(n14836), .A2(n11055), .ZN(n16130) );
  XNOR2_X1 U13881 ( .A(n9721), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14826) );
  INV_X1 U13882 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14893) );
  NAND2_X1 U13883 ( .A1(n9721), .A2(n14893), .ZN(n14839) );
  NAND2_X1 U13884 ( .A1(n14826), .A2(n14839), .ZN(n11056) );
  AOI21_X1 U13885 ( .B1(n14825), .B2(n16130), .A(n11056), .ZN(n16128) );
  INV_X1 U13886 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11057) );
  NAND2_X1 U13887 ( .A1(n9721), .A2(n11057), .ZN(n11058) );
  AND2_X1 U13888 ( .A1(n16128), .A2(n11058), .ZN(n11059) );
  NOR2_X1 U13889 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14850) );
  NAND4_X1 U13890 ( .A1(n14850), .A2(n16198), .A3(n15055), .A4(n16214), .ZN(
        n11060) );
  NAND2_X1 U13891 ( .A1(n14734), .A2(n11060), .ZN(n14837) );
  NAND2_X1 U13892 ( .A1(n14836), .A2(n14837), .ZN(n14840) );
  NOR2_X1 U13893 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11061) );
  NOR2_X1 U13894 ( .A1(n9721), .A2(n11061), .ZN(n11062) );
  NOR2_X1 U13895 ( .A1(n14840), .A2(n11062), .ZN(n11063) );
  XNOR2_X1 U13896 ( .A(n9721), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14821) );
  AND2_X1 U13897 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14904) );
  NAND2_X1 U13898 ( .A1(n14794), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11066) );
  INV_X1 U13899 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14894) );
  INV_X1 U13900 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15020) );
  INV_X1 U13901 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15014) );
  INV_X1 U13902 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15024) );
  NAND4_X1 U13903 ( .A1(n14894), .A2(n15020), .A3(n15014), .A4(n15024), .ZN(
        n11065) );
  NOR2_X1 U13904 ( .A1(n11064), .A2(n11065), .ZN(n14795) );
  AND2_X1 U13905 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14963) );
  NAND2_X1 U13906 ( .A1(n14963), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14897) );
  NAND2_X1 U13907 ( .A1(n14752), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11067) );
  AOI21_X2 U13908 ( .B1(n14765), .B2(n14897), .A(n11067), .ZN(n11069) );
  INV_X1 U13909 ( .A(n11069), .ZN(n14745) );
  INV_X1 U13910 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15002) );
  INV_X1 U13911 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14993) );
  INV_X1 U13912 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14962) );
  AND3_X1 U13913 ( .A1(n15002), .A2(n14993), .A3(n14962), .ZN(n14753) );
  INV_X1 U13914 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14740) );
  INV_X1 U13915 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14958) );
  AND2_X1 U13916 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14912) );
  AND3_X2 U13917 ( .A1(n14724), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n9721), .ZN(n14714) );
  NAND2_X1 U13918 ( .A1(n10331), .A2(n10430), .ZN(n11072) );
  XNOR2_X1 U13919 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11086) );
  NAND2_X1 U13920 ( .A1(n20573), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11090) );
  NAND2_X1 U13921 ( .A1(n11086), .A2(n11087), .ZN(n11077) );
  NAND2_X1 U13922 ( .A1(n20541), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11076) );
  NAND2_X1 U13923 ( .A1(n11077), .A2(n11076), .ZN(n11100) );
  XNOR2_X1 U13924 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11099) );
  NAND2_X1 U13925 ( .A1(n11100), .A2(n11099), .ZN(n11079) );
  NAND2_X1 U13926 ( .A1(n20459), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11078) );
  NAND2_X1 U13927 ( .A1(n11079), .A2(n11078), .ZN(n11085) );
  XNOR2_X1 U13928 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11084) );
  NAND2_X1 U13929 ( .A1(n11085), .A2(n11084), .ZN(n11081) );
  NAND2_X1 U13930 ( .A1(n21022), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11080) );
  NAND2_X1 U13931 ( .A1(n11081), .A2(n11080), .ZN(n11113) );
  NOR2_X1 U13932 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10603), .ZN(
        n11082) );
  NAND2_X1 U13933 ( .A1(n11111), .A2(n12865), .ZN(n11124) );
  NAND2_X1 U13934 ( .A1(n12865), .A2(n11089), .ZN(n11122) );
  XNOR2_X1 U13935 ( .A(n11085), .B(n11084), .ZN(n12861) );
  XNOR2_X1 U13936 ( .A(n11087), .B(n11086), .ZN(n12860) );
  INV_X1 U13937 ( .A(n11098), .ZN(n11088) );
  NOR2_X1 U13938 ( .A1(n12860), .A2(n11088), .ZN(n11096) );
  OAI21_X1 U13939 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20573), .A(
        n11090), .ZN(n11092) );
  NOR2_X1 U13940 ( .A1(n11106), .A2(n11092), .ZN(n11095) );
  NAND2_X1 U13941 ( .A1(n11149), .A2(n20135), .ZN(n11091) );
  NAND2_X1 U13942 ( .A1(n11091), .A2(n13165), .ZN(n11105) );
  INV_X1 U13943 ( .A(n11092), .ZN(n11093) );
  OAI211_X1 U13944 ( .C1(n10430), .C2(n10422), .A(n11105), .B(n11093), .ZN(
        n11094) );
  OAI21_X1 U13945 ( .B1(n11111), .B2(n11095), .A(n11094), .ZN(n11097) );
  NAND2_X1 U13946 ( .A1(n11096), .A2(n11097), .ZN(n11104) );
  OAI211_X1 U13947 ( .C1(n11098), .C2(n11097), .A(n12860), .B(n11117), .ZN(
        n11103) );
  XNOR2_X1 U13948 ( .A(n11100), .B(n11099), .ZN(n12862) );
  NAND2_X1 U13949 ( .A1(n11115), .A2(n12862), .ZN(n11101) );
  OAI211_X1 U13950 ( .C1(n11106), .C2(n12862), .A(n11101), .B(n11105), .ZN(
        n11102) );
  NAND3_X1 U13951 ( .A1(n11104), .A2(n11103), .A3(n11102), .ZN(n11108) );
  AOI22_X1 U13952 ( .A1(n11109), .A2(n12861), .B1(n11108), .B2(n11107), .ZN(
        n11110) );
  AOI21_X1 U13953 ( .B1(n11111), .B2(n12861), .A(n11110), .ZN(n11119) );
  INV_X1 U13954 ( .A(n12863), .ZN(n11114) );
  NOR2_X1 U13955 ( .A1(n11115), .A2(n11114), .ZN(n11118) );
  NAND2_X1 U13956 ( .A1(n11115), .A2(n12863), .ZN(n11116) );
  OAI22_X1 U13957 ( .A1(n11119), .A2(n11118), .B1(n11117), .B2(n11116), .ZN(
        n11120) );
  AOI21_X1 U13958 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20815), .A(
        n11120), .ZN(n11121) );
  NAND2_X1 U13959 ( .A1(n11122), .A2(n11121), .ZN(n11123) );
  OR2_X1 U13960 ( .A1(n16052), .A2(n20815), .ZN(n19964) );
  NAND2_X1 U13961 ( .A1(n11126), .A2(n11125), .ZN(n11133) );
  INV_X1 U13962 ( .A(n20661), .ZN(n20653) );
  NAND2_X1 U13963 ( .A1(n20653), .A2(n11129), .ZN(n20818) );
  NAND2_X1 U13964 ( .A1(n20818), .A2(n20815), .ZN(n11127) );
  NAND2_X1 U13965 ( .A1(n20815), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16045) );
  INV_X1 U13966 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20812) );
  NAND2_X1 U13967 ( .A1(n20812), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11128) );
  AND2_X1 U13968 ( .A1(n16045), .A2(n11128), .ZN(n13041) );
  NAND2_X1 U13969 ( .A1(n14383), .A2(n16151), .ZN(n11130) );
  INV_X1 U13970 ( .A(n16200), .ZN(n16171) );
  NAND2_X1 U13971 ( .A1(n16171), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14925) );
  OAI211_X1 U13972 ( .C1(n14818), .C2(n20950), .A(n11130), .B(n14925), .ZN(
        n11131) );
  INV_X1 U13973 ( .A(n11131), .ZN(n11132) );
  NAND3_X1 U13974 ( .A1(n11134), .A2(n11133), .A3(n11132), .ZN(P1_U2969) );
  INV_X1 U13975 ( .A(n14729), .ZN(n14644) );
  OAI21_X1 U13976 ( .B1(n11074), .B2(n13583), .A(n11137), .ZN(n11138) );
  NOR2_X1 U13977 ( .A1(n11139), .A2(n11138), .ZN(n11143) );
  OAI21_X1 U13978 ( .B1(n10387), .B2(n21125), .A(n10389), .ZN(n11140) );
  OAI211_X1 U13979 ( .C1(n11071), .C2(n11233), .A(n11143), .B(n11142), .ZN(
        n13158) );
  INV_X1 U13980 ( .A(n11146), .ZN(n11147) );
  NAND3_X1 U13981 ( .A1(n11145), .A2(n11147), .A3(n13160), .ZN(n11148) );
  OR2_X1 U13982 ( .A1(n10424), .A2(n13165), .ZN(n13141) );
  INV_X1 U13983 ( .A(n16055), .ZN(n13201) );
  NAND2_X1 U13984 ( .A1(n13190), .A2(n13201), .ZN(n13209) );
  INV_X1 U13985 ( .A(n10389), .ZN(n14071) );
  NAND4_X1 U13986 ( .A1(n14071), .A2(n11149), .A3(n10421), .A4(n21125), .ZN(
        n11150) );
  NOR2_X1 U13987 ( .A1(n11150), .A2(n10429), .ZN(n13054) );
  NAND2_X1 U13988 ( .A1(n13054), .A2(n13587), .ZN(n11151) );
  NAND2_X1 U13989 ( .A1(n13209), .A2(n11151), .ZN(n11152) );
  INV_X1 U13990 ( .A(n11246), .ZN(n14058) );
  OR2_X1 U13991 ( .A1(n11243), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n11157) );
  INV_X1 U13992 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11153) );
  NAND2_X1 U13993 ( .A1(n11194), .A2(n11153), .ZN(n11155) );
  INV_X1 U13995 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13068) );
  NAND2_X1 U13996 ( .A1(n13587), .A2(n13068), .ZN(n11154) );
  NAND3_X1 U13997 ( .A1(n11155), .A2(n11233), .A3(n11154), .ZN(n11156) );
  INV_X1 U13998 ( .A(n11163), .ZN(n11194) );
  NAND2_X1 U13999 ( .A1(n11194), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11159) );
  INV_X1 U14000 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13613) );
  NAND2_X1 U14001 ( .A1(n11233), .A2(n13613), .ZN(n11158) );
  NAND2_X1 U14002 ( .A1(n11159), .A2(n11158), .ZN(n13011) );
  XNOR2_X1 U14003 ( .A(n11160), .B(n13011), .ZN(n13590) );
  INV_X1 U14004 ( .A(n11160), .ZN(n11161) );
  AOI21_X1 U14005 ( .B1(n13590), .B2(n13587), .A(n11161), .ZN(n13135) );
  MUX2_X1 U14006 ( .A(n11243), .B(n11194), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n11166) );
  INV_X1 U14007 ( .A(n11162), .ZN(n11163) );
  NAND2_X1 U14008 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14358), .ZN(
        n11164) );
  AND2_X1 U14009 ( .A1(n11196), .A2(n11164), .ZN(n11165) );
  NAND2_X1 U14010 ( .A1(n11166), .A2(n11165), .ZN(n13134) );
  MUX2_X1 U14011 ( .A(n11229), .B(n11246), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n11169) );
  OR2_X1 U14012 ( .A1(n11167), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11168) );
  AND2_X1 U14013 ( .A1(n11169), .A2(n11168), .ZN(n13259) );
  MUX2_X1 U14014 ( .A(n11243), .B(n11194), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n11171) );
  NAND2_X1 U14015 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n14358), .ZN(
        n11170) );
  INV_X1 U14016 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n13417) );
  NAND2_X1 U14017 ( .A1(n13587), .A2(n13417), .ZN(n11173) );
  NAND2_X1 U14018 ( .A1(n11224), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11172) );
  NAND3_X1 U14019 ( .A1(n11194), .A2(n11173), .A3(n11172), .ZN(n11174) );
  OAI21_X1 U14020 ( .B1(n11229), .B2(P1_EBX_REG_5__SCAN_IN), .A(n11174), .ZN(
        n13415) );
  MUX2_X1 U14021 ( .A(n11243), .B(n11194), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n11177) );
  NAND2_X1 U14022 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14358), .ZN(
        n11175) );
  AND2_X1 U14023 ( .A1(n11196), .A2(n11175), .ZN(n11176) );
  NAND2_X1 U14024 ( .A1(n11177), .A2(n11176), .ZN(n13510) );
  INV_X1 U14025 ( .A(n11229), .ZN(n11232) );
  INV_X1 U14026 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20001) );
  NAND2_X1 U14027 ( .A1(n11232), .A2(n20001), .ZN(n11181) );
  NAND2_X1 U14028 ( .A1(n13587), .A2(n20001), .ZN(n11179) );
  NAND2_X1 U14029 ( .A1(n11224), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11178) );
  NAND3_X1 U14030 ( .A1(n11194), .A2(n11179), .A3(n11178), .ZN(n11180) );
  MUX2_X1 U14031 ( .A(n11243), .B(n11194), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n11183) );
  NAND2_X1 U14032 ( .A1(n14358), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11182) );
  INV_X1 U14033 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n13794) );
  NAND2_X1 U14034 ( .A1(n13587), .A2(n13794), .ZN(n11185) );
  NAND2_X1 U14035 ( .A1(n11224), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11184) );
  NAND3_X1 U14036 ( .A1(n11194), .A2(n11185), .A3(n11184), .ZN(n11186) );
  OAI21_X1 U14037 ( .B1(n11229), .B2(P1_EBX_REG_9__SCAN_IN), .A(n11186), .ZN(
        n13790) );
  OR2_X1 U14038 ( .A1(n11243), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n11190) );
  NAND2_X1 U14039 ( .A1(n11194), .A2(n16234), .ZN(n11188) );
  INV_X1 U14040 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n16109) );
  NAND2_X1 U14041 ( .A1(n13587), .A2(n16109), .ZN(n11187) );
  NAND3_X1 U14042 ( .A1(n11188), .A2(n11224), .A3(n11187), .ZN(n11189) );
  NAND2_X1 U14043 ( .A1(n11190), .A2(n11189), .ZN(n13926) );
  NAND2_X1 U14044 ( .A1(n13927), .A2(n13926), .ZN(n13955) );
  MUX2_X1 U14045 ( .A(n11229), .B(n11233), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n11191) );
  OAI21_X1 U14046 ( .B1(n11167), .B2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11191), .ZN(n13956) );
  MUX2_X1 U14047 ( .A(n11229), .B(n11233), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n11192) );
  OAI21_X1 U14048 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n11167), .A(
        n11192), .ZN(n11193) );
  INV_X1 U14049 ( .A(n11193), .ZN(n14632) );
  MUX2_X1 U14050 ( .A(n11243), .B(n11194), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n11198) );
  NAND2_X1 U14051 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14358), .ZN(
        n11195) );
  AND2_X1 U14052 ( .A1(n11196), .A2(n11195), .ZN(n11197) );
  NAND2_X1 U14053 ( .A1(n11198), .A2(n11197), .ZN(n16100) );
  OR2_X1 U14054 ( .A1(n11243), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n11202) );
  NAND2_X1 U14055 ( .A1(n11194), .A2(n16198), .ZN(n11200) );
  INV_X1 U14056 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14625) );
  NAND2_X1 U14057 ( .A1(n13587), .A2(n14625), .ZN(n11199) );
  NAND3_X1 U14058 ( .A1(n11200), .A2(n11224), .A3(n11199), .ZN(n11201) );
  MUX2_X1 U14059 ( .A(n11229), .B(n11233), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n11203) );
  OAI21_X1 U14060 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n11167), .A(
        n11203), .ZN(n14548) );
  INV_X1 U14061 ( .A(n14548), .ZN(n11204) );
  OR2_X1 U14062 ( .A1(n11243), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n11209) );
  INV_X1 U14063 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14892) );
  NAND2_X1 U14064 ( .A1(n11194), .A2(n14892), .ZN(n11207) );
  INV_X1 U14065 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n11205) );
  NAND2_X1 U14066 ( .A1(n13587), .A2(n11205), .ZN(n11206) );
  NAND3_X1 U14067 ( .A1(n11207), .A2(n11246), .A3(n11206), .ZN(n11208) );
  MUX2_X1 U14068 ( .A(n11229), .B(n11224), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n11211) );
  OR2_X1 U14069 ( .A1(n11167), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11210) );
  NAND2_X1 U14070 ( .A1(n11211), .A2(n11210), .ZN(n14617) );
  NOR2_X1 U14071 ( .A1(n14614), .A2(n14617), .ZN(n11212) );
  OR2_X1 U14072 ( .A1(n11243), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n11216) );
  NAND2_X1 U14073 ( .A1(n11194), .A2(n14894), .ZN(n11214) );
  INV_X1 U14074 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14608) );
  NAND2_X1 U14075 ( .A1(n13587), .A2(n14608), .ZN(n11213) );
  NAND3_X1 U14076 ( .A1(n11214), .A2(n11233), .A3(n11213), .ZN(n11215) );
  AND2_X1 U14077 ( .A1(n11216), .A2(n11215), .ZN(n14526) );
  MUX2_X1 U14078 ( .A(n11229), .B(n11224), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n11217) );
  OAI21_X1 U14079 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n11167), .A(
        n11217), .ZN(n14517) );
  MUX2_X1 U14080 ( .A(n11243), .B(n11194), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n11219) );
  NAND2_X1 U14081 ( .A1(n14358), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11218) );
  NAND2_X1 U14082 ( .A1(n11219), .A2(n11218), .ZN(n14498) );
  MUX2_X1 U14083 ( .A(n11229), .B(n11233), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n11221) );
  OR2_X1 U14084 ( .A1(n11167), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11220) );
  NAND2_X1 U14085 ( .A1(n11221), .A2(n11220), .ZN(n14489) );
  MUX2_X1 U14086 ( .A(n11243), .B(n11194), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n11223) );
  NAND2_X1 U14087 ( .A1(n14358), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11222) );
  AND2_X1 U14088 ( .A1(n11223), .A2(n11222), .ZN(n14477) );
  MUX2_X1 U14089 ( .A(n11229), .B(n11224), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n11225) );
  OAI21_X1 U14090 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n11167), .A(
        n11225), .ZN(n14465) );
  OR2_X1 U14091 ( .A1(n11243), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n11228) );
  NAND2_X1 U14092 ( .A1(n11194), .A2(n14993), .ZN(n11226) );
  OAI211_X1 U14093 ( .C1(n14358), .C2(P1_EBX_REG_24__SCAN_IN), .A(n11224), .B(
        n11226), .ZN(n11227) );
  AND2_X1 U14094 ( .A1(n11228), .A2(n11227), .ZN(n14451) );
  MUX2_X1 U14095 ( .A(n11229), .B(n11224), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n11231) );
  OR2_X1 U14096 ( .A1(n11167), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11230) );
  AND2_X1 U14097 ( .A1(n11231), .A2(n11230), .ZN(n14432) );
  INV_X1 U14098 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14598) );
  NAND2_X1 U14099 ( .A1(n11232), .A2(n14598), .ZN(n11237) );
  NAND2_X1 U14100 ( .A1(n13587), .A2(n14598), .ZN(n11235) );
  NAND2_X1 U14101 ( .A1(n11233), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11234) );
  NAND3_X1 U14102 ( .A1(n11194), .A2(n11235), .A3(n11234), .ZN(n11236) );
  AND2_X1 U14103 ( .A1(n11237), .A2(n11236), .ZN(n14406) );
  OR2_X1 U14104 ( .A1(n11243), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n11242) );
  INV_X1 U14105 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14967) );
  NAND2_X1 U14106 ( .A1(n11194), .A2(n14967), .ZN(n11240) );
  INV_X1 U14107 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n11238) );
  NAND2_X1 U14108 ( .A1(n13587), .A2(n11238), .ZN(n11239) );
  NAND3_X1 U14109 ( .A1(n11240), .A2(n11224), .A3(n11239), .ZN(n11241) );
  NAND2_X1 U14110 ( .A1(n11242), .A2(n11241), .ZN(n14422) );
  OR2_X1 U14111 ( .A1(n11243), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n11249) );
  NAND2_X1 U14112 ( .A1(n11194), .A2(n14740), .ZN(n11247) );
  INV_X1 U14113 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n11244) );
  NAND2_X1 U14114 ( .A1(n13587), .A2(n11244), .ZN(n11245) );
  NAND3_X1 U14115 ( .A1(n11247), .A2(n11246), .A3(n11245), .ZN(n11248) );
  NAND2_X1 U14116 ( .A1(n11249), .A2(n11248), .ZN(n14395) );
  OR2_X1 U14117 ( .A1(n11167), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11250) );
  INV_X1 U14118 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n11252) );
  NAND2_X1 U14119 ( .A1(n13587), .A2(n11252), .ZN(n11251) );
  NAND2_X1 U14120 ( .A1(n11250), .A2(n11251), .ZN(n14059) );
  MUX2_X1 U14121 ( .A(n14059), .B(n11251), .S(n14058), .Z(n14056) );
  XNOR2_X1 U14122 ( .A(n14396), .B(n14056), .ZN(n14932) );
  INV_X1 U14123 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11462) );
  AND2_X4 U14124 ( .A1(n11509), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14127) );
  AND2_X4 U14125 ( .A1(n11509), .A2(n13290), .ZN(n11500) );
  AOI22_X1 U14126 ( .A1(n11353), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11500), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11259) );
  AND3_X4 U14127 ( .A1(n11515), .A2(n11658), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11514) );
  BUF_X2 U14128 ( .A(n11334), .Z(n14292) );
  AOI22_X1 U14129 ( .A1(n14127), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14140), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11263) );
  AOI22_X1 U14130 ( .A1(n11514), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14292), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11262) );
  AOI22_X1 U14131 ( .A1(n11500), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11261) );
  AOI22_X1 U14132 ( .A1(n11353), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11498), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11260) );
  NAND4_X1 U14133 ( .A1(n11263), .A2(n11262), .A3(n11261), .A4(n11260), .ZN(
        n11264) );
  INV_X1 U14134 ( .A(n11379), .ZN(n11278) );
  AOI22_X1 U14135 ( .A1(n14127), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14140), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11269) );
  AOI22_X1 U14136 ( .A1(n11514), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14292), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11268) );
  AOI22_X1 U14137 ( .A1(n11353), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11498), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11267) );
  AOI22_X1 U14138 ( .A1(n11500), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11266) );
  NAND4_X1 U14139 ( .A1(n11269), .A2(n11268), .A3(n11267), .A4(n11266), .ZN(
        n11270) );
  NAND2_X1 U14140 ( .A1(n11270), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11277) );
  AOI22_X1 U14141 ( .A1(n11514), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11354), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11274) );
  AOI22_X1 U14142 ( .A1(n14127), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14140), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11273) );
  AOI22_X1 U14143 ( .A1(n11500), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11272) );
  AOI22_X1 U14144 ( .A1(n11353), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11498), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11271) );
  NAND4_X1 U14145 ( .A1(n11274), .A2(n11273), .A3(n11272), .A4(n11271), .ZN(
        n11275) );
  NAND2_X1 U14146 ( .A1(n11275), .A2(n20841), .ZN(n11276) );
  AOI22_X1 U14147 ( .A1(n11353), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11498), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11280) );
  AOI22_X1 U14148 ( .A1(n11500), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11279) );
  AOI22_X1 U14149 ( .A1(n14127), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14140), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11282) );
  AOI22_X1 U14150 ( .A1(n11514), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11354), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11281) );
  AOI22_X1 U14151 ( .A1(n11353), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11498), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11290) );
  AOI22_X1 U14152 ( .A1(n14127), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14140), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11289) );
  AOI22_X1 U14153 ( .A1(n11500), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11288) );
  INV_X1 U14154 ( .A(n11285), .ZN(n11286) );
  NOR2_X1 U14155 ( .A1(n11286), .A2(n20841), .ZN(n11287) );
  NAND4_X1 U14156 ( .A1(n11290), .A2(n11289), .A3(n11288), .A4(n11287), .ZN(
        n11291) );
  AOI22_X1 U14157 ( .A1(n11353), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11500), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11296) );
  AOI22_X1 U14158 ( .A1(n14127), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14140), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11295) );
  AOI22_X1 U14159 ( .A1(n11514), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14292), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11294) );
  AOI22_X1 U14160 ( .A1(n11355), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11498), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11293) );
  NAND4_X1 U14161 ( .A1(n11296), .A2(n11295), .A3(n11294), .A4(n11293), .ZN(
        n11297) );
  NAND2_X1 U14162 ( .A1(n11297), .A2(n20841), .ZN(n11304) );
  AOI22_X1 U14163 ( .A1(n14140), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11498), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11299) );
  AOI22_X1 U14164 ( .A1(n11500), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11298) );
  NAND4_X1 U14165 ( .A1(n11301), .A2(n11300), .A3(n11299), .A4(n11298), .ZN(
        n11302) );
  NAND2_X1 U14166 ( .A1(n11302), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11303) );
  INV_X1 U14167 ( .A(n11308), .ZN(n11305) );
  NAND2_X1 U14168 ( .A1(n11381), .A2(n11366), .ZN(n11364) );
  INV_X1 U14169 ( .A(n11366), .ZN(n11307) );
  NAND2_X1 U14170 ( .A1(n11307), .A2(n12954), .ZN(n11915) );
  NAND3_X1 U14171 ( .A1(n11364), .A2(n11915), .A3(n13939), .ZN(n11922) );
  AOI22_X1 U14172 ( .A1(n14127), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14140), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11313) );
  AOI22_X1 U14173 ( .A1(n11514), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14292), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11312) );
  AOI22_X1 U14174 ( .A1(n11500), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11311) );
  AOI22_X1 U14175 ( .A1(n11353), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11498), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11310) );
  NAND4_X1 U14176 ( .A1(n11313), .A2(n11312), .A3(n11311), .A4(n11310), .ZN(
        n11314) );
  AOI22_X1 U14177 ( .A1(n14127), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14140), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11318) );
  AOI22_X1 U14178 ( .A1(n11514), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14292), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11317) );
  AOI22_X1 U14179 ( .A1(n11353), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11498), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11316) );
  AOI22_X1 U14180 ( .A1(n11500), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11315) );
  NAND4_X1 U14181 ( .A1(n11318), .A2(n11317), .A3(n11316), .A4(n11315), .ZN(
        n11319) );
  AOI22_X1 U14182 ( .A1(n11514), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14292), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U14183 ( .A1(n11500), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11323) );
  AOI22_X1 U14184 ( .A1(n14127), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14140), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11322) );
  NAND4_X1 U14185 ( .A1(n11325), .A2(n11324), .A3(n11323), .A4(n11322), .ZN(
        n11326) );
  NAND2_X1 U14186 ( .A1(n11326), .A2(n20841), .ZN(n11333) );
  AOI22_X1 U14187 ( .A1(n14127), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11498), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11329) );
  AOI22_X1 U14188 ( .A1(n11514), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14292), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11328) );
  AOI22_X1 U14189 ( .A1(n11353), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11500), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11327) );
  NAND4_X1 U14190 ( .A1(n11330), .A2(n11329), .A3(n11328), .A4(n11327), .ZN(
        n11331) );
  NAND2_X1 U14191 ( .A1(n11331), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11332) );
  AOI22_X1 U14192 ( .A1(n11514), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11334), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11337) );
  AOI22_X1 U14193 ( .A1(n11500), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U14194 ( .A1(n11353), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11498), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11335) );
  NAND4_X1 U14195 ( .A1(n11338), .A2(n11337), .A3(n11336), .A4(n11335), .ZN(
        n11339) );
  NAND2_X1 U14196 ( .A1(n11339), .A2(n20841), .ZN(n11346) );
  AOI22_X1 U14197 ( .A1(n11514), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14292), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14198 ( .A1(n14127), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14140), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14199 ( .A1(n11500), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U14200 ( .A1(n11353), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11498), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11340) );
  NAND4_X1 U14201 ( .A1(n11343), .A2(n11342), .A3(n11341), .A4(n11340), .ZN(
        n11344) );
  NAND2_X1 U14202 ( .A1(n11344), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11345) );
  INV_X1 U14203 ( .A(n13635), .ZN(n11679) );
  INV_X1 U14204 ( .A(n11370), .ZN(n11348) );
  NAND2_X1 U14205 ( .A1(n12358), .A2(n11379), .ZN(n11391) );
  NAND2_X1 U14206 ( .A1(n11348), .A2(n11391), .ZN(n11365) );
  NAND2_X1 U14207 ( .A1(n11386), .A2(n12350), .ZN(n11363) );
  AOI22_X1 U14208 ( .A1(n11500), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14140), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U14209 ( .A1(n11355), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11498), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11349) );
  AOI22_X1 U14210 ( .A1(n11353), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14127), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U14211 ( .A1(n11514), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11354), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11351) );
  NAND3_X1 U14212 ( .A1(n10161), .A2(n11352), .A3(n11351), .ZN(n11362) );
  AOI22_X1 U14213 ( .A1(n11353), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14140), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U14214 ( .A1(n11514), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11354), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14215 ( .A1(n11500), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11498), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14216 ( .A1(n14127), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11356) );
  NAND3_X1 U14217 ( .A1(n11365), .A2(n9783), .A3(n11364), .ZN(n11369) );
  INV_X1 U14218 ( .A(n11380), .ZN(n11367) );
  NAND2_X1 U14219 ( .A1(n11368), .A2(n11370), .ZN(n11377) );
  NAND3_X1 U14220 ( .A1(n11372), .A2(n11370), .A3(n9720), .ZN(n11946) );
  BUF_X4 U14221 ( .A(n11371), .Z(n19944) );
  NAND3_X1 U14222 ( .A1(n11946), .A2(n13682), .A3(n19944), .ZN(n11375) );
  NOR2_X1 U14223 ( .A1(n11915), .A2(n12358), .ZN(n11373) );
  AND2_X2 U14224 ( .A1(n11373), .A2(n11372), .ZN(n11395) );
  INV_X1 U14225 ( .A(n11395), .ZN(n11374) );
  INV_X1 U14226 ( .A(n11895), .ZN(n11376) );
  NAND2_X1 U14227 ( .A1(n11440), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11384) );
  INV_X1 U14228 ( .A(n11377), .ZN(n11378) );
  NAND2_X1 U14229 ( .A1(n11378), .A2(n19943), .ZN(n11912) );
  INV_X1 U14230 ( .A(n11385), .ZN(n11382) );
  NAND2_X1 U14231 ( .A1(n11395), .A2(n12359), .ZN(n12742) );
  NOR2_X1 U14232 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13348) );
  AOI22_X1 U14233 ( .A1(n15928), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n13348), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11383) );
  NAND2_X1 U14234 ( .A1(n11384), .A2(n11383), .ZN(n11422) );
  INV_X1 U14235 ( .A(n11386), .ZN(n12098) );
  NAND2_X1 U14236 ( .A1(n12098), .A2(n12350), .ZN(n11390) );
  INV_X1 U14237 ( .A(n11915), .ZN(n11388) );
  NAND2_X1 U14238 ( .A1(n11390), .A2(n11389), .ZN(n11393) );
  INV_X1 U14239 ( .A(n11391), .ZN(n11392) );
  AND2_X1 U14240 ( .A1(n14263), .A2(n12359), .ZN(n11937) );
  INV_X1 U14241 ( .A(n13349), .ZN(n11394) );
  NAND2_X1 U14242 ( .A1(n11395), .A2(n11396), .ZN(n11401) );
  NAND2_X1 U14243 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11398) );
  XNOR2_X1 U14244 ( .A(n11422), .B(n11423), .ZN(n11459) );
  INV_X1 U14245 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15923) );
  INV_X1 U14246 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n11406) );
  INV_X1 U14247 ( .A(n13348), .ZN(n11417) );
  NAND2_X1 U14248 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11402) );
  NAND2_X1 U14249 ( .A1(n11417), .A2(n11402), .ZN(n11403) );
  AOI21_X1 U14250 ( .B1(n12012), .B2(P2_EBX_REG_0__SCAN_IN), .A(n11403), .ZN(
        n11404) );
  OAI211_X1 U14251 ( .C1(n11401), .C2(n11406), .A(n11405), .B(n11404), .ZN(
        n11407) );
  INV_X1 U14252 ( .A(n11407), .ZN(n11414) );
  NAND2_X1 U14253 ( .A1(n11409), .A2(n11408), .ZN(n12347) );
  INV_X1 U14254 ( .A(n11410), .ZN(n11411) );
  NAND2_X1 U14255 ( .A1(n12347), .A2(n11411), .ZN(n11412) );
  NAND2_X1 U14256 ( .A1(n11412), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11413) );
  INV_X1 U14257 ( .A(n11416), .ZN(n11419) );
  NOR2_X1 U14258 ( .A1(n11417), .A2(n19931), .ZN(n11418) );
  AOI21_X1 U14259 ( .B1(n11419), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11418), 
        .ZN(n11420) );
  NAND2_X1 U14260 ( .A1(n11421), .A2(n11420), .ZN(n11451) );
  NAND2_X1 U14261 ( .A1(n11450), .A2(n11451), .ZN(n11457) );
  NAND2_X1 U14262 ( .A1(n11459), .A2(n11457), .ZN(n11454) );
  INV_X1 U14263 ( .A(n11422), .ZN(n11424) );
  NAND2_X1 U14264 ( .A1(n11424), .A2(n11423), .ZN(n11425) );
  AND2_X2 U14265 ( .A1(n11426), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11443) );
  AOI22_X1 U14266 ( .A1(n12012), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11427) );
  INV_X1 U14267 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n11428) );
  NAND2_X1 U14268 ( .A1(n11440), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11434) );
  AOI21_X1 U14269 ( .B1(n16510), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11433) );
  NAND2_X1 U14270 ( .A1(n11434), .A2(n11433), .ZN(n11436) );
  NAND2_X1 U14271 ( .A1(n11436), .A2(n11435), .ZN(n11437) );
  NAND2_X1 U14272 ( .A1(n11449), .A2(n11448), .ZN(n11439) );
  NAND2_X1 U14273 ( .A1(n11440), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11442) );
  NAND2_X1 U14274 ( .A1(n13348), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11441) );
  INV_X1 U14275 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n11446) );
  NAND2_X1 U14276 ( .A1(n12076), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n11445) );
  NAND2_X1 U14277 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11444) );
  OAI211_X1 U14278 ( .C1(n11401), .C2(n11446), .A(n11445), .B(n11444), .ZN(
        n11447) );
  XNOR2_X1 U14279 ( .A(n11449), .B(n11448), .ZN(n12930) );
  INV_X1 U14280 ( .A(n11458), .ZN(n11455) );
  OR2_X1 U14281 ( .A1(n11455), .A2(n11454), .ZN(n11486) );
  INV_X1 U14282 ( .A(n12982), .ZN(n11456) );
  BUF_X1 U14283 ( .A(n11459), .Z(n11465) );
  INV_X1 U14284 ( .A(n11465), .ZN(n11460) );
  NAND2_X1 U14285 ( .A1(n12816), .A2(n11460), .ZN(n11483) );
  INV_X1 U14286 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11461) );
  OAI22_X1 U14287 ( .A1(n11462), .A2(n19399), .B1(n19462), .B2(n11461), .ZN(
        n11468) );
  INV_X1 U14288 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14174) );
  INV_X1 U14289 ( .A(n19295), .ZN(n11463) );
  XNOR2_X2 U14290 ( .A(n11465), .B(n11464), .ZN(n15917) );
  INV_X1 U14291 ( .A(n12816), .ZN(n12889) );
  NAND2_X1 U14292 ( .A1(n15917), .A2(n12889), .ZN(n11482) );
  INV_X1 U14293 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13728) );
  OAI22_X1 U14294 ( .A1(n14174), .A2(n19349), .B1(n19605), .B2(n13728), .ZN(
        n11467) );
  NOR2_X1 U14295 ( .A1(n11468), .A2(n11467), .ZN(n11497) );
  INV_X1 U14296 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11469) );
  INV_X1 U14297 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12828) );
  OAI22_X1 U14298 ( .A1(n11469), .A2(n19425), .B1(n19300), .B2(n12828), .ZN(
        n11473) );
  INV_X1 U14299 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11471) );
  INV_X1 U14300 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12169) );
  OAI22_X1 U14301 ( .A1(n11612), .A2(n11471), .B1(n19537), .B2(n12169), .ZN(
        n11472) );
  NOR2_X1 U14302 ( .A1(n11473), .A2(n11472), .ZN(n11496) );
  INV_X1 U14303 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11477) );
  NAND2_X1 U14304 ( .A1(n19295), .A2(n12982), .ZN(n11489) );
  INV_X1 U14305 ( .A(n11489), .ZN(n11474) );
  INV_X1 U14306 ( .A(n11616), .ZN(n11475) );
  NAND2_X1 U14307 ( .A1(n11475), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11476) );
  OAI211_X1 U14308 ( .C1(n19627), .C2(n11477), .A(n11476), .B(n19944), .ZN(
        n11481) );
  INV_X1 U14309 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13731) );
  INV_X1 U14310 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11479) );
  OAI22_X1 U14311 ( .A1(n13731), .A2(n13931), .B1(n11608), .B2(n11479), .ZN(
        n11480) );
  NOR2_X1 U14312 ( .A1(n11481), .A2(n11480), .ZN(n11495) );
  INV_X1 U14313 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11485) );
  INV_X1 U14314 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14181) );
  OAI22_X1 U14315 ( .A1(n11485), .A2(n11615), .B1(n19572), .B2(n14181), .ZN(
        n11493) );
  INV_X1 U14316 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11491) );
  INV_X1 U14317 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11490) );
  OAI22_X1 U14318 ( .A1(n11491), .A2(n13709), .B1(n11603), .B2(n11490), .ZN(
        n11492) );
  NOR2_X1 U14319 ( .A1(n11493), .A2(n11492), .ZN(n11494) );
  NAND4_X1 U14320 ( .A1(n11497), .A2(n11496), .A3(n11495), .A4(n11494), .ZN(
        n11550) );
  INV_X1 U14321 ( .A(n11498), .ZN(n11499) );
  AND2_X2 U14322 ( .A1(n14128), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14161) );
  AND2_X2 U14323 ( .A1(n14311), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12262) );
  AOI22_X1 U14324 ( .A1(n12262), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U14325 ( .A1(n11588), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12292), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11502) );
  NAND3_X1 U14326 ( .A1(n11503), .A2(n11502), .A3(n11501), .ZN(n11506) );
  INV_X1 U14327 ( .A(n11355), .ZN(n13266) );
  AND2_X2 U14328 ( .A1(n14325), .A2(n20841), .ZN(n14156) );
  AOI22_X1 U14329 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11504) );
  INV_X1 U14330 ( .A(n11504), .ZN(n11505) );
  NOR2_X1 U14331 ( .A1(n11506), .A2(n11505), .ZN(n11507) );
  NAND2_X1 U14332 ( .A1(n11508), .A2(n11507), .ZN(n11522) );
  AND2_X1 U14333 ( .A1(n11509), .A2(n14129), .ZN(n11528) );
  NOR2_X1 U14334 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U14335 ( .A1(n11528), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11520) );
  AND2_X1 U14336 ( .A1(n11511), .A2(n14129), .ZN(n11537) );
  AND2_X1 U14337 ( .A1(n14129), .A2(n11512), .ZN(n11513) );
  AOI22_X1 U14338 ( .A1(n11537), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11513), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11519) );
  AND2_X2 U14339 ( .A1(n14312), .A2(n20841), .ZN(n14162) );
  INV_X2 U14340 ( .A(n14310), .ZN(n11516) );
  AND2_X2 U14341 ( .A1(n11516), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11529) );
  AOI22_X1 U14342 ( .A1(n14162), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11518) );
  AND2_X2 U14343 ( .A1(n11516), .A2(n20841), .ZN(n11523) );
  AOI22_X1 U14344 ( .A1(n14155), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11523), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11517) );
  NAND4_X1 U14345 ( .A1(n11520), .A2(n11519), .A3(n11518), .A4(n11517), .ZN(
        n11521) );
  AOI22_X1 U14346 ( .A1(n14162), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n11523), .ZN(n11527) );
  AOI22_X1 U14347 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11571), .B1(
        n12262), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14348 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n14161), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11525) );
  AOI22_X1 U14349 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11588), .B1(
        n11575), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11524) );
  NAND4_X1 U14350 ( .A1(n11527), .A2(n11526), .A3(n11525), .A4(n11524), .ZN(
        n11535) );
  AOI22_X1 U14351 ( .A1(n11537), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11513), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14352 ( .A1(n11528), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U14353 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n14155), .B1(
        n13998), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U14354 ( .A1(n12292), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11530) );
  NAND4_X1 U14355 ( .A1(n11533), .A2(n11532), .A3(n11531), .A4(n11530), .ZN(
        n11534) );
  NOR2_X1 U14356 ( .A1(n12880), .A2(n12112), .ZN(n11536) );
  NAND2_X1 U14357 ( .A1(n14263), .A2(n11536), .ZN(n11950) );
  AOI22_X1 U14358 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n11529), .B1(
        n13998), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11539) );
  AOI22_X1 U14359 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n11528), .B1(
        n11537), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14360 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11588), .B1(
        n11575), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11547) );
  INV_X1 U14361 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11542) );
  NAND2_X1 U14362 ( .A1(n14163), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11541) );
  NAND2_X1 U14363 ( .A1(n11513), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11540) );
  OAI211_X1 U14364 ( .C1(n14153), .C2(n11542), .A(n11541), .B(n11540), .ZN(
        n11543) );
  INV_X1 U14365 ( .A(n11543), .ZN(n11546) );
  AOI22_X1 U14366 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n14161), .B1(
        n14155), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U14367 ( .A1(n14162), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11544) );
  NAND4_X1 U14368 ( .A1(n11547), .A2(n11546), .A3(n11545), .A4(n11544), .ZN(
        n11548) );
  NAND2_X1 U14369 ( .A1(n11950), .A2(n12117), .ZN(n11549) );
  NAND2_X1 U14370 ( .A1(n11550), .A2(n11549), .ZN(n11683) );
  INV_X1 U14371 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14009) );
  INV_X1 U14372 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14006) );
  OAI22_X1 U14373 ( .A1(n14009), .A2(n13931), .B1(n19605), .B2(n14006), .ZN(
        n11554) );
  INV_X1 U14374 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11552) );
  INV_X1 U14375 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11551) );
  NOR2_X1 U14376 ( .A1(n11554), .A2(n11553), .ZN(n11570) );
  INV_X1 U14377 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14003) );
  INV_X1 U14378 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12202) );
  OAI22_X1 U14379 ( .A1(n14003), .A2(n11615), .B1(n11616), .B2(n12202), .ZN(
        n11557) );
  INV_X1 U14380 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11555) );
  INV_X1 U14381 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14227) );
  OAI22_X1 U14382 ( .A1(n13709), .A2(n11555), .B1(n19572), .B2(n14227), .ZN(
        n11556) );
  NOR2_X1 U14383 ( .A1(n11557), .A2(n11556), .ZN(n11569) );
  INV_X1 U14384 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11558) );
  INV_X1 U14385 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12206) );
  OAI22_X1 U14386 ( .A1(n11558), .A2(n19399), .B1(n19300), .B2(n12206), .ZN(
        n11561) );
  INV_X1 U14387 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11559) );
  INV_X1 U14388 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14220) );
  OAI22_X1 U14389 ( .A1(n11559), .A2(n19462), .B1(n19349), .B2(n14220), .ZN(
        n11560) );
  NOR2_X1 U14390 ( .A1(n11561), .A2(n11560), .ZN(n11568) );
  INV_X1 U14391 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11563) );
  INV_X1 U14392 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11562) );
  OAI22_X1 U14393 ( .A1(n11612), .A2(n11563), .B1(n11603), .B2(n11562), .ZN(
        n11566) );
  INV_X1 U14394 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11564) );
  INV_X1 U14395 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12203) );
  OAI22_X1 U14396 ( .A1(n11564), .A2(n19425), .B1(n19537), .B2(n12203), .ZN(
        n11565) );
  NOR2_X1 U14397 ( .A1(n11566), .A2(n11565), .ZN(n11567) );
  NAND4_X1 U14398 ( .A1(n11570), .A2(n11569), .A3(n11568), .A4(n11567), .ZN(
        n11587) );
  AOI22_X1 U14399 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n11571), .B1(
        n12262), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11579) );
  NAND2_X1 U14400 ( .A1(n11513), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11573) );
  NAND2_X1 U14401 ( .A1(n11537), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11572) );
  OAI211_X1 U14402 ( .C1(n14153), .C2(n12206), .A(n11573), .B(n11572), .ZN(
        n11574) );
  INV_X1 U14403 ( .A(n11574), .ZN(n11578) );
  AOI22_X1 U14404 ( .A1(n11588), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__3__SCAN_IN), .B2(n14155), .ZN(n11577) );
  AOI22_X1 U14405 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11576) );
  NAND4_X1 U14406 ( .A1(n11579), .A2(n11578), .A3(n11577), .A4(n11576), .ZN(
        n11585) );
  AOI22_X1 U14407 ( .A1(n14162), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14161), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14408 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11523), .B1(
        n13998), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14409 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n11528), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11581) );
  NAND2_X1 U14410 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11580) );
  NAND4_X1 U14411 ( .A1(n11583), .A2(n11582), .A3(n11581), .A4(n11580), .ZN(
        n11584) );
  INV_X1 U14412 ( .A(n11674), .ZN(n12125) );
  NAND2_X1 U14413 ( .A1(n12125), .A2(n14263), .ZN(n11586) );
  INV_X1 U14414 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n20934) );
  AOI22_X1 U14415 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11588), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U14416 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12262), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11594) );
  INV_X1 U14417 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12220) );
  NAND2_X1 U14418 ( .A1(n11513), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11590) );
  NAND2_X1 U14419 ( .A1(n11537), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11589) );
  OAI211_X1 U14420 ( .C1(n14153), .C2(n12220), .A(n11590), .B(n11589), .ZN(
        n11591) );
  INV_X1 U14421 ( .A(n11591), .ZN(n11593) );
  AOI22_X1 U14422 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14155), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11592) );
  NAND4_X1 U14423 ( .A1(n11595), .A2(n11594), .A3(n11593), .A4(n11592), .ZN(
        n11601) );
  AOI22_X1 U14424 ( .A1(n14162), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14161), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U14425 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11529), .B1(
        n13998), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U14426 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11528), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11597) );
  NAND2_X1 U14427 ( .A1(n11523), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11596) );
  NAND4_X1 U14428 ( .A1(n11599), .A2(n11598), .A3(n11597), .A4(n11596), .ZN(
        n11600) );
  INV_X1 U14429 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11602) );
  INV_X1 U14430 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14274) );
  OAI22_X1 U14431 ( .A1(n11602), .A2(n13709), .B1(n19572), .B2(n14274), .ZN(
        n11607) );
  INV_X1 U14432 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11605) );
  INV_X1 U14433 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11604) );
  OAI22_X1 U14434 ( .A1(n11605), .A2(n19399), .B1(n11603), .B2(n11604), .ZN(
        n11606) );
  NOR2_X1 U14435 ( .A1(n11607), .A2(n11606), .ZN(n11626) );
  INV_X1 U14436 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14267) );
  INV_X1 U14437 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13002) );
  OAI22_X1 U14438 ( .A1(n14267), .A2(n19349), .B1(n19300), .B2(n13002), .ZN(
        n11611) );
  INV_X1 U14439 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14104) );
  INV_X1 U14440 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11609) );
  OAI22_X1 U14441 ( .A1(n14104), .A2(n13931), .B1(n11608), .B2(n11609), .ZN(
        n11610) );
  NOR2_X1 U14442 ( .A1(n11611), .A2(n11610), .ZN(n11625) );
  INV_X1 U14443 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11614) );
  INV_X1 U14444 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11613) );
  OAI22_X1 U14445 ( .A1(n11614), .A2(n19425), .B1(n11612), .B2(n11613), .ZN(
        n11618) );
  INV_X1 U14446 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14094) );
  INV_X1 U14447 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12241) );
  OAI22_X1 U14448 ( .A1(n14094), .A2(n11615), .B1(n11616), .B2(n12241), .ZN(
        n11617) );
  NOR2_X1 U14449 ( .A1(n11618), .A2(n11617), .ZN(n11624) );
  INV_X1 U14450 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11619) );
  INV_X1 U14451 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12242) );
  OAI22_X1 U14452 ( .A1(n11619), .A2(n19462), .B1(n19537), .B2(n12242), .ZN(
        n11622) );
  INV_X1 U14453 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11620) );
  INV_X1 U14454 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14100) );
  OAI22_X1 U14455 ( .A1(n11620), .A2(n19627), .B1(n19605), .B2(n14100), .ZN(
        n11621) );
  NOR2_X1 U14456 ( .A1(n11622), .A2(n11621), .ZN(n11623) );
  NAND4_X1 U14457 ( .A1(n11626), .A2(n11625), .A3(n11624), .A4(n11623), .ZN(
        n11641) );
  AOI22_X1 U14458 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11588), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11633) );
  AOI22_X1 U14459 ( .A1(n12262), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11632) );
  NAND2_X1 U14460 ( .A1(n11513), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11628) );
  NAND2_X1 U14461 ( .A1(n11537), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11627) );
  OAI211_X1 U14462 ( .C1(n14153), .C2(n13002), .A(n11628), .B(n11627), .ZN(
        n11629) );
  INV_X1 U14463 ( .A(n11629), .ZN(n11631) );
  AOI22_X1 U14464 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14155), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11630) );
  NAND4_X1 U14465 ( .A1(n11633), .A2(n11632), .A3(n11631), .A4(n11630), .ZN(
        n11639) );
  AOI22_X1 U14466 ( .A1(n14162), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14161), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11637) );
  AOI22_X1 U14467 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13998), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U14468 ( .A1(n11528), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11635) );
  NAND2_X1 U14469 ( .A1(n11523), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11634) );
  NAND4_X1 U14470 ( .A1(n11637), .A2(n11636), .A3(n11635), .A4(n11634), .ZN(
        n11638) );
  INV_X1 U14471 ( .A(n11680), .ZN(n12089) );
  NAND2_X1 U14472 ( .A1(n12089), .A2(n14263), .ZN(n11640) );
  NAND2_X1 U14473 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11645) );
  NAND2_X1 U14474 ( .A1(n14162), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11644) );
  NAND2_X1 U14475 ( .A1(n11588), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11643) );
  NAND2_X1 U14476 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11642) );
  AOI22_X1 U14477 ( .A1(n11571), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14161), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11656) );
  NAND2_X1 U14478 ( .A1(n12262), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11649) );
  AOI22_X1 U14479 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n11537), .B1(
        n11513), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11648) );
  NAND2_X1 U14480 ( .A1(n12292), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11647) );
  NAND2_X1 U14481 ( .A1(n14155), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11646) );
  AOI22_X1 U14482 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n11528), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11653) );
  NAND2_X1 U14483 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11652) );
  NAND2_X1 U14484 ( .A1(n13998), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11651) );
  NAND2_X1 U14485 ( .A1(n11523), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11650) );
  NAND2_X1 U14486 ( .A1(n11960), .A2(n12139), .ZN(n11681) );
  NAND2_X1 U14487 ( .A1(n19922), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11660) );
  NAND2_X1 U14488 ( .A1(n11256), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11659) );
  NAND2_X1 U14489 ( .A1(n11660), .A2(n11659), .ZN(n11881) );
  NAND2_X1 U14490 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19931), .ZN(
        n11880) );
  NAND2_X1 U14491 ( .A1(n13290), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11661) );
  NAND2_X1 U14492 ( .A1(n11672), .A2(n11661), .ZN(n11663) );
  NAND2_X1 U14493 ( .A1(n11662), .A2(n11663), .ZN(n11666) );
  INV_X1 U14494 ( .A(n11663), .ZN(n11664) );
  INV_X1 U14495 ( .A(n11900), .ZN(n11667) );
  INV_X1 U14496 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n11670) );
  INV_X1 U14497 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n12824) );
  NAND2_X1 U14498 ( .A1(n11670), .A2(n12824), .ZN(n11671) );
  MUX2_X1 U14499 ( .A(n12112), .B(n11671), .S(n19325), .Z(n11694) );
  XNOR2_X1 U14500 ( .A(n11675), .B(n11676), .ZN(n11890) );
  MUX2_X1 U14501 ( .A(n11674), .B(n11890), .S(n13635), .Z(n11933) );
  INV_X1 U14502 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n21011) );
  MUX2_X1 U14503 ( .A(n11933), .B(n21011), .S(n19325), .Z(n11688) );
  NAND3_X1 U14504 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n11878), .A3(
        n20966), .ZN(n11891) );
  MUX2_X1 U14505 ( .A(n11891), .B(n11955), .S(n11679), .Z(n11932) );
  INV_X1 U14506 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n19163) );
  MUX2_X1 U14507 ( .A(n11932), .B(n19163), .S(n19325), .Z(n11700) );
  INV_X1 U14508 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n19108) );
  MUX2_X1 U14509 ( .A(n11680), .B(n19108), .S(n19325), .Z(n11755) );
  XNOR2_X1 U14510 ( .A(n11756), .B(n11755), .ZN(n19106) );
  INV_X1 U14511 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n20980) );
  INV_X1 U14512 ( .A(n11682), .ZN(n11684) );
  NAND2_X1 U14513 ( .A1(n11684), .A2(n11683), .ZN(n11685) );
  INV_X1 U14514 ( .A(n11701), .ZN(n11686) );
  OAI21_X1 U14515 ( .B1(n11688), .B2(n11687), .A(n11686), .ZN(n13641) );
  OAI21_X2 U14516 ( .B1(n11947), .B2(n11763), .A(n13641), .ZN(n13357) );
  OAI21_X1 U14517 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19931), .A(
        n11880), .ZN(n11905) );
  MUX2_X1 U14518 ( .A(n12880), .B(n11905), .S(n13635), .Z(n11931) );
  AND2_X1 U14519 ( .A1(n19325), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n11691) );
  INV_X1 U14520 ( .A(n11691), .ZN(n11690) );
  OAI21_X1 U14521 ( .B1(n11931), .B2(n19325), .A(n11690), .ZN(n19124) );
  NAND2_X1 U14522 ( .A1(n19124), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12877) );
  NAND2_X1 U14523 ( .A1(n11691), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n11692) );
  NAND2_X1 U14524 ( .A1(n11694), .A2(n11692), .ZN(n15381) );
  NOR2_X1 U14525 ( .A1(n12877), .A2(n15381), .ZN(n11693) );
  INV_X1 U14526 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15914) );
  XNOR2_X1 U14527 ( .A(n15381), .B(n12877), .ZN(n15622) );
  NOR2_X1 U14528 ( .A1(n15914), .A2(n15622), .ZN(n15621) );
  NOR2_X1 U14529 ( .A1(n11693), .A2(n15621), .ZN(n12904) );
  XNOR2_X1 U14530 ( .A(n11695), .B(n11694), .ZN(n15370) );
  NAND2_X1 U14531 ( .A1(n12904), .A2(n15370), .ZN(n11696) );
  NAND2_X1 U14532 ( .A1(n11696), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11697) );
  OR2_X1 U14533 ( .A1(n12904), .A2(n15370), .ZN(n12902) );
  NAND2_X1 U14534 ( .A1(n11697), .A2(n12902), .ZN(n13355) );
  OAI21_X1 U14535 ( .B1(n13357), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n13355), .ZN(n11699) );
  NAND2_X1 U14536 ( .A1(n13357), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11698) );
  NAND2_X1 U14537 ( .A1(n11699), .A2(n11698), .ZN(n13515) );
  XNOR2_X1 U14538 ( .A(n11701), .B(n11700), .ZN(n11702) );
  XNOR2_X1 U14539 ( .A(n11702), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13514) );
  NAND2_X1 U14540 ( .A1(n13515), .A2(n13514), .ZN(n11704) );
  INV_X1 U14541 ( .A(n11702), .ZN(n15357) );
  NAND2_X1 U14542 ( .A1(n15357), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11703) );
  NAND2_X1 U14543 ( .A1(n11704), .A2(n11703), .ZN(n13687) );
  NAND2_X1 U14544 ( .A1(n13686), .A2(n13687), .ZN(n11707) );
  NAND2_X1 U14545 ( .A1(n11705), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11706) );
  NAND2_X1 U14546 ( .A1(n11707), .A2(n11706), .ZN(n13766) );
  INV_X1 U14547 ( .A(n11958), .ZN(n11709) );
  NAND2_X1 U14548 ( .A1(n11709), .A2(n11708), .ZN(n11970) );
  INV_X1 U14549 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11711) );
  INV_X1 U14550 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11710) );
  OAI22_X1 U14551 ( .A1(n11711), .A2(n11615), .B1(n11616), .B2(n11710), .ZN(
        n11715) );
  INV_X1 U14552 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11713) );
  INV_X1 U14553 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11712) );
  OAI22_X1 U14554 ( .A1(n11713), .A2(n13709), .B1(n19572), .B2(n11712), .ZN(
        n11714) );
  NOR2_X1 U14555 ( .A1(n11715), .A2(n11714), .ZN(n11733) );
  INV_X1 U14556 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11717) );
  INV_X1 U14557 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11716) );
  OAI22_X1 U14558 ( .A1(n11717), .A2(n11612), .B1(n11603), .B2(n11716), .ZN(
        n11719) );
  INV_X1 U14559 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14285) );
  INV_X1 U14560 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12263) );
  OAI22_X1 U14561 ( .A1(n14285), .A2(n19425), .B1(n19537), .B2(n12263), .ZN(
        n11718) );
  NOR2_X1 U14562 ( .A1(n11719), .A2(n11718), .ZN(n11732) );
  INV_X1 U14563 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11721) );
  INV_X1 U14564 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11720) );
  OAI22_X1 U14565 ( .A1(n11721), .A2(n19399), .B1(n19300), .B2(n11720), .ZN(
        n11725) );
  INV_X1 U14566 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11723) );
  INV_X1 U14567 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11722) );
  OAI22_X1 U14568 ( .A1(n11723), .A2(n19349), .B1(n19462), .B2(n11722), .ZN(
        n11724) );
  NOR2_X1 U14569 ( .A1(n11725), .A2(n11724), .ZN(n11731) );
  INV_X1 U14570 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14113) );
  INV_X1 U14571 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11726) );
  OAI22_X1 U14572 ( .A1(n14113), .A2(n13931), .B1(n19605), .B2(n11726), .ZN(
        n11729) );
  INV_X1 U14573 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11727) );
  INV_X1 U14574 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14295) );
  OAI22_X1 U14575 ( .A1(n11727), .A2(n19627), .B1(n11608), .B2(n14295), .ZN(
        n11728) );
  NOR2_X1 U14576 ( .A1(n11729), .A2(n11728), .ZN(n11730) );
  NAND4_X1 U14577 ( .A1(n11733), .A2(n11732), .A3(n11731), .A4(n11730), .ZN(
        n11754) );
  NAND2_X1 U14578 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11735) );
  NAND2_X1 U14579 ( .A1(n11588), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11734) );
  AND2_X1 U14580 ( .A1(n11735), .A2(n11734), .ZN(n11743) );
  AOI22_X1 U14581 ( .A1(n14162), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11742) );
  NAND2_X1 U14582 ( .A1(n14155), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11737) );
  NAND2_X1 U14583 ( .A1(n14163), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11736) );
  OAI211_X1 U14584 ( .C1(n11738), .C2(n14285), .A(n11737), .B(n11736), .ZN(
        n11739) );
  INV_X1 U14585 ( .A(n11739), .ZN(n11741) );
  AOI22_X1 U14586 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12292), .B1(
        n14161), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11740) );
  NAND4_X1 U14587 ( .A1(n11743), .A2(n11742), .A3(n11741), .A4(n11740), .ZN(
        n11752) );
  AOI22_X1 U14588 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11523), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11750) );
  NAND2_X1 U14589 ( .A1(n9741), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11746) );
  NAND2_X1 U14590 ( .A1(n11528), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11745) );
  NAND2_X1 U14591 ( .A1(n11537), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11744) );
  AND3_X1 U14592 ( .A1(n11746), .A2(n11745), .A3(n11744), .ZN(n11749) );
  NAND2_X1 U14593 ( .A1(n12262), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11748) );
  NAND2_X1 U14594 ( .A1(n11571), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11747) );
  NAND4_X1 U14595 ( .A1(n11750), .A2(n11749), .A3(n11748), .A4(n11747), .ZN(
        n11751) );
  NAND2_X1 U14596 ( .A1(n12135), .A2(n14263), .ZN(n11753) );
  XNOR2_X1 U14597 ( .A(n11970), .B(n11971), .ZN(n11961) );
  NAND2_X1 U14598 ( .A1(n11961), .A2(n12139), .ZN(n11757) );
  MUX2_X1 U14599 ( .A(n12135), .B(P2_EBX_REG_6__SCAN_IN), .S(n19325), .Z(
        n11761) );
  XNOR2_X1 U14600 ( .A(n11762), .B(n11761), .ZN(n19092) );
  NAND2_X1 U14601 ( .A1(n11757), .A2(n19092), .ZN(n11758) );
  INV_X1 U14602 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16471) );
  NAND2_X1 U14603 ( .A1(n13766), .A2(n13767), .ZN(n11760) );
  NAND2_X1 U14604 ( .A1(n11758), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11759) );
  INV_X1 U14605 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12996) );
  MUX2_X1 U14606 ( .A(n11763), .B(n12996), .S(n19325), .Z(n11768) );
  INV_X1 U14607 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n11764) );
  NAND2_X1 U14608 ( .A1(n11771), .A2(n11764), .ZN(n11765) );
  NAND2_X1 U14609 ( .A1(n19325), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11766) );
  NOR2_X1 U14610 ( .A1(n11771), .A2(n11766), .ZN(n11767) );
  OR2_X1 U14611 ( .A1(n11775), .A2(n11767), .ZN(n15345) );
  OR2_X1 U14612 ( .A1(n15345), .A2(n12139), .ZN(n11772) );
  INV_X1 U14613 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16472) );
  NOR2_X1 U14614 ( .A1(n11772), .A2(n16472), .ZN(n16399) );
  NOR2_X1 U14615 ( .A1(n11769), .A2(n11768), .ZN(n11770) );
  OR2_X1 U14616 ( .A1(n11771), .A2(n11770), .ZN(n19082) );
  INV_X1 U14617 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16482) );
  NOR2_X1 U14618 ( .A1(n19082), .A2(n16482), .ZN(n13910) );
  NAND2_X1 U14619 ( .A1(n11772), .A2(n16472), .ZN(n16400) );
  NAND2_X1 U14620 ( .A1(n19082), .A2(n16482), .ZN(n16396) );
  AND2_X1 U14621 ( .A1(n16400), .A2(n16396), .ZN(n11773) );
  AND2_X1 U14622 ( .A1(n19325), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11774) );
  XNOR2_X1 U14623 ( .A(n11775), .B(n11774), .ZN(n19071) );
  NAND2_X1 U14624 ( .A1(n19071), .A2(n11763), .ZN(n11786) );
  INV_X1 U14625 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15820) );
  AND2_X1 U14626 ( .A1(n11786), .A2(n15820), .ZN(n15898) );
  INV_X1 U14627 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n21042) );
  INV_X1 U14628 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n11776) );
  INV_X1 U14629 ( .A(n11851), .ZN(n11780) );
  NAND2_X1 U14630 ( .A1(n19325), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11777) );
  NOR2_X1 U14631 ( .A1(n11778), .A2(n11777), .ZN(n11779) );
  OR3_X1 U14632 ( .A1(n11782), .A2(n11780), .A3(n11779), .ZN(n19058) );
  INV_X1 U14633 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16380) );
  OAI21_X1 U14634 ( .B1(n19058), .B2(n12139), .A(n16380), .ZN(n16374) );
  INV_X1 U14635 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n11781) );
  OR3_X1 U14636 ( .A1(n11782), .A2(n9720), .A3(n11781), .ZN(n11784) );
  INV_X1 U14637 ( .A(n11791), .ZN(n11783) );
  AOI21_X1 U14638 ( .B1(n15323), .B2(n11763), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15883) );
  AND2_X1 U14639 ( .A1(n11763), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11785) );
  NAND2_X1 U14640 ( .A1(n15323), .A2(n11785), .ZN(n15881) );
  OR2_X1 U14641 ( .A1(n11786), .A2(n15820), .ZN(n15897) );
  INV_X1 U14642 ( .A(n19058), .ZN(n11788) );
  AND2_X1 U14643 ( .A1(n11763), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11787) );
  NAND2_X1 U14644 ( .A1(n11788), .A2(n11787), .ZN(n16373) );
  AND3_X1 U14645 ( .A1(n15881), .A2(n15897), .A3(n16373), .ZN(n11789) );
  NAND2_X1 U14646 ( .A1(n19325), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11790) );
  NAND2_X1 U14647 ( .A1(n11791), .A2(n11790), .ZN(n11800) );
  NAND3_X1 U14648 ( .A1(n19325), .A2(n11792), .A3(P2_EBX_REG_12__SCAN_IN), 
        .ZN(n11793) );
  NAND2_X1 U14649 ( .A1(n11800), .A2(n11793), .ZN(n19049) );
  INV_X1 U14650 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11794) );
  NOR2_X1 U14651 ( .A1(n11795), .A2(n11794), .ZN(n15873) );
  NAND2_X1 U14652 ( .A1(n11795), .A2(n11794), .ZN(n15871) );
  OAI21_X1 U14653 ( .B1(n15870), .B2(n15873), .A(n15871), .ZN(n15841) );
  INV_X1 U14654 ( .A(n15841), .ZN(n11798) );
  AND2_X1 U14655 ( .A1(n19325), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11799) );
  INV_X1 U14656 ( .A(n11799), .ZN(n11796) );
  XNOR2_X1 U14657 ( .A(n11800), .B(n11796), .ZN(n19037) );
  NAND2_X1 U14658 ( .A1(n19037), .A2(n11763), .ZN(n11832) );
  INV_X1 U14659 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15846) );
  AND2_X1 U14660 ( .A1(n11832), .A2(n15846), .ZN(n15839) );
  AND2_X1 U14661 ( .A1(n19325), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11821) );
  NAND2_X1 U14662 ( .A1(n19325), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11813) );
  AND2_X1 U14663 ( .A1(n19325), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11808) );
  AND2_X1 U14664 ( .A1(n19325), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11805) );
  INV_X1 U14665 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n16293) );
  NAND3_X1 U14666 ( .A1(n11840), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n19325), 
        .ZN(n11801) );
  OAI211_X1 U14667 ( .C1(n11840), .C2(P2_EBX_REG_21__SCAN_IN), .A(n11801), .B(
        n11851), .ZN(n15278) );
  OR2_X1 U14668 ( .A1(n15278), .A2(n12139), .ZN(n11802) );
  INV_X1 U14669 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11836) );
  NAND2_X1 U14670 ( .A1(n11802), .A2(n11836), .ZN(n15567) );
  INV_X1 U14671 ( .A(n11807), .ZN(n11804) );
  NAND2_X1 U14672 ( .A1(n19325), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11803) );
  XNOR2_X1 U14673 ( .A(n11804), .B(n11803), .ZN(n18978) );
  NAND2_X1 U14674 ( .A1(n18978), .A2(n11763), .ZN(n11834) );
  INV_X1 U14675 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15761) );
  NAND2_X1 U14676 ( .A1(n11834), .A2(n15761), .ZN(n15753) );
  AND2_X1 U14677 ( .A1(n11811), .A2(n11805), .ZN(n11806) );
  OR2_X1 U14678 ( .A1(n11807), .A2(n11806), .ZN(n18994) );
  NOR2_X1 U14679 ( .A1(n18994), .A2(n12139), .ZN(n11826) );
  NOR2_X1 U14680 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n11826), .ZN(
        n15583) );
  NAND2_X1 U14681 ( .A1(n11809), .A2(n11808), .ZN(n11810) );
  AND2_X1 U14682 ( .A1(n11811), .A2(n11810), .ZN(n15279) );
  NOR2_X1 U14683 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n11827), .ZN(
        n16335) );
  NOR2_X1 U14684 ( .A1(n15583), .A2(n16335), .ZN(n15755) );
  AND2_X1 U14685 ( .A1(n15753), .A2(n15755), .ZN(n15574) );
  XNOR2_X1 U14686 ( .A(n11812), .B(n10021), .ZN(n19006) );
  NAND2_X1 U14687 ( .A1(n19006), .A2(n11763), .ZN(n11814) );
  INV_X1 U14688 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21013) );
  NAND2_X1 U14689 ( .A1(n11814), .A2(n21013), .ZN(n15594) );
  NAND3_X1 U14690 ( .A1(n11815), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n19325), 
        .ZN(n11816) );
  NAND3_X1 U14691 ( .A1(n11817), .A2(n11851), .A3(n11816), .ZN(n15312) );
  OR2_X1 U14692 ( .A1(n15312), .A2(n12139), .ZN(n11818) );
  XNOR2_X1 U14693 ( .A(n11818), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15602) );
  XNOR2_X1 U14694 ( .A(n11819), .B(n9818), .ZN(n19018) );
  NAND2_X1 U14695 ( .A1(n19018), .A2(n11763), .ZN(n11820) );
  INV_X1 U14696 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16446) );
  NAND2_X1 U14697 ( .A1(n11820), .A2(n16446), .ZN(n15612) );
  INV_X1 U14698 ( .A(n11821), .ZN(n11822) );
  XNOR2_X1 U14699 ( .A(n11823), .B(n11822), .ZN(n19027) );
  NAND2_X1 U14700 ( .A1(n19027), .A2(n11763), .ZN(n11824) );
  INV_X1 U14701 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15834) );
  NAND2_X1 U14702 ( .A1(n11824), .A2(n15834), .ZN(n15814) );
  AND4_X1 U14703 ( .A1(n15594), .A2(n15602), .A3(n15612), .A4(n15814), .ZN(
        n11825) );
  NAND3_X1 U14704 ( .A1(n15567), .A2(n15574), .A3(n11825), .ZN(n11839) );
  NAND2_X1 U14705 ( .A1(n11826), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15585) );
  NAND2_X1 U14706 ( .A1(n11827), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16337) );
  AND2_X1 U14707 ( .A1(n15585), .A2(n16337), .ZN(n15573) );
  INV_X1 U14708 ( .A(n19006), .ZN(n11828) );
  INV_X1 U14709 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11829) );
  OR3_X1 U14710 ( .A1(n15312), .A2(n12139), .A3(n11829), .ZN(n15571) );
  INV_X1 U14711 ( .A(n19018), .ZN(n11830) );
  AND2_X1 U14712 ( .A1(n11763), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11831) );
  NAND2_X1 U14713 ( .A1(n19027), .A2(n11831), .ZN(n15813) );
  OR2_X1 U14714 ( .A1(n11832), .A2(n15846), .ZN(n15838) );
  AND4_X1 U14715 ( .A1(n15571), .A2(n15611), .A3(n15813), .A4(n15838), .ZN(
        n11833) );
  AND2_X1 U14716 ( .A1(n15593), .A2(n11833), .ZN(n11837) );
  INV_X1 U14717 ( .A(n11834), .ZN(n11835) );
  NAND2_X1 U14718 ( .A1(n11835), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15754) );
  OR3_X1 U14719 ( .A1(n15278), .A2(n12139), .A3(n11836), .ZN(n15566) );
  AND4_X1 U14720 ( .A1(n15573), .A2(n11837), .A3(n15754), .A4(n15566), .ZN(
        n11838) );
  AND2_X1 U14721 ( .A1(n19325), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11841) );
  AND2_X1 U14722 ( .A1(n11841), .A2(n10164), .ZN(n11842) );
  OR2_X1 U14723 ( .A1(n11846), .A2(n11842), .ZN(n15263) );
  OR2_X1 U14724 ( .A1(n15263), .A2(n12139), .ZN(n11843) );
  NAND2_X1 U14725 ( .A1(n11843), .A2(n15735), .ZN(n15729) );
  NAND2_X1 U14726 ( .A1(n11763), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11844) );
  OR2_X1 U14727 ( .A1(n15263), .A2(n11844), .ZN(n15728) );
  NAND2_X1 U14728 ( .A1(n19325), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11845) );
  NOR2_X1 U14729 ( .A1(n11846), .A2(n11845), .ZN(n11847) );
  XNOR2_X1 U14730 ( .A(n11848), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15558) );
  NAND2_X1 U14731 ( .A1(n11763), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11849) );
  NOR2_X1 U14732 ( .A1(n15249), .A2(n11849), .ZN(n11850) );
  INV_X1 U14733 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15705) );
  NOR2_X1 U14734 ( .A1(n10158), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15546) );
  INV_X1 U14735 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n15223) );
  INV_X1 U14736 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n15189) );
  NOR3_X1 U14737 ( .A1(n11852), .A2(n15189), .A3(n9720), .ZN(n11853) );
  NOR2_X1 U14738 ( .A1(n15093), .A2(n11853), .ZN(n11854) );
  INV_X1 U14739 ( .A(n11854), .ZN(n15200) );
  NOR2_X1 U14740 ( .A1(n15200), .A2(n12139), .ZN(n11855) );
  NAND3_X1 U14741 ( .A1(n11854), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n11763), .ZN(n11866) );
  OAI21_X1 U14742 ( .B1(n11855), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11866), .ZN(n15537) );
  NAND2_X1 U14743 ( .A1(n19325), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11856) );
  NAND2_X1 U14744 ( .A1(n11857), .A2(n10015), .ZN(n11858) );
  NAND2_X1 U14745 ( .A1(n11859), .A2(n11858), .ZN(n15184) );
  NOR2_X1 U14746 ( .A1(n15184), .A2(n12139), .ZN(n15518) );
  AND2_X1 U14747 ( .A1(n19325), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11860) );
  AOI21_X1 U14748 ( .B1(n11860), .B2(n11859), .A(n11872), .ZN(n15168) );
  NAND2_X1 U14749 ( .A1(n15168), .A2(n11763), .ZN(n15520) );
  INV_X1 U14750 ( .A(n15520), .ZN(n11861) );
  OAI21_X1 U14751 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n11861), .ZN(n11862) );
  NAND2_X1 U14752 ( .A1(n11863), .A2(n11862), .ZN(n11865) );
  INV_X1 U14753 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15519) );
  NAND2_X1 U14754 ( .A1(n15520), .A2(n15519), .ZN(n11864) );
  NAND2_X1 U14755 ( .A1(n11865), .A2(n11864), .ZN(n11868) );
  NAND2_X1 U14756 ( .A1(n10158), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15547) );
  NAND2_X1 U14757 ( .A1(n11866), .A2(n15547), .ZN(n15514) );
  INV_X1 U14758 ( .A(n15514), .ZN(n11867) );
  NAND2_X1 U14759 ( .A1(n11868), .A2(n11867), .ZN(n15504) );
  NAND2_X1 U14760 ( .A1(n19325), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11871) );
  INV_X1 U14761 ( .A(n11872), .ZN(n11869) );
  XOR2_X1 U14762 ( .A(n11871), .B(n11869), .Z(n11870) );
  INV_X1 U14763 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15642) );
  OAI21_X1 U14764 ( .B1(n11870), .B2(n12139), .A(n15642), .ZN(n15503) );
  NAND2_X1 U14765 ( .A1(n15504), .A2(n15503), .ZN(n15482) );
  INV_X1 U14766 ( .A(n11870), .ZN(n16277) );
  NAND3_X1 U14767 ( .A1(n16277), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11763), .ZN(n15502) );
  NAND2_X1 U14768 ( .A1(n15482), .A2(n15502), .ZN(n11876) );
  NAND2_X1 U14769 ( .A1(n19325), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11873) );
  AOI21_X1 U14770 ( .B1(n11874), .B2(n11763), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15481) );
  INV_X1 U14771 ( .A(n11874), .ZN(n15152) );
  INV_X1 U14772 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n20856) );
  NOR2_X1 U14773 ( .A1(n15481), .A2(n9803), .ZN(n11875) );
  XNOR2_X1 U14774 ( .A(n11876), .B(n11875), .ZN(n15501) );
  INV_X1 U14775 ( .A(n11903), .ZN(n11936) );
  NAND2_X1 U14776 ( .A1(n11895), .A2(n19944), .ZN(n11879) );
  MUX2_X1 U14777 ( .A(n11879), .B(n13635), .S(n11900), .Z(n11889) );
  NOR2_X1 U14778 ( .A1(n11881), .A2(n11905), .ZN(n11887) );
  INV_X1 U14779 ( .A(n11905), .ZN(n11884) );
  NAND2_X1 U14780 ( .A1(n11881), .A2(n11880), .ZN(n11928) );
  NAND2_X1 U14781 ( .A1(n11882), .A2(n11928), .ZN(n11901) );
  INV_X1 U14782 ( .A(n11901), .ZN(n11883) );
  OAI211_X1 U14783 ( .C1(n19944), .C2(n11884), .A(n19943), .B(n11883), .ZN(
        n11886) );
  NAND3_X1 U14784 ( .A1(n14263), .A2(n19943), .A3(n11900), .ZN(n11885) );
  OAI211_X1 U14785 ( .C1(n13635), .C2(n11887), .A(n11886), .B(n11885), .ZN(
        n11888) );
  NAND2_X1 U14786 ( .A1(n11889), .A2(n11888), .ZN(n11892) );
  MUX2_X1 U14787 ( .A(n13635), .B(n11892), .S(n11899), .Z(n11893) );
  NAND2_X1 U14788 ( .A1(n11936), .A2(n11893), .ZN(n11894) );
  MUX2_X1 U14789 ( .A(n11894), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n16510), .Z(n11897) );
  NAND2_X1 U14790 ( .A1(n11903), .A2(n11376), .ZN(n11896) );
  NAND2_X1 U14791 ( .A1(n13330), .A2(n19944), .ZN(n13282) );
  INV_X1 U14792 ( .A(n13682), .ZN(n12360) );
  NAND2_X1 U14793 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n16075) );
  INV_X1 U14794 ( .A(n16075), .ZN(n19952) );
  NOR2_X1 U14795 ( .A1(n18956), .A2(n19838), .ZN(n19831) );
  NAND2_X1 U14796 ( .A1(n18956), .A2(n19838), .ZN(n19833) );
  INV_X1 U14797 ( .A(n19833), .ZN(n19820) );
  NOR3_X1 U14798 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19831), .A3(n19820), 
        .ZN(n19825) );
  INV_X1 U14799 ( .A(n19825), .ZN(n19942) );
  NOR2_X1 U14800 ( .A1(n19952), .A2(n19942), .ZN(n13346) );
  NAND2_X1 U14801 ( .A1(n12360), .A2(n13346), .ZN(n11943) );
  AOI21_X1 U14802 ( .B1(n11897), .B2(n19943), .A(n13939), .ZN(n11898) );
  NAND2_X1 U14803 ( .A1(n13282), .A2(n11898), .ZN(n11942) );
  NAND2_X1 U14804 ( .A1(n11900), .A2(n11899), .ZN(n11904) );
  NOR2_X1 U14805 ( .A1(n11901), .A2(n11904), .ZN(n11902) );
  OR2_X1 U14806 ( .A1(n11903), .A2(n11902), .ZN(n12949) );
  INV_X1 U14807 ( .A(n12949), .ZN(n13322) );
  OAI21_X1 U14808 ( .B1(n11905), .B2(n11904), .A(n13322), .ZN(n11906) );
  INV_X1 U14809 ( .A(n11906), .ZN(n11908) );
  INV_X1 U14810 ( .A(n13272), .ZN(n11907) );
  NAND2_X1 U14811 ( .A1(n11907), .A2(n20966), .ZN(n15977) );
  INV_X1 U14812 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12750) );
  OAI21_X1 U14813 ( .B1(n12262), .B2(n15977), .A(n12750), .ZN(n19927) );
  MUX2_X1 U14814 ( .A(n11908), .B(n19927), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n16507) );
  NOR2_X1 U14815 ( .A1(n11946), .A2(n14263), .ZN(n11909) );
  NAND2_X1 U14816 ( .A1(n16507), .A2(n11909), .ZN(n11940) );
  NAND2_X1 U14817 ( .A1(n11395), .A2(n13346), .ZN(n11910) );
  OR2_X1 U14818 ( .A1(n12949), .A2(n11910), .ZN(n11924) );
  OAI21_X1 U14819 ( .B1(n11914), .B2(n12360), .A(n11913), .ZN(n11921) );
  NAND2_X1 U14820 ( .A1(n11915), .A2(n11364), .ZN(n11916) );
  NAND2_X1 U14821 ( .A1(n11916), .A2(n12957), .ZN(n11917) );
  NAND2_X1 U14822 ( .A1(n11917), .A2(n11937), .ZN(n12349) );
  NAND2_X1 U14823 ( .A1(n14263), .A2(n12358), .ZN(n12370) );
  NAND2_X1 U14824 ( .A1(n12370), .A2(n19943), .ZN(n11918) );
  NAND3_X1 U14825 ( .A1(n11918), .A2(n12350), .A3(n12957), .ZN(n11919) );
  NAND2_X1 U14826 ( .A1(n11919), .A2(n13682), .ZN(n11920) );
  NAND4_X1 U14827 ( .A1(n11922), .A2(n11921), .A3(n12349), .A4(n11920), .ZN(
        n12371) );
  INV_X1 U14828 ( .A(n12371), .ZN(n11923) );
  NAND2_X1 U14829 ( .A1(n11924), .A2(n11923), .ZN(n13278) );
  MUX2_X1 U14830 ( .A(n11395), .B(n12360), .S(n14263), .Z(n11925) );
  NAND2_X1 U14831 ( .A1(n11925), .A2(n16075), .ZN(n11926) );
  NOR2_X1 U14832 ( .A1(n12949), .A2(n11926), .ZN(n11927) );
  NOR2_X1 U14833 ( .A1(n13278), .A2(n11927), .ZN(n11939) );
  INV_X1 U14834 ( .A(n11928), .ZN(n11930) );
  OAI21_X1 U14835 ( .B1(n11931), .B2(n11930), .A(n11929), .ZN(n11934) );
  NAND3_X1 U14836 ( .A1(n11934), .A2(n11933), .A3(n11932), .ZN(n11935) );
  AND2_X1 U14837 ( .A1(n11936), .A2(n11935), .ZN(n13324) );
  INV_X1 U14838 ( .A(n11937), .ZN(n11938) );
  NOR2_X1 U14839 ( .A1(n11946), .A2(n11938), .ZN(n13320) );
  NAND2_X1 U14840 ( .A1(n13324), .A2(n13320), .ZN(n13335) );
  AND3_X1 U14841 ( .A1(n11940), .A2(n11939), .A3(n13335), .ZN(n11941) );
  OAI211_X1 U14842 ( .C1(n13282), .C2(n11943), .A(n11942), .B(n11941), .ZN(
        n11945) );
  NAND2_X1 U14843 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12874), .ZN(n13637) );
  INV_X1 U14844 ( .A(n13637), .ZN(n11944) );
  OR2_X1 U14845 ( .A1(n11946), .A2(n13635), .ZN(n13334) );
  INV_X1 U14846 ( .A(n11947), .ZN(n13368) );
  INV_X1 U14847 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12905) );
  NAND2_X1 U14848 ( .A1(n12880), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12879) );
  NOR2_X1 U14849 ( .A1(n12112), .A2(n12879), .ZN(n11949) );
  AND2_X1 U14850 ( .A1(n12880), .A2(n15923), .ZN(n11948) );
  XNOR2_X1 U14851 ( .A(n11948), .B(n12112), .ZN(n15625) );
  NOR2_X1 U14852 ( .A1(n15914), .A2(n15625), .ZN(n15624) );
  NOR2_X1 U14853 ( .A1(n11949), .A2(n15624), .ZN(n11951) );
  XNOR2_X1 U14854 ( .A(n11950), .B(n12117), .ZN(n12900) );
  NAND2_X1 U14855 ( .A1(n9794), .A2(n12900), .ZN(n12899) );
  OR2_X1 U14856 ( .A1(n11951), .A2(n12905), .ZN(n11952) );
  NAND2_X1 U14857 ( .A1(n12899), .A2(n11952), .ZN(n11953) );
  INV_X1 U14858 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13363) );
  XNOR2_X1 U14859 ( .A(n11953), .B(n13363), .ZN(n13367) );
  NAND2_X1 U14860 ( .A1(n11953), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11954) );
  NAND2_X1 U14861 ( .A1(n13366), .A2(n11954), .ZN(n13519) );
  INV_X1 U14862 ( .A(n11955), .ZN(n12131) );
  NAND2_X1 U14863 ( .A1(n11956), .A2(n12131), .ZN(n11957) );
  NAND2_X1 U14864 ( .A1(n11958), .A2(n11957), .ZN(n13517) );
  INV_X1 U14865 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13516) );
  INV_X1 U14866 ( .A(n11960), .ZN(n11959) );
  NAND2_X1 U14867 ( .A1(n11959), .A2(n20980), .ZN(n13688) );
  NAND2_X1 U14868 ( .A1(n11960), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13689) );
  NAND2_X1 U14869 ( .A1(n13692), .A2(n13689), .ZN(n11967) );
  INV_X1 U14870 ( .A(n11966), .ZN(n11965) );
  OR2_X1 U14871 ( .A1(n13689), .A2(n11971), .ZN(n11964) );
  NAND2_X1 U14872 ( .A1(n13765), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11969) );
  NAND2_X1 U14873 ( .A1(n11967), .A2(n11966), .ZN(n11968) );
  XNOR2_X1 U14874 ( .A(n11976), .B(n12139), .ZN(n13906) );
  INV_X1 U14875 ( .A(n13906), .ZN(n11973) );
  NAND2_X1 U14876 ( .A1(n11973), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11974) );
  XNOR2_X1 U14877 ( .A(n11975), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16393) );
  INV_X1 U14878 ( .A(n11976), .ZN(n11977) );
  NAND3_X1 U14879 ( .A1(n11977), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n11763), .ZN(n11978) );
  NAND2_X2 U14880 ( .A1(n11979), .A2(n11978), .ZN(n15598) );
  AND2_X1 U14881 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15888) );
  AND2_X1 U14882 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15599) );
  NAND2_X1 U14883 ( .A1(n15888), .A2(n15599), .ZN(n15830) );
  NAND2_X1 U14884 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11980) );
  NOR2_X1 U14885 ( .A1(n15830), .A2(n11980), .ZN(n15796) );
  NAND2_X1 U14886 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15790) );
  NOR2_X1 U14887 ( .A1(n15790), .A2(n21013), .ZN(n11981) );
  NAND2_X1 U14888 ( .A1(n15796), .A2(n11981), .ZN(n16432) );
  INV_X1 U14889 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16441) );
  NOR2_X1 U14890 ( .A1(n16432), .A2(n16441), .ZN(n15767) );
  AND2_X1 U14891 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15769) );
  INV_X1 U14892 ( .A(n15769), .ZN(n15746) );
  AND2_X1 U14893 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15721) );
  INV_X1 U14894 ( .A(n15721), .ZN(n12390) );
  INV_X1 U14895 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11982) );
  INV_X1 U14896 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15538) );
  NAND2_X1 U14897 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12380) );
  AND2_X2 U14898 ( .A1(n12372), .A2(n13320), .ZN(n16460) );
  NAND2_X1 U14899 ( .A1(n11984), .A2(n11983), .ZN(n11989) );
  INV_X1 U14900 ( .A(n11985), .ZN(n11987) );
  OR2_X1 U14901 ( .A1(n11987), .A2(n11986), .ZN(n11988) );
  NAND2_X1 U14902 ( .A1(n11989), .A2(n11988), .ZN(n13521) );
  INV_X1 U14903 ( .A(n13521), .ZN(n11995) );
  INV_X1 U14904 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11992) );
  NAND2_X1 U14905 ( .A1(n12012), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11991) );
  NAND2_X1 U14906 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11990) );
  OAI211_X1 U14907 ( .C1(n15099), .C2(n11992), .A(n11991), .B(n11990), .ZN(
        n11993) );
  AOI21_X1 U14908 ( .B1(n11443), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n11993), .ZN(n13520) );
  NAND2_X1 U14909 ( .A1(n11995), .A2(n11994), .ZN(n13523) );
  INV_X1 U14910 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n11998) );
  NAND2_X1 U14911 ( .A1(n12012), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11997) );
  NAND2_X1 U14912 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11996) );
  OAI211_X1 U14913 ( .C1(n15099), .C2(n11998), .A(n11997), .B(n11996), .ZN(
        n11999) );
  AOI21_X1 U14914 ( .B1(n11443), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11999), .ZN(n13007) );
  AOI22_X1 U14915 ( .A1(n12076), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12001) );
  NAND2_X1 U14916 ( .A1(n12003), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12000) );
  OAI211_X1 U14917 ( .C1(n12002), .C2(n16471), .A(n12001), .B(n12000), .ZN(
        n13000) );
  NAND2_X1 U14918 ( .A1(n12999), .A2(n13000), .ZN(n12993) );
  INV_X1 U14919 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n12005) );
  AOI22_X1 U14920 ( .A1(n12076), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12004) );
  OAI21_X1 U14921 ( .B1(n15099), .B2(n12005), .A(n12004), .ZN(n12006) );
  AOI21_X1 U14922 ( .B1(n15101), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n12006), .ZN(n12995) );
  INV_X1 U14923 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n15340) );
  NAND2_X1 U14924 ( .A1(n15101), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12008) );
  AOI22_X1 U14925 ( .A1(n12076), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12007) );
  OAI211_X1 U14926 ( .C1(n15099), .C2(n15340), .A(n12008), .B(n12007), .ZN(
        n15330) );
  INV_X1 U14927 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U14928 ( .A1(n12076), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12009) );
  OAI21_X1 U14929 ( .B1(n15099), .B2(n12010), .A(n12009), .ZN(n12011) );
  AOI21_X1 U14930 ( .B1(n15101), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n12011), .ZN(n13028) );
  NAND2_X1 U14931 ( .A1(n15101), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12018) );
  INV_X1 U14932 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n12015) );
  NAND2_X1 U14933 ( .A1(n12012), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12014) );
  NAND2_X1 U14934 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12013) );
  OAI211_X1 U14935 ( .C1(n15099), .C2(n12015), .A(n12014), .B(n12013), .ZN(
        n12016) );
  INV_X1 U14936 ( .A(n12016), .ZN(n12017) );
  NAND2_X1 U14937 ( .A1(n12018), .A2(n12017), .ZN(n16377) );
  INV_X1 U14938 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n12021) );
  NAND2_X1 U14939 ( .A1(n15101), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12020) );
  AOI22_X1 U14940 ( .A1(n12076), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n12019) );
  OAI211_X1 U14941 ( .C1(n15099), .C2(n12021), .A(n12020), .B(n12019), .ZN(
        n13223) );
  INV_X1 U14942 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n12024) );
  NAND2_X1 U14943 ( .A1(n15101), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12023) );
  AOI22_X1 U14944 ( .A1(n12076), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n12022) );
  OAI211_X1 U14945 ( .C1(n15099), .C2(n12024), .A(n12023), .B(n12022), .ZN(
        n15864) );
  INV_X1 U14946 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n15847) );
  NAND2_X1 U14947 ( .A1(n12076), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12026) );
  NAND2_X1 U14948 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12025) );
  OAI211_X1 U14949 ( .C1(n15099), .C2(n15847), .A(n12026), .B(n12025), .ZN(
        n12027) );
  AOI21_X1 U14950 ( .B1(n15101), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n12027), .ZN(n13376) );
  NAND2_X1 U14951 ( .A1(n15101), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12033) );
  INV_X1 U14952 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n12030) );
  NAND2_X1 U14953 ( .A1(n12076), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12029) );
  NAND2_X1 U14954 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12028) );
  OAI211_X1 U14955 ( .C1(n15099), .C2(n12030), .A(n12029), .B(n12028), .ZN(
        n12031) );
  INV_X1 U14956 ( .A(n12031), .ZN(n12032) );
  NAND2_X1 U14957 ( .A1(n12033), .A2(n12032), .ZN(n15827) );
  INV_X1 U14958 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n15617) );
  NAND2_X1 U14959 ( .A1(n12076), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12035) );
  NAND2_X1 U14960 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12034) );
  OAI211_X1 U14961 ( .C1(n15099), .C2(n15617), .A(n12035), .B(n12034), .ZN(
        n12036) );
  AOI21_X1 U14962 ( .B1(n15101), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n12036), .ZN(n13623) );
  INV_X1 U14963 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19856) );
  NAND2_X1 U14964 ( .A1(n12076), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12038) );
  NAND2_X1 U14965 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12037) );
  OAI211_X1 U14966 ( .C1(n15099), .C2(n19856), .A(n12038), .B(n12037), .ZN(
        n12039) );
  AOI21_X1 U14967 ( .B1(n15101), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n12039), .ZN(n15304) );
  INV_X1 U14968 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19858) );
  NAND2_X1 U14969 ( .A1(n15101), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12041) );
  AOI22_X1 U14970 ( .A1(n12076), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n12040) );
  OAI211_X1 U14971 ( .C1(n15099), .C2(n19858), .A(n12041), .B(n12040), .ZN(
        n13727) );
  INV_X1 U14972 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15287) );
  NAND2_X1 U14973 ( .A1(n12076), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12043) );
  NAND2_X1 U14974 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12042) );
  OAI211_X1 U14975 ( .C1(n15099), .C2(n15287), .A(n12043), .B(n12042), .ZN(
        n12044) );
  AOI21_X1 U14976 ( .B1(n15101), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n12044), .ZN(n15289) );
  INV_X1 U14977 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n12047) );
  NAND2_X1 U14978 ( .A1(n12076), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12046) );
  NAND2_X1 U14979 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12045) );
  OAI211_X1 U14980 ( .C1(n15099), .C2(n12047), .A(n12046), .B(n12045), .ZN(
        n12048) );
  AOI21_X1 U14981 ( .B1(n15101), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n12048), .ZN(n15430) );
  INV_X1 U14982 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n18980) );
  NAND2_X1 U14983 ( .A1(n15101), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12051) );
  AOI22_X1 U14984 ( .A1(n12076), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n12050) );
  OAI211_X1 U14985 ( .C1(n15099), .C2(n18980), .A(n12051), .B(n12050), .ZN(
        n15762) );
  INV_X1 U14986 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20953) );
  NAND2_X1 U14987 ( .A1(n15101), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12053) );
  AOI22_X1 U14988 ( .A1(n12076), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n12052) );
  OAI211_X1 U14989 ( .C1(n15099), .C2(n20953), .A(n12053), .B(n12052), .ZN(
        n15270) );
  INV_X1 U14990 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n12056) );
  NAND2_X1 U14991 ( .A1(n12076), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12055) );
  NAND2_X1 U14992 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12054) );
  OAI211_X1 U14993 ( .C1(n15099), .C2(n12056), .A(n12055), .B(n12054), .ZN(
        n12057) );
  AOI21_X1 U14994 ( .B1(n15101), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n12057), .ZN(n15256) );
  INV_X1 U14995 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n12060) );
  NAND2_X1 U14996 ( .A1(n12076), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12059) );
  NAND2_X1 U14997 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12058) );
  OAI211_X1 U14998 ( .C1(n15099), .C2(n12060), .A(n12059), .B(n12058), .ZN(
        n12061) );
  AOI21_X1 U14999 ( .B1(n15101), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n12061), .ZN(n15237) );
  INV_X1 U15000 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n12064) );
  NAND2_X1 U15001 ( .A1(n12076), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12063) );
  NAND2_X1 U15002 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12062) );
  OAI211_X1 U15003 ( .C1(n15099), .C2(n12064), .A(n12063), .B(n12062), .ZN(
        n12065) );
  AOI21_X1 U15004 ( .B1(n15101), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n12065), .ZN(n15226) );
  INV_X1 U15005 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19867) );
  NAND2_X1 U15006 ( .A1(n11443), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12067) );
  AOI22_X1 U15007 ( .A1(n12076), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n12066) );
  OAI211_X1 U15008 ( .C1(n15099), .C2(n19867), .A(n12067), .B(n12066), .ZN(
        n15206) );
  NAND2_X1 U15009 ( .A1(n15228), .A2(n15206), .ZN(n15208) );
  INV_X1 U15010 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19869) );
  NAND2_X1 U15011 ( .A1(n12076), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12069) );
  NAND2_X1 U15012 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12068) );
  OAI211_X1 U15013 ( .C1(n15099), .C2(n19869), .A(n12069), .B(n12068), .ZN(
        n12070) );
  AOI21_X1 U15014 ( .B1(n15101), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12070), .ZN(n15192) );
  INV_X1 U15015 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19871) );
  NAND2_X1 U15016 ( .A1(n12076), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12072) );
  NAND2_X1 U15017 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12071) );
  OAI211_X1 U15018 ( .C1(n15099), .C2(n19871), .A(n12072), .B(n12071), .ZN(
        n12073) );
  AOI21_X1 U15019 ( .B1(n15101), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n12073), .ZN(n15170) );
  INV_X1 U15020 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n12332) );
  NAND2_X1 U15021 ( .A1(n11443), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12075) );
  AOI22_X1 U15022 ( .A1(n12076), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12074) );
  OAI211_X1 U15023 ( .C1(n15099), .C2(n12332), .A(n12075), .B(n12074), .ZN(
        n15158) );
  INV_X1 U15024 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19873) );
  NAND2_X1 U15025 ( .A1(n11443), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12078) );
  AOI22_X1 U15026 ( .A1(n12076), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12077) );
  OAI211_X1 U15027 ( .C1(n15099), .C2(n19873), .A(n12078), .B(n12077), .ZN(
        n15388) );
  INV_X1 U15028 ( .A(n15390), .ZN(n12084) );
  INV_X1 U15029 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n12346) );
  NAND2_X1 U15030 ( .A1(n12076), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12080) );
  NAND2_X1 U15031 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12079) );
  OAI211_X1 U15032 ( .C1(n15099), .C2(n12346), .A(n12080), .B(n12079), .ZN(
        n12081) );
  AOI21_X1 U15033 ( .B1(n15101), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12081), .ZN(n12082) );
  INV_X1 U15034 ( .A(n12082), .ZN(n12083) );
  NAND2_X1 U15035 ( .A1(n15928), .A2(n14263), .ZN(n12085) );
  NAND2_X1 U15036 ( .A1(n12085), .A2(n11416), .ZN(n12086) );
  NAND2_X1 U15037 ( .A1(n12372), .A2(n12086), .ZN(n16466) );
  NOR2_X1 U15038 ( .A1(n12957), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12087) );
  INV_X1 U15039 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n12094) );
  NAND2_X1 U15040 ( .A1(n9719), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12093) );
  NOR2_X1 U15041 ( .A1(n12089), .A2(n19325), .ZN(n12090) );
  MUX2_X1 U15042 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n12090), .S(
        n14263), .Z(n12091) );
  NAND2_X1 U15043 ( .A1(n12091), .A2(n19757), .ZN(n12092) );
  OAI211_X1 U15044 ( .C1(n12338), .C2(n12094), .A(n12093), .B(n12092), .ZN(
        n13693) );
  INV_X1 U15045 ( .A(n12880), .ZN(n12097) );
  NOR2_X1 U15046 ( .A1(n19944), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12095) );
  INV_X1 U15047 ( .A(n12304), .ZN(n12096) );
  NAND2_X1 U15048 ( .A1(n12097), .A2(n12096), .ZN(n12102) );
  AND2_X2 U15049 ( .A1(n19944), .A2(n19757), .ZN(n12142) );
  NAND2_X1 U15050 ( .A1(n12098), .A2(n12142), .ZN(n12115) );
  OAI22_X1 U15051 ( .A1(n12957), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n19931), 
        .B2(n19757), .ZN(n12099) );
  INV_X1 U15052 ( .A(n12099), .ZN(n12100) );
  AND2_X1 U15053 ( .A1(n12115), .A2(n12100), .ZN(n12101) );
  NAND2_X1 U15054 ( .A1(n12107), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12106) );
  INV_X1 U15055 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12966) );
  NAND2_X1 U15056 ( .A1(n19944), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12103) );
  OAI211_X1 U15057 ( .C1(n12957), .C2(n12966), .A(n19757), .B(n12103), .ZN(
        n12104) );
  INV_X1 U15058 ( .A(n12104), .ZN(n12105) );
  NAND2_X1 U15059 ( .A1(n12106), .A2(n12105), .ZN(n12961) );
  INV_X1 U15060 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19839) );
  NAND2_X1 U15061 ( .A1(n12107), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U15062 ( .A1(n12087), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12142), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12108) );
  NAND2_X1 U15063 ( .A1(n12109), .A2(n12108), .ZN(n12114) );
  AND2_X1 U15064 ( .A1(n12957), .A2(n19757), .ZN(n12110) );
  AOI22_X1 U15065 ( .A1(n11386), .A2(n12110), .B1(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12111) );
  OAI21_X1 U15066 ( .B1(n12112), .B2(n12304), .A(n12111), .ZN(n13031) );
  NAND2_X1 U15067 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12116) );
  OAI211_X1 U15068 ( .C1(n12304), .C2(n12117), .A(n12116), .B(n12115), .ZN(
        n12120) );
  NAND2_X1 U15069 ( .A1(n9719), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12119) );
  INV_X2 U15070 ( .A(n12338), .ZN(n12312) );
  AOI22_X1 U15071 ( .A1(n12312), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12142), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12118) );
  NAND2_X1 U15072 ( .A1(n12119), .A2(n12118), .ZN(n12890) );
  NOR2_X1 U15073 ( .A1(n12891), .A2(n12890), .ZN(n12892) );
  NOR2_X1 U15074 ( .A1(n12121), .A2(n12120), .ZN(n12122) );
  AOI22_X1 U15075 ( .A1(n12142), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12124) );
  NAND2_X1 U15076 ( .A1(n12312), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12123) );
  OAI211_X1 U15077 ( .C1(n12304), .C2(n12125), .A(n12124), .B(n12123), .ZN(
        n12126) );
  INV_X1 U15078 ( .A(n12126), .ZN(n12128) );
  NAND2_X1 U15079 ( .A1(n9719), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12127) );
  NAND2_X1 U15080 ( .A1(n12128), .A2(n12127), .ZN(n13359) );
  NAND2_X1 U15081 ( .A1(n13358), .A2(n13359), .ZN(n13527) );
  NAND2_X1 U15082 ( .A1(n12142), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12130) );
  NAND2_X1 U15083 ( .A1(n12312), .A2(P2_EAX_REG_4__SCAN_IN), .ZN(n12129) );
  OAI211_X1 U15084 ( .C1(n12304), .C2(n12131), .A(n12130), .B(n12129), .ZN(
        n12132) );
  INV_X1 U15085 ( .A(n12132), .ZN(n12134) );
  NAND2_X1 U15086 ( .A1(n9719), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12133) );
  NOR2_X1 U15087 ( .A1(n12304), .A2(n12135), .ZN(n12136) );
  AOI21_X1 U15088 ( .B1(n13693), .B2(n13694), .A(n12136), .ZN(n13775) );
  NAND2_X1 U15089 ( .A1(n9719), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U15090 ( .A1(n12312), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12142), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12137) );
  NAND2_X1 U15091 ( .A1(n12138), .A2(n12137), .ZN(n13774) );
  INV_X1 U15092 ( .A(n13774), .ZN(n12141) );
  OR2_X1 U15093 ( .A1(n12304), .A2(n12139), .ZN(n12140) );
  NAND2_X1 U15094 ( .A1(n9719), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n12144) );
  AOI22_X1 U15095 ( .A1(n12312), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n12142), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12143) );
  NAND2_X1 U15096 ( .A1(n12144), .A2(n12143), .ZN(n16477) );
  AOI22_X1 U15097 ( .A1(n14162), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12262), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15098 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11523), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12147) );
  AOI22_X1 U15099 ( .A1(n11528), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12146) );
  NAND2_X1 U15100 ( .A1(n9741), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12145) );
  NAND4_X1 U15101 ( .A1(n12148), .A2(n12147), .A3(n12146), .A4(n12145), .ZN(
        n12158) );
  AOI22_X1 U15102 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11588), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12156) );
  INV_X1 U15103 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12151) );
  NAND2_X1 U15104 ( .A1(n11513), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12150) );
  NAND2_X1 U15105 ( .A1(n11537), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12149) );
  OAI211_X1 U15106 ( .C1(n14153), .C2(n12151), .A(n12150), .B(n12149), .ZN(
        n12152) );
  INV_X1 U15107 ( .A(n12152), .ZN(n12155) );
  AOI22_X1 U15108 ( .A1(n14161), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14155), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U15109 ( .A1(n11571), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12153) );
  NAND4_X1 U15110 ( .A1(n12156), .A2(n12155), .A3(n12154), .A4(n12153), .ZN(
        n12157) );
  INV_X1 U15111 ( .A(n13023), .ZN(n19158) );
  NAND2_X1 U15112 ( .A1(n12312), .A2(P2_EAX_REG_8__SCAN_IN), .ZN(n12160) );
  NAND2_X1 U15113 ( .A1(n12142), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12159) );
  OAI211_X1 U15114 ( .C1(n12304), .C2(n19158), .A(n12160), .B(n12159), .ZN(
        n12161) );
  INV_X1 U15115 ( .A(n12161), .ZN(n12163) );
  NAND2_X1 U15116 ( .A1(n9719), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U15117 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11528), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12167) );
  NAND2_X1 U15118 ( .A1(n9741), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12166) );
  NAND2_X1 U15119 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12165) );
  NAND2_X1 U15120 ( .A1(n11523), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12164) );
  NAND4_X1 U15121 ( .A1(n12167), .A2(n12166), .A3(n12165), .A4(n12164), .ZN(
        n12171) );
  INV_X1 U15122 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12168) );
  OAI22_X1 U15123 ( .A1(n14096), .A2(n12169), .B1(n14095), .B2(n12168), .ZN(
        n12170) );
  NOR2_X1 U15124 ( .A1(n12171), .A2(n12170), .ZN(n12179) );
  OAI22_X1 U15125 ( .A1(n14181), .A2(n14101), .B1(n14099), .B2(n12828), .ZN(
        n12175) );
  NAND2_X1 U15126 ( .A1(n11513), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12173) );
  NAND2_X1 U15127 ( .A1(n11537), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12172) );
  OAI211_X1 U15128 ( .C1(n14153), .C2(n14174), .A(n12173), .B(n12172), .ZN(
        n12174) );
  NOR2_X1 U15129 ( .A1(n12175), .A2(n12174), .ZN(n12178) );
  AOI22_X1 U15130 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11588), .B1(
        n11575), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12177) );
  AOI22_X1 U15131 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11571), .B1(
        n12262), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12176) );
  NAND4_X1 U15132 ( .A1(n12179), .A2(n12178), .A3(n12177), .A4(n12176), .ZN(
        n13026) );
  INV_X1 U15133 ( .A(n13026), .ZN(n13025) );
  NAND2_X1 U15134 ( .A1(n9719), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15135 ( .A1(n12312), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12142), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12180) );
  OAI211_X1 U15136 ( .C1(n13025), .C2(n12304), .A(n12181), .B(n12180), .ZN(
        n15901) );
  AOI22_X1 U15137 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n14162), .B1(
        n12262), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12185) );
  AOI22_X1 U15138 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11523), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U15139 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n11537), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12183) );
  NAND2_X1 U15140 ( .A1(n9741), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12182) );
  NAND4_X1 U15141 ( .A1(n12185), .A2(n12184), .A3(n12183), .A4(n12182), .ZN(
        n12195) );
  AOI22_X1 U15142 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n11575), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12193) );
  INV_X1 U15143 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12188) );
  INV_X1 U15144 ( .A(n14163), .ZN(n12217) );
  INV_X1 U15145 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13985) );
  OR2_X1 U15146 ( .A1(n12217), .A2(n13985), .ZN(n12187) );
  NAND2_X1 U15147 ( .A1(n11513), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12186) );
  OAI211_X1 U15148 ( .C1(n14153), .C2(n12188), .A(n12187), .B(n12186), .ZN(
        n12189) );
  INV_X1 U15149 ( .A(n12189), .ZN(n12192) );
  AOI22_X1 U15150 ( .A1(n11588), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n14155), .ZN(n12191) );
  AOI22_X1 U15151 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n14161), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12190) );
  NAND4_X1 U15152 ( .A1(n12193), .A2(n12192), .A3(n12191), .A4(n12190), .ZN(
        n12194) );
  INV_X1 U15153 ( .A(n19150), .ZN(n13221) );
  AOI22_X1 U15154 ( .A1(n12312), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12142), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12196) );
  OAI21_X1 U15155 ( .B1(n13221), .B2(n12304), .A(n12196), .ZN(n12197) );
  AOI21_X1 U15156 ( .B1(n9719), .B2(P2_REIP_REG_10__SCAN_IN), .A(n12197), .ZN(
        n16453) );
  NOR2_X2 U15157 ( .A1(n15902), .A2(n16453), .ZN(n15317) );
  AOI22_X1 U15158 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n11528), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12201) );
  NAND2_X1 U15159 ( .A1(n13998), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12200) );
  NAND2_X1 U15160 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12199) );
  NAND2_X1 U15161 ( .A1(n11523), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12198) );
  NAND4_X1 U15162 ( .A1(n12201), .A2(n12200), .A3(n12199), .A4(n12198), .ZN(
        n12205) );
  OAI22_X1 U15163 ( .A1(n14096), .A2(n12203), .B1(n14095), .B2(n12202), .ZN(
        n12204) );
  NOR2_X1 U15164 ( .A1(n12205), .A2(n12204), .ZN(n12214) );
  OAI22_X1 U15165 ( .A1(n14227), .A2(n14101), .B1(n14099), .B2(n12206), .ZN(
        n12210) );
  NAND2_X1 U15166 ( .A1(n11513), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n12208) );
  NAND2_X1 U15167 ( .A1(n11537), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12207) );
  OAI211_X1 U15168 ( .C1(n14153), .C2(n14220), .A(n12208), .B(n12207), .ZN(
        n12209) );
  NOR2_X1 U15169 ( .A1(n12210), .A2(n12209), .ZN(n12213) );
  AOI22_X1 U15170 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11588), .B1(
        n11575), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15171 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n11571), .B1(
        n12262), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12211) );
  NAND4_X1 U15172 ( .A1(n12214), .A2(n12213), .A3(n12212), .A4(n12211), .ZN(
        n13218) );
  INV_X1 U15173 ( .A(n13218), .ZN(n13220) );
  NAND2_X1 U15174 ( .A1(n9719), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15175 ( .A1(n12312), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12142), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12215) );
  OAI211_X1 U15176 ( .C1(n13220), .C2(n12304), .A(n12216), .B(n12215), .ZN(
        n15318) );
  NAND2_X1 U15177 ( .A1(n15317), .A2(n15318), .ZN(n15319) );
  AOI22_X1 U15178 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11588), .B1(
        n11575), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12225) );
  INV_X1 U15179 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14077) );
  OR2_X1 U15180 ( .A1(n12217), .A2(n14077), .ZN(n12219) );
  NAND2_X1 U15181 ( .A1(n11513), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12218) );
  OAI211_X1 U15182 ( .C1(n14099), .C2(n12220), .A(n12219), .B(n12218), .ZN(
        n12221) );
  INV_X1 U15183 ( .A(n12221), .ZN(n12224) );
  AOI22_X1 U15184 ( .A1(n11571), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n12292), .ZN(n12223) );
  AOI22_X1 U15185 ( .A1(n14162), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12222) );
  NAND4_X1 U15186 ( .A1(n12225), .A2(n12224), .A3(n12223), .A4(n12222), .ZN(
        n12231) );
  AOI22_X1 U15187 ( .A1(n12262), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14161), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12229) );
  AOI22_X1 U15188 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11529), .B1(
        n11523), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15189 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11537), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12227) );
  NAND2_X1 U15190 ( .A1(n13998), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12226) );
  NAND4_X1 U15191 ( .A1(n12229), .A2(n12228), .A3(n12227), .A4(n12226), .ZN(
        n12230) );
  NAND2_X1 U15192 ( .A1(n12312), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n12233) );
  NAND2_X1 U15193 ( .A1(n12142), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12232) );
  OAI211_X1 U15194 ( .C1(n12304), .C2(n9816), .A(n12233), .B(n12232), .ZN(
        n12234) );
  INV_X1 U15195 ( .A(n12234), .ZN(n12236) );
  NAND2_X1 U15196 ( .A1(n9719), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12235) );
  NOR2_X2 U15197 ( .A1(n15319), .A2(n15868), .ZN(n15850) );
  AOI22_X1 U15198 ( .A1(n11528), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12240) );
  NAND2_X1 U15199 ( .A1(n9741), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12239) );
  NAND2_X1 U15200 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12238) );
  NAND2_X1 U15201 ( .A1(n11523), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12237) );
  NAND4_X1 U15202 ( .A1(n12240), .A2(n12239), .A3(n12238), .A4(n12237), .ZN(
        n12244) );
  OAI22_X1 U15203 ( .A1(n14096), .A2(n12242), .B1(n14095), .B2(n12241), .ZN(
        n12243) );
  NOR2_X1 U15204 ( .A1(n12244), .A2(n12243), .ZN(n12255) );
  NAND2_X1 U15205 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12248) );
  NAND2_X1 U15206 ( .A1(n11588), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12247) );
  NAND2_X1 U15207 ( .A1(n12262), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12246) );
  NAND2_X1 U15208 ( .A1(n11571), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12245) );
  AND4_X1 U15209 ( .A1(n12248), .A2(n12247), .A3(n12246), .A4(n12245), .ZN(
        n12254) );
  OAI22_X1 U15210 ( .A1(n14101), .A2(n14274), .B1(n14099), .B2(n13002), .ZN(
        n12252) );
  NAND2_X1 U15211 ( .A1(n11513), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n12250) );
  NAND2_X1 U15212 ( .A1(n11537), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12249) );
  OAI211_X1 U15213 ( .C1(n14153), .C2(n14267), .A(n12250), .B(n12249), .ZN(
        n12251) );
  NOR2_X1 U15214 ( .A1(n12252), .A2(n12251), .ZN(n12253) );
  NAND2_X1 U15215 ( .A1(n9719), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12257) );
  AOI22_X1 U15216 ( .A1(n12312), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12142), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12256) );
  OAI211_X1 U15217 ( .C1(n13372), .C2(n12304), .A(n12257), .B(n12256), .ZN(
        n15851) );
  NAND2_X1 U15218 ( .A1(n15850), .A2(n15851), .ZN(n15824) );
  INV_X1 U15219 ( .A(n15824), .ZN(n12284) );
  AOI22_X1 U15220 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11537), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12261) );
  NAND2_X1 U15221 ( .A1(n13998), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12260) );
  NAND2_X1 U15222 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12259) );
  NAND2_X1 U15223 ( .A1(n11523), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12258) );
  NAND4_X1 U15224 ( .A1(n12261), .A2(n12260), .A3(n12259), .A4(n12258), .ZN(
        n12266) );
  INV_X1 U15225 ( .A(n12262), .ZN(n12264) );
  OAI22_X1 U15226 ( .A1(n14295), .A2(n12264), .B1(n14096), .B2(n12263), .ZN(
        n12265) );
  NOR2_X1 U15227 ( .A1(n12266), .A2(n12265), .ZN(n12278) );
  NAND2_X1 U15228 ( .A1(n11588), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12270) );
  NAND2_X1 U15229 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12269) );
  NAND2_X1 U15230 ( .A1(n11571), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12268) );
  NAND2_X1 U15231 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12267) );
  NAND4_X1 U15232 ( .A1(n12270), .A2(n12269), .A3(n12268), .A4(n12267), .ZN(
        n12276) );
  AOI22_X1 U15233 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11513), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12274) );
  NAND2_X1 U15234 ( .A1(n12292), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12273) );
  NAND2_X1 U15235 ( .A1(n14161), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12272) );
  NAND2_X1 U15236 ( .A1(n14155), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12271) );
  NAND4_X1 U15237 ( .A1(n12274), .A2(n12273), .A3(n12272), .A4(n12271), .ZN(
        n12275) );
  NOR2_X1 U15238 ( .A1(n12276), .A2(n12275), .ZN(n12277) );
  NAND2_X1 U15239 ( .A1(n12312), .A2(P2_EAX_REG_14__SCAN_IN), .ZN(n12280) );
  NAND2_X1 U15240 ( .A1(n12142), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12279) );
  OAI211_X1 U15241 ( .C1(n12304), .C2(n19143), .A(n12280), .B(n12279), .ZN(
        n12281) );
  INV_X1 U15242 ( .A(n12281), .ZN(n12283) );
  NAND2_X1 U15243 ( .A1(n9719), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12282) );
  NAND2_X1 U15244 ( .A1(n12283), .A2(n12282), .ZN(n15823) );
  AOI22_X1 U15245 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11528), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12288) );
  NAND2_X1 U15246 ( .A1(n13998), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12287) );
  NAND2_X1 U15247 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12286) );
  NAND2_X1 U15248 ( .A1(n11523), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12285) );
  NAND4_X1 U15249 ( .A1(n12288), .A2(n12287), .A3(n12286), .A4(n12285), .ZN(
        n12291) );
  INV_X1 U15250 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n19564) );
  INV_X1 U15251 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12289) );
  OAI22_X1 U15252 ( .A1(n14096), .A2(n19564), .B1(n14095), .B2(n12289), .ZN(
        n12290) );
  NOR2_X1 U15253 ( .A1(n12291), .A2(n12290), .ZN(n12300) );
  AOI22_X1 U15254 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n11537), .B1(
        n11513), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12296) );
  NAND2_X1 U15255 ( .A1(n12292), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12295) );
  NAND2_X1 U15256 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12294) );
  NAND2_X1 U15257 ( .A1(n14155), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12293) );
  AND4_X1 U15258 ( .A1(n12296), .A2(n12295), .A3(n12294), .A4(n12293), .ZN(
        n12299) );
  AOI22_X1 U15259 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11588), .B1(
        n11575), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15260 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n12262), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12297) );
  NAND4_X1 U15261 ( .A1(n12300), .A2(n12299), .A3(n12298), .A4(n12297), .ZN(
        n13622) );
  INV_X1 U15262 ( .A(n13622), .ZN(n12303) );
  NAND2_X1 U15263 ( .A1(n12312), .A2(P2_EAX_REG_15__SCAN_IN), .ZN(n12302) );
  NAND2_X1 U15264 ( .A1(n12142), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12301) );
  OAI211_X1 U15265 ( .C1(n12304), .C2(n12303), .A(n12302), .B(n12301), .ZN(
        n12305) );
  INV_X1 U15266 ( .A(n12305), .ZN(n12307) );
  NAND2_X1 U15267 ( .A1(n9719), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12306) );
  NAND2_X1 U15268 ( .A1(n9719), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U15269 ( .A1(n12312), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12142), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12308) );
  NAND2_X1 U15270 ( .A1(n9719), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U15271 ( .A1(n12312), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12142), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12310) );
  NAND2_X1 U15272 ( .A1(n12311), .A2(n12310), .ZN(n13959) );
  NAND2_X1 U15273 ( .A1(n9719), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12314) );
  AOI22_X1 U15274 ( .A1(n12312), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12142), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12313) );
  AND2_X1 U15275 ( .A1(n12314), .A2(n12313), .ZN(n15283) );
  NAND2_X1 U15276 ( .A1(n9719), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12316) );
  AOI22_X1 U15277 ( .A1(n12312), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12142), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12315) );
  NAND2_X1 U15278 ( .A1(n12316), .A2(n12315), .ZN(n14020) );
  NAND2_X1 U15279 ( .A1(n14019), .A2(n14020), .ZN(n14021) );
  NAND2_X1 U15280 ( .A1(n9719), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12318) );
  AOI22_X1 U15281 ( .A1(n12312), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12142), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12317) );
  AND2_X1 U15282 ( .A1(n12318), .A2(n12317), .ZN(n15766) );
  NOR2_X2 U15283 ( .A1(n14021), .A2(n15766), .ZN(n15765) );
  NAND2_X1 U15284 ( .A1(n9719), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12320) );
  AOI22_X1 U15285 ( .A1(n12312), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12142), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12319) );
  NAND2_X1 U15286 ( .A1(n12320), .A2(n12319), .ZN(n15272) );
  NAND2_X1 U15287 ( .A1(n9719), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12322) );
  AOI22_X1 U15288 ( .A1(n12312), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12142), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12321) );
  NAND2_X1 U15289 ( .A1(n12322), .A2(n12321), .ZN(n15260) );
  INV_X1 U15290 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n12839) );
  INV_X1 U15291 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15722) );
  INV_X1 U15292 ( .A(n12142), .ZN(n12336) );
  OAI22_X1 U15293 ( .A1(n12338), .A2(n12839), .B1(n15722), .B2(n12336), .ZN(
        n12323) );
  AOI21_X1 U15294 ( .B1(n9719), .B2(P2_REIP_REG_23__SCAN_IN), .A(n12323), .ZN(
        n15241) );
  NAND2_X1 U15295 ( .A1(n9719), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12325) );
  AOI22_X1 U15296 ( .A1(n12312), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12142), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12324) );
  AND2_X1 U15297 ( .A1(n12325), .A2(n12324), .ZN(n15229) );
  OR2_X1 U15298 ( .A1(n12333), .A2(n19867), .ZN(n12327) );
  AOI22_X1 U15299 ( .A1(n12312), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12142), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12326) );
  NAND2_X1 U15300 ( .A1(n12327), .A2(n12326), .ZN(n15209) );
  OR2_X1 U15301 ( .A1(n12333), .A2(n19869), .ZN(n12329) );
  AOI22_X1 U15302 ( .A1(n12312), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12142), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12328) );
  NAND2_X1 U15303 ( .A1(n12329), .A2(n12328), .ZN(n15194) );
  INV_X1 U15304 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n12848) );
  INV_X1 U15305 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15669) );
  OAI22_X1 U15306 ( .A1(n12338), .A2(n12848), .B1(n15669), .B2(n12336), .ZN(
        n12330) );
  AOI21_X1 U15307 ( .B1(n9719), .B2(P2_REIP_REG_27__SCAN_IN), .A(n12330), .ZN(
        n15172) );
  AOI22_X1 U15308 ( .A1(n12312), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12142), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12331) );
  OAI21_X1 U15309 ( .B1(n12333), .B2(n12332), .A(n12331), .ZN(n15160) );
  INV_X1 U15310 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14348) );
  OAI22_X1 U15311 ( .A1(n12338), .A2(n14348), .B1(n15642), .B2(n12336), .ZN(
        n12334) );
  AOI21_X1 U15312 ( .B1(n9719), .B2(P2_REIP_REG_29__SCAN_IN), .A(n12334), .ZN(
        n14346) );
  INV_X1 U15313 ( .A(n14346), .ZN(n12335) );
  INV_X1 U15314 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12337) );
  OAI22_X1 U15315 ( .A1(n12338), .A2(n12337), .B1(n20856), .B2(n12336), .ZN(
        n12339) );
  AOI21_X1 U15316 ( .B1(n9719), .B2(P2_REIP_REG_30__SCAN_IN), .A(n12339), .ZN(
        n12340) );
  OR2_X2 U15317 ( .A1(n9775), .A2(n12340), .ZN(n15138) );
  NAND2_X1 U15318 ( .A1(n9775), .A2(n12340), .ZN(n12341) );
  INV_X1 U15319 ( .A(n14337), .ZN(n15148) );
  AND2_X1 U15320 ( .A1(n12342), .A2(n12343), .ZN(n13326) );
  INV_X1 U15321 ( .A(n13326), .ZN(n13268) );
  NAND2_X1 U15322 ( .A1(n12742), .A2(n11913), .ZN(n12947) );
  NAND2_X1 U15323 ( .A1(n12947), .A2(n19944), .ZN(n12344) );
  NAND2_X1 U15324 ( .A1(n13268), .A2(n12344), .ZN(n12345) );
  NOR2_X1 U15325 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15937) );
  INV_X1 U15326 ( .A(n15937), .ZN(n19889) );
  NOR2_X1 U15327 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19889), .ZN(n12743) );
  AND2_X2 U15328 ( .A1(n12743), .A2(n16510), .ZN(n19276) );
  NOR2_X1 U15329 ( .A1(n9725), .A2(n12346), .ZN(n15494) );
  INV_X1 U15330 ( .A(n12347), .ZN(n12366) );
  NAND2_X1 U15331 ( .A1(n12348), .A2(n19944), .ZN(n13297) );
  NAND2_X1 U15332 ( .A1(n13297), .A2(n12349), .ZN(n12351) );
  NAND2_X1 U15333 ( .A1(n12351), .A2(n12350), .ZN(n12364) );
  NOR2_X1 U15334 ( .A1(n12353), .A2(n12352), .ZN(n12354) );
  NAND2_X1 U15335 ( .A1(n12355), .A2(n12354), .ZN(n12952) );
  INV_X1 U15336 ( .A(n12357), .ZN(n12745) );
  OAI21_X1 U15337 ( .B1(n12365), .B2(n12358), .A(n12745), .ZN(n12362) );
  NAND2_X1 U15338 ( .A1(n12360), .A2(n12359), .ZN(n12361) );
  AND4_X1 U15339 ( .A1(n12952), .A2(n12356), .A3(n12362), .A4(n12361), .ZN(
        n12363) );
  NAND2_X1 U15340 ( .A1(n12364), .A2(n12363), .ZN(n12814) );
  AOI21_X1 U15341 ( .B1(n12366), .B2(n12365), .A(n12814), .ZN(n13264) );
  NAND2_X1 U15342 ( .A1(n13264), .A2(n12367), .ZN(n12368) );
  NAND2_X1 U15343 ( .A1(n12372), .A2(n12368), .ZN(n15798) );
  NOR2_X1 U15344 ( .A1(n15923), .A2(n15914), .ZN(n15918) );
  INV_X1 U15345 ( .A(n12372), .ZN(n12369) );
  NAND2_X1 U15346 ( .A1(n12369), .A2(n9725), .ZN(n16490) );
  OAI21_X1 U15347 ( .B1(n15798), .B2(n15918), .A(n16490), .ZN(n12896) );
  NOR2_X1 U15348 ( .A1(n15798), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12895) );
  NAND2_X1 U15349 ( .A1(n12372), .A2(n12951), .ZN(n15793) );
  NOR2_X1 U15350 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n15918), .ZN(
        n12383) );
  INV_X1 U15351 ( .A(n12383), .ZN(n12909) );
  NOR2_X1 U15352 ( .A1(n15793), .A2(n12909), .ZN(n12373) );
  AND4_X1 U15353 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13770) );
  AND3_X1 U15354 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n13770), .ZN(n12386) );
  NOR2_X1 U15355 ( .A1(n16491), .A2(n12386), .ZN(n12374) );
  NOR2_X1 U15356 ( .A1(n13361), .A2(n12374), .ZN(n15887) );
  NAND2_X1 U15357 ( .A1(n15887), .A2(n16491), .ZN(n15695) );
  NAND3_X1 U15358 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15767), .A3(
        n15769), .ZN(n12389) );
  INV_X1 U15359 ( .A(n12389), .ZN(n12375) );
  NAND2_X1 U15360 ( .A1(n15887), .A2(n12375), .ZN(n12376) );
  NAND2_X1 U15361 ( .A1(n15695), .A2(n12376), .ZN(n15734) );
  OAI21_X1 U15362 ( .B1(n16491), .B2(n15721), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12377) );
  INV_X1 U15363 ( .A(n12377), .ZN(n12378) );
  NAND2_X1 U15364 ( .A1(n15734), .A2(n12378), .ZN(n15709) );
  NAND2_X1 U15365 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12391) );
  OAI21_X1 U15366 ( .B1(n15709), .B2(n12391), .A(n15695), .ZN(n12379) );
  NAND2_X1 U15367 ( .A1(n12379), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15667) );
  OR2_X1 U15368 ( .A1(n15667), .A2(n12380), .ZN(n15631) );
  NAND3_X1 U15369 ( .A1(n15631), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15695), .ZN(n12381) );
  OAI211_X1 U15370 ( .C1(n15497), .C2(n16466), .A(n12382), .B(n12381), .ZN(
        n12393) );
  NOR2_X1 U15371 ( .A1(n15793), .A2(n12383), .ZN(n12385) );
  INV_X1 U15372 ( .A(n15798), .ZN(n12384) );
  OR2_X1 U15373 ( .A1(n12385), .A2(n12384), .ZN(n12388) );
  AOI21_X1 U15374 ( .B1(n15918), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n12385), .ZN(n13362) );
  INV_X1 U15375 ( .A(n13362), .ZN(n13524) );
  AND2_X1 U15376 ( .A1(n13524), .A2(n12386), .ZN(n12387) );
  NOR2_X1 U15377 ( .A1(n12390), .A2(n15736), .ZN(n15710) );
  NAND2_X1 U15378 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15710), .ZN(
        n15698) );
  NOR2_X1 U15379 ( .A1(n15698), .A2(n12391), .ZN(n15641) );
  NAND3_X1 U15380 ( .A1(n15641), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15644) );
  NOR3_X1 U15381 ( .A1(n15644), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15642), .ZN(n12392) );
  OAI21_X1 U15382 ( .B1(n15501), .B2(n16498), .A(n12396), .ZN(P2_U3016) );
  AOI22_X1 U15383 ( .A1(n17256), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12401) );
  AOI22_X1 U15384 ( .A1(n15950), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12400) );
  INV_X2 U15385 ( .A(n9769), .ZN(n15951) );
  AOI22_X1 U15386 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15951), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15387 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15952), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12398) );
  NAND4_X1 U15388 ( .A1(n12401), .A2(n12400), .A3(n12399), .A4(n12398), .ZN(
        n12413) );
  INV_X2 U15389 ( .A(n13871), .ZN(n17286) );
  INV_X2 U15390 ( .A(n14035), .ZN(n15949) );
  AOI22_X1 U15391 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15949), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12411) );
  AOI22_X1 U15392 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12410) );
  AOI22_X1 U15393 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12409) );
  INV_X2 U15394 ( .A(n17075), .ZN(n17300) );
  AOI22_X1 U15395 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12408) );
  NAND4_X1 U15396 ( .A1(n12411), .A2(n12410), .A3(n12409), .A4(n12408), .ZN(
        n12412) );
  AOI22_X1 U15397 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U15398 ( .A1(n17256), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12416) );
  AOI22_X1 U15399 ( .A1(n15950), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17220), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12415) );
  AOI22_X1 U15400 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15949), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12414) );
  NAND4_X1 U15401 ( .A1(n12417), .A2(n12416), .A3(n12415), .A4(n12414), .ZN(
        n12424) );
  AOI22_X1 U15402 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15951), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12422) );
  INV_X2 U15403 ( .A(n17006), .ZN(n17254) );
  AOI22_X1 U15404 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U15405 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9718), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12420) );
  AOI22_X1 U15406 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12419) );
  NAND4_X1 U15407 ( .A1(n12422), .A2(n12421), .A3(n12420), .A4(n12419), .ZN(
        n12423) );
  INV_X4 U15408 ( .A(n13859), .ZN(n17289) );
  AOI22_X1 U15409 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12428) );
  AOI22_X1 U15410 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12427) );
  AOI22_X1 U15411 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15951), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12426) );
  AOI22_X1 U15412 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15952), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12425) );
  NAND4_X1 U15413 ( .A1(n12428), .A2(n12427), .A3(n12426), .A4(n12425), .ZN(
        n12434) );
  AOI22_X1 U15414 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U15415 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12431) );
  AOI22_X1 U15416 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12430) );
  AOI22_X1 U15417 ( .A1(n15950), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15949), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12429) );
  NAND4_X1 U15418 ( .A1(n12432), .A2(n12431), .A3(n12430), .A4(n12429), .ZN(
        n12433) );
  AOI22_X1 U15419 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U15420 ( .A1(n17268), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15951), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U15421 ( .A1(n15950), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U15422 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12435) );
  AOI22_X1 U15423 ( .A1(n13891), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12442) );
  AOI22_X1 U15424 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12441) );
  AOI22_X1 U15425 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15949), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12443) );
  OAI21_X1 U15426 ( .B1(n17006), .B2(n17329), .A(n12443), .ZN(n12444) );
  INV_X1 U15427 ( .A(n12444), .ZN(n12445) );
  NAND3_X1 U15428 ( .A1(n10154), .A2(n10155), .A3(n12445), .ZN(n17479) );
  AOI22_X1 U15429 ( .A1(n12450), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17269), .ZN(n12448) );
  AOI22_X1 U15430 ( .A1(n12405), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15951), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12447) );
  AOI22_X1 U15431 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n15949), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n12556), .ZN(n12449) );
  NAND2_X1 U15432 ( .A1(n17479), .A2(n12477), .ZN(n12476) );
  NOR2_X1 U15433 ( .A1(n17472), .A2(n12476), .ZN(n12475) );
  AOI22_X1 U15434 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12460) );
  AOI22_X1 U15435 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12459) );
  INV_X1 U15436 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17320) );
  AOI22_X1 U15437 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15949), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12451) );
  OAI21_X1 U15438 ( .B1(n17006), .B2(n17320), .A(n12451), .ZN(n12457) );
  AOI22_X1 U15439 ( .A1(n15950), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U15440 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U15441 ( .A1(n17287), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U15442 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15952), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12452) );
  NAND4_X1 U15443 ( .A1(n12455), .A2(n12454), .A3(n12453), .A4(n12452), .ZN(
        n12456) );
  AOI211_X1 U15444 ( .C1(n17157), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n12457), .B(n12456), .ZN(n12458) );
  NAND3_X1 U15445 ( .A1(n12460), .A2(n12459), .A3(n12458), .ZN(n12652) );
  NAND2_X1 U15446 ( .A1(n12475), .A2(n12652), .ZN(n12474) );
  AOI22_X1 U15447 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12470) );
  AOI22_X1 U15448 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12469) );
  INV_X1 U15449 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17312) );
  AOI22_X1 U15450 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15949), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12461) );
  OAI21_X1 U15451 ( .B1(n17006), .B2(n17312), .A(n12461), .ZN(n12467) );
  AOI22_X1 U15452 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12465) );
  AOI22_X1 U15453 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U15454 ( .A1(n15950), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15951), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12463) );
  INV_X1 U15455 ( .A(n9771), .ZN(n17293) );
  AOI22_X1 U15456 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12462) );
  NAND4_X1 U15457 ( .A1(n12465), .A2(n12464), .A3(n12463), .A4(n12462), .ZN(
        n12466) );
  AOI211_X1 U15458 ( .C1(n17268), .C2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n12467), .B(n12466), .ZN(n12468) );
  NAND3_X1 U15459 ( .A1(n12470), .A2(n12469), .A3(n12468), .ZN(n12653) );
  INV_X1 U15460 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16066) );
  NAND2_X1 U15461 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16066), .ZN(
        n12471) );
  OAI21_X1 U15462 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n17868), .A(
        n12471), .ZN(n12523) );
  INV_X1 U15463 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18892) );
  NAND2_X1 U15464 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18892), .ZN(
        n12517) );
  INV_X1 U15465 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17988) );
  NAND2_X1 U15466 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15999) );
  INV_X1 U15467 ( .A(n15999), .ZN(n17974) );
  INV_X1 U15468 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18006) );
  NOR2_X1 U15469 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18101) );
  INV_X1 U15470 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12505) );
  INV_X1 U15471 ( .A(n12653), .ZN(n17461) );
  XNOR2_X1 U15472 ( .A(n17461), .B(n12472), .ZN(n12473) );
  NAND2_X1 U15473 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12473), .ZN(
        n12499) );
  INV_X1 U15474 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18201) );
  XNOR2_X1 U15475 ( .A(n18201), .B(n12473), .ZN(n17900) );
  XOR2_X1 U15476 ( .A(n17464), .B(n12474), .Z(n12495) );
  INV_X1 U15477 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18217) );
  INV_X1 U15478 ( .A(n12652), .ZN(n17468) );
  XNOR2_X1 U15479 ( .A(n17468), .B(n12475), .ZN(n12493) );
  XNOR2_X1 U15480 ( .A(n18217), .B(n12493), .ZN(n17921) );
  INV_X1 U15481 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18245) );
  XOR2_X1 U15482 ( .A(n17472), .B(n12476), .Z(n17937) );
  INV_X1 U15483 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18254) );
  OR2_X1 U15484 ( .A1(n18254), .A2(n12478), .ZN(n12491) );
  XNOR2_X1 U15485 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12478), .ZN(
        n17950) );
  NAND2_X1 U15486 ( .A1(n17491), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12490) );
  AOI22_X1 U15487 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U15488 ( .A1(n13891), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U15489 ( .A1(n15950), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12481) );
  AOI22_X1 U15490 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12480) );
  NAND4_X1 U15491 ( .A1(n12483), .A2(n12482), .A3(n12481), .A4(n12480), .ZN(
        n12489) );
  INV_X2 U15492 ( .A(n9769), .ZN(n17287) );
  AOI22_X1 U15493 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12487) );
  AOI22_X1 U15494 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12418), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12486) );
  AOI22_X1 U15495 ( .A1(n12405), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12485) );
  AOI22_X1 U15496 ( .A1(n15949), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12484) );
  NAND4_X1 U15497 ( .A1(n12487), .A2(n12486), .A3(n12485), .A4(n12484), .ZN(
        n12488) );
  INV_X1 U15498 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18911) );
  NOR2_X1 U15499 ( .A1(n17967), .A2(n18911), .ZN(n17966) );
  NAND2_X1 U15500 ( .A1(n17958), .A2(n17966), .ZN(n17957) );
  NAND2_X1 U15501 ( .A1(n12490), .A2(n17957), .ZN(n17949) );
  NAND2_X1 U15502 ( .A1(n17950), .A2(n17949), .ZN(n17948) );
  NAND2_X1 U15503 ( .A1(n12491), .A2(n17948), .ZN(n17938) );
  NAND2_X1 U15504 ( .A1(n17937), .A2(n17938), .ZN(n17936) );
  NOR2_X1 U15505 ( .A1(n17937), .A2(n17938), .ZN(n12492) );
  AOI21_X2 U15506 ( .B1(n18245), .B2(n17936), .A(n12492), .ZN(n17920) );
  NAND2_X1 U15507 ( .A1(n17921), .A2(n17920), .ZN(n17919) );
  NAND2_X1 U15508 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12493), .ZN(
        n12494) );
  NAND2_X1 U15509 ( .A1(n12495), .A2(n12497), .ZN(n12498) );
  NAND2_X1 U15510 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17913), .ZN(
        n17912) );
  AOI21_X1 U15511 ( .B1(n17458), .B2(n12500), .A(n17795), .ZN(n12502) );
  NAND2_X1 U15512 ( .A1(n12502), .A2(n12501), .ZN(n12503) );
  INV_X1 U15513 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18143) );
  INV_X1 U15514 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18117) );
  INV_X1 U15515 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17852) );
  NAND2_X1 U15516 ( .A1(n18176), .A2(n17852), .ZN(n17848) );
  INV_X1 U15517 ( .A(n17848), .ZN(n12504) );
  INV_X1 U15518 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18093) );
  NOR2_X1 U15519 ( .A1(n18176), .A2(n17852), .ZN(n18160) );
  NAND2_X1 U15520 ( .A1(n18160), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18144) );
  NOR2_X1 U15521 ( .A1(n18144), .A2(n18143), .ZN(n18100) );
  NAND3_X1 U15522 ( .A1(n18100), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18118) );
  INV_X1 U15523 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18103) );
  NOR2_X1 U15524 ( .A1(n18118), .A2(n18103), .ZN(n15997) );
  INV_X1 U15525 ( .A(n15997), .ZN(n18080) );
  NAND2_X2 U15526 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n12506), .ZN(
        n17833) );
  NOR2_X2 U15527 ( .A1(n18080), .A2(n17833), .ZN(n18036) );
  INV_X1 U15528 ( .A(n18036), .ZN(n17762) );
  INV_X1 U15529 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n20847) );
  NAND2_X1 U15530 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18071) );
  INV_X1 U15531 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17737) );
  INV_X1 U15532 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18031) );
  NOR2_X1 U15533 ( .A1(n17737), .A2(n18031), .ZN(n18033) );
  NAND3_X1 U15534 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n18033), .ZN(n16013) );
  NOR2_X1 U15535 ( .A1(n18071), .A2(n16013), .ZN(n16518) );
  NAND3_X1 U15536 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n16518), .ZN(n12680) );
  INV_X1 U15537 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17749) );
  NAND2_X1 U15538 ( .A1(n17749), .A2(n17868), .ZN(n17744) );
  NOR2_X1 U15539 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17744), .ZN(
        n12509) );
  NAND2_X1 U15540 ( .A1(n12509), .A2(n18031), .ZN(n17707) );
  NOR2_X1 U15541 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17707), .ZN(
        n17685) );
  INV_X1 U15542 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18012) );
  INV_X1 U15543 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n20842) );
  INV_X1 U15544 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18018) );
  INV_X1 U15545 ( .A(n17667), .ZN(n17652) );
  MUX2_X1 U15546 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17652), .S(
        n17868), .Z(n12512) );
  INV_X1 U15547 ( .A(n16013), .ZN(n16570) );
  OR2_X1 U15548 ( .A1(n18071), .A2(n17762), .ZN(n17706) );
  NAND2_X1 U15549 ( .A1(n12510), .A2(n17706), .ZN(n17746) );
  NAND2_X1 U15550 ( .A1(n16570), .A2(n17746), .ZN(n17686) );
  NAND3_X1 U15551 ( .A1(n17673), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n17667), .ZN(n12513) );
  INV_X1 U15552 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17995) );
  NAND2_X1 U15553 ( .A1(n17795), .A2(n12513), .ZN(n17651) );
  NAND2_X1 U15554 ( .A1(n17795), .A2(n17625), .ZN(n16565) );
  AND2_X2 U15555 ( .A1(n12514), .A2(n17988), .ZN(n17626) );
  INV_X1 U15556 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17613) );
  NAND2_X1 U15557 ( .A1(n17626), .A2(n17613), .ZN(n12515) );
  NOR2_X1 U15558 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17868), .ZN(
        n16560) );
  AOI22_X1 U15559 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17868), .B1(
        n12517), .B2(n12516), .ZN(n12522) );
  NOR2_X1 U15560 ( .A1(n17795), .A2(n12518), .ZN(n16061) );
  INV_X1 U15561 ( .A(n16060), .ZN(n12519) );
  OAI22_X1 U15562 ( .A1(n18892), .A2(n16061), .B1(n16066), .B2(n12519), .ZN(
        n12520) );
  NAND2_X1 U15563 ( .A1(n12523), .A2(n12520), .ZN(n12521) );
  OAI21_X1 U15564 ( .B1(n12523), .B2(n12522), .A(n12521), .ZN(n16555) );
  AOI22_X1 U15565 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18754), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18908), .ZN(n12640) );
  OAI21_X1 U15566 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18900), .A(
        n12525), .ZN(n12526) );
  OAI22_X1 U15567 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18762), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12526), .ZN(n12532) );
  NOR2_X1 U15568 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18762), .ZN(
        n12527) );
  NAND2_X1 U15569 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12526), .ZN(
        n12531) );
  AOI22_X1 U15570 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12532), .B1(
        n12527), .B2(n12531), .ZN(n12535) );
  AOI21_X1 U15571 ( .B1(n18914), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n12639), .ZN(n12643) );
  AND2_X1 U15572 ( .A1(n12640), .A2(n12643), .ZN(n12534) );
  OAI21_X1 U15573 ( .B1(n12530), .B2(n12529), .A(n12535), .ZN(n12528) );
  INV_X1 U15574 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18780) );
  OAI22_X1 U15575 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18780), .B1(
        n12533), .B2(n12532), .ZN(n12641) );
  AOI211_X1 U15576 ( .C1(n12535), .C2(n12534), .A(n12644), .B(n12641), .ZN(
        n18769) );
  AOI22_X1 U15577 ( .A1(n17287), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12539) );
  AOI22_X1 U15578 ( .A1(n17256), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12538) );
  AOI22_X1 U15579 ( .A1(n15949), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12537) );
  AOI22_X1 U15580 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15952), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12536) );
  NAND4_X1 U15581 ( .A1(n12539), .A2(n12538), .A3(n12537), .A4(n12536), .ZN(
        n12545) );
  AOI22_X1 U15582 ( .A1(n13891), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12543) );
  AOI22_X1 U15584 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17220), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12542) );
  AOI22_X1 U15585 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12541) );
  AOI22_X1 U15586 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12540) );
  NAND4_X1 U15587 ( .A1(n12543), .A2(n12542), .A3(n12541), .A4(n12540), .ZN(
        n12544) );
  AOI22_X1 U15588 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U15589 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12554) );
  AOI22_X1 U15590 ( .A1(n17256), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12546) );
  OAI21_X1 U15591 ( .B1(n14035), .B2(n21100), .A(n12546), .ZN(n12552) );
  AOI22_X1 U15592 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12550) );
  AOI22_X1 U15593 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12549) );
  AOI22_X1 U15594 ( .A1(n17287), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12548) );
  AOI22_X1 U15595 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15952), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12547) );
  NAND4_X1 U15596 ( .A1(n12550), .A2(n12549), .A3(n12548), .A4(n12547), .ZN(
        n12551) );
  NAND2_X1 U15597 ( .A1(n18305), .A2(n17494), .ZN(n12633) );
  NAND2_X1 U15598 ( .A1(n12633), .A2(n12627), .ZN(n18947) );
  AOI22_X1 U15599 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17291), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12560) );
  AOI22_X1 U15600 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12559) );
  AOI22_X1 U15601 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12558) );
  AOI22_X1 U15602 ( .A1(n13891), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15952), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12557) );
  NAND4_X1 U15603 ( .A1(n12560), .A2(n12559), .A3(n12558), .A4(n12557), .ZN(
        n12566) );
  AOI22_X1 U15604 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U15605 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12563) );
  AOI22_X1 U15606 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12562) );
  INV_X1 U15607 ( .A(n14035), .ZN(n12577) );
  AOI22_X1 U15608 ( .A1(n17256), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12561) );
  NAND4_X1 U15609 ( .A1(n12564), .A2(n12563), .A3(n12562), .A4(n12561), .ZN(
        n12565) );
  AOI22_X1 U15610 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12570) );
  AOI22_X1 U15611 ( .A1(n13891), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12569) );
  AOI22_X1 U15612 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12568) );
  AOI22_X1 U15613 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12567) );
  NAND4_X1 U15614 ( .A1(n12570), .A2(n12569), .A3(n12568), .A4(n12567), .ZN(
        n12576) );
  AOI22_X1 U15615 ( .A1(n17268), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12574) );
  AOI22_X1 U15616 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12573) );
  AOI22_X1 U15617 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17291), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12572) );
  AOI22_X1 U15618 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12571) );
  NAND4_X1 U15619 ( .A1(n12574), .A2(n12573), .A3(n12572), .A4(n12571), .ZN(
        n12575) );
  AOI22_X1 U15620 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12586) );
  AOI22_X1 U15621 ( .A1(n13891), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U15622 ( .A1(n17190), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12578) );
  OAI21_X1 U15623 ( .B1(n9772), .B2(n17329), .A(n12578), .ZN(n12584) );
  AOI22_X1 U15624 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(n9726), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12583) );
  AOI22_X1 U15625 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12579), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12582) );
  AOI22_X1 U15626 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12581) );
  AOI22_X1 U15627 ( .A1(n17287), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15952), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12580) );
  AOI22_X1 U15628 ( .A1(n17256), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12596) );
  AOI22_X1 U15629 ( .A1(n17292), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U15630 ( .A1(n17287), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12418), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12587) );
  OAI21_X1 U15631 ( .B1(n9772), .B2(n17320), .A(n12587), .ZN(n12593) );
  AOI22_X1 U15632 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U15633 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12590) );
  AOI22_X1 U15634 ( .A1(n13891), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15949), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U15635 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15952), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12588) );
  NAND4_X1 U15636 ( .A1(n12591), .A2(n12590), .A3(n12589), .A4(n12588), .ZN(
        n12592) );
  AOI211_X1 U15637 ( .C1(n17291), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n12593), .B(n12592), .ZN(n12594) );
  NAND3_X1 U15638 ( .A1(n12596), .A2(n12595), .A3(n12594), .ZN(n13822) );
  NOR3_X1 U15639 ( .A1(n17341), .A2(n13822), .A3(n12647), .ZN(n12620) );
  NOR2_X1 U15640 ( .A1(n15987), .A2(n12620), .ZN(n12634) );
  AOI22_X1 U15641 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12607) );
  AOI22_X1 U15642 ( .A1(n17256), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15949), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12606) );
  AOI22_X1 U15643 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12597) );
  OAI21_X1 U15644 ( .B1(n12446), .B2(n20889), .A(n12597), .ZN(n12604) );
  AOI22_X1 U15645 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12602) );
  AOI22_X1 U15646 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12601) );
  AOI22_X1 U15647 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12600) );
  AOI22_X1 U15648 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12599) );
  NAND4_X1 U15649 ( .A1(n12602), .A2(n12601), .A3(n12600), .A4(n12599), .ZN(
        n12603) );
  AOI22_X1 U15650 ( .A1(n17268), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12617) );
  AOI22_X1 U15651 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12616) );
  INV_X1 U15652 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n21060) );
  AOI22_X1 U15653 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15949), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12608) );
  OAI21_X1 U15654 ( .B1(n12446), .B2(n21060), .A(n12608), .ZN(n12614) );
  AOI22_X1 U15655 ( .A1(n17190), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9718), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12612) );
  AOI22_X1 U15656 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12611) );
  AOI22_X1 U15657 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13891), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12610) );
  AOI22_X1 U15658 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15952), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12609) );
  NAND4_X1 U15659 ( .A1(n12612), .A2(n12611), .A3(n12610), .A4(n12609), .ZN(
        n12613) );
  AOI211_X1 U15660 ( .C1(n17256), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n12614), .B(n12613), .ZN(n12615) );
  NAND3_X1 U15661 ( .A1(n12617), .A2(n12616), .A3(n12615), .ZN(n12635) );
  NAND2_X1 U15662 ( .A1(n17392), .A2(n12635), .ZN(n12618) );
  NAND3_X1 U15663 ( .A1(n18326), .A2(n12646), .A3(n13822), .ZN(n13823) );
  NAND2_X1 U15664 ( .A1(n17341), .A2(n17347), .ZN(n12629) );
  INV_X1 U15665 ( .A(n13822), .ZN(n18318) );
  NAND2_X1 U15666 ( .A1(n15987), .A2(n17341), .ZN(n15989) );
  INV_X1 U15667 ( .A(n15989), .ZN(n12619) );
  OAI21_X1 U15668 ( .B1(n12620), .B2(n12619), .A(n18932), .ZN(n12621) );
  OAI211_X1 U15669 ( .C1(n12629), .C2(n18318), .A(n17392), .B(n12621), .ZN(
        n12626) );
  NAND2_X1 U15670 ( .A1(n18932), .A2(n17392), .ZN(n12630) );
  NOR4_X1 U15671 ( .A1(n13822), .A2(n12635), .A3(n12630), .A4(n12629), .ZN(
        n12636) );
  NAND2_X1 U15672 ( .A1(n12647), .A2(n12636), .ZN(n15969) );
  OAI21_X1 U15673 ( .B1(n12622), .B2(n12626), .A(n15969), .ZN(n16668) );
  INV_X1 U15674 ( .A(n16668), .ZN(n16662) );
  NAND2_X1 U15675 ( .A1(n17554), .A2(n17494), .ZN(n13826) );
  INV_X1 U15676 ( .A(n12635), .ZN(n18314) );
  NAND2_X1 U15677 ( .A1(n18309), .A2(n18314), .ZN(n12637) );
  NOR2_X1 U15678 ( .A1(n17554), .A2(n12630), .ZN(n12623) );
  INV_X1 U15679 ( .A(n12626), .ZN(n12632) );
  AOI22_X1 U15680 ( .A1(n18314), .A2(n12630), .B1(n12629), .B2(n12628), .ZN(
        n12631) );
  NAND2_X1 U15681 ( .A1(n18326), .A2(n17347), .ZN(n16080) );
  NOR2_X1 U15682 ( .A1(n16080), .A2(n12633), .ZN(n15967) );
  NAND2_X1 U15683 ( .A1(n12636), .A2(n12638), .ZN(n15974) );
  NAND2_X1 U15684 ( .A1(n12715), .A2(n15974), .ZN(n18282) );
  INV_X1 U15685 ( .A(n12637), .ZN(n16010) );
  INV_X1 U15686 ( .A(n12638), .ZN(n16011) );
  XOR2_X1 U15687 ( .A(n12640), .B(n12639), .Z(n12642) );
  INV_X1 U15688 ( .A(n18772), .ZN(n15986) );
  AOI21_X1 U15689 ( .B1(n12644), .B2(n12643), .A(n15986), .ZN(n18773) );
  NAND2_X1 U15690 ( .A1(n12646), .A2(n12645), .ZN(n15968) );
  NOR2_X1 U15691 ( .A1(n18305), .A2(n12647), .ZN(n15985) );
  NAND2_X1 U15692 ( .A1(n15985), .A2(n17341), .ZN(n15982) );
  INV_X1 U15693 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18945) );
  NAND2_X1 U15694 ( .A1(n18893), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18796) );
  NAND2_X1 U15695 ( .A1(n16555), .A2(n17861), .ZN(n12689) );
  NOR2_X1 U15696 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18946) );
  INV_X1 U15697 ( .A(n18946), .ZN(n18896) );
  NAND2_X1 U15698 ( .A1(n18945), .A2(n18887), .ZN(n16664) );
  NAND2_X1 U15699 ( .A1(n18896), .A2(n16664), .ZN(n14045) );
  INV_X1 U15700 ( .A(n14045), .ZN(n18929) );
  NAND2_X1 U15701 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17872) );
  NAND2_X1 U15702 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17926) );
  NAND2_X1 U15703 ( .A1(n17871), .A2(n17829), .ZN(n17801) );
  NAND2_X1 U15704 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17803) );
  NAND2_X1 U15705 ( .A1(n17789), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12724) );
  NAND2_X1 U15706 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17765) );
  NAND2_X1 U15707 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17731) );
  NAND2_X1 U15708 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17695) );
  NAND2_X1 U15709 ( .A1(n17676), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17655) );
  NAND2_X1 U15710 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17656) );
  INV_X1 U15711 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17607) );
  INV_X1 U15712 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16726) );
  INV_X1 U15713 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16719) );
  NAND2_X1 U15714 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16535), .ZN(
        n16520) );
  XOR2_X2 U15715 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n16520), .Z(
        n16933) );
  INV_X1 U15716 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18874) );
  INV_X1 U15717 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18935) );
  NOR2_X1 U15718 ( .A1(n18874), .A2(n18280), .ZN(n16548) );
  NAND2_X1 U15719 ( .A1(n9828), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12648) );
  NOR2_X1 U15720 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18945), .ZN(n17690) );
  NOR2_X1 U15721 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18887), .ZN(
        n18909) );
  NOR2_X1 U15722 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18938) );
  AOI21_X1 U15723 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(
        P3_STATE2_REG_2__SCAN_IN), .A(n18938), .ZN(n18800) );
  NOR3_X2 U15724 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n16666), .ZN(n18641) );
  INV_X2 U15725 ( .A(n18313), .ZN(n18678) );
  OR2_X1 U15726 ( .A1(n12648), .A2(n17802), .ZN(n16523) );
  INV_X1 U15727 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16688) );
  XOR2_X1 U15728 ( .A(n16688), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n12650) );
  NOR2_X1 U15729 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17750), .ZN(
        n16537) );
  INV_X1 U15730 ( .A(n16536), .ZN(n16684) );
  NAND2_X1 U15731 ( .A1(n18678), .A2(n12648), .ZN(n12649) );
  OAI211_X1 U15732 ( .C1(n16684), .C2(n18804), .A(n12649), .B(n17968), .ZN(
        n16538) );
  NOR2_X1 U15733 ( .A1(n16537), .A2(n16538), .ZN(n16522) );
  OAI22_X1 U15734 ( .A1(n16523), .A2(n12650), .B1(n16522), .B2(n16688), .ZN(
        n12651) );
  AOI211_X1 U15735 ( .C1(n17730), .C2(n9959), .A(n16548), .B(n12651), .ZN(
        n12687) );
  NOR2_X1 U15736 ( .A1(n17967), .A2(n17491), .ZN(n12660) );
  NOR2_X1 U15737 ( .A1(n12660), .A2(n17479), .ZN(n12658) );
  NOR2_X1 U15738 ( .A1(n12658), .A2(n17472), .ZN(n12668) );
  NAND2_X1 U15739 ( .A1(n12668), .A2(n12652), .ZN(n12656) );
  NOR2_X1 U15740 ( .A1(n17464), .A2(n12656), .ZN(n12655) );
  NAND2_X1 U15741 ( .A1(n12655), .A2(n12653), .ZN(n12654) );
  NOR2_X1 U15742 ( .A1(n17458), .A2(n12654), .ZN(n12678) );
  INV_X1 U15743 ( .A(n17458), .ZN(n16006) );
  XNOR2_X1 U15744 ( .A(n12654), .B(n16006), .ZN(n17890) );
  XNOR2_X1 U15745 ( .A(n12655), .B(n17461), .ZN(n12671) );
  XOR2_X1 U15746 ( .A(n12656), .B(n17464), .Z(n12657) );
  NAND2_X1 U15747 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12657), .ZN(
        n12670) );
  INV_X1 U15748 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18222) );
  XNOR2_X1 U15749 ( .A(n18222), .B(n12657), .ZN(n17910) );
  XOR2_X1 U15750 ( .A(n17472), .B(n12658), .Z(n12659) );
  NAND2_X1 U15751 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12659), .ZN(
        n12666) );
  XNOR2_X1 U15752 ( .A(n18245), .B(n12659), .ZN(n17935) );
  XOR2_X1 U15753 ( .A(n17479), .B(n12660), .Z(n12664) );
  OR2_X1 U15754 ( .A1(n18254), .A2(n12664), .ZN(n12665) );
  INV_X1 U15755 ( .A(n17967), .ZN(n12663) );
  AOI21_X1 U15756 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12477), .A(
        n12663), .ZN(n12662) );
  NOR2_X1 U15757 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12477), .ZN(
        n12661) );
  AOI221_X1 U15758 ( .B1(n12663), .B2(n12477), .C1(n12662), .C2(n18911), .A(
        n12661), .ZN(n17947) );
  XNOR2_X1 U15759 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12664), .ZN(
        n17946) );
  NAND2_X1 U15760 ( .A1(n17947), .A2(n17946), .ZN(n17945) );
  NAND2_X1 U15761 ( .A1(n12665), .A2(n17945), .ZN(n17934) );
  NAND2_X1 U15762 ( .A1(n17935), .A2(n17934), .ZN(n17933) );
  NAND2_X1 U15763 ( .A1(n12666), .A2(n17933), .ZN(n12667) );
  NAND2_X1 U15764 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12667), .ZN(
        n12669) );
  XOR2_X1 U15765 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n12667), .Z(
        n17924) );
  XNOR2_X1 U15766 ( .A(n12668), .B(n17468), .ZN(n17923) );
  NAND2_X1 U15767 ( .A1(n17924), .A2(n17923), .ZN(n17922) );
  NAND2_X1 U15768 ( .A1(n12669), .A2(n17922), .ZN(n17909) );
  NAND2_X1 U15769 ( .A1(n17910), .A2(n17909), .ZN(n17908) );
  NAND2_X1 U15770 ( .A1(n12670), .A2(n17908), .ZN(n12672) );
  NAND2_X1 U15771 ( .A1(n12671), .A2(n12672), .ZN(n12673) );
  XOR2_X1 U15772 ( .A(n12672), .B(n12671), .Z(n17897) );
  NAND2_X1 U15773 ( .A1(n17897), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17896) );
  INV_X1 U15774 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18203) );
  NAND2_X1 U15775 ( .A1(n12678), .A2(n12674), .ZN(n12679) );
  INV_X1 U15776 ( .A(n12674), .ZN(n12677) );
  NAND2_X1 U15777 ( .A1(n17890), .A2(n17889), .ZN(n12676) );
  NAND2_X1 U15778 ( .A1(n12678), .A2(n12677), .ZN(n12675) );
  OAI211_X1 U15779 ( .C1(n12678), .C2(n12677), .A(n12676), .B(n12675), .ZN(
        n17866) );
  NAND2_X1 U15780 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17866), .ZN(
        n17865) );
  NAND2_X1 U15781 ( .A1(n15997), .A2(n17777), .ZN(n18104) );
  NAND2_X1 U15782 ( .A1(n18008), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17650) );
  NAND2_X1 U15783 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16533) );
  INV_X1 U15784 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16015) );
  NOR2_X1 U15785 ( .A1(n16533), .A2(n16015), .ZN(n16527) );
  NAND3_X1 U15786 ( .A1(n17978), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n16527), .ZN(n12681) );
  XOR2_X1 U15787 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12681), .Z(
        n16558) );
  NAND3_X1 U15788 ( .A1(n16527), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n18892), .ZN(n16552) );
  INV_X1 U15789 ( .A(n17666), .ZN(n18010) );
  NOR2_X1 U15790 ( .A1(n18018), .A2(n18010), .ZN(n17649) );
  NAND2_X1 U15791 ( .A1(n17974), .A2(n17649), .ZN(n17981) );
  INV_X1 U15792 ( .A(n17981), .ZN(n17612) );
  NAND2_X1 U15793 ( .A1(n16527), .A2(n17612), .ZN(n16005) );
  OAI21_X1 U15794 ( .B1(n16066), .B2(n16005), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12683) );
  OAI21_X1 U15795 ( .B1(n16552), .B2(n17981), .A(n12683), .ZN(n16550) );
  NOR2_X2 U15796 ( .A1(n16006), .A2(n17971), .ZN(n17881) );
  INV_X1 U15797 ( .A(n12685), .ZN(n12686) );
  AND2_X1 U15798 ( .A1(n12687), .A2(n12686), .ZN(n12688) );
  NOR4_X1 U15799 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n12693) );
  NOR4_X1 U15800 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n12692) );
  NOR4_X1 U15801 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12691) );
  NOR4_X1 U15802 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n12690) );
  AND4_X1 U15803 ( .A1(n12693), .A2(n12692), .A3(n12691), .A4(n12690), .ZN(
        n12698) );
  NOR4_X1 U15804 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_7__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n12696) );
  NOR4_X1 U15805 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n12695) );
  NOR4_X1 U15806 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n12694) );
  INV_X1 U15807 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20738) );
  AND4_X1 U15808 ( .A1(n12696), .A2(n12695), .A3(n12694), .A4(n20738), .ZN(
        n12697) );
  NAND2_X1 U15809 ( .A1(n12698), .A2(n12697), .ZN(n12699) );
  AND2_X2 U15810 ( .A1(n12699), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20130)
         );
  INV_X1 U15811 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20808) );
  NOR3_X1 U15812 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20808), .ZN(n12701) );
  NOR4_X1 U15813 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12700) );
  NAND4_X1 U15814 ( .A1(n20130), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12701), .A4(
        n12700), .ZN(U214) );
  NOR4_X1 U15815 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12705) );
  NOR4_X1 U15816 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12704) );
  NOR4_X1 U15817 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12703) );
  NOR4_X1 U15818 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12702) );
  NAND4_X1 U15819 ( .A1(n12705), .A2(n12704), .A3(n12703), .A4(n12702), .ZN(
        n12710) );
  NOR4_X1 U15820 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n12708) );
  NOR4_X1 U15821 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12707) );
  NOR4_X1 U15822 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12706) );
  INV_X1 U15823 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19842) );
  NAND4_X1 U15824 ( .A1(n12708), .A2(n12707), .A3(n12706), .A4(n19842), .ZN(
        n12709) );
  OAI21_X1 U15825 ( .B1(n12710), .B2(n12709), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12711) );
  INV_X1 U15826 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19933) );
  NOR2_X1 U15827 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(n19933), .ZN(n12713) );
  NOR4_X1 U15828 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .A3(P2_BE_N_REG_3__SCAN_IN), .A4(P2_D_C_N_REG_SCAN_IN), .ZN(n12712) );
  INV_X1 U15829 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n20917) );
  NAND4_X1 U15830 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(n12713), .A3(n12712), .A4(
        n20917), .ZN(n12714) );
  NOR2_X1 U15831 ( .A1(n13962), .A2(n12714), .ZN(n16578) );
  NAND2_X1 U15832 ( .A1(n16578), .A2(U214), .ZN(U212) );
  NOR2_X1 U15833 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12714), .ZN(n16651)
         );
  NOR3_X1 U15834 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17020) );
  INV_X1 U15835 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17319) );
  NAND2_X1 U15836 ( .A1(n17020), .A2(n17319), .ZN(n17014) );
  NOR2_X1 U15837 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17014), .ZN(n16993) );
  NAND2_X1 U15838 ( .A1(n16993), .A2(n17307), .ZN(n16988) );
  INV_X1 U15839 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17310) );
  NAND2_X1 U15840 ( .A1(n16969), .A2(n17310), .ZN(n16964) );
  INV_X1 U15841 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16930) );
  NAND2_X1 U15842 ( .A1(n16942), .A2(n16930), .ZN(n16929) );
  INV_X1 U15843 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n20906) );
  NAND2_X1 U15844 ( .A1(n16922), .A2(n20906), .ZN(n16914) );
  INV_X1 U15845 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16890) );
  NAND2_X1 U15846 ( .A1(n16895), .A2(n16890), .ZN(n16889) );
  INV_X1 U15847 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16862) );
  NAND2_X1 U15848 ( .A1(n16871), .A2(n16862), .ZN(n16861) );
  INV_X1 U15849 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16840) );
  NAND2_X1 U15850 ( .A1(n16848), .A2(n16840), .ZN(n16839) );
  INV_X1 U15851 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16823) );
  NAND2_X1 U15852 ( .A1(n16824), .A2(n16823), .ZN(n16820) );
  INV_X1 U15853 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17141) );
  NAND2_X1 U15854 ( .A1(n16804), .A2(n17141), .ZN(n16797) );
  NOR2_X1 U15855 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16797), .ZN(n16782) );
  INV_X1 U15856 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16773) );
  NAND2_X1 U15857 ( .A1(n16782), .A2(n16773), .ZN(n16772) );
  NOR2_X1 U15858 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16772), .ZN(n16743) );
  INV_X1 U15859 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16754) );
  NAND2_X1 U15860 ( .A1(n16743), .A2(n16754), .ZN(n12718) );
  NOR2_X1 U15861 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n12718), .ZN(n16739) );
  NAND2_X1 U15862 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18927) );
  INV_X1 U15863 ( .A(n12715), .ZN(n18733) );
  INV_X1 U15864 ( .A(n12716), .ZN(n17552) );
  NAND2_X1 U15865 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n17554), .ZN(n12717) );
  AOI211_X4 U15866 ( .C1(n16666), .C2(n18927), .A(n12734), .B(n12717), .ZN(
        n17015) );
  AOI211_X1 U15867 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n12718), .A(n16739), .B(
        n17049), .ZN(n12740) );
  INV_X1 U15868 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18867) );
  INV_X1 U15869 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18818) );
  INV_X2 U15870 ( .A(n18943), .ZN(n18942) );
  NAND2_X2 U15871 ( .A1(n18942), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18876) );
  OAI211_X1 U15872 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18818), .B(n18876), .ZN(n15983) );
  INV_X1 U15873 ( .A(n15983), .ZN(n18931) );
  OAI211_X1 U15874 ( .C1(n18931), .C2(n17554), .A(n18927), .B(n16666), .ZN(
        n18785) );
  INV_X1 U15875 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18865) );
  INV_X1 U15876 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18860) );
  INV_X1 U15877 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18847) );
  INV_X1 U15878 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18844) );
  INV_X1 U15879 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18832) );
  INV_X1 U15880 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18829) );
  INV_X1 U15881 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18825) );
  NAND2_X1 U15882 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17030) );
  NOR2_X1 U15883 ( .A1(n18825), .A2(n17030), .ZN(n17002) );
  NAND2_X1 U15884 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17002), .ZN(n16985) );
  NOR2_X1 U15885 ( .A1(n18829), .A2(n16985), .ZN(n16956) );
  NAND2_X1 U15886 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16956), .ZN(n16967) );
  NOR2_X1 U15887 ( .A1(n18832), .A2(n16967), .ZN(n16950) );
  NAND2_X1 U15888 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16950), .ZN(n16921) );
  INV_X1 U15889 ( .A(n16921), .ZN(n16948) );
  INV_X1 U15890 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18838) );
  INV_X1 U15891 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18836) );
  NOR2_X1 U15892 ( .A1(n18838), .A2(n18836), .ZN(n16908) );
  AND3_X1 U15893 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16948), .A3(n16908), 
        .ZN(n16902) );
  NAND2_X1 U15894 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16902), .ZN(n16870) );
  NOR3_X1 U15895 ( .A1(n18847), .A2(n18844), .A3(n16870), .ZN(n16785) );
  INV_X1 U15896 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n21058) );
  INV_X1 U15897 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n20997) );
  INV_X1 U15898 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18852) );
  NAND2_X1 U15899 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16837) );
  NOR2_X1 U15900 ( .A1(n18852), .A2(n16837), .ZN(n16811) );
  NAND2_X1 U15901 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16811), .ZN(n16812) );
  NOR2_X1 U15902 ( .A1(n20997), .A2(n16812), .ZN(n16801) );
  NAND2_X1 U15903 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16801), .ZN(n16786) );
  NOR2_X1 U15904 ( .A1(n21058), .A2(n16786), .ZN(n16779) );
  NAND3_X1 U15905 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16785), .A3(n16779), 
        .ZN(n16777) );
  NOR2_X1 U15906 ( .A1(n18860), .A2(n16777), .ZN(n16761) );
  NAND2_X1 U15907 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16761), .ZN(n16747) );
  NOR2_X1 U15908 ( .A1(n18865), .A2(n16747), .ZN(n12719) );
  NAND2_X1 U15909 ( .A1(n17031), .A2(n12719), .ZN(n16686) );
  NOR4_X4 U15910 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n18893), .ZN(n16974) );
  NOR2_X1 U15911 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18887), .ZN(n18794) );
  INV_X1 U15912 ( .A(n18794), .ZN(n18637) );
  NOR2_X1 U15913 ( .A1(n18796), .A2(n18637), .ZN(n18789) );
  NOR4_X2 U15914 ( .A1(n18125), .A2(n18948), .A3(n16974), .A4(n18789), .ZN(
        n17045) );
  OAI221_X1 U15915 ( .B1(n17041), .B2(P3_REIP_REG_26__SCAN_IN), .C1(n17041), 
        .C2(n12719), .A(n17053), .ZN(n16736) );
  INV_X1 U15916 ( .A(n16736), .ZN(n12720) );
  AOI21_X1 U15917 ( .B1(n18867), .B2(n16686), .A(n12720), .ZN(n12739) );
  INV_X1 U15918 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17636) );
  INV_X1 U15919 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17961) );
  INV_X1 U15920 ( .A(n12721), .ZN(n17637) );
  NOR2_X1 U15921 ( .A1(n17961), .A2(n17637), .ZN(n17605) );
  INV_X1 U15922 ( .A(n17605), .ZN(n12722) );
  NOR2_X1 U15923 ( .A1(n17636), .A2(n12722), .ZN(n16682) );
  AOI21_X1 U15924 ( .B1(n17636), .B2(n12722), .A(n16682), .ZN(n17639) );
  INV_X1 U15925 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16748) );
  INV_X1 U15926 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16768) );
  NAND2_X1 U15927 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17676), .ZN(
        n12730) );
  NOR2_X1 U15928 ( .A1(n16768), .A2(n12730), .ZN(n12732) );
  NAND2_X1 U15929 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n12732), .ZN(
        n12723) );
  AOI21_X1 U15930 ( .B1(n16748), .B2(n12723), .A(n17605), .ZN(n17648) );
  AOI21_X1 U15931 ( .B1(n16768), .B2(n12730), .A(n12732), .ZN(n17677) );
  INV_X1 U15932 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17704) );
  INV_X1 U15933 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n20989) );
  NAND2_X1 U15934 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17720), .ZN(
        n17689) );
  NOR2_X1 U15935 ( .A1(n20989), .A2(n17689), .ZN(n12729) );
  XNOR2_X1 U15936 ( .A(n17704), .B(n12729), .ZN(n17712) );
  INV_X1 U15937 ( .A(n17765), .ZN(n12725) );
  NOR2_X1 U15938 ( .A1(n17961), .A2(n12724), .ZN(n17764) );
  NAND2_X1 U15939 ( .A1(n12725), .A2(n17764), .ZN(n16835) );
  NOR2_X1 U15940 ( .A1(n9958), .A2(n16835), .ZN(n17728) );
  NAND2_X1 U15941 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17728), .ZN(
        n16825) );
  INV_X1 U15942 ( .A(n16825), .ZN(n12727) );
  NAND2_X1 U15943 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17764), .ZN(
        n16858) );
  NOR2_X1 U15944 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16858), .ZN(
        n16857) );
  OAI21_X1 U15945 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n12727), .A(
        n17689), .ZN(n12728) );
  INV_X1 U15946 ( .A(n12728), .ZN(n17729) );
  AOI21_X1 U15947 ( .B1(n20989), .B2(n17689), .A(n12729), .ZN(n17721) );
  NOR2_X1 U15948 ( .A1(n16790), .A2(n16933), .ZN(n16781) );
  INV_X1 U15949 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17698) );
  NAND2_X1 U15950 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12729), .ZN(
        n12731) );
  INV_X1 U15951 ( .A(n12730), .ZN(n17646) );
  AOI21_X1 U15952 ( .B1(n17698), .B2(n12731), .A(n17646), .ZN(n17693) );
  NOR2_X1 U15953 ( .A1(n16780), .A2(n16933), .ZN(n16767) );
  XOR2_X1 U15954 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n12732), .Z(
        n17660) );
  NOR2_X1 U15955 ( .A1(n17648), .A2(n16745), .ZN(n16744) );
  NOR2_X1 U15956 ( .A1(n16744), .A2(n16933), .ZN(n12733) );
  INV_X1 U15957 ( .A(n16974), .ZN(n18799) );
  AOI211_X1 U15958 ( .C1(n17639), .C2(n12733), .A(n16683), .B(n18799), .ZN(
        n12738) );
  INV_X1 U15959 ( .A(n18785), .ZN(n12735) );
  AOI211_X4 U15960 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n17554), .A(n12735), .B(
        n12734), .ZN(n17019) );
  INV_X1 U15961 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n12736) );
  OAI22_X1 U15962 ( .A1(n17636), .A2(n17035), .B1(n17050), .B2(n12736), .ZN(
        n12737) );
  OR4_X1 U15963 ( .A1(n12740), .A2(n12739), .A3(n12738), .A4(n12737), .ZN(
        P3_U2645) );
  INV_X1 U15964 ( .A(n15925), .ZN(n16516) );
  INV_X1 U15965 ( .A(n12752), .ZN(n12741) );
  INV_X1 U15966 ( .A(n11913), .ZN(n13332) );
  NAND2_X1 U15967 ( .A1(n12741), .A2(n13332), .ZN(n19130) );
  INV_X1 U15968 ( .A(n19130), .ZN(n12744) );
  INV_X1 U15969 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n21023) );
  NOR2_X1 U15970 ( .A1(n12752), .A2(n12742), .ZN(n13646) );
  NOR2_X1 U15971 ( .A1(n13646), .A2(n12743), .ZN(n12746) );
  OAI21_X1 U15972 ( .B1(n12744), .B2(n21023), .A(n12746), .ZN(P2_U2814) );
  NOR2_X1 U15973 ( .A1(n12744), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n12747)
         );
  AOI22_X1 U15974 ( .A1(n12747), .A2(n12746), .B1(n12745), .B2(n19953), .ZN(
        P2_U3612) );
  AND2_X1 U15975 ( .A1(n12357), .A2(n16075), .ZN(n12946) );
  NOR4_X1 U15976 ( .A1(n12949), .A2(n13321), .A3(n12946), .A4(n13346), .ZN(
        n13331) );
  NOR2_X1 U15977 ( .A1(n13331), .A2(n16516), .ZN(n19934) );
  NAND2_X1 U15978 ( .A1(n16507), .A2(n19937), .ZN(n12748) );
  NAND2_X1 U15979 ( .A1(n12748), .A2(n13335), .ZN(n12749) );
  NAND2_X1 U15980 ( .A1(n12749), .A2(n15925), .ZN(n12884) );
  OAI21_X1 U15981 ( .B1(n19934), .B2(n12750), .A(n12884), .ZN(P2_U2819) );
  INV_X1 U15982 ( .A(n13349), .ZN(n12751) );
  NOR2_X4 U15983 ( .A1(n12752), .A2(n12751), .ZN(n19272) );
  NAND2_X1 U15984 ( .A1(n13646), .A2(n16075), .ZN(n12753) );
  AND2_X2 U15985 ( .A1(n12835), .A2(n12753), .ZN(n19273) );
  AOI22_X1 U15986 ( .A1(n19273), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n19272), .ZN(n12756) );
  NOR2_X2 U15987 ( .A1(n12753), .A2(n14263), .ZN(n12806) );
  NAND2_X1 U15988 ( .A1(n13962), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12755) );
  INV_X1 U15989 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n21045) );
  OR2_X1 U15990 ( .A1(n13962), .A2(n21045), .ZN(n12754) );
  NAND2_X1 U15991 ( .A1(n12755), .A2(n12754), .ZN(n19197) );
  NAND2_X1 U15992 ( .A1(n12806), .A2(n19197), .ZN(n12758) );
  NAND2_X1 U15993 ( .A1(n12756), .A2(n12758), .ZN(P2_U2961) );
  INV_X1 U15994 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19252) );
  NAND2_X1 U15995 ( .A1(n19273), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n12757) );
  OAI211_X1 U15996 ( .C1(n19252), .C2(n12835), .A(n12758), .B(n12757), .ZN(
        P2_U2976) );
  NAND2_X1 U15997 ( .A1(n13962), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12760) );
  INV_X1 U15998 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14050) );
  OR2_X1 U15999 ( .A1(n13962), .A2(n14050), .ZN(n12759) );
  NAND2_X1 U16000 ( .A1(n12760), .A2(n12759), .ZN(n19184) );
  NAND2_X1 U16001 ( .A1(n12806), .A2(n19184), .ZN(n12771) );
  NAND2_X1 U16002 ( .A1(n19273), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12761) );
  OAI211_X1 U16003 ( .C1(n12337), .C2(n12835), .A(n12771), .B(n12761), .ZN(
        P2_U2966) );
  INV_X1 U16004 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n20992) );
  MUX2_X1 U16005 ( .A(BUF1_REG_8__SCAN_IN), .B(BUF2_REG_8__SCAN_IN), .S(n13962), .Z(n19200) );
  NAND2_X1 U16006 ( .A1(n12806), .A2(n19200), .ZN(n12767) );
  NAND2_X1 U16007 ( .A1(n19273), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n12762) );
  OAI211_X1 U16008 ( .C1(n20992), .C2(n12835), .A(n12767), .B(n12762), .ZN(
        P2_U2975) );
  INV_X1 U16009 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n12843) );
  NAND2_X1 U16010 ( .A1(n13962), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12764) );
  INV_X1 U16011 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16608) );
  OR2_X1 U16012 ( .A1(n13962), .A2(n16608), .ZN(n12763) );
  NAND2_X1 U16013 ( .A1(n12764), .A2(n12763), .ZN(n19194) );
  NAND2_X1 U16014 ( .A1(n12806), .A2(n19194), .ZN(n12769) );
  NAND2_X1 U16015 ( .A1(n19273), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12765) );
  OAI211_X1 U16016 ( .C1(n12843), .C2(n12835), .A(n12769), .B(n12765), .ZN(
        P2_U2962) );
  INV_X1 U16017 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n12850) );
  NAND2_X1 U16018 ( .A1(n19273), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12766) );
  OAI211_X1 U16019 ( .C1(n12850), .C2(n12835), .A(n12767), .B(n12766), .ZN(
        P2_U2960) );
  INV_X1 U16020 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19250) );
  NAND2_X1 U16021 ( .A1(n19273), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12768) );
  OAI211_X1 U16022 ( .C1(n19250), .C2(n12835), .A(n12769), .B(n12768), .ZN(
        P2_U2977) );
  INV_X1 U16023 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19244) );
  NAND2_X1 U16024 ( .A1(n19273), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n12770) );
  OAI211_X1 U16025 ( .C1(n19244), .C2(n12835), .A(n12771), .B(n12770), .ZN(
        P2_U2981) );
  INV_X1 U16026 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n20977) );
  MUX2_X1 U16027 ( .A(BUF1_REG_12__SCAN_IN), .B(BUF2_REG_12__SCAN_IN), .S(
        n13962), .Z(n19189) );
  NAND2_X1 U16028 ( .A1(n12806), .A2(n19189), .ZN(n19274) );
  NAND2_X1 U16029 ( .A1(n19273), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12772) );
  OAI211_X1 U16030 ( .C1(n20977), .C2(n12835), .A(n19274), .B(n12772), .ZN(
        P2_U2964) );
  AOI22_X1 U16031 ( .A1(n19273), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19272), .ZN(n12776) );
  INV_X1 U16032 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14639) );
  OR2_X1 U16033 ( .A1(n13962), .A2(n14639), .ZN(n12774) );
  NAND2_X1 U16034 ( .A1(n13962), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12773) );
  AND2_X1 U16035 ( .A1(n12774), .A2(n12773), .ZN(n19187) );
  INV_X1 U16036 ( .A(n19187), .ZN(n12775) );
  NAND2_X1 U16037 ( .A1(n12806), .A2(n12775), .ZN(n12793) );
  NAND2_X1 U16038 ( .A1(n12776), .A2(n12793), .ZN(P2_U2965) );
  AOI22_X1 U16039 ( .A1(n19273), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19272), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12777) );
  INV_X1 U16040 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16618) );
  INV_X1 U16041 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18308) );
  AOI22_X1 U16042 ( .A1(n13961), .A2(n16618), .B1(n18308), .B2(n13962), .ZN(
        n16311) );
  NAND2_X1 U16043 ( .A1(n12806), .A2(n16311), .ZN(n12787) );
  NAND2_X1 U16044 ( .A1(n12777), .A2(n12787), .ZN(P2_U2969) );
  AOI22_X1 U16045 ( .A1(n19273), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19272), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12778) );
  AOI22_X1 U16046 ( .A1(n13961), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13962), .ZN(n19344) );
  INV_X1 U16047 ( .A(n19344), .ZN(n15467) );
  NAND2_X1 U16048 ( .A1(n12806), .A2(n15467), .ZN(n12795) );
  NAND2_X1 U16049 ( .A1(n12778), .A2(n12795), .ZN(P2_U2959) );
  AOI22_X1 U16050 ( .A1(n19273), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19272), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12779) );
  AOI22_X1 U16051 ( .A1(n13961), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13962), .ZN(n19326) );
  INV_X1 U16052 ( .A(n19326), .ZN(n19208) );
  NAND2_X1 U16053 ( .A1(n12806), .A2(n19208), .ZN(n12785) );
  NAND2_X1 U16054 ( .A1(n12779), .A2(n12785), .ZN(P2_U2972) );
  AOI22_X1 U16055 ( .A1(n19273), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n19272), .ZN(n12783) );
  INV_X1 U16056 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n12780) );
  OR2_X1 U16057 ( .A1(n13962), .A2(n12780), .ZN(n12782) );
  NAND2_X1 U16058 ( .A1(n13962), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12781) );
  AND2_X1 U16059 ( .A1(n12782), .A2(n12781), .ZN(n19192) );
  INV_X1 U16060 ( .A(n19192), .ZN(n15441) );
  NAND2_X1 U16061 ( .A1(n12806), .A2(n15441), .ZN(n12789) );
  NAND2_X1 U16062 ( .A1(n12783), .A2(n12789), .ZN(P2_U2963) );
  AOI22_X1 U16063 ( .A1(n19273), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19272), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12784) );
  AOI22_X1 U16064 ( .A1(n13961), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13962), .ZN(n19320) );
  INV_X1 U16065 ( .A(n19320), .ZN(n14023) );
  NAND2_X1 U16066 ( .A1(n12806), .A2(n14023), .ZN(n12802) );
  NAND2_X1 U16067 ( .A1(n12784), .A2(n12802), .ZN(P2_U2955) );
  AOI22_X1 U16068 ( .A1(n19273), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19272), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12786) );
  NAND2_X1 U16069 ( .A1(n12786), .A2(n12785), .ZN(P2_U2957) );
  AOI22_X1 U16070 ( .A1(n19273), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19272), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n12788) );
  NAND2_X1 U16071 ( .A1(n12788), .A2(n12787), .ZN(P2_U2954) );
  AOI22_X1 U16072 ( .A1(n19273), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n19272), .ZN(n12790) );
  NAND2_X1 U16073 ( .A1(n12790), .A2(n12789), .ZN(P2_U2978) );
  AOI22_X1 U16074 ( .A1(n19273), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19272), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12791) );
  OAI22_X1 U16075 ( .A1(n13962), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13961), .ZN(n19223) );
  INV_X1 U16076 ( .A(n19223), .ZN(n16304) );
  NAND2_X1 U16077 ( .A1(n12806), .A2(n16304), .ZN(n12804) );
  NAND2_X1 U16078 ( .A1(n12791), .A2(n12804), .ZN(P2_U2971) );
  AOI22_X1 U16079 ( .A1(n19273), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_17__SCAN_IN), .B2(n19272), .ZN(n12792) );
  AOI22_X1 U16080 ( .A1(n13961), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13962), .ZN(n19313) );
  INV_X1 U16081 ( .A(n19313), .ZN(n13964) );
  NAND2_X1 U16082 ( .A1(n12806), .A2(n13964), .ZN(n12800) );
  NAND2_X1 U16083 ( .A1(n12792), .A2(n12800), .ZN(P2_U2953) );
  AOI22_X1 U16084 ( .A1(n19273), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n19272), .ZN(n12794) );
  NAND2_X1 U16085 ( .A1(n12794), .A2(n12793), .ZN(P2_U2980) );
  AOI22_X1 U16086 ( .A1(n19273), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19272), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n12796) );
  NAND2_X1 U16087 ( .A1(n12796), .A2(n12795), .ZN(P2_U2974) );
  AOI22_X1 U16088 ( .A1(n19273), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19272), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12797) );
  OAI22_X1 U16089 ( .A1(n13962), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13961), .ZN(n19331) );
  INV_X1 U16090 ( .A(n19331), .ZN(n16298) );
  NAND2_X1 U16091 ( .A1(n12806), .A2(n16298), .ZN(n12798) );
  NAND2_X1 U16092 ( .A1(n12797), .A2(n12798), .ZN(P2_U2973) );
  AOI22_X1 U16093 ( .A1(n19273), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n19272), .ZN(n12799) );
  NAND2_X1 U16094 ( .A1(n12799), .A2(n12798), .ZN(P2_U2958) );
  AOI22_X1 U16095 ( .A1(n19273), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19272), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12801) );
  NAND2_X1 U16096 ( .A1(n12801), .A2(n12800), .ZN(P2_U2968) );
  AOI22_X1 U16097 ( .A1(n19273), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19272), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n12803) );
  NAND2_X1 U16098 ( .A1(n12803), .A2(n12802), .ZN(P2_U2970) );
  AOI22_X1 U16099 ( .A1(n19273), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n19272), .ZN(n12805) );
  NAND2_X1 U16100 ( .A1(n12805), .A2(n12804), .ZN(P2_U2956) );
  INV_X1 U16101 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n12807) );
  INV_X1 U16102 ( .A(n19273), .ZN(n12811) );
  INV_X1 U16103 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n12975) );
  INV_X1 U16104 ( .A(n12806), .ZN(n12810) );
  INV_X1 U16105 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16625) );
  INV_X1 U16106 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18296) );
  AOI22_X1 U16107 ( .A1(n13961), .A2(n16625), .B1(n18296), .B2(n13962), .ZN(
        n19171) );
  INV_X1 U16108 ( .A(n19171), .ZN(n13678) );
  OAI222_X1 U16109 ( .A1(n12807), .A2(n12811), .B1(n12835), .B2(n12975), .C1(
        n12810), .C2(n13678), .ZN(P2_U2952) );
  INV_X1 U16110 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n12808) );
  OAI222_X1 U16111 ( .A1(n12808), .A2(n12811), .B1(n12810), .B2(n13678), .C1(
        n12835), .C2(n12966), .ZN(P2_U2967) );
  INV_X1 U16112 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12812) );
  AOI22_X1 U16113 ( .A1(n13961), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13962), .ZN(n19181) );
  INV_X1 U16114 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12809) );
  OAI222_X1 U16115 ( .A1(n12812), .A2(n12811), .B1(n12810), .B2(n19181), .C1(
        n12809), .C2(n12835), .ZN(P2_U2982) );
  INV_X1 U16116 ( .A(n13330), .ZN(n12813) );
  NAND2_X1 U16117 ( .A1(n12813), .A2(n13326), .ZN(n13280) );
  NAND2_X1 U16118 ( .A1(n13280), .A2(n13265), .ZN(n12815) );
  NAND2_X1 U16119 ( .A1(n15348), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12817) );
  NOR2_X2 U16120 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19894) );
  AOI22_X1 U16121 ( .A1(n12986), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19894), .B2(n19931), .ZN(n12818) );
  NOR2_X1 U16122 ( .A1(n15348), .A2(n16510), .ZN(n12827) );
  AOI21_X1 U16123 ( .B1(n19944), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12820) );
  AND2_X1 U16124 ( .A1(n12827), .A2(n12820), .ZN(n12821) );
  NAND2_X1 U16125 ( .A1(n19164), .A2(n12957), .ZN(n19165) );
  NAND2_X1 U16126 ( .A1(n13708), .A2(n19151), .ZN(n12823) );
  NAND2_X1 U16127 ( .A1(n19164), .A2(n12816), .ZN(n12822) );
  OAI211_X1 U16128 ( .C1(n19164), .C2(n12824), .A(n12823), .B(n12822), .ZN(
        P2_U2887) );
  NAND2_X1 U16129 ( .A1(n12986), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12825) );
  NAND2_X1 U16130 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19922), .ZN(
        n19566) );
  NAND2_X1 U16131 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19931), .ZN(
        n19598) );
  NAND2_X1 U16132 ( .A1(n19566), .A2(n19598), .ZN(n13669) );
  NAND2_X1 U16133 ( .A1(n19894), .A2(n13669), .ZN(n19601) );
  NAND2_X1 U16134 ( .A1(n12825), .A2(n19601), .ZN(n12826) );
  INV_X1 U16135 ( .A(n14258), .ZN(n14236) );
  XNOR2_X1 U16136 ( .A(n12829), .B(n12926), .ZN(n12831) );
  NAND2_X1 U16137 ( .A1(n12830), .A2(n12831), .ZN(n12929) );
  OR2_X1 U16138 ( .A1(n12831), .A2(n12830), .ZN(n12832) );
  NOR2_X1 U16139 ( .A1(n19164), .A2(n11670), .ZN(n12833) );
  AOI21_X1 U16140 ( .B1(n19164), .B2(n15917), .A(n12833), .ZN(n12834) );
  OAI21_X1 U16141 ( .B1(n19915), .B2(n19165), .A(n12834), .ZN(P2_U2886) );
  NAND2_X1 U16142 ( .A1(n13332), .A2(n15925), .ZN(n12836) );
  OAI21_X1 U16143 ( .B1(n13282), .B2(n12836), .A(n12835), .ZN(n12837) );
  NAND2_X1 U16144 ( .A1(n19259), .A2(n11376), .ZN(n12978) );
  NOR2_X1 U16145 ( .A1(n19685), .A2(n12874), .ZN(n19928) );
  INV_X1 U16146 ( .A(n19928), .ZN(n13352) );
  NOR2_X1 U16147 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13352), .ZN(n12976) );
  INV_X1 U16148 ( .A(n12976), .ZN(n19951) );
  AOI22_X1 U16149 ( .A1(n19269), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n12970), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12838) );
  OAI21_X1 U16150 ( .B1(n12839), .B2(n12978), .A(n12838), .ZN(P2_U2928) );
  INV_X1 U16151 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n12841) );
  AOI22_X1 U16152 ( .A1(n12976), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n12970), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12840) );
  OAI21_X1 U16153 ( .B1(n12841), .B2(n12978), .A(n12840), .ZN(P2_U2926) );
  AOI22_X1 U16154 ( .A1(n19269), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n12970), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12842) );
  OAI21_X1 U16155 ( .B1(n12843), .B2(n12978), .A(n12842), .ZN(P2_U2925) );
  INV_X1 U16156 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n12845) );
  AOI22_X1 U16157 ( .A1(n12976), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n12970), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n12844) );
  OAI21_X1 U16158 ( .B1(n12845), .B2(n12978), .A(n12844), .ZN(P2_U2929) );
  AOI22_X1 U16159 ( .A1(n19269), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n12970), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12846) );
  OAI21_X1 U16160 ( .B1(n14348), .B2(n12978), .A(n12846), .ZN(P2_U2922) );
  AOI22_X1 U16161 ( .A1(n12976), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n12970), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12847) );
  OAI21_X1 U16162 ( .B1(n12848), .B2(n12978), .A(n12847), .ZN(P2_U2924) );
  AOI22_X1 U16163 ( .A1(n19269), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n12970), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12849) );
  OAI21_X1 U16164 ( .B1(n12850), .B2(n12978), .A(n12849), .ZN(P2_U2927) );
  INV_X1 U16165 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n12852) );
  AOI22_X1 U16166 ( .A1(n12976), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n12970), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12851) );
  OAI21_X1 U16167 ( .B1(n12852), .B2(n12978), .A(n12851), .ZN(P2_U2930) );
  INV_X1 U16168 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n12854) );
  AOI22_X1 U16169 ( .A1(n12976), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n12970), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12853) );
  OAI21_X1 U16170 ( .B1(n12854), .B2(n12978), .A(n12853), .ZN(P2_U2932) );
  AOI22_X1 U16171 ( .A1(n12976), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n12970), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12855) );
  OAI21_X1 U16172 ( .B1(n20977), .B2(n12978), .A(n12855), .ZN(P2_U2923) );
  INV_X1 U16173 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n12857) );
  AOI22_X1 U16174 ( .A1(n12976), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n12970), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12856) );
  OAI21_X1 U16175 ( .B1(n12857), .B2(n12978), .A(n12856), .ZN(P2_U2931) );
  INV_X1 U16176 ( .A(n12859), .ZN(n12867) );
  NOR4_X1 U16177 ( .A1(n12863), .A2(n12862), .A3(n12861), .A4(n12860), .ZN(
        n12864) );
  OR2_X1 U16178 ( .A1(n12865), .A2(n12864), .ZN(n13052) );
  NOR2_X1 U16179 ( .A1(n13052), .A2(n19964), .ZN(n12866) );
  NAND2_X1 U16180 ( .A1(n12867), .A2(n12866), .ZN(n14353) );
  INV_X1 U16181 ( .A(n12868), .ZN(n12869) );
  INV_X1 U16182 ( .A(n20817), .ZN(n12872) );
  NAND2_X1 U16183 ( .A1(n20661), .A2(n20714), .ZN(n19967) );
  INV_X1 U16184 ( .A(n19967), .ZN(n12870) );
  OAI21_X1 U16185 ( .B1(n12870), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n12872), 
        .ZN(n12871) );
  OAI21_X1 U16186 ( .B1(n12873), .B2(n12872), .A(n12871), .ZN(P1_U3487) );
  AOI21_X1 U16187 ( .B1(n19685), .B2(n12874), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19947) );
  NAND2_X1 U16188 ( .A1(n13352), .A2(n19947), .ZN(n12875) );
  INV_X1 U16189 ( .A(n12884), .ZN(n12878) );
  NAND2_X1 U16190 ( .A1(n12878), .A2(n19944), .ZN(n16421) );
  OAI21_X1 U16191 ( .B1(n19124), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12877), .ZN(n16497) );
  INV_X1 U16192 ( .A(n16497), .ZN(n12882) );
  OAI21_X1 U16193 ( .B1(n12880), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12879), .ZN(n16502) );
  NAND2_X1 U16194 ( .A1(n19276), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n16500) );
  OAI21_X1 U16195 ( .B1(n16418), .B2(n16502), .A(n16500), .ZN(n12881) );
  AOI21_X1 U16196 ( .B1(n19285), .B2(n12882), .A(n12881), .ZN(n12888) );
  OR2_X1 U16197 ( .A1(n19894), .A2(n15937), .ZN(n19913) );
  NAND2_X1 U16198 ( .A1(n19913), .A2(n16510), .ZN(n12883) );
  INV_X1 U16199 ( .A(n12981), .ZN(n12886) );
  NAND2_X1 U16200 ( .A1(n19941), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12885) );
  NAND2_X1 U16201 ( .A1(n12886), .A2(n12885), .ZN(n13779) );
  OAI21_X1 U16202 ( .B1(n19284), .B2(n13779), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12887) );
  OAI211_X1 U16203 ( .C1(n13674), .C2(n12889), .A(n12888), .B(n12887), .ZN(
        P2_U3014) );
  NAND2_X1 U16204 ( .A1(n12891), .A2(n12890), .ZN(n12894) );
  INV_X1 U16205 ( .A(n12892), .ZN(n12893) );
  AND2_X1 U16206 ( .A1(n12894), .A2(n12893), .ZN(n19905) );
  AND2_X1 U16207 ( .A1(n19276), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n19287) );
  AOI21_X1 U16208 ( .B1(n12895), .B2(n15918), .A(n19287), .ZN(n12898) );
  NAND2_X1 U16209 ( .A1(n12896), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12897) );
  OAI211_X1 U16210 ( .C1(n19905), .C2(n16479), .A(n12898), .B(n12897), .ZN(
        n12911) );
  NAND2_X1 U16211 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n15918), .ZN(
        n12908) );
  OAI21_X1 U16212 ( .B1(n9794), .B2(n12900), .A(n12899), .ZN(n12901) );
  INV_X1 U16213 ( .A(n12901), .ZN(n19289) );
  INV_X1 U16214 ( .A(n12902), .ZN(n12903) );
  AOI21_X1 U16215 ( .B1(n12904), .B2(n15370), .A(n12903), .ZN(n12906) );
  XNOR2_X1 U16216 ( .A(n12906), .B(n12905), .ZN(n19286) );
  AOI22_X1 U16217 ( .A1(n16460), .A2(n19289), .B1(n16485), .B2(n19286), .ZN(
        n12907) );
  OAI221_X1 U16218 ( .B1(n15793), .B2(n12909), .C1(n15793), .C2(n12908), .A(
        n12907), .ZN(n12910) );
  AOI211_X1 U16219 ( .C1(n16494), .C2(n19295), .A(n12911), .B(n12910), .ZN(
        n12912) );
  INV_X1 U16220 ( .A(n12912), .ZN(P2_U3044) );
  INV_X1 U16221 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n20868) );
  OAI21_X1 U16222 ( .B1(n12859), .B2(n13052), .A(n12868), .ZN(n12914) );
  OR2_X1 U16223 ( .A1(n16055), .A2(n13055), .ZN(n12913) );
  AND2_X1 U16224 ( .A1(n12914), .A2(n12913), .ZN(n19963) );
  INV_X1 U16225 ( .A(n12915), .ZN(n12917) );
  INV_X1 U16226 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n12916) );
  NAND2_X1 U16227 ( .A1(n12917), .A2(n12916), .ZN(n16072) );
  INV_X1 U16228 ( .A(n16072), .ZN(n13072) );
  OR2_X1 U16229 ( .A1(n12918), .A2(n13072), .ZN(n12919) );
  NAND2_X1 U16230 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20819) );
  NAND2_X1 U16231 ( .A1(n12919), .A2(n20819), .ZN(n20810) );
  AND2_X1 U16232 ( .A1(n19963), .A2(n20810), .ZN(n16039) );
  NOR2_X1 U16233 ( .A1(n16039), .A2(n19964), .ZN(n19972) );
  NAND2_X1 U16234 ( .A1(n10422), .A2(n13579), .ZN(n12920) );
  NAND2_X1 U16235 ( .A1(n13144), .A2(n12920), .ZN(n13156) );
  INV_X1 U16236 ( .A(n13156), .ZN(n12921) );
  MUX2_X1 U16237 ( .A(n13190), .B(n12921), .S(n13201), .Z(n12923) );
  INV_X1 U16238 ( .A(n13052), .ZN(n13147) );
  OAI22_X1 U16239 ( .A1(n12859), .A2(n13147), .B1(n12868), .B2(n16055), .ZN(
        n12922) );
  NOR2_X1 U16240 ( .A1(n12923), .A2(n12922), .ZN(n16041) );
  INV_X1 U16241 ( .A(n16041), .ZN(n12924) );
  NAND2_X1 U16242 ( .A1(n12924), .A2(n19972), .ZN(n12925) );
  OAI21_X1 U16243 ( .B1(n20868), .B2(n19972), .A(n12925), .ZN(P1_U3484) );
  INV_X1 U16244 ( .A(n12829), .ZN(n12927) );
  NAND2_X1 U16245 ( .A1(n12927), .A2(n12926), .ZN(n12928) );
  NAND2_X1 U16246 ( .A1(n12929), .A2(n12928), .ZN(n12941) );
  INV_X1 U16247 ( .A(n12941), .ZN(n12940) );
  NAND2_X1 U16248 ( .A1(n12930), .A2(n12981), .ZN(n12935) );
  INV_X1 U16249 ( .A(n19894), .ZN(n19719) );
  NOR2_X1 U16250 ( .A1(n19912), .A2(n19922), .ZN(n19714) );
  INV_X1 U16251 ( .A(n12983), .ZN(n12932) );
  NAND2_X1 U16252 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19629) );
  NAND2_X1 U16253 ( .A1(n19629), .A2(n19912), .ZN(n12931) );
  NAND2_X1 U16254 ( .A1(n12932), .A2(n12931), .ZN(n13670) );
  NOR2_X1 U16255 ( .A1(n19719), .A2(n13670), .ZN(n12933) );
  AOI21_X1 U16256 ( .B1(n12986), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12933), .ZN(n12934) );
  NAND2_X1 U16257 ( .A1(n12979), .A2(n12938), .ZN(n12942) );
  INV_X1 U16258 ( .A(n12942), .ZN(n12939) );
  NAND2_X1 U16259 ( .A1(n12940), .A2(n12939), .ZN(n12980) );
  NAND2_X1 U16260 ( .A1(n12942), .A2(n12941), .ZN(n12943) );
  MUX2_X1 U16261 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n19295), .S(n19164), .Z(
        n12944) );
  AOI21_X1 U16262 ( .B1(n19907), .B2(n19151), .A(n12944), .ZN(n12945) );
  INV_X1 U16263 ( .A(n12945), .ZN(P2_U2885) );
  NAND2_X1 U16264 ( .A1(n12947), .A2(n12946), .ZN(n12948) );
  NOR2_X1 U16265 ( .A1(n12949), .A2(n12948), .ZN(n12950) );
  AOI21_X1 U16266 ( .B1(n13330), .B2(n12951), .A(n12950), .ZN(n13281) );
  NAND2_X1 U16267 ( .A1(n13281), .A2(n12952), .ZN(n12953) );
  INV_X1 U16268 ( .A(n12957), .ZN(n19341) );
  NOR2_X1 U16269 ( .A1(n19341), .A2(n12955), .ZN(n12956) );
  NAND2_X1 U16270 ( .A1(n19205), .A2(n12956), .ZN(n13963) );
  INV_X1 U16271 ( .A(n13963), .ZN(n12959) );
  AND2_X1 U16272 ( .A1(n19325), .A2(n12957), .ZN(n12958) );
  NAND2_X1 U16273 ( .A1(n19205), .A2(n19341), .ZN(n19180) );
  INV_X1 U16274 ( .A(n12113), .ZN(n12965) );
  INV_X1 U16275 ( .A(n12960), .ZN(n12963) );
  INV_X1 U16276 ( .A(n12961), .ZN(n12962) );
  NAND2_X1 U16277 ( .A1(n12963), .A2(n12962), .ZN(n12964) );
  NAND2_X1 U16278 ( .A1(n12965), .A2(n12964), .ZN(n16492) );
  OAI22_X1 U16279 ( .A1(n19180), .A2(n16492), .B1(n19205), .B2(n12966), .ZN(
        n12968) );
  NAND2_X1 U16280 ( .A1(n19205), .A2(n12098), .ZN(n19236) );
  NOR2_X1 U16281 ( .A1(n19925), .A2(n16492), .ZN(n19235) );
  AOI211_X1 U16282 ( .C1(n19925), .C2(n16492), .A(n19236), .B(n19235), .ZN(
        n12967) );
  AOI211_X1 U16283 ( .C1(n19171), .C2(n19207), .A(n12968), .B(n12967), .ZN(
        n12969) );
  INV_X1 U16284 ( .A(n12969), .ZN(P2_U2919) );
  AOI22_X1 U16285 ( .A1(n19269), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19268), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12971) );
  OAI21_X1 U16286 ( .B1(n12337), .B2(n12978), .A(n12971), .ZN(P2_U2921) );
  INV_X1 U16287 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n12973) );
  AOI22_X1 U16288 ( .A1(n12976), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19268), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12972) );
  OAI21_X1 U16289 ( .B1(n12973), .B2(n12978), .A(n12972), .ZN(P2_U2933) );
  AOI22_X1 U16290 ( .A1(n12976), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19268), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n12974) );
  OAI21_X1 U16291 ( .B1(n12975), .B2(n12978), .A(n12974), .ZN(P2_U2935) );
  INV_X1 U16292 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n20858) );
  AOI22_X1 U16293 ( .A1(n12976), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19268), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n12977) );
  OAI21_X1 U16294 ( .B1(n20858), .B2(n12978), .A(n12977), .ZN(P2_U2934) );
  NAND2_X1 U16295 ( .A1(n12980), .A2(n12979), .ZN(n13017) );
  AND2_X1 U16296 ( .A1(n14258), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12988) );
  OAI21_X1 U16297 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12983), .A(
        n19894), .ZN(n12984) );
  NOR2_X1 U16298 ( .A1(n12984), .A2(n19810), .ZN(n12985) );
  AOI21_X1 U16299 ( .B1(n12986), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12985), .ZN(n12987) );
  NAND2_X1 U16300 ( .A1(n12991), .A2(n12988), .ZN(n15353) );
  OAI21_X1 U16301 ( .B1(n12988), .B2(n12991), .A(n15353), .ZN(n12989) );
  INV_X1 U16302 ( .A(n12989), .ZN(n13016) );
  NAND2_X1 U16303 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12991), .ZN(
        n13018) );
  NAND2_X1 U16304 ( .A1(n15350), .A2(n13018), .ZN(n13001) );
  AND2_X1 U16305 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12992) );
  NAND2_X1 U16306 ( .A1(n13001), .A2(n13015), .ZN(n13003) );
  XOR2_X1 U16307 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n13003), .Z(n12998)
         );
  AOI21_X1 U16308 ( .B1(n12995), .B2(n12993), .A(n12994), .ZN(n16484) );
  INV_X1 U16309 ( .A(n16484), .ZN(n19086) );
  MUX2_X1 U16310 ( .A(n12996), .B(n19086), .S(n19164), .Z(n12997) );
  OAI21_X1 U16311 ( .B1(n12998), .B2(n19165), .A(n12997), .ZN(P2_U2880) );
  OAI21_X1 U16312 ( .B1(n12999), .B2(n13000), .A(n12993), .ZN(n19101) );
  NAND2_X1 U16313 ( .A1(n13001), .A2(n15351), .ZN(n15356) );
  NOR2_X1 U16314 ( .A1(n15356), .A2(n13002), .ZN(n13004) );
  OAI211_X1 U16315 ( .C1(n13004), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n19151), .B(n13003), .ZN(n13006) );
  NAND2_X1 U16316 ( .A1(n19161), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13005) );
  OAI211_X1 U16317 ( .C1(n19101), .C2(n19161), .A(n13006), .B(n13005), .ZN(
        P2_U2881) );
  XOR2_X1 U16318 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n15356), .Z(n13010)
         );
  AND2_X1 U16319 ( .A1(n13523), .A2(n13007), .ZN(n13008) );
  OR2_X1 U16320 ( .A1(n12999), .A2(n13008), .ZN(n13699) );
  MUX2_X1 U16321 ( .A(n13699), .B(n19108), .S(n19161), .Z(n13009) );
  OAI21_X1 U16322 ( .B1(n13010), .B2(n19165), .A(n13009), .ZN(P2_U2882) );
  OR2_X1 U16323 ( .A1(n11167), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13012) );
  NAND2_X1 U16324 ( .A1(n13012), .A2(n13011), .ZN(n20114) );
  XNOR2_X1 U16325 ( .A(n13014), .B(n13013), .ZN(n13618) );
  OAI222_X1 U16326 ( .A1(n20114), .A2(n14636), .B1(n13613), .B2(n16118), .C1(
        n14638), .C2(n13618), .ZN(P1_U2872) );
  NAND3_X1 U16327 ( .A1(n13017), .A2(n13016), .A3(n13020), .ZN(n13022) );
  INV_X1 U16328 ( .A(n13018), .ZN(n13019) );
  NAND2_X1 U16329 ( .A1(n13022), .A2(n13021), .ZN(n19155) );
  NAND2_X1 U16330 ( .A1(n19155), .A2(n13023), .ZN(n13024) );
  INV_X1 U16331 ( .A(n13024), .ZN(n19156) );
  OAI211_X1 U16332 ( .C1(n19156), .C2(n13026), .A(n19151), .B(n13219), .ZN(
        n13030) );
  AOI21_X1 U16333 ( .B1(n13028), .B2(n15331), .A(n13027), .ZN(n19073) );
  NAND2_X1 U16334 ( .A1(n19164), .A2(n19073), .ZN(n13029) );
  OAI211_X1 U16335 ( .C1(n19164), .C2(n21042), .A(n13030), .B(n13029), .ZN(
        P2_U2878) );
  XNOR2_X1 U16336 ( .A(n19210), .B(n19905), .ZN(n13036) );
  XNOR2_X1 U16337 ( .A(n13032), .B(n13031), .ZN(n19920) );
  INV_X1 U16338 ( .A(n19920), .ZN(n15384) );
  NAND2_X1 U16339 ( .A1(n19915), .A2(n15384), .ZN(n13033) );
  OAI21_X1 U16340 ( .B1(n19915), .B2(n15384), .A(n13033), .ZN(n19234) );
  NOR2_X1 U16341 ( .A1(n19234), .A2(n19235), .ZN(n19233) );
  INV_X1 U16342 ( .A(n13033), .ZN(n13034) );
  NOR2_X1 U16343 ( .A1(n19233), .A2(n13034), .ZN(n13035) );
  NOR2_X1 U16344 ( .A1(n13035), .A2(n13036), .ZN(n19209) );
  AOI21_X1 U16345 ( .B1(n13036), .B2(n13035), .A(n19209), .ZN(n13040) );
  AOI22_X1 U16346 ( .A1(n19207), .A2(n16311), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19231), .ZN(n13039) );
  INV_X1 U16347 ( .A(n19905), .ZN(n13037) );
  NAND2_X1 U16348 ( .A1(n13037), .A2(n19232), .ZN(n13038) );
  OAI211_X1 U16349 ( .C1(n13040), .C2(n19236), .A(n13039), .B(n13038), .ZN(
        P2_U2917) );
  NAND2_X1 U16350 ( .A1(n14818), .A2(n13041), .ZN(n13042) );
  AOI22_X1 U16351 ( .A1(n13042), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n16171), .B2(P1_REIP_REG_0__SCAN_IN), .ZN(n13047) );
  OR2_X1 U16352 ( .A1(n13043), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13044) );
  AND2_X1 U16353 ( .A1(n13045), .A2(n13044), .ZN(n20118) );
  NAND2_X1 U16354 ( .A1(n20118), .A2(n11125), .ZN(n13046) );
  OAI211_X1 U16355 ( .C1(n13618), .C2(n20129), .A(n13047), .B(n13046), .ZN(
        P1_U2999) );
  INV_X1 U16356 ( .A(n16425), .ZN(n13360) );
  NOR2_X1 U16357 ( .A1(n13360), .A2(n19161), .ZN(n13050) );
  AOI21_X1 U16358 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n19161), .A(n13050), .ZN(
        n13051) );
  OAI21_X1 U16359 ( .B1(n19567), .B2(n19165), .A(n13051), .ZN(P2_U2884) );
  INV_X1 U16360 ( .A(n20819), .ZN(n20724) );
  NOR2_X1 U16361 ( .A1(n13052), .A2(n20724), .ZN(n13053) );
  NAND2_X1 U16362 ( .A1(n16256), .A2(n13053), .ZN(n13206) );
  NAND2_X1 U16363 ( .A1(n13054), .A2(n13055), .ZN(n13059) );
  NAND2_X1 U16364 ( .A1(n13144), .A2(n13055), .ZN(n13200) );
  NAND2_X1 U16365 ( .A1(n13587), .A2(n20819), .ZN(n13056) );
  OR2_X1 U16366 ( .A1(n11145), .A2(n13056), .ZN(n13057) );
  NAND2_X1 U16367 ( .A1(n13200), .A2(n13057), .ZN(n13058) );
  NAND2_X1 U16368 ( .A1(n13058), .A2(n16055), .ZN(n13203) );
  NAND3_X1 U16369 ( .A1(n13206), .A2(n13059), .A3(n13203), .ZN(n13060) );
  NOR2_X1 U16370 ( .A1(n13061), .A2(n13062), .ZN(n13065) );
  OAI21_X1 U16371 ( .B1(n13064), .B2(n13063), .A(n13132), .ZN(n13603) );
  INV_X2 U16372 ( .A(n14679), .ZN(n14661) );
  INV_X1 U16373 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n13100) );
  INV_X1 U16374 ( .A(n20130), .ZN(n20128) );
  NAND2_X1 U16375 ( .A1(n20128), .A2(DATAI_1_), .ZN(n13067) );
  NAND2_X1 U16376 ( .A1(n20130), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13066) );
  AND2_X1 U16377 ( .A1(n13067), .A2(n13066), .ZN(n20151) );
  OAI222_X1 U16378 ( .A1(n14712), .A2(n13603), .B1(n14661), .B2(n13100), .C1(
        n14711), .C2(n20151), .ZN(P1_U2903) );
  INV_X1 U16379 ( .A(n13603), .ZN(n13497) );
  XNOR2_X1 U16380 ( .A(n13590), .B(n14358), .ZN(n13172) );
  OAI22_X1 U16381 ( .A1(n14636), .A2(n13172), .B1(n13068), .B2(n16118), .ZN(
        n13069) );
  AOI21_X1 U16382 ( .B1(n13497), .B2(n16116), .A(n13069), .ZN(n13070) );
  INV_X1 U16383 ( .A(n13070), .ZN(P1_U2871) );
  INV_X1 U16384 ( .A(P1_UWORD_REG_13__SCAN_IN), .ZN(n13077) );
  NOR2_X1 U16385 ( .A1(n20811), .A2(n20714), .ZN(n16263) );
  INV_X1 U16386 ( .A(n16263), .ZN(n13490) );
  NOR2_X1 U16387 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13490), .ZN(n20820) );
  INV_X1 U16388 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13076) );
  INV_X1 U16389 ( .A(n13073), .ZN(n13074) );
  INV_X1 U16390 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13075) );
  OAI222_X1 U16391 ( .A1(n13077), .A2(n13442), .B1(n13409), .B2(n13076), .C1(
        n13387), .C2(n13075), .ZN(P1_U2907) );
  INV_X1 U16392 ( .A(P1_UWORD_REG_14__SCAN_IN), .ZN(n13080) );
  INV_X1 U16393 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13079) );
  INV_X1 U16394 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13078) );
  OAI222_X1 U16395 ( .A1(n13080), .A2(n13442), .B1(n13409), .B2(n13079), .C1(
        n13387), .C2(n13078), .ZN(P1_U2906) );
  INV_X1 U16396 ( .A(P1_UWORD_REG_11__SCAN_IN), .ZN(n13083) );
  INV_X1 U16397 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13082) );
  INV_X1 U16398 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13081) );
  OAI222_X1 U16399 ( .A1(n13083), .A2(n13442), .B1(n13409), .B2(n13082), .C1(
        n13387), .C2(n13081), .ZN(P1_U2909) );
  INV_X1 U16400 ( .A(P1_UWORD_REG_10__SCAN_IN), .ZN(n13086) );
  INV_X1 U16401 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13085) );
  INV_X1 U16402 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13084) );
  OAI222_X1 U16403 ( .A1(n13086), .A2(n13442), .B1(n13409), .B2(n13085), .C1(
        n13387), .C2(n13084), .ZN(P1_U2910) );
  INV_X1 U16404 ( .A(P1_UWORD_REG_9__SCAN_IN), .ZN(n13089) );
  INV_X1 U16405 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13088) );
  INV_X1 U16406 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13087) );
  OAI222_X1 U16407 ( .A1(n13089), .A2(n13442), .B1(n13409), .B2(n13088), .C1(
        n13387), .C2(n13087), .ZN(P1_U2911) );
  INV_X1 U16408 ( .A(P1_UWORD_REG_8__SCAN_IN), .ZN(n13092) );
  INV_X1 U16409 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13091) );
  INV_X1 U16410 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13090) );
  OAI222_X1 U16411 ( .A1(n13092), .A2(n13442), .B1(n13409), .B2(n13091), .C1(
        n13387), .C2(n13090), .ZN(P1_U2912) );
  INV_X1 U16412 ( .A(P1_UWORD_REG_12__SCAN_IN), .ZN(n13095) );
  INV_X1 U16413 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13094) );
  INV_X1 U16414 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13093) );
  OAI222_X1 U16415 ( .A1(n13095), .A2(n13442), .B1(n13409), .B2(n13094), .C1(
        n13387), .C2(n13093), .ZN(P1_U2908) );
  INV_X1 U16416 ( .A(P1_LWORD_REG_6__SCAN_IN), .ZN(n13098) );
  INV_X1 U16417 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n13097) );
  OAI222_X1 U16418 ( .A1(n13098), .A2(n13442), .B1(n10644), .B2(n13445), .C1(
        n13097), .C2(n13387), .ZN(P1_U2930) );
  INV_X1 U16419 ( .A(P1_LWORD_REG_1__SCAN_IN), .ZN(n13101) );
  INV_X1 U16420 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n13099) );
  OAI222_X1 U16421 ( .A1(n13101), .A2(n13442), .B1(n13100), .B2(n13445), .C1(
        n13099), .C2(n13387), .ZN(P1_U2935) );
  INV_X1 U16422 ( .A(P1_LWORD_REG_4__SCAN_IN), .ZN(n13103) );
  INV_X1 U16423 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n13455) );
  INV_X1 U16424 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n13102) );
  OAI222_X1 U16425 ( .A1(n13103), .A2(n13442), .B1(n13455), .B2(n13445), .C1(
        n13102), .C2(n13387), .ZN(P1_U2932) );
  INV_X1 U16426 ( .A(P1_LWORD_REG_5__SCAN_IN), .ZN(n13105) );
  INV_X1 U16427 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13447) );
  INV_X1 U16428 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n13104) );
  OAI222_X1 U16429 ( .A1(n13105), .A2(n13442), .B1(n13447), .B2(n13445), .C1(
        n13104), .C2(n13387), .ZN(P1_U2931) );
  INV_X1 U16430 ( .A(P1_LWORD_REG_2__SCAN_IN), .ZN(n13107) );
  INV_X1 U16431 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n13139) );
  INV_X1 U16432 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n13106) );
  OAI222_X1 U16433 ( .A1(n13107), .A2(n13442), .B1(n13139), .B2(n13445), .C1(
        n13106), .C2(n13387), .ZN(P1_U2934) );
  INV_X1 U16434 ( .A(P1_LWORD_REG_3__SCAN_IN), .ZN(n13109) );
  INV_X1 U16435 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n13263) );
  INV_X1 U16436 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n13108) );
  OAI222_X1 U16437 ( .A1(n13109), .A2(n13442), .B1(n13263), .B2(n13445), .C1(
        n13108), .C2(n13387), .ZN(P1_U2933) );
  AND2_X1 U16438 ( .A1(n13166), .A2(n20724), .ZN(n13110) );
  NOR2_X2 U16439 ( .A1(n13252), .A2(n13165), .ZN(n20071) );
  INV_X1 U16440 ( .A(DATAI_11_), .ZN(n13112) );
  NAND2_X1 U16441 ( .A1(n20130), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13111) );
  OAI21_X1 U16442 ( .B1(n20130), .B2(n13112), .A(n13111), .ZN(n14649) );
  NAND2_X1 U16443 ( .A1(n20071), .A2(n14649), .ZN(n13231) );
  AOI22_X1 U16444 ( .A1(n20083), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n13252), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n13113) );
  NAND2_X1 U16445 ( .A1(n13231), .A2(n13113), .ZN(P1_U2963) );
  INV_X1 U16446 ( .A(DATAI_4_), .ZN(n13115) );
  NAND2_X1 U16447 ( .A1(n20130), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13114) );
  OAI21_X1 U16448 ( .B1(n20130), .B2(n13115), .A(n13114), .ZN(n14680) );
  NAND2_X1 U16449 ( .A1(n20071), .A2(n14680), .ZN(n13241) );
  AOI22_X1 U16450 ( .A1(n20083), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n13252), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13116) );
  NAND2_X1 U16451 ( .A1(n13241), .A2(n13116), .ZN(P1_U2956) );
  NAND2_X1 U16452 ( .A1(n20128), .A2(DATAI_5_), .ZN(n13118) );
  NAND2_X1 U16453 ( .A1(n20130), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13117) );
  AND2_X1 U16454 ( .A1(n13118), .A2(n13117), .ZN(n20165) );
  INV_X1 U16455 ( .A(n20165), .ZN(n13119) );
  NAND2_X1 U16456 ( .A1(n20071), .A2(n13119), .ZN(n13235) );
  AOI22_X1 U16457 ( .A1(n20083), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n13252), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13120) );
  NAND2_X1 U16458 ( .A1(n13235), .A2(n13120), .ZN(P1_U2957) );
  NAND2_X1 U16459 ( .A1(n20128), .A2(DATAI_7_), .ZN(n13122) );
  NAND2_X1 U16460 ( .A1(n20130), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13121) );
  AND2_X1 U16461 ( .A1(n13122), .A2(n13121), .ZN(n20174) );
  INV_X1 U16462 ( .A(n20174), .ZN(n13123) );
  NAND2_X1 U16463 ( .A1(n20071), .A2(n13123), .ZN(n13239) );
  AOI22_X1 U16464 ( .A1(n20083), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n13252), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13124) );
  NAND2_X1 U16465 ( .A1(n13239), .A2(n13124), .ZN(P1_U2959) );
  NAND2_X1 U16466 ( .A1(n20128), .A2(DATAI_3_), .ZN(n13126) );
  NAND2_X1 U16467 ( .A1(n20130), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13125) );
  AND2_X1 U16468 ( .A1(n13126), .A2(n13125), .ZN(n20158) );
  INV_X1 U16469 ( .A(n20158), .ZN(n13127) );
  NAND2_X1 U16470 ( .A1(n20071), .A2(n13127), .ZN(n13243) );
  AOI22_X1 U16471 ( .A1(n20083), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n13252), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13128) );
  NAND2_X1 U16472 ( .A1(n13243), .A2(n13128), .ZN(P1_U2955) );
  INV_X1 U16473 ( .A(DATAI_6_), .ZN(n13130) );
  NAND2_X1 U16474 ( .A1(n20130), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13129) );
  OAI21_X1 U16475 ( .B1(n20130), .B2(n13130), .A(n13129), .ZN(n14669) );
  NAND2_X1 U16476 ( .A1(n20071), .A2(n14669), .ZN(n13237) );
  AOI22_X1 U16477 ( .A1(n20083), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n13252), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13131) );
  NAND2_X1 U16478 ( .A1(n13237), .A2(n13131), .ZN(P1_U2958) );
  OAI21_X1 U16479 ( .B1(n9822), .B2(n10555), .A(n13133), .ZN(n14594) );
  INV_X1 U16480 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n20831) );
  NOR2_X1 U16481 ( .A1(n13135), .A2(n13134), .ZN(n13136) );
  OR2_X1 U16482 ( .A1(n13260), .A2(n13136), .ZN(n20106) );
  OAI222_X1 U16483 ( .A1(n14594), .A2(n14638), .B1(n16118), .B2(n20831), .C1(
        n20106), .C2(n14636), .ZN(P1_U2870) );
  NAND2_X1 U16484 ( .A1(n20128), .A2(DATAI_2_), .ZN(n13138) );
  NAND2_X1 U16485 ( .A1(n20130), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13137) );
  AND2_X1 U16486 ( .A1(n13138), .A2(n13137), .ZN(n20154) );
  OAI222_X1 U16487 ( .A1(n14712), .A2(n14594), .B1(n14661), .B2(n13139), .C1(
        n14711), .C2(n20154), .ZN(P1_U2902) );
  XNOR2_X1 U16488 ( .A(n13140), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13499) );
  AND2_X1 U16489 ( .A1(n13141), .A2(n20135), .ZN(n13142) );
  NAND2_X1 U16490 ( .A1(n13143), .A2(n13142), .ZN(n13184) );
  NAND2_X1 U16491 ( .A1(n13144), .A2(n13184), .ZN(n13145) );
  NAND2_X1 U16492 ( .A1(n12859), .A2(n13145), .ZN(n13199) );
  NAND2_X1 U16493 ( .A1(n13147), .A2(n13146), .ZN(n13151) );
  NAND2_X1 U16494 ( .A1(n13165), .A2(n16072), .ZN(n13585) );
  NAND2_X1 U16495 ( .A1(n13585), .A2(n20819), .ZN(n13148) );
  OAI211_X1 U16496 ( .C1(n11145), .C2(n13148), .A(n20135), .B(n14049), .ZN(
        n13149) );
  NAND2_X1 U16497 ( .A1(n13149), .A2(n16055), .ZN(n13150) );
  MUX2_X1 U16498 ( .A(n13151), .B(n13150), .S(n10387), .Z(n13153) );
  OR3_X1 U16499 ( .A1(n10331), .A2(n13165), .A3(n16055), .ZN(n13152) );
  NAND3_X1 U16500 ( .A1(n13199), .A2(n13153), .A3(n13152), .ZN(n13154) );
  OAI211_X1 U16501 ( .C1(n10421), .C2(n13167), .A(n13155), .B(n13156), .ZN(
        n13157) );
  INV_X1 U16502 ( .A(n13158), .ZN(n13163) );
  OAI21_X1 U16503 ( .B1(n13160), .B2(n20135), .A(n13159), .ZN(n13161) );
  INV_X1 U16504 ( .A(n13161), .ZN(n13162) );
  NAND4_X1 U16505 ( .A1(n13163), .A2(n13162), .A3(n13185), .A4(n13184), .ZN(
        n13164) );
  NOR2_X1 U16506 ( .A1(n16207), .A2(n15035), .ZN(n20119) );
  NOR2_X1 U16507 ( .A1(n12859), .A2(n13165), .ZN(n16019) );
  NAND2_X1 U16508 ( .A1(n13169), .A2(n16019), .ZN(n15051) );
  AND2_X1 U16509 ( .A1(n20119), .A2(n15051), .ZN(n15043) );
  NOR2_X1 U16510 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20122), .ZN(
        n13549) );
  NOR2_X1 U16511 ( .A1(n15043), .A2(n13549), .ZN(n13174) );
  OR2_X1 U16512 ( .A1(n11145), .A2(n13166), .ZN(n16048) );
  OAI21_X1 U16513 ( .B1(n13167), .B2(n20161), .A(n16048), .ZN(n13168) );
  INV_X1 U16514 ( .A(n13169), .ZN(n13170) );
  NAND2_X1 U16515 ( .A1(n13170), .A2(n16200), .ZN(n15037) );
  OAI21_X1 U16516 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n20119), .A(
        n15037), .ZN(n20121) );
  AOI22_X1 U16517 ( .A1(n16171), .A2(P1_REIP_REG_1__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20121), .ZN(n13171) );
  OAI21_X1 U16518 ( .B1(n20107), .B2(n13172), .A(n13171), .ZN(n13173) );
  AOI21_X1 U16519 ( .B1(n13174), .B2(n11153), .A(n13173), .ZN(n13175) );
  OAI21_X1 U16520 ( .B1(n13499), .B2(n20091), .A(n13175), .ZN(P1_U3030) );
  INV_X1 U16521 ( .A(n20083), .ZN(n13228) );
  INV_X1 U16522 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13180) );
  INV_X1 U16523 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13443) );
  INV_X1 U16524 ( .A(n20071), .ZN(n13178) );
  INV_X1 U16525 ( .A(DATAI_15_), .ZN(n13177) );
  INV_X1 U16526 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13176) );
  MUX2_X1 U16527 ( .A(n13177), .B(n13176), .S(n20130), .Z(n14706) );
  OAI222_X1 U16528 ( .A1(n13228), .A2(n13180), .B1(n13443), .B2(n13179), .C1(
        n13178), .C2(n14706), .ZN(P1_U2967) );
  INV_X1 U16529 ( .A(n13183), .ZN(n13186) );
  NAND3_X1 U16530 ( .A1(n13186), .A2(n13185), .A3(n13184), .ZN(n13187) );
  NOR2_X1 U16531 ( .A1(n13187), .A2(n16256), .ZN(n15073) );
  XNOR2_X1 U16532 ( .A(n13188), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13196) );
  NOR2_X1 U16533 ( .A1(n10429), .A2(n13196), .ZN(n13191) );
  INV_X1 U16534 ( .A(n13200), .ZN(n13189) );
  OR2_X1 U16535 ( .A1(n13190), .A2(n13189), .ZN(n13459) );
  AOI22_X1 U16536 ( .A1(n15073), .A2(n13191), .B1(n13459), .B2(n13196), .ZN(
        n13194) );
  NAND2_X1 U16537 ( .A1(n16019), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13192) );
  NAND2_X1 U16538 ( .A1(n16019), .A2(n10455), .ZN(n15078) );
  MUX2_X1 U16539 ( .A(n13192), .B(n15078), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13193) );
  OAI211_X1 U16540 ( .C1(n13182), .C2(n15073), .A(n13194), .B(n13193), .ZN(
        n13470) );
  INV_X1 U16541 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20100) );
  NOR2_X1 U16542 ( .A1(n20714), .A2(n20100), .ZN(n15083) );
  INV_X1 U16543 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13195) );
  AOI22_X1 U16544 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n11153), .B2(n13195), .ZN(
        n15081) );
  INV_X1 U16545 ( .A(n13196), .ZN(n13197) );
  AOI222_X1 U16546 ( .A1(n13470), .A2(n16255), .B1(n15083), .B2(n15081), .C1(
        n13482), .C2(n13197), .ZN(n13211) );
  INV_X1 U16547 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20547) );
  OR2_X1 U16548 ( .A1(n13583), .A2(n10423), .ZN(n13198) );
  AND2_X1 U16549 ( .A1(n13199), .A2(n13198), .ZN(n13208) );
  NAND2_X1 U16550 ( .A1(n13200), .A2(n11145), .ZN(n13205) );
  NOR3_X1 U16551 ( .A1(n13201), .A2(n20724), .A3(n16072), .ZN(n16044) );
  INV_X1 U16552 ( .A(n16044), .ZN(n13202) );
  NAND2_X1 U16553 ( .A1(n13203), .A2(n13202), .ZN(n13204) );
  OAI21_X1 U16554 ( .B1(n16019), .B2(n13205), .A(n13204), .ZN(n13207) );
  NAND4_X1 U16555 ( .A1(n13209), .A2(n13208), .A3(n13207), .A4(n13206), .ZN(
        n13475) );
  NAND2_X1 U16556 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16263), .ZN(n16267) );
  INV_X1 U16557 ( .A(n16267), .ZN(n13481) );
  AOI22_X1 U16558 ( .A1(n13210), .A2(n13475), .B1(P1_FLUSH_REG_SCAN_IN), .B2(
        n13481), .ZN(n16259) );
  OAI21_X1 U16559 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n20547), .A(n16259), 
        .ZN(n16257) );
  MUX2_X1 U16560 ( .A(n10094), .B(n13211), .S(n16257), .Z(n13212) );
  INV_X1 U16561 ( .A(n13212), .ZN(P1_U3472) );
  INV_X1 U16562 ( .A(n16255), .ZN(n15090) );
  INV_X1 U16563 ( .A(n16019), .ZN(n13462) );
  OAI21_X1 U16564 ( .B1(n15090), .B2(n13462), .A(n16257), .ZN(n13216) );
  INV_X1 U16565 ( .A(n15073), .ZN(n13465) );
  NOR2_X1 U16566 ( .A1(n10331), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13213) );
  AOI21_X1 U16567 ( .B1(n10552), .B2(n13465), .A(n13213), .ZN(n16021) );
  AOI22_X1 U16568 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20100), .B1(n10173), 
        .B2(n13482), .ZN(n13214) );
  OAI21_X1 U16569 ( .B1(n16021), .B2(n15090), .A(n13214), .ZN(n13215) );
  AOI22_X1 U16570 ( .A1(n13216), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n16257), .B2(n13215), .ZN(n13217) );
  INV_X1 U16571 ( .A(n13217), .ZN(P1_U3474) );
  OAI21_X1 U16572 ( .B1(n13219), .B2(n13221), .A(n13220), .ZN(n13222) );
  NAND3_X1 U16573 ( .A1(n10149), .A2(n19151), .A3(n13222), .ZN(n13226) );
  NOR2_X1 U16574 ( .A1(n16379), .A2(n13223), .ZN(n13224) );
  OR2_X1 U16575 ( .A1(n15865), .A2(n13224), .ZN(n15321) );
  INV_X1 U16576 ( .A(n15321), .ZN(n16367) );
  NAND2_X1 U16577 ( .A1(n19164), .A2(n16367), .ZN(n13225) );
  OAI211_X1 U16578 ( .C1(n19164), .C2(n11781), .A(n13226), .B(n13225), .ZN(
        P2_U2876) );
  INV_X1 U16579 ( .A(n20154), .ZN(n13227) );
  NAND2_X1 U16580 ( .A1(n20071), .A2(n13227), .ZN(n13255) );
  AOI22_X1 U16581 ( .A1(n13253), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n13252), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13229) );
  NAND2_X1 U16582 ( .A1(n13255), .A2(n13229), .ZN(P1_U2954) );
  AOI22_X1 U16583 ( .A1(n13253), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n13252), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13230) );
  NAND2_X1 U16584 ( .A1(n13231), .A2(n13230), .ZN(P1_U2948) );
  INV_X1 U16585 ( .A(n20151), .ZN(n13232) );
  NAND2_X1 U16586 ( .A1(n20071), .A2(n13232), .ZN(n13249) );
  AOI22_X1 U16587 ( .A1(n13253), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n13252), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13233) );
  NAND2_X1 U16588 ( .A1(n13249), .A2(n13233), .ZN(P1_U2938) );
  AOI22_X1 U16589 ( .A1(n13253), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n13252), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13234) );
  NAND2_X1 U16590 ( .A1(n13235), .A2(n13234), .ZN(P1_U2942) );
  AOI22_X1 U16591 ( .A1(n13253), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n13252), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13236) );
  NAND2_X1 U16592 ( .A1(n13237), .A2(n13236), .ZN(P1_U2943) );
  AOI22_X1 U16593 ( .A1(n13253), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n13252), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13238) );
  NAND2_X1 U16594 ( .A1(n13239), .A2(n13238), .ZN(P1_U2944) );
  AOI22_X1 U16595 ( .A1(n13253), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n13252), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13240) );
  NAND2_X1 U16596 ( .A1(n13241), .A2(n13240), .ZN(P1_U2941) );
  AOI22_X1 U16597 ( .A1(n13253), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n13252), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13242) );
  NAND2_X1 U16598 ( .A1(n13243), .A2(n13242), .ZN(P1_U2940) );
  NAND2_X1 U16599 ( .A1(n20128), .A2(DATAI_0_), .ZN(n13245) );
  NAND2_X1 U16600 ( .A1(n20130), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13244) );
  AND2_X1 U16601 ( .A1(n13245), .A2(n13244), .ZN(n20142) );
  INV_X1 U16602 ( .A(n20142), .ZN(n13246) );
  NAND2_X1 U16603 ( .A1(n20071), .A2(n13246), .ZN(n13251) );
  AOI22_X1 U16604 ( .A1(n13253), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n13252), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13247) );
  NAND2_X1 U16605 ( .A1(n13251), .A2(n13247), .ZN(P1_U2952) );
  AOI22_X1 U16606 ( .A1(n13253), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n13252), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13248) );
  NAND2_X1 U16607 ( .A1(n13249), .A2(n13248), .ZN(P1_U2953) );
  AOI22_X1 U16608 ( .A1(n13253), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n13252), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13250) );
  NAND2_X1 U16609 ( .A1(n13251), .A2(n13250), .ZN(P1_U2937) );
  AOI22_X1 U16610 ( .A1(n13253), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n13252), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13254) );
  NAND2_X1 U16611 ( .A1(n13255), .A2(n13254), .ZN(P1_U2939) );
  OAI21_X1 U16612 ( .B1(n13256), .B2(n13258), .A(n13257), .ZN(n13502) );
  INV_X1 U16613 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13262) );
  OR2_X1 U16614 ( .A1(n13260), .A2(n13259), .ZN(n13261) );
  AND2_X1 U16615 ( .A1(n13451), .A2(n13261), .ZN(n20088) );
  INV_X1 U16616 ( .A(n20088), .ZN(n14577) );
  OAI222_X1 U16617 ( .A1(n13502), .A2(n14638), .B1(n13262), .B2(n16118), .C1(
        n14577), .C2(n14636), .ZN(P1_U2869) );
  OAI222_X1 U16618 ( .A1(n14712), .A2(n13502), .B1(n14661), .B2(n13263), .C1(
        n14711), .C2(n20158), .ZN(P1_U2901) );
  INV_X1 U16619 ( .A(n13264), .ZN(n13301) );
  NAND2_X1 U16620 ( .A1(n13265), .A2(n11416), .ZN(n13288) );
  OAI21_X1 U16621 ( .B1(n14325), .B2(n20841), .A(n14101), .ZN(n13267) );
  NAND2_X1 U16622 ( .A1(n13288), .A2(n13267), .ZN(n13276) );
  NAND2_X1 U16623 ( .A1(n13268), .A2(n13329), .ZN(n13292) );
  INV_X1 U16624 ( .A(n11512), .ZN(n13269) );
  NAND2_X1 U16625 ( .A1(n13269), .A2(n13290), .ZN(n13289) );
  XNOR2_X1 U16626 ( .A(n13289), .B(n20841), .ZN(n13270) );
  NAND2_X1 U16627 ( .A1(n13292), .A2(n13270), .ZN(n13275) );
  AOI21_X1 U16628 ( .B1(n21077), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13271) );
  NOR2_X1 U16629 ( .A1(n13272), .A2(n13271), .ZN(n13273) );
  NAND2_X1 U16630 ( .A1(n15928), .A2(n13273), .ZN(n13274) );
  NAND3_X1 U16631 ( .A1(n13276), .A2(n13275), .A3(n13274), .ZN(n13277) );
  AOI21_X1 U16632 ( .B1(n16425), .B2(n13301), .A(n13277), .ZN(n15947) );
  INV_X1 U16633 ( .A(n13278), .ZN(n13279) );
  AND3_X1 U16634 ( .A1(n13281), .A2(n13280), .A3(n13279), .ZN(n13285) );
  INV_X1 U16635 ( .A(n13282), .ZN(n13283) );
  NAND3_X1 U16636 ( .A1(n13283), .A2(n13332), .A3(n13346), .ZN(n13284) );
  INV_X1 U16637 ( .A(n13319), .ZN(n15926) );
  NAND2_X1 U16638 ( .A1(n15947), .A2(n15926), .ZN(n13287) );
  NAND2_X1 U16639 ( .A1(n13319), .A2(n20841), .ZN(n13286) );
  NAND2_X1 U16640 ( .A1(n13287), .A2(n13286), .ZN(n13318) );
  INV_X1 U16641 ( .A(n13288), .ZN(n13296) );
  NAND2_X1 U16642 ( .A1(n13266), .A2(n13289), .ZN(n13295) );
  NAND2_X1 U16643 ( .A1(n19295), .A2(n13301), .ZN(n13294) );
  XNOR2_X1 U16644 ( .A(n13290), .B(n21077), .ZN(n13291) );
  AOI22_X1 U16645 ( .A1(n13292), .A2(n13295), .B1(n13291), .B2(n15928), .ZN(
        n13293) );
  OAI211_X1 U16646 ( .C1(n13296), .C2(n13295), .A(n13294), .B(n13293), .ZN(
        n15942) );
  MUX2_X1 U16647 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n15942), .S(
        n15926), .Z(n13341) );
  INV_X1 U16648 ( .A(n12342), .ZN(n13298) );
  NAND2_X1 U16649 ( .A1(n13298), .A2(n13297), .ZN(n13305) );
  AND2_X1 U16650 ( .A1(n13305), .A2(n11515), .ZN(n13299) );
  AOI21_X1 U16651 ( .B1(n12816), .B2(n13301), .A(n13299), .ZN(n15924) );
  AOI21_X1 U16652 ( .B1(n15928), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n19931), .ZN(n13300) );
  AND2_X1 U16653 ( .A1(n15924), .A2(n13300), .ZN(n13308) );
  NOR2_X1 U16654 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n13308), .ZN(
        n13310) );
  NAND2_X1 U16655 ( .A1(n15917), .A2(n13301), .ZN(n13307) );
  INV_X1 U16656 ( .A(n11511), .ZN(n13303) );
  INV_X1 U16657 ( .A(n11509), .ZN(n13302) );
  NAND2_X1 U16658 ( .A1(n13303), .A2(n13302), .ZN(n13304) );
  AOI22_X1 U16659 ( .A1(n13305), .A2(n13304), .B1(n11256), .B2(n15928), .ZN(
        n13306) );
  NAND2_X1 U16660 ( .A1(n13307), .A2(n13306), .ZN(n15938) );
  INV_X1 U16661 ( .A(n13308), .ZN(n13309) );
  OAI22_X1 U16662 ( .A1(n13310), .A2(n15938), .B1(n19922), .B2(n13309), .ZN(
        n13311) );
  AOI211_X1 U16663 ( .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n15947), .A(
        n13319), .B(n13311), .ZN(n13313) );
  INV_X1 U16664 ( .A(n13313), .ZN(n13312) );
  AOI21_X1 U16665 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n13312), .A(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13314) );
  AOI22_X1 U16666 ( .A1(n13341), .A2(n13314), .B1(n13313), .B2(n19912), .ZN(
        n13315) );
  OAI21_X1 U16667 ( .B1(n13318), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n13315), .ZN(n13317) );
  INV_X1 U16668 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n13316) );
  NAND2_X1 U16669 ( .A1(n13317), .A2(n13316), .ZN(n13344) );
  INV_X1 U16670 ( .A(n13318), .ZN(n13342) );
  NAND2_X1 U16671 ( .A1(n13319), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13339) );
  INV_X1 U16672 ( .A(n13320), .ZN(n13323) );
  OAI22_X1 U16673 ( .A1(n13324), .A2(n13323), .B1(n13322), .B2(n13321), .ZN(
        n13325) );
  INV_X1 U16674 ( .A(n13325), .ZN(n13328) );
  NAND2_X1 U16675 ( .A1(n13330), .A2(n13326), .ZN(n13327) );
  OAI211_X1 U16676 ( .C1(n13330), .C2(n13329), .A(n13328), .B(n13327), .ZN(
        n19935) );
  OAI21_X1 U16677 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n13331), .ZN(n13336) );
  NAND3_X1 U16678 ( .A1(n13332), .A2(n14263), .A3(n15977), .ZN(n13333) );
  NAND4_X1 U16679 ( .A1(n13336), .A2(n13335), .A3(n13334), .A4(n13333), .ZN(
        n13337) );
  NOR2_X1 U16680 ( .A1(n19935), .A2(n13337), .ZN(n13338) );
  NAND2_X1 U16681 ( .A1(n13339), .A2(n13338), .ZN(n13340) );
  AOI21_X1 U16682 ( .B1(n13342), .B2(n13341), .A(n13340), .ZN(n13343) );
  NAND2_X1 U16683 ( .A1(n16517), .A2(n12874), .ZN(n13345) );
  NAND2_X1 U16684 ( .A1(n13345), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13351) );
  INV_X1 U16685 ( .A(n13346), .ZN(n13347) );
  NOR2_X1 U16686 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13347), .ZN(n13642) );
  OR2_X1 U16687 ( .A1(n13348), .A2(n19685), .ZN(n19955) );
  AOI21_X1 U16688 ( .B1(n13349), .B2(n13642), .A(n19955), .ZN(n13350) );
  OAI21_X1 U16689 ( .B1(n16509), .B2(n16510), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13354) );
  NOR2_X1 U16690 ( .A1(n16510), .A2(n13352), .ZN(n16506) );
  INV_X1 U16691 ( .A(n16506), .ZN(n13353) );
  NAND2_X1 U16692 ( .A1(n13354), .A2(n13353), .ZN(P2_U3593) );
  XNOR2_X1 U16693 ( .A(n13355), .B(n13363), .ZN(n13356) );
  XNOR2_X1 U16694 ( .A(n13357), .B(n13356), .ZN(n16422) );
  XNOR2_X1 U16695 ( .A(n13358), .B(n13359), .ZN(n19900) );
  INV_X1 U16696 ( .A(n19900), .ZN(n19224) );
  OAI22_X1 U16697 ( .A1(n13360), .A2(n16466), .B1(n11446), .B2(n9725), .ZN(
        n13365) );
  INV_X1 U16698 ( .A(n13361), .ZN(n13769) );
  INV_X1 U16699 ( .A(n16491), .ZN(n16431) );
  NAND2_X1 U16700 ( .A1(n13363), .A2(n16431), .ZN(n13525) );
  OAI22_X1 U16701 ( .A1(n13769), .A2(n13363), .B1(n13362), .B2(n13525), .ZN(
        n13364) );
  AOI211_X1 U16702 ( .C1(n16493), .C2(n19224), .A(n13365), .B(n13364), .ZN(
        n13370) );
  INV_X1 U16703 ( .A(n13366), .ZN(n16419) );
  NOR2_X1 U16704 ( .A1(n13368), .A2(n13367), .ZN(n16420) );
  OR3_X1 U16705 ( .A1(n16419), .A2(n16420), .A3(n16503), .ZN(n13369) );
  OAI211_X1 U16706 ( .C1(n16422), .C2(n16498), .A(n13370), .B(n13369), .ZN(
        P2_U3043) );
  INV_X1 U16707 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n13433) );
  OAI222_X1 U16708 ( .A1(n14711), .A2(n20142), .B1(n14712), .B2(n13618), .C1(
        n13433), .C2(n14661), .ZN(P1_U2904) );
  INV_X1 U16709 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n13381) );
  OAI211_X1 U16710 ( .C1(n13374), .C2(n13373), .A(n19151), .B(n13375), .ZN(
        n13380) );
  NAND2_X1 U16711 ( .A1(n13376), .A2(n15866), .ZN(n13378) );
  INV_X1 U16712 ( .A(n15826), .ZN(n13377) );
  NAND2_X1 U16713 ( .A1(n19164), .A2(n19045), .ZN(n13379) );
  OAI211_X1 U16714 ( .C1(n19164), .C2(n13381), .A(n13380), .B(n13379), .ZN(
        P2_U2874) );
  NAND2_X1 U16715 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15937), .ZN(n18955) );
  INV_X1 U16716 ( .A(n18955), .ZN(n13382) );
  AOI21_X1 U16717 ( .B1(n13382), .B2(n16075), .A(n15925), .ZN(n13386) );
  NOR2_X1 U16718 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n16510), .ZN(n13383) );
  OAI211_X1 U16719 ( .C1(n16509), .C2(n13383), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n19952), .ZN(n13385) );
  NOR4_X1 U16720 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n12874), .ZN(n13384) );
  OAI211_X1 U16721 ( .C1(n16509), .C2(n13386), .A(n13385), .B(n19090), .ZN(
        P2_U3177) );
  INV_X1 U16722 ( .A(P1_UWORD_REG_5__SCAN_IN), .ZN(n13389) );
  INV_X1 U16723 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n13388) );
  OAI222_X1 U16724 ( .A1(n13389), .A2(n13442), .B1(n13409), .B2(n14674), .C1(
        n13387), .C2(n13388), .ZN(P1_U2915) );
  INV_X1 U16725 ( .A(P1_UWORD_REG_7__SCAN_IN), .ZN(n13392) );
  INV_X1 U16726 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13391) );
  INV_X1 U16727 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n13390) );
  OAI222_X1 U16728 ( .A1(n13392), .A2(n13442), .B1(n13409), .B2(n13391), .C1(
        n13387), .C2(n13390), .ZN(P1_U2913) );
  INV_X1 U16729 ( .A(P1_UWORD_REG_3__SCAN_IN), .ZN(n13394) );
  INV_X1 U16730 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n13393) );
  OAI222_X1 U16731 ( .A1(n13394), .A2(n13442), .B1(n13409), .B2(n14687), .C1(
        n13387), .C2(n13393), .ZN(P1_U2917) );
  INV_X1 U16732 ( .A(P1_UWORD_REG_6__SCAN_IN), .ZN(n13397) );
  INV_X1 U16733 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13396) );
  INV_X1 U16734 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n13395) );
  OAI222_X1 U16735 ( .A1(n13397), .A2(n13442), .B1(n13409), .B2(n13396), .C1(
        n13387), .C2(n13395), .ZN(P1_U2914) );
  INV_X1 U16736 ( .A(P1_UWORD_REG_0__SCAN_IN), .ZN(n13400) );
  INV_X1 U16737 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13399) );
  INV_X1 U16738 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n13398) );
  OAI222_X1 U16739 ( .A1(n13400), .A2(n13442), .B1(n13409), .B2(n13399), .C1(
        n13387), .C2(n13398), .ZN(P1_U2920) );
  INV_X1 U16740 ( .A(P1_UWORD_REG_4__SCAN_IN), .ZN(n13403) );
  INV_X1 U16741 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13402) );
  INV_X1 U16742 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n13401) );
  OAI222_X1 U16743 ( .A1(n13403), .A2(n13442), .B1(n13409), .B2(n13402), .C1(
        n13387), .C2(n13401), .ZN(P1_U2916) );
  INV_X1 U16744 ( .A(P1_UWORD_REG_2__SCAN_IN), .ZN(n13406) );
  INV_X1 U16745 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13405) );
  INV_X1 U16746 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n13404) );
  OAI222_X1 U16747 ( .A1(n13406), .A2(n13442), .B1(n13409), .B2(n13405), .C1(
        n13387), .C2(n13404), .ZN(P1_U2918) );
  INV_X1 U16748 ( .A(P1_UWORD_REG_1__SCAN_IN), .ZN(n13410) );
  INV_X1 U16749 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13408) );
  INV_X1 U16750 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n13407) );
  OAI222_X1 U16751 ( .A1(n13410), .A2(n13442), .B1(n13409), .B2(n13408), .C1(
        n13387), .C2(n13407), .ZN(P1_U2919) );
  AND2_X1 U16752 ( .A1(n13411), .A2(n13412), .ZN(n13414) );
  OR2_X1 U16753 ( .A1(n13414), .A2(n9727), .ZN(n13538) );
  AOI21_X1 U16754 ( .B1(n13415), .B2(n13453), .A(n13511), .ZN(n20023) );
  INV_X1 U16755 ( .A(n20023), .ZN(n13416) );
  OAI222_X1 U16756 ( .A1(n13538), .A2(n14638), .B1(n13417), .B2(n16118), .C1(
        n14636), .C2(n13416), .ZN(P1_U2867) );
  INV_X1 U16757 ( .A(P1_LWORD_REG_12__SCAN_IN), .ZN(n13420) );
  INV_X1 U16758 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n13419) );
  INV_X1 U16759 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n13418) );
  OAI222_X1 U16760 ( .A1(n13420), .A2(n13442), .B1(n13445), .B2(n13419), .C1(
        n13418), .C2(n13387), .ZN(P1_U2924) );
  INV_X1 U16761 ( .A(P1_LWORD_REG_14__SCAN_IN), .ZN(n13423) );
  INV_X1 U16762 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n13422) );
  INV_X1 U16763 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n13421) );
  OAI222_X1 U16764 ( .A1(n13423), .A2(n13442), .B1(n13445), .B2(n13422), .C1(
        n13421), .C2(n13387), .ZN(P1_U2922) );
  INV_X1 U16765 ( .A(P1_LWORD_REG_8__SCAN_IN), .ZN(n13426) );
  INV_X1 U16766 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13425) );
  INV_X1 U16767 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n13424) );
  OAI222_X1 U16768 ( .A1(n13426), .A2(n13442), .B1(n13445), .B2(n13425), .C1(
        n13424), .C2(n13387), .ZN(P1_U2928) );
  INV_X1 U16769 ( .A(P1_LWORD_REG_7__SCAN_IN), .ZN(n13428) );
  INV_X1 U16770 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n13427) );
  OAI222_X1 U16771 ( .A1(n13428), .A2(n13442), .B1(n10656), .B2(n13445), .C1(
        n13427), .C2(n13387), .ZN(P1_U2929) );
  INV_X1 U16772 ( .A(P1_LWORD_REG_13__SCAN_IN), .ZN(n13431) );
  INV_X1 U16773 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n13430) );
  INV_X1 U16774 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n13429) );
  OAI222_X1 U16775 ( .A1(n13431), .A2(n13442), .B1(n13445), .B2(n13430), .C1(
        n13429), .C2(n13387), .ZN(P1_U2923) );
  INV_X1 U16776 ( .A(P1_LWORD_REG_0__SCAN_IN), .ZN(n13434) );
  INV_X1 U16777 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n13432) );
  OAI222_X1 U16778 ( .A1(n13434), .A2(n13442), .B1(n13433), .B2(n13445), .C1(
        n13432), .C2(n13387), .ZN(P1_U2936) );
  INV_X1 U16779 ( .A(P1_LWORD_REG_9__SCAN_IN), .ZN(n13437) );
  INV_X1 U16780 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n13436) );
  INV_X1 U16781 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n13435) );
  OAI222_X1 U16782 ( .A1(n13437), .A2(n13442), .B1(n13445), .B2(n13436), .C1(
        n13435), .C2(n13387), .ZN(P1_U2927) );
  INV_X1 U16783 ( .A(P1_LWORD_REG_10__SCAN_IN), .ZN(n13440) );
  INV_X1 U16784 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13439) );
  INV_X1 U16785 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n13438) );
  OAI222_X1 U16786 ( .A1(n13440), .A2(n13442), .B1(n13445), .B2(n13439), .C1(
        n13438), .C2(n13387), .ZN(P1_U2926) );
  INV_X1 U16787 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n13441) );
  OAI222_X1 U16788 ( .A1(n13443), .A2(n13442), .B1(n13180), .B2(n13445), .C1(
        n13441), .C2(n13387), .ZN(P1_U2921) );
  INV_X1 U16789 ( .A(P1_LWORD_REG_11__SCAN_IN), .ZN(n13446) );
  INV_X1 U16790 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n13982) );
  INV_X1 U16791 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n13444) );
  OAI222_X1 U16792 ( .A1(n13446), .A2(n13442), .B1(n13982), .B2(n13445), .C1(
        n13444), .C2(n13387), .ZN(P1_U2925) );
  OAI222_X1 U16793 ( .A1(n14712), .A2(n13538), .B1(n14661), .B2(n13447), .C1(
        n14711), .C2(n20165), .ZN(P1_U2899) );
  INV_X1 U16794 ( .A(n13411), .ZN(n13448) );
  AOI21_X1 U16795 ( .B1(n13449), .B2(n13257), .A(n13448), .ZN(n20049) );
  INV_X1 U16796 ( .A(n20049), .ZN(n13456) );
  INV_X1 U16797 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13454) );
  NAND2_X1 U16798 ( .A1(n13451), .A2(n13450), .ZN(n13452) );
  NAND2_X1 U16799 ( .A1(n13453), .A2(n13452), .ZN(n20052) );
  OAI222_X1 U16800 ( .A1(n13456), .A2(n14638), .B1(n13454), .B2(n16118), .C1(
        n14636), .C2(n20052), .ZN(P1_U2868) );
  INV_X1 U16801 ( .A(n14680), .ZN(n20162) );
  OAI222_X1 U16802 ( .A1(n14712), .A2(n13456), .B1(n14661), .B2(n13455), .C1(
        n14711), .C2(n20162), .ZN(P1_U2900) );
  INV_X1 U16803 ( .A(n20406), .ZN(n15071) );
  INV_X1 U16804 ( .A(n15078), .ZN(n13468) );
  AOI21_X1 U16805 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n13457), .A(
        n13458), .ZN(n13463) );
  MUX2_X1 U16806 ( .A(n13458), .B(n10575), .S(n13188), .Z(n13460) );
  OAI21_X1 U16807 ( .B1(n13457), .B2(n13460), .A(n13459), .ZN(n13461) );
  OAI21_X1 U16808 ( .B1(n13463), .B2(n13462), .A(n13461), .ZN(n13467) );
  AOI21_X1 U16809 ( .B1(n13188), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10575), .ZN(n13464) );
  NOR2_X1 U16810 ( .A1(n9723), .A2(n13464), .ZN(n15088) );
  NOR3_X1 U16811 ( .A1(n13465), .A2(n15088), .A3(n10429), .ZN(n13466) );
  AOI211_X1 U16812 ( .C1(n13468), .C2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13467), .B(n13466), .ZN(n13469) );
  OAI21_X1 U16813 ( .B1(n15071), .B2(n15073), .A(n13469), .ZN(n15087) );
  MUX2_X1 U16814 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15087), .S(
        n13475), .Z(n16033) );
  NOR2_X1 U16815 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20714), .ZN(n13480) );
  AOI22_X1 U16816 ( .A1(n20714), .A2(n16033), .B1(n13480), .B2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13472) );
  MUX2_X1 U16817 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13470), .S(
        n13475), .Z(n16028) );
  AOI22_X1 U16818 ( .A1(n16028), .A2(n20714), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n13480), .ZN(n13471) );
  INV_X1 U16819 ( .A(n13475), .ZN(n16022) );
  INV_X1 U16820 ( .A(n20285), .ZN(n20545) );
  OR2_X1 U16821 ( .A1(n13476), .A2(n20545), .ZN(n13477) );
  XNOR2_X1 U16822 ( .A(n13477), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20036) );
  AOI21_X1 U16823 ( .B1(n20036), .B2(n16256), .A(n16022), .ZN(n13478) );
  AOI211_X1 U16824 ( .C1(n10603), .C2(n16022), .A(P1_STATE2_REG_1__SCAN_IN), 
        .B(n13478), .ZN(n13479) );
  AOI21_X1 U16825 ( .B1(n13480), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13479), .ZN(n16035) );
  OAI21_X1 U16826 ( .B1(n16034), .B2(n13474), .A(n16035), .ZN(n13491) );
  OAI21_X1 U16827 ( .B1(n13491), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13481), .ZN(
        n13484) );
  NAND2_X1 U16828 ( .A1(n20811), .A2(n20714), .ZN(n20814) );
  NAND2_X1 U16829 ( .A1(n13484), .A2(n20291), .ZN(n20126) );
  AND2_X1 U16830 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20547), .ZN(n15070) );
  NOR2_X1 U16831 ( .A1(n13182), .A2(n15070), .ZN(n13488) );
  NAND2_X1 U16832 ( .A1(n20208), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20249) );
  AND2_X1 U16833 ( .A1(n20249), .A2(n20661), .ZN(n20658) );
  NOR2_X1 U16834 ( .A1(n20249), .A2(n20653), .ZN(n13486) );
  MUX2_X1 U16835 ( .A(n20658), .B(n13486), .S(n13485), .Z(n13487) );
  OAI21_X1 U16836 ( .B1(n13488), .B2(n13487), .A(n20126), .ZN(n13489) );
  OAI21_X1 U16837 ( .B1(n20126), .B2(n20459), .A(n13489), .ZN(P1_U3476) );
  OR2_X1 U16838 ( .A1(n13491), .A2(n13490), .ZN(n16050) );
  INV_X1 U16839 ( .A(n16050), .ZN(n13493) );
  INV_X1 U16840 ( .A(n10552), .ZN(n20246) );
  OAI22_X1 U16841 ( .A1(n20207), .A2(n20653), .B1(n20246), .B2(n15070), .ZN(
        n13492) );
  OAI21_X1 U16842 ( .B1(n13493), .B2(n13492), .A(n20126), .ZN(n13494) );
  OAI21_X1 U16843 ( .B1(n20126), .B2(n20573), .A(n13494), .ZN(P1_U3478) );
  AOI22_X1 U16844 ( .A1(n16135), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n16171), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13495) );
  OAI21_X1 U16845 ( .B1(n16127), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13495), .ZN(n13496) );
  AOI21_X1 U16846 ( .B1(n13497), .B2(n16152), .A(n13496), .ZN(n13498) );
  OAI21_X1 U16847 ( .B1(n13499), .B2(n19970), .A(n13498), .ZN(P1_U2998) );
  XNOR2_X1 U16848 ( .A(n13500), .B(n13501), .ZN(n20092) );
  INV_X1 U16849 ( .A(n13502), .ZN(n14582) );
  INV_X1 U16850 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20739) );
  NOR2_X1 U16851 ( .A1(n16200), .A2(n20739), .ZN(n20087) );
  AOI21_X1 U16852 ( .B1(n16135), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20087), .ZN(n13503) );
  OAI21_X1 U16853 ( .B1(n16127), .B2(n14572), .A(n13503), .ZN(n13504) );
  AOI21_X1 U16854 ( .B1(n14582), .B2(n16152), .A(n13504), .ZN(n13505) );
  OAI21_X1 U16855 ( .B1(n20092), .B2(n19970), .A(n13505), .ZN(P1_U2996) );
  INV_X1 U16856 ( .A(n13506), .ZN(n13509) );
  INV_X1 U16857 ( .A(n9727), .ZN(n13508) );
  INV_X1 U16858 ( .A(n13507), .ZN(n13608) );
  AOI21_X1 U16859 ( .B1(n13509), .B2(n13508), .A(n13608), .ZN(n20019) );
  INV_X1 U16860 ( .A(n20019), .ZN(n13542) );
  INV_X1 U16861 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n13513) );
  NOR2_X1 U16862 ( .A1(n13511), .A2(n13510), .ZN(n13512) );
  OR2_X1 U16863 ( .A1(n13610), .A2(n13512), .ZN(n20014) );
  OAI222_X1 U16864 ( .A1(n13542), .A2(n14638), .B1(n13513), .B2(n16118), .C1(
        n14636), .C2(n20014), .ZN(P1_U2866) );
  XOR2_X1 U16865 ( .A(n13515), .B(n13514), .Z(n19278) );
  INV_X1 U16866 ( .A(n19278), .ZN(n13535) );
  XNOR2_X1 U16867 ( .A(n13517), .B(n13516), .ZN(n13518) );
  XNOR2_X1 U16868 ( .A(n13519), .B(n13518), .ZN(n19280) );
  NAND2_X1 U16869 ( .A1(n13521), .A2(n13520), .ZN(n13522) );
  NAND2_X1 U16870 ( .A1(n13523), .A2(n13522), .ZN(n19277) );
  NAND3_X1 U16871 ( .A1(n16431), .A2(n13524), .A3(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13526) );
  INV_X1 U16872 ( .A(n13526), .ZN(n13695) );
  OAI211_X1 U16873 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n13526), .A(
        n13769), .B(n13525), .ZN(n13697) );
  OAI21_X1 U16874 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13695), .A(
        n13697), .ZN(n13532) );
  NAND2_X1 U16875 ( .A1(n13528), .A2(n13527), .ZN(n13530) );
  INV_X1 U16876 ( .A(n13694), .ZN(n13529) );
  NAND2_X1 U16877 ( .A1(n13530), .A2(n13529), .ZN(n15360) );
  INV_X1 U16878 ( .A(n15360), .ZN(n19216) );
  AOI22_X1 U16879 ( .A1(n16493), .A2(n19216), .B1(n19276), .B2(
        P2_REIP_REG_4__SCAN_IN), .ZN(n13531) );
  OAI211_X1 U16880 ( .C1(n16466), .C2(n19277), .A(n13532), .B(n13531), .ZN(
        n13533) );
  AOI21_X1 U16881 ( .B1(n19280), .B2(n16460), .A(n13533), .ZN(n13534) );
  OAI21_X1 U16882 ( .B1(n13535), .B2(n16498), .A(n13534), .ZN(P2_U3042) );
  XNOR2_X1 U16883 ( .A(n13537), .B(n13536), .ZN(n13565) );
  INV_X1 U16884 ( .A(n13538), .ZN(n20033) );
  INV_X1 U16885 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20742) );
  NOR2_X1 U16886 ( .A1(n16200), .A2(n20742), .ZN(n13562) );
  AOI21_X1 U16887 ( .B1(n16135), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n13562), .ZN(n13539) );
  OAI21_X1 U16888 ( .B1(n16127), .B2(n20029), .A(n13539), .ZN(n13540) );
  AOI21_X1 U16889 ( .B1(n20033), .B2(n16152), .A(n13540), .ZN(n13541) );
  OAI21_X1 U16890 ( .B1(n13565), .B2(n19970), .A(n13541), .ZN(P1_U2994) );
  INV_X1 U16891 ( .A(n14669), .ZN(n20168) );
  OAI222_X1 U16892 ( .A1(n14712), .A2(n13542), .B1(n14661), .B2(n10644), .C1(
        n14711), .C2(n20168), .ZN(P1_U2898) );
  XNOR2_X1 U16893 ( .A(n13543), .B(n13544), .ZN(n13557) );
  INV_X1 U16894 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n13545) );
  OR2_X1 U16895 ( .A1(n16200), .A2(n13545), .ZN(n13552) );
  NAND2_X1 U16896 ( .A1(n16135), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13546) );
  OAI211_X1 U16897 ( .C1(n16127), .C2(n20035), .A(n13552), .B(n13546), .ZN(
        n13547) );
  AOI21_X1 U16898 ( .B1(n20049), .B2(n16152), .A(n13547), .ZN(n13548) );
  OAI21_X1 U16899 ( .B1(n19970), .B2(n13557), .A(n13548), .ZN(P1_U2995) );
  AOI21_X1 U16900 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20101) );
  NOR2_X1 U16901 ( .A1(n16201), .A2(n13549), .ZN(n14888) );
  NAND2_X1 U16902 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14888), .ZN(
        n20113) );
  NOR2_X1 U16903 ( .A1(n16207), .A2(n16209), .ZN(n13657) );
  NOR2_X1 U16904 ( .A1(n20101), .A2(n13657), .ZN(n20086) );
  INV_X1 U16905 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20095) );
  NOR2_X1 U16906 ( .A1(n21014), .A2(n20095), .ZN(n14884) );
  AOI21_X1 U16907 ( .B1(n21014), .B2(n20095), .A(n14884), .ZN(n13555) );
  NAND2_X1 U16908 ( .A1(n15035), .A2(n20100), .ZN(n13550) );
  OAI21_X1 U16909 ( .B1(n11153), .B2(n10996), .A(n20099), .ZN(n13559) );
  NAND2_X1 U16910 ( .A1(n20097), .A2(n13559), .ZN(n16227) );
  AND2_X1 U16911 ( .A1(n16207), .A2(n20101), .ZN(n13551) );
  NOR2_X1 U16912 ( .A1(n16227), .A2(n13551), .ZN(n20096) );
  NOR2_X1 U16913 ( .A1(n20096), .A2(n21014), .ZN(n13554) );
  OAI21_X1 U16914 ( .B1(n20052), .B2(n20107), .A(n13552), .ZN(n13553) );
  AOI211_X1 U16915 ( .C1(n20086), .C2(n13555), .A(n13554), .B(n13553), .ZN(
        n13556) );
  OAI21_X1 U16916 ( .B1(n20091), .B2(n13557), .A(n13556), .ZN(P1_U3027) );
  INV_X1 U16917 ( .A(n14884), .ZN(n13561) );
  NOR3_X1 U16918 ( .A1(n13561), .A2(n13558), .A3(n20101), .ZN(n14889) );
  INV_X1 U16919 ( .A(n16207), .ZN(n20104) );
  OAI21_X1 U16920 ( .B1(n14889), .B2(n20104), .A(n20097), .ZN(n16204) );
  INV_X1 U16921 ( .A(n16204), .ZN(n13560) );
  OAI211_X1 U16922 ( .C1(n16201), .C2(n14884), .A(n13560), .B(n13559), .ZN(
        n13659) );
  NOR2_X1 U16923 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13561), .ZN(
        n13660) );
  AOI22_X1 U16924 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13659), .B1(
        n13660), .B2(n20086), .ZN(n13564) );
  AOI21_X1 U16925 ( .B1(n20023), .B2(n20116), .A(n13562), .ZN(n13563) );
  OAI211_X1 U16926 ( .C1(n20091), .C2(n13565), .A(n13564), .B(n13563), .ZN(
        P1_U3026) );
  XOR2_X1 U16927 ( .A(n13567), .B(n13566), .Z(n20110) );
  NAND2_X1 U16928 ( .A1(n20110), .A2(n11125), .ZN(n13571) );
  INV_X1 U16929 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20737) );
  OR2_X1 U16930 ( .A1(n16200), .A2(n20737), .ZN(n20105) );
  INV_X1 U16931 ( .A(n20105), .ZN(n13569) );
  NOR2_X1 U16932 ( .A1(n16127), .A2(n14584), .ZN(n13568) );
  AOI211_X1 U16933 ( .C1(n16135), .C2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13569), .B(n13568), .ZN(n13570) );
  OAI211_X1 U16934 ( .C1(n20129), .C2(n14594), .A(n13571), .B(n13570), .ZN(
        P1_U2997) );
  AND2_X1 U16935 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20815), .ZN(n13572) );
  NOR2_X1 U16936 ( .A1(n20547), .A2(n20814), .ZN(n16056) );
  AOI22_X1 U16937 ( .A1(n10960), .A2(n13572), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n16056), .ZN(n13573) );
  NAND2_X1 U16938 ( .A1(n16200), .A2(n13573), .ZN(n13574) );
  INV_X1 U16939 ( .A(n13597), .ZN(n13578) );
  INV_X1 U16940 ( .A(n13575), .ZN(n13576) );
  NAND2_X1 U16941 ( .A1(n13576), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13577) );
  INV_X1 U16942 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14369) );
  NAND2_X1 U16943 ( .A1(n14585), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13580) );
  OAI21_X1 U16944 ( .B1(n13579), .B2(n13578), .A(n14571), .ZN(n20048) );
  INV_X1 U16945 ( .A(n20048), .ZN(n14595) );
  INV_X1 U16946 ( .A(n13580), .ZN(n13581) );
  AND2_X2 U16947 ( .A1(n14719), .A2(n13581), .ZN(n20039) );
  INV_X1 U16948 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13601) );
  INV_X1 U16949 ( .A(n13583), .ZN(n13584) );
  AND2_X1 U16950 ( .A1(n13597), .A2(n13584), .ZN(n20037) );
  INV_X1 U16951 ( .A(n20037), .ZN(n13593) );
  AND2_X1 U16952 ( .A1(n20819), .A2(n20812), .ZN(n13588) );
  NAND2_X1 U16953 ( .A1(n13585), .A2(n13588), .ZN(n13595) );
  NOR2_X1 U16954 ( .A1(n13595), .A2(n10430), .ZN(n13586) );
  INV_X1 U16955 ( .A(n14590), .ZN(n14578) );
  INV_X1 U16956 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20734) );
  AOI22_X1 U16957 ( .A1(n14578), .A2(n20734), .B1(n20042), .B2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13592) );
  NAND2_X1 U16958 ( .A1(n13587), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13594) );
  NOR2_X1 U16959 ( .A1(n13594), .A2(n13588), .ZN(n13589) );
  NAND2_X1 U16960 ( .A1(n20024), .A2(n13590), .ZN(n13591) );
  OAI211_X1 U16961 ( .C1(n20464), .C2(n13593), .A(n13592), .B(n13591), .ZN(
        n13600) );
  AND3_X1 U16962 ( .A1(n13595), .A2(n20135), .A3(n13594), .ZN(n13596) );
  AND2_X2 U16963 ( .A1(n13597), .A2(n13596), .ZN(n20041) );
  INV_X1 U16964 ( .A(n14585), .ZN(n14479) );
  AOI22_X1 U16965 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(n20041), .B1(n14479), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n13598) );
  INV_X1 U16966 ( .A(n13598), .ZN(n13599) );
  AOI211_X1 U16967 ( .C1(n20039), .C2(n13601), .A(n13600), .B(n13599), .ZN(
        n13602) );
  OAI21_X1 U16968 ( .B1(n14595), .B2(n13603), .A(n13602), .ZN(P1_U2839) );
  INV_X1 U16969 ( .A(n13604), .ZN(n13607) );
  INV_X1 U16970 ( .A(n13606), .ZN(n13805) );
  OAI21_X1 U16971 ( .B1(n13608), .B2(n13607), .A(n13805), .ZN(n20006) );
  OAI21_X1 U16972 ( .B1(n13610), .B2(n13609), .A(n13813), .ZN(n13611) );
  INV_X1 U16973 ( .A(n13611), .ZN(n20005) );
  AOI22_X1 U16974 ( .A1(n20005), .A2(n16115), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n14623), .ZN(n13612) );
  OAI21_X1 U16975 ( .B1(n20006), .B2(n14628), .A(n13612), .ZN(P1_U2865) );
  NAND2_X1 U16976 ( .A1(n14590), .A2(n14585), .ZN(n19996) );
  INV_X1 U16977 ( .A(n19996), .ZN(n16095) );
  INV_X1 U16978 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n20125) );
  NOR2_X1 U16979 ( .A1(n16095), .A2(n20125), .ZN(n13615) );
  OAI22_X1 U16980 ( .A1(n13613), .A2(n20000), .B1(n20053), .B2(n20114), .ZN(
        n13614) );
  AOI211_X1 U16981 ( .C1(n20037), .C2(n10552), .A(n13615), .B(n13614), .ZN(
        n13617) );
  OAI21_X1 U16982 ( .B1(n20039), .B2(n20042), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13616) );
  OAI211_X1 U16983 ( .C1(n14595), .C2(n13618), .A(n13617), .B(n13616), .ZN(
        P1_U2840) );
  INV_X1 U16984 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n13627) );
  OAI211_X1 U16985 ( .C1(n13620), .C2(n13622), .A(n13621), .B(n19151), .ZN(
        n13626) );
  INV_X1 U16986 ( .A(n15829), .ZN(n13624) );
  OAI21_X1 U16987 ( .B1(n13624), .B2(n10123), .A(n15305), .ZN(n19020) );
  INV_X1 U16988 ( .A(n19020), .ZN(n16448) );
  NAND2_X1 U16989 ( .A1(n19164), .A2(n16448), .ZN(n13625) );
  OAI211_X1 U16990 ( .C1(n19164), .C2(n13627), .A(n13626), .B(n13625), .ZN(
        P2_U2872) );
  AOI21_X1 U16991 ( .B1(n16429), .B2(n13630), .A(n15113), .ZN(n16416) );
  INV_X1 U16992 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13629) );
  INV_X1 U16993 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15559) );
  INV_X1 U16994 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15577) );
  INV_X1 U16995 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18993) );
  INV_X1 U16996 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15109) );
  INV_X1 U16997 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15616) );
  INV_X1 U16998 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15210) );
  INV_X1 U16999 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16272) );
  NAND2_X1 U17000 ( .A1(n15103), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13628) );
  OAI22_X1 U17001 ( .A1(n16510), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19138) );
  INV_X1 U17002 ( .A(n19138), .ZN(n15378) );
  AOI22_X1 U17003 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15914), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16510), .ZN(n15377) );
  NOR2_X1 U17004 ( .A1(n15378), .A2(n15377), .ZN(n15376) );
  OAI21_X1 U17005 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n13630), .ZN(n19292) );
  NAND2_X1 U17006 ( .A1(n15376), .A2(n19292), .ZN(n15111) );
  NAND2_X1 U17007 ( .A1(n9740), .A2(n15111), .ZN(n13631) );
  XNOR2_X1 U17008 ( .A(n16416), .B(n13631), .ZN(n13653) );
  NOR2_X1 U17009 ( .A1(n19567), .A2(n19130), .ZN(n13652) );
  NOR2_X1 U17010 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19952), .ZN(n13644) );
  INV_X1 U17011 ( .A(n13644), .ZN(n13633) );
  NOR2_X1 U17012 ( .A1(n13635), .A2(n13633), .ZN(n13632) );
  NAND2_X1 U17013 ( .A1(n19953), .A2(n13632), .ZN(n19085) );
  NAND2_X1 U17014 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13633), .ZN(n13634) );
  NOR2_X1 U17015 ( .A1(n13635), .A2(n13634), .ZN(n13636) );
  NOR3_X1 U17016 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13637), .A3(n19757), 
        .ZN(n16504) );
  INV_X1 U17017 ( .A(n16504), .ZN(n13638) );
  NAND2_X1 U17018 ( .A1(n19090), .A2(n13638), .ZN(n13639) );
  OR2_X1 U17019 ( .A1(n19276), .A2(n13639), .ZN(n13640) );
  OAI22_X1 U17020 ( .A1(n19107), .A2(n13641), .B1(n11446), .B2(n19129), .ZN(
        n13649) );
  INV_X1 U17021 ( .A(n13642), .ZN(n13643) );
  NAND2_X1 U17022 ( .A1(n19272), .A2(n13643), .ZN(n15140) );
  NOR2_X1 U17023 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13644), .ZN(n13645) );
  NAND2_X1 U17024 ( .A1(n13646), .A2(n13645), .ZN(n13647) );
  INV_X1 U17025 ( .A(n9717), .ZN(n18992) );
  OAI22_X1 U17026 ( .A1(n19109), .A2(n21011), .B1(n16429), .B2(n18992), .ZN(
        n13648) );
  AOI211_X1 U17027 ( .C1(n19133), .C2(n16425), .A(n13649), .B(n13648), .ZN(
        n13650) );
  OAI21_X1 U17028 ( .B1(n19900), .B2(n19121), .A(n13650), .ZN(n13651) );
  AOI211_X1 U17029 ( .C1(n13653), .C2(n19117), .A(n13652), .B(n13651), .ZN(
        n13654) );
  INV_X1 U17030 ( .A(n13654), .ZN(P2_U2852) );
  XOR2_X1 U17031 ( .A(n13656), .B(n13655), .Z(n13668) );
  INV_X1 U17032 ( .A(n14889), .ZN(n16228) );
  INV_X1 U17033 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n13658) );
  OR2_X1 U17034 ( .A1(n16200), .A2(n13658), .ZN(n13665) );
  OAI21_X1 U17035 ( .B1(n20014), .B2(n20107), .A(n13665), .ZN(n13662) );
  AOI21_X1 U17036 ( .B1(n16209), .B2(n13660), .A(n13659), .ZN(n13918) );
  NOR2_X1 U17037 ( .A1(n13918), .A2(n14886), .ZN(n13661) );
  AOI211_X1 U17038 ( .C1(n16231), .C2(n14886), .A(n13662), .B(n13661), .ZN(
        n13663) );
  OAI21_X1 U17039 ( .B1(n13668), .B2(n20091), .A(n13663), .ZN(P1_U3025) );
  NAND2_X1 U17040 ( .A1(n16135), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13664) );
  OAI211_X1 U17041 ( .C1(n16127), .C2(n20012), .A(n13665), .B(n13664), .ZN(
        n13666) );
  AOI21_X1 U17042 ( .B1(n20019), .B2(n16152), .A(n13666), .ZN(n13667) );
  OAI21_X1 U17043 ( .B1(n13668), .B2(n19970), .A(n13667), .ZN(P1_U2993) );
  OAI222_X1 U17044 ( .A1(n14712), .A2(n20006), .B1(n14661), .B2(n10656), .C1(
        n14711), .C2(n20174), .ZN(P1_U2897) );
  NOR2_X2 U17045 ( .A1(n19687), .A2(n19713), .ZN(n19708) );
  NOR2_X2 U17046 ( .A1(n19683), .A2(n19888), .ZN(n19678) );
  OAI21_X1 U17047 ( .B1(n19708), .B2(n19678), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13673) );
  NOR2_X1 U17048 ( .A1(n13670), .A2(n13669), .ZN(n19426) );
  NAND2_X1 U17049 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19426), .ZN(
        n13677) );
  NAND2_X1 U17050 ( .A1(n11603), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13671) );
  NAND3_X1 U17051 ( .A1(n19922), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19689) );
  NOR2_X1 U17052 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19689), .ZN(
        n19676) );
  AOI21_X1 U17053 ( .B1(n13671), .B2(n19757), .A(n19676), .ZN(n13672) );
  INV_X1 U17054 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14141) );
  INV_X1 U17055 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16587) );
  INV_X1 U17056 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n17382) );
  OAI22_X2 U17057 ( .A1(n16587), .A2(n19338), .B1(n17382), .B2(n19336), .ZN(
        n19767) );
  AOI22_X1 U17058 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19335), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19334), .ZN(n19770) );
  INV_X1 U17059 ( .A(n19770), .ZN(n19637) );
  AOI22_X1 U17060 ( .A1(n19678), .A2(n19767), .B1(n19708), .B2(n19637), .ZN(
        n13680) );
  INV_X1 U17061 ( .A(n11603), .ZN(n13675) );
  OAI21_X1 U17062 ( .B1(n13675), .B2(n19676), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13676) );
  OAI21_X1 U17063 ( .B1(n13677), .B2(n19719), .A(n13676), .ZN(n19677) );
  NOR2_X2 U17064 ( .A1(n13678), .A2(n19343), .ZN(n19760) );
  AOI22_X1 U17065 ( .A1(n19677), .A2(n19760), .B1(n19759), .B2(n19676), .ZN(
        n13679) );
  OAI211_X1 U17066 ( .C1(n19682), .C2(n14141), .A(n13680), .B(n13679), .ZN(
        P2_U3144) );
  INV_X1 U17067 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13685) );
  INV_X1 U17068 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20859) );
  INV_X1 U17069 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n17370) );
  OAI22_X2 U17070 ( .A1(n20859), .A2(n19338), .B1(n17370), .B2(n19336), .ZN(
        n19779) );
  AOI22_X1 U17071 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19335), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19334), .ZN(n19782) );
  INV_X1 U17072 ( .A(n19782), .ZN(n19643) );
  AOI22_X1 U17073 ( .A1(n19678), .A2(n19779), .B1(n19708), .B2(n19643), .ZN(
        n13684) );
  INV_X1 U17074 ( .A(n16311), .ZN(n13681) );
  NOR2_X2 U17075 ( .A1(n13681), .A2(n19343), .ZN(n19778) );
  NOR2_X2 U17076 ( .A1(n13682), .A2(n19340), .ZN(n19777) );
  AOI22_X1 U17077 ( .A1(n19677), .A2(n19778), .B1(n19676), .B2(n19777), .ZN(
        n13683) );
  OAI211_X1 U17078 ( .C1(n19682), .C2(n13685), .A(n13684), .B(n13683), .ZN(
        P2_U3146) );
  XNOR2_X1 U17079 ( .A(n13686), .B(n13687), .ZN(n16411) );
  INV_X1 U17080 ( .A(n13689), .ZN(n13691) );
  AND2_X1 U17081 ( .A1(n13689), .A2(n13688), .ZN(n13690) );
  INV_X1 U17082 ( .A(n16410), .ZN(n13703) );
  XNOR2_X1 U17083 ( .A(n13694), .B(n13693), .ZN(n19214) );
  NAND2_X1 U17084 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13695), .ZN(
        n16470) );
  INV_X1 U17085 ( .A(n16470), .ZN(n13698) );
  NOR2_X1 U17086 ( .A1(n11998), .A2(n9725), .ZN(n13696) );
  AOI221_X1 U17087 ( .B1(n13698), .B2(n20980), .C1(n13697), .C2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n13696), .ZN(n13701) );
  INV_X1 U17088 ( .A(n13699), .ZN(n19116) );
  NAND2_X1 U17089 ( .A1(n19116), .A2(n16494), .ZN(n13700) );
  OAI211_X1 U17090 ( .C1(n19214), .C2(n16479), .A(n13701), .B(n13700), .ZN(
        n13702) );
  AOI21_X1 U17091 ( .B1(n13703), .B2(n16460), .A(n13702), .ZN(n13704) );
  OAI21_X1 U17092 ( .B1(n16498), .B2(n16411), .A(n13704), .ZN(P2_U3041) );
  NAND2_X1 U17093 ( .A1(n19567), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19896) );
  NAND2_X1 U17094 ( .A1(n19714), .A2(n19903), .ZN(n13712) );
  OAI21_X1 U17095 ( .B1(n19896), .B2(n19712), .A(n13712), .ZN(n13707) );
  NAND2_X1 U17096 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19903), .ZN(
        n19490) );
  NOR2_X1 U17097 ( .A1(n19629), .A2(n19490), .ZN(n19533) );
  INV_X1 U17098 ( .A(n19533), .ZN(n13705) );
  OAI211_X1 U17099 ( .C1(n13709), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19719), 
        .B(n13705), .ZN(n13706) );
  NAND3_X1 U17100 ( .A1(n13707), .A2(n19765), .A3(n13706), .ZN(n19526) );
  INV_X1 U17101 ( .A(n19526), .ZN(n13718) );
  INV_X1 U17102 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14134) );
  NAND2_X1 U17103 ( .A1(n19567), .A2(n19925), .ZN(n19427) );
  AOI22_X1 U17104 ( .A1(n19492), .A2(n19767), .B1(n19560), .B2(n19637), .ZN(
        n13714) );
  INV_X1 U17105 ( .A(n13709), .ZN(n13710) );
  OAI21_X1 U17106 ( .B1(n13710), .B2(n19533), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13711) );
  OAI21_X1 U17107 ( .B1(n13712), .B2(n19719), .A(n13711), .ZN(n19525) );
  AOI22_X1 U17108 ( .A1(n19525), .A2(n19760), .B1(n19759), .B2(n19533), .ZN(
        n13713) );
  OAI211_X1 U17109 ( .C1(n13718), .C2(n14134), .A(n13714), .B(n13713), .ZN(
        P2_U3104) );
  INV_X1 U17110 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13717) );
  AOI22_X1 U17111 ( .A1(n19492), .A2(n19779), .B1(n19560), .B2(n19643), .ZN(
        n13716) );
  AOI22_X1 U17112 ( .A1(n19525), .A2(n19778), .B1(n19777), .B2(n19533), .ZN(
        n13715) );
  OAI211_X1 U17113 ( .C1(n13718), .C2(n13717), .A(n13716), .B(n13715), .ZN(
        P2_U3106) );
  OAI21_X1 U17114 ( .B1(n13721), .B2(n13720), .A(n13719), .ZN(n16252) );
  NAND2_X1 U17115 ( .A1(n16252), .A2(n11125), .ZN(n13725) );
  INV_X1 U17116 ( .A(n20002), .ZN(n13723) );
  INV_X1 U17117 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20745) );
  OR2_X1 U17118 ( .A1(n16200), .A2(n20745), .ZN(n16248) );
  OAI21_X1 U17119 ( .B1(n14818), .B2(n19998), .A(n16248), .ZN(n13722) );
  AOI21_X1 U17120 ( .B1(n13723), .B2(n16151), .A(n13722), .ZN(n13724) );
  OAI211_X1 U17121 ( .C1(n20129), .C2(n20006), .A(n13725), .B(n13724), .ZN(
        P1_U2992) );
  OAI21_X1 U17122 ( .B1(n15303), .B2(n13727), .A(n13726), .ZN(n19009) );
  AOI22_X1 U17123 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11575), .B1(
        n11588), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13736) );
  AOI22_X1 U17124 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12262), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13735) );
  OAI22_X1 U17125 ( .A1(n13728), .A2(n14101), .B1(n14099), .B2(n14174), .ZN(
        n13733) );
  NAND2_X1 U17126 ( .A1(n11513), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13730) );
  NAND2_X1 U17127 ( .A1(n11537), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n13729) );
  OAI211_X1 U17128 ( .C1(n14153), .C2(n13731), .A(n13730), .B(n13729), .ZN(
        n13732) );
  NOR2_X1 U17129 ( .A1(n13733), .A2(n13732), .ZN(n13734) );
  NAND3_X1 U17130 ( .A1(n13736), .A2(n13735), .A3(n13734), .ZN(n13742) );
  AOI22_X1 U17131 ( .A1(n14162), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14161), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13740) );
  AOI22_X1 U17132 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n11529), .B1(
        n13998), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13739) );
  AOI22_X1 U17133 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11528), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13738) );
  NAND2_X1 U17134 ( .A1(n11523), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13737) );
  NAND4_X1 U17135 ( .A1(n13740), .A2(n13739), .A3(n13738), .A4(n13737), .ZN(
        n13741) );
  NOR2_X1 U17136 ( .A1(n13742), .A2(n13741), .ZN(n13762) );
  AOI22_X1 U17137 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11588), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13750) );
  AOI22_X1 U17138 ( .A1(n12262), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13749) );
  INV_X1 U17139 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13944) );
  NAND2_X1 U17140 ( .A1(n11513), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13745) );
  NAND2_X1 U17141 ( .A1(n11537), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n13744) );
  OAI211_X1 U17142 ( .C1(n14153), .C2(n13944), .A(n13745), .B(n13744), .ZN(
        n13746) );
  INV_X1 U17143 ( .A(n13746), .ZN(n13748) );
  AOI22_X1 U17144 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14155), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13747) );
  NAND4_X1 U17145 ( .A1(n13750), .A2(n13749), .A3(n13748), .A4(n13747), .ZN(
        n13756) );
  AOI22_X1 U17146 ( .A1(n14162), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14161), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13754) );
  AOI22_X1 U17147 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9741), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13753) );
  AOI22_X1 U17148 ( .A1(n11528), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13752) );
  NAND2_X1 U17149 ( .A1(n11523), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13751) );
  NAND4_X1 U17150 ( .A1(n13754), .A2(n13753), .A3(n13752), .A4(n13751), .ZN(
        n13755) );
  NOR2_X1 U17151 ( .A1(n13756), .A2(n13755), .ZN(n19140) );
  INV_X1 U17152 ( .A(n19140), .ZN(n13757) );
  INV_X1 U17153 ( .A(n13762), .ZN(n13759) );
  INV_X1 U17154 ( .A(n13760), .ZN(n13761) );
  AOI21_X1 U17155 ( .B1(n13762), .B2(n13758), .A(n13761), .ZN(n13969) );
  NAND2_X1 U17156 ( .A1(n13969), .A2(n19151), .ZN(n13764) );
  NAND2_X1 U17157 ( .A1(n19161), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13763) );
  OAI211_X1 U17158 ( .C1(n19009), .C2(n19161), .A(n13764), .B(n13763), .ZN(
        P2_U2870) );
  XNOR2_X1 U17159 ( .A(n13765), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13785) );
  XOR2_X1 U17160 ( .A(n13768), .B(n13767), .Z(n13783) );
  NOR2_X1 U17161 ( .A1(n20980), .A2(n16470), .ZN(n13772) );
  OAI21_X1 U17162 ( .B1(n16491), .B2(n13770), .A(n13769), .ZN(n16481) );
  INV_X1 U17163 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19845) );
  NOR2_X1 U17164 ( .A1(n19845), .A2(n9725), .ZN(n13771) );
  AOI221_X1 U17165 ( .B1(n13772), .B2(n16471), .C1(n16481), .C2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n13771), .ZN(n13773) );
  INV_X1 U17166 ( .A(n13773), .ZN(n13777) );
  XOR2_X1 U17167 ( .A(n13775), .B(n13774), .Z(n19206) );
  OAI22_X1 U17168 ( .A1(n19101), .A2(n16466), .B1(n16479), .B2(n19206), .ZN(
        n13776) );
  AOI211_X1 U17169 ( .C1(n13783), .C2(n16485), .A(n13777), .B(n13776), .ZN(
        n13778) );
  OAI21_X1 U17170 ( .B1(n13785), .B2(n16503), .A(n13778), .ZN(P2_U3040) );
  OAI21_X1 U17171 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n15110), .A(
        n13912), .ZN(n19099) );
  OAI22_X1 U17172 ( .A1(n19845), .A2(n9725), .B1(n19291), .B2(n19099), .ZN(
        n13780) );
  AOI21_X1 U17173 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19284), .A(
        n13780), .ZN(n13781) );
  OAI21_X1 U17174 ( .B1(n19101), .B2(n13674), .A(n13781), .ZN(n13782) );
  AOI21_X1 U17175 ( .B1(n13783), .B2(n19285), .A(n13782), .ZN(n13784) );
  OAI21_X1 U17176 ( .B1(n13785), .B2(n16418), .A(n13784), .ZN(P2_U3008) );
  AND2_X1 U17177 ( .A1(n13786), .A2(n13787), .ZN(n13789) );
  OR2_X1 U17178 ( .A1(n13789), .A2(n13788), .ZN(n13951) );
  AOI21_X1 U17179 ( .B1(n13790), .B2(n13811), .A(n13927), .ZN(n16241) );
  AOI22_X1 U17180 ( .A1(n16241), .A2(n16115), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n14623), .ZN(n13791) );
  OAI21_X1 U17181 ( .B1(n13951), .B2(n14628), .A(n13791), .ZN(P1_U2863) );
  INV_X1 U17182 ( .A(n13947), .ZN(n13799) );
  NAND4_X1 U17183 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n14361)
         );
  NAND4_X1 U17184 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n14362)
         );
  NOR2_X1 U17185 ( .A1(n14361), .A2(n20028), .ZN(n14501) );
  INV_X1 U17186 ( .A(n14501), .ZN(n14560) );
  INV_X1 U17187 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20748) );
  NAND3_X1 U17188 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n13792) );
  NOR2_X1 U17189 ( .A1(n14479), .A2(n13792), .ZN(n20040) );
  NAND2_X1 U17190 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20040), .ZN(n19997) );
  NAND2_X1 U17191 ( .A1(n19996), .A2(n19997), .ZN(n20045) );
  INV_X1 U17192 ( .A(n20045), .ZN(n13793) );
  AOI21_X1 U17193 ( .B1(n14361), .B2(n19996), .A(n13793), .ZN(n19995) );
  OAI22_X1 U17194 ( .A1(n13795), .A2(n19999), .B1(n13794), .B2(n20000), .ZN(
        n13796) );
  AOI211_X1 U17195 ( .C1(n20024), .C2(n16241), .A(n19987), .B(n13796), .ZN(
        n13797) );
  OAI221_X1 U17196 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n14560), .C1(n20748), 
        .C2(n19995), .A(n13797), .ZN(n13798) );
  AOI21_X1 U17197 ( .B1(n20039), .B2(n13799), .A(n13798), .ZN(n13800) );
  OAI21_X1 U17198 ( .B1(n13951), .B2(n14571), .A(n13800), .ZN(P1_U2831) );
  NAND2_X1 U17199 ( .A1(n10162), .A2(n13802), .ZN(n13803) );
  XNOR2_X1 U17200 ( .A(n13801), .B(n13803), .ZN(n13924) );
  INV_X1 U17201 ( .A(n13786), .ZN(n13804) );
  AOI21_X1 U17202 ( .B1(n13806), .B2(n13805), .A(n13804), .ZN(n19993) );
  AOI22_X1 U17203 ( .A1(n16135), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16171), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13807) );
  OAI21_X1 U17204 ( .B1(n16127), .B2(n13808), .A(n13807), .ZN(n13809) );
  AOI21_X1 U17205 ( .B1(n19993), .B2(n16152), .A(n13809), .ZN(n13810) );
  OAI21_X1 U17206 ( .B1(n13924), .B2(n19970), .A(n13810), .ZN(P1_U2991) );
  INV_X1 U17207 ( .A(n19993), .ZN(n13817) );
  INV_X1 U17208 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13815) );
  INV_X1 U17209 ( .A(n13811), .ZN(n13812) );
  AOI21_X1 U17210 ( .B1(n13814), .B2(n13813), .A(n13812), .ZN(n13922) );
  INV_X1 U17211 ( .A(n13922), .ZN(n19990) );
  OAI222_X1 U17212 ( .A1(n13817), .A2(n14638), .B1(n13815), .B2(n16118), .C1(
        n14636), .C2(n19990), .ZN(P1_U2864) );
  INV_X1 U17213 ( .A(DATAI_8_), .ZN(n13816) );
  INV_X1 U17214 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16611) );
  MUX2_X1 U17215 ( .A(n13816), .B(n16611), .S(n20130), .Z(n20054) );
  OAI222_X1 U17216 ( .A1(n13817), .A2(n14712), .B1(n13425), .B2(n14661), .C1(
        n14711), .C2(n20054), .ZN(P1_U2896) );
  INV_X1 U17217 ( .A(DATAI_9_), .ZN(n13818) );
  MUX2_X1 U17218 ( .A(n13818), .B(n21045), .S(n20130), .Z(n20057) );
  OAI222_X1 U17219 ( .A1(n13951), .A2(n14712), .B1(n13436), .B2(n14661), .C1(
        n14711), .C2(n20057), .ZN(P1_U2895) );
  OAI21_X1 U17220 ( .B1(n13788), .B2(n13820), .A(n13819), .ZN(n13925) );
  INV_X1 U17221 ( .A(DATAI_10_), .ZN(n13821) );
  MUX2_X1 U17222 ( .A(n13821), .B(n16608), .S(n20130), .Z(n20060) );
  OAI222_X1 U17223 ( .A1(n13925), .A2(n14712), .B1(n13439), .B2(n14661), .C1(
        n14711), .C2(n20060), .ZN(P1_U2894) );
  NOR2_X1 U17224 ( .A1(n13822), .A2(n17392), .ZN(n13824) );
  INV_X1 U17225 ( .A(n18769), .ZN(n15988) );
  INV_X1 U17226 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n13827) );
  INV_X1 U17227 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n20981) );
  INV_X1 U17228 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17323) );
  NAND2_X1 U17229 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17327) );
  OR4_X1 U17230 ( .A1(n20981), .A2(n17319), .A3(n17323), .A4(n17327), .ZN(
        n17284) );
  INV_X1 U17231 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17311) );
  NOR3_X1 U17232 ( .A1(n17310), .A2(n17311), .A3(n17307), .ZN(n17285) );
  NAND3_X1 U17233 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17316), .A3(n17285), .ZN(
        n17281) );
  NAND2_X1 U17234 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17253), .ZN(n17250) );
  AND4_X1 U17235 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(P3_EBX_REG_13__SCAN_IN), .A4(P3_EBX_REG_12__SCAN_IN), .ZN(n14028)
         );
  AND2_X1 U17236 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(P3_EBX_REG_16__SCAN_IN), 
        .ZN(n17182) );
  NAND4_X1 U17237 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17237), .A3(n14028), 
        .A4(n17182), .ZN(n17170) );
  NOR2_X1 U17238 ( .A1(n17392), .A2(n17154), .ZN(n17142) );
  NAND2_X1 U17239 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17142), .ZN(n17130) );
  NAND2_X1 U17240 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17107), .ZN(n17098) );
  AND2_X1 U17241 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17093) );
  NAND2_X1 U17242 ( .A1(n18332), .A2(n17334), .ZN(n17340) );
  OAI22_X1 U17243 ( .A1(n17338), .A2(n17103), .B1(n17093), .B2(n17340), .ZN(
        n17091) );
  AOI22_X1 U17244 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15951), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13831) );
  AOI22_X1 U17245 ( .A1(n17256), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13830) );
  AOI22_X1 U17246 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13829) );
  AOI22_X1 U17247 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15952), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13828) );
  NAND4_X1 U17248 ( .A1(n13831), .A2(n13830), .A3(n13829), .A4(n13828), .ZN(
        n13837) );
  AOI22_X1 U17249 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13835) );
  AOI22_X1 U17250 ( .A1(n15949), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13834) );
  AOI22_X1 U17251 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13833) );
  AOI22_X1 U17252 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13891), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13832) );
  NAND4_X1 U17253 ( .A1(n13835), .A2(n13834), .A3(n13833), .A4(n13832), .ZN(
        n13836) );
  NOR2_X1 U17254 ( .A1(n13837), .A2(n13836), .ZN(n13902) );
  AOI22_X1 U17255 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15951), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13841) );
  AOI22_X1 U17256 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13840) );
  AOI22_X1 U17257 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13839) );
  AOI22_X1 U17258 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13838) );
  NAND4_X1 U17259 ( .A1(n13841), .A2(n13840), .A3(n13839), .A4(n13838), .ZN(
        n13847) );
  AOI22_X1 U17260 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15949), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13845) );
  AOI22_X1 U17261 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17288), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13844) );
  AOI22_X1 U17262 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13843) );
  AOI22_X1 U17263 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13842) );
  NAND4_X1 U17264 ( .A1(n13845), .A2(n13844), .A3(n13843), .A4(n13842), .ZN(
        n13846) );
  NOR2_X1 U17265 ( .A1(n13847), .A2(n13846), .ZN(n17100) );
  AOI22_X1 U17266 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17287), .ZN(n13851) );
  AOI22_X1 U17267 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13850) );
  AOI22_X1 U17268 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17254), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17274), .ZN(n13849) );
  AOI22_X1 U17269 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n9722), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17269), .ZN(n13848) );
  NAND4_X1 U17270 ( .A1(n13851), .A2(n13850), .A3(n13849), .A4(n13848), .ZN(
        n13857) );
  AOI22_X1 U17271 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13855) );
  AOI22_X1 U17272 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n9726), .ZN(n13854) );
  AOI22_X1 U17273 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17268), .B1(
        n13891), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13853) );
  AOI22_X1 U17274 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17286), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n15949), .ZN(n13852) );
  NAND4_X1 U17275 ( .A1(n13855), .A2(n13854), .A3(n13853), .A4(n13852), .ZN(
        n13856) );
  NOR2_X1 U17276 ( .A1(n13857), .A2(n13856), .ZN(n17109) );
  AOI22_X1 U17277 ( .A1(n17287), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13869) );
  AOI22_X1 U17278 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13868) );
  AOI22_X1 U17279 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15949), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13858) );
  OAI21_X1 U17280 ( .B1(n13859), .B2(n21100), .A(n13858), .ZN(n13866) );
  AOI22_X1 U17281 ( .A1(n13891), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13864) );
  AOI22_X1 U17282 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13863) );
  AOI22_X1 U17283 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13862) );
  AOI22_X1 U17284 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13861) );
  NAND4_X1 U17285 ( .A1(n13864), .A2(n13863), .A3(n13862), .A4(n13861), .ZN(
        n13865) );
  AOI211_X1 U17286 ( .C1(n17254), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n13866), .B(n13865), .ZN(n13867) );
  NAND3_X1 U17287 ( .A1(n13869), .A2(n13868), .A3(n13867), .ZN(n17115) );
  AOI22_X1 U17288 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13880) );
  AOI22_X1 U17289 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13879) );
  AOI22_X1 U17290 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13870) );
  OAI21_X1 U17291 ( .B1(n13871), .B2(n20889), .A(n13870), .ZN(n13877) );
  AOI22_X1 U17292 ( .A1(n15950), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15951), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13875) );
  AOI22_X1 U17293 ( .A1(n15949), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13874) );
  AOI22_X1 U17294 ( .A1(n13891), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13873) );
  AOI22_X1 U17295 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15952), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13872) );
  NAND4_X1 U17296 ( .A1(n13875), .A2(n13874), .A3(n13873), .A4(n13872), .ZN(
        n13876) );
  AOI211_X1 U17297 ( .C1(n9722), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n13877), .B(n13876), .ZN(n13878) );
  NAND3_X1 U17298 ( .A1(n13880), .A2(n13879), .A3(n13878), .ZN(n17116) );
  NAND2_X1 U17299 ( .A1(n17115), .A2(n17116), .ZN(n17114) );
  NOR2_X1 U17300 ( .A1(n17109), .A2(n17114), .ZN(n17108) );
  AOI22_X1 U17301 ( .A1(n12577), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13890) );
  AOI22_X1 U17302 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13889) );
  AOI22_X1 U17303 ( .A1(n17256), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13881) );
  OAI21_X1 U17304 ( .B1(n17075), .B2(n17329), .A(n13881), .ZN(n13887) );
  AOI22_X1 U17305 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15951), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13885) );
  AOI22_X1 U17306 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13884) );
  AOI22_X1 U17307 ( .A1(n15950), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13883) );
  AOI22_X1 U17308 ( .A1(n13891), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15952), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13882) );
  NAND4_X1 U17309 ( .A1(n13885), .A2(n13884), .A3(n13883), .A4(n13882), .ZN(
        n13886) );
  AOI211_X1 U17310 ( .C1(n9722), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n13887), .B(n13886), .ZN(n13888) );
  NAND3_X1 U17311 ( .A1(n13890), .A2(n13889), .A3(n13888), .ZN(n17105) );
  NAND2_X1 U17312 ( .A1(n17108), .A2(n17105), .ZN(n17104) );
  NOR2_X1 U17313 ( .A1(n17100), .A2(n17104), .ZN(n17099) );
  AOI22_X1 U17314 ( .A1(n13891), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13901) );
  AOI22_X1 U17315 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13900) );
  AOI22_X1 U17316 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13892) );
  OAI21_X1 U17317 ( .B1(n17075), .B2(n17320), .A(n13892), .ZN(n13898) );
  AOI22_X1 U17318 ( .A1(n15950), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15949), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13896) );
  AOI22_X1 U17319 ( .A1(n17256), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15951), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13895) );
  AOI22_X1 U17320 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13894) );
  AOI22_X1 U17321 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15952), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13893) );
  NAND4_X1 U17322 ( .A1(n13896), .A2(n13895), .A3(n13894), .A4(n13893), .ZN(
        n13897) );
  AOI211_X1 U17323 ( .C1(n9722), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n13898), .B(n13897), .ZN(n13899) );
  NAND3_X1 U17324 ( .A1(n13901), .A2(n13900), .A3(n13899), .ZN(n17096) );
  NAND2_X1 U17325 ( .A1(n17099), .A2(n17096), .ZN(n17095) );
  NOR2_X1 U17326 ( .A1(n13902), .A2(n17095), .ZN(n17090) );
  AOI21_X1 U17327 ( .B1(n13902), .B2(n17095), .A(n17090), .ZN(n17357) );
  AOI22_X1 U17328 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17091), .B1(n17357), 
        .B2(n17338), .ZN(n13905) );
  INV_X1 U17329 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n13903) );
  NAND3_X1 U17330 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n13903), .A3(n17103), 
        .ZN(n13904) );
  NAND2_X1 U17331 ( .A1(n13905), .A2(n13904), .ZN(P3_U2675) );
  XNOR2_X1 U17332 ( .A(n13906), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13907) );
  XNOR2_X1 U17333 ( .A(n13908), .B(n13907), .ZN(n16489) );
  INV_X1 U17334 ( .A(n13910), .ZN(n16397) );
  NAND2_X1 U17335 ( .A1(n16397), .A2(n16396), .ZN(n13911) );
  XNOR2_X1 U17336 ( .A(n13909), .B(n13911), .ZN(n16486) );
  OAI22_X1 U17337 ( .A1(n16428), .A2(n13913), .B1(n12005), .B2(n9725), .ZN(
        n13916) );
  AOI21_X1 U17338 ( .B1(n13913), .B2(n13912), .A(n15115), .ZN(n19080) );
  INV_X1 U17339 ( .A(n19080), .ZN(n13914) );
  OAI22_X1 U17340 ( .A1(n19291), .A2(n13914), .B1(n13674), .B2(n19086), .ZN(
        n13915) );
  AOI211_X1 U17341 ( .C1(n16486), .C2(n19285), .A(n13916), .B(n13915), .ZN(
        n13917) );
  OAI21_X1 U17342 ( .B1(n16489), .B2(n16418), .A(n13917), .ZN(P2_U3007) );
  INV_X1 U17343 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20746) );
  OAI21_X1 U17344 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15043), .A(
        n13918), .ZN(n16247) );
  INV_X1 U17345 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14887) );
  NAND2_X1 U17346 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16231), .ZN(
        n16250) );
  AOI221_X1 U17347 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n14887), .C2(n11040), .A(
        n16250), .ZN(n13919) );
  AOI21_X1 U17348 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16247), .A(
        n13919), .ZN(n13920) );
  OAI21_X1 U17349 ( .B1(n16200), .B2(n20746), .A(n13920), .ZN(n13921) );
  AOI21_X1 U17350 ( .B1(n13922), .B2(n20116), .A(n13921), .ZN(n13923) );
  OAI21_X1 U17351 ( .B1(n13924), .B2(n20091), .A(n13923), .ZN(P1_U3023) );
  INV_X1 U17352 ( .A(n13925), .ZN(n16153) );
  OR2_X1 U17353 ( .A1(n13927), .A2(n13926), .ZN(n13928) );
  NAND2_X1 U17354 ( .A1(n13955), .A2(n13928), .ZN(n16235) );
  OAI22_X1 U17355 ( .A1(n16235), .A2(n14636), .B1(n16109), .B2(n16118), .ZN(
        n13929) );
  AOI21_X1 U17356 ( .B1(n16153), .B2(n16116), .A(n13929), .ZN(n13930) );
  INV_X1 U17357 ( .A(n13930), .ZN(P1_U2862) );
  INV_X1 U17358 ( .A(n13931), .ZN(n13935) );
  NAND2_X1 U17359 ( .A1(n19903), .A2(n19912), .ZN(n19395) );
  NOR2_X1 U17360 ( .A1(n19598), .A2(n19395), .ZN(n19389) );
  AOI21_X1 U17361 ( .B1(n13935), .B2(n19757), .A(n19389), .ZN(n13933) );
  NOR2_X2 U17362 ( .A1(n19568), .A2(n19458), .ZN(n19391) );
  NOR2_X1 U17363 ( .A1(n19601), .A2(n19395), .ZN(n13936) );
  AOI221_X1 U17364 ( .B1(n19391), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19412), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n13936), .ZN(n13932) );
  MUX2_X1 U17365 ( .A(n13933), .B(n13932), .S(n19894), .Z(n13934) );
  INV_X1 U17366 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n17361) );
  INV_X1 U17367 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16583) );
  OAI22_X2 U17368 ( .A1(n17361), .A2(n19336), .B1(n16583), .B2(n19338), .ZN(
        n19738) );
  AOI22_X1 U17369 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19335), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19334), .ZN(n19741) );
  INV_X1 U17370 ( .A(n19741), .ZN(n19791) );
  AOI22_X1 U17371 ( .A1(n19391), .A2(n19738), .B1(n19412), .B2(n19791), .ZN(
        n13941) );
  OAI21_X1 U17372 ( .B1(n13935), .B2(n19389), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13938) );
  INV_X1 U17373 ( .A(n13936), .ZN(n13937) );
  NAND2_X1 U17374 ( .A1(n13938), .A2(n13937), .ZN(n19390) );
  NOR2_X2 U17375 ( .A1(n19223), .A2(n19343), .ZN(n19790) );
  NOR2_X2 U17376 ( .A1(n13939), .A2(n19340), .ZN(n19789) );
  AOI22_X1 U17377 ( .A1(n19390), .A2(n19790), .B1(n19389), .B2(n19789), .ZN(
        n13940) );
  OAI211_X1 U17378 ( .C1(n19394), .C2(n14077), .A(n13941), .B(n13940), .ZN(
        P2_U3068) );
  AOI22_X1 U17379 ( .A1(n19391), .A2(n19767), .B1(n19412), .B2(n19637), .ZN(
        n13943) );
  AOI22_X1 U17380 ( .A1(n19390), .A2(n19760), .B1(n19759), .B2(n19389), .ZN(
        n13942) );
  OAI211_X1 U17381 ( .C1(n19394), .C2(n13944), .A(n13943), .B(n13942), .ZN(
        P2_U3064) );
  XNOR2_X1 U17382 ( .A(n9721), .B(n16233), .ZN(n13945) );
  XNOR2_X1 U17383 ( .A(n13946), .B(n13945), .ZN(n16243) );
  NAND2_X1 U17384 ( .A1(n16243), .A2(n11125), .ZN(n13950) );
  NOR2_X1 U17385 ( .A1(n16200), .A2(n20748), .ZN(n16240) );
  NOR2_X1 U17386 ( .A1(n16127), .A2(n13947), .ZN(n13948) );
  AOI211_X1 U17387 ( .C1(n16135), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16240), .B(n13948), .ZN(n13949) );
  OAI211_X1 U17388 ( .C1(n20129), .C2(n13951), .A(n13950), .B(n13949), .ZN(
        P1_U2990) );
  OAI21_X1 U17389 ( .B1(n13952), .B2(n13954), .A(n13953), .ZN(n14882) );
  AOI21_X1 U17390 ( .B1(n13956), .B2(n13955), .A(n9951), .ZN(n16220) );
  AOI22_X1 U17391 ( .A1(n16220), .A2(n16115), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n14623), .ZN(n13957) );
  OAI21_X1 U17392 ( .B1(n14882), .B2(n14628), .A(n13957), .ZN(P1_U2861) );
  INV_X1 U17393 ( .A(n19236), .ZN(n19219) );
  OR2_X1 U17394 ( .A1(n9808), .A2(n13959), .ZN(n13960) );
  AND2_X1 U17395 ( .A1(n13958), .A2(n13960), .ZN(n19010) );
  INV_X1 U17396 ( .A(n19010), .ZN(n13967) );
  NOR2_X2 U17397 ( .A1(n13963), .A2(n13961), .ZN(n19174) );
  NOR2_X2 U17398 ( .A1(n13963), .A2(n13962), .ZN(n19173) );
  AOI22_X1 U17399 ( .A1(n19174), .A2(BUF2_REG_17__SCAN_IN), .B1(n19173), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n13966) );
  AOI22_X1 U17400 ( .A1(n19172), .A2(n13964), .B1(n19231), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n13965) );
  OAI211_X1 U17401 ( .C1(n19180), .C2(n13967), .A(n13966), .B(n13965), .ZN(
        n13968) );
  AOI21_X1 U17402 ( .B1(n13969), .B2(n19219), .A(n13968), .ZN(n13970) );
  INV_X1 U17403 ( .A(n13970), .ZN(P2_U2902) );
  INV_X1 U17404 ( .A(n14878), .ZN(n13979) );
  AOI22_X1 U17405 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(n20041), .B1(n20024), 
        .B2(n16220), .ZN(n13971) );
  OAI211_X1 U17406 ( .C1(n19999), .C2(n13972), .A(n13971), .B(n20043), .ZN(
        n13978) );
  NAND2_X1 U17407 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n13974) );
  NOR2_X1 U17408 ( .A1(n13974), .A2(n14560), .ZN(n13976) );
  INV_X1 U17409 ( .A(n19995), .ZN(n13973) );
  AOI21_X1 U17410 ( .B1(n13974), .B2(n19996), .A(n13973), .ZN(n16114) );
  INV_X1 U17411 ( .A(n16114), .ZN(n13975) );
  MUX2_X1 U17412 ( .A(n13976), .B(n13975), .S(P1_REIP_REG_11__SCAN_IN), .Z(
        n13977) );
  AOI211_X1 U17413 ( .C1(n20039), .C2(n13979), .A(n13978), .B(n13977), .ZN(
        n13980) );
  OAI21_X1 U17414 ( .B1(n14571), .B2(n14882), .A(n13980), .ZN(P1_U2829) );
  INV_X1 U17415 ( .A(n14649), .ZN(n13981) );
  OAI222_X1 U17416 ( .A1(n14712), .A2(n14882), .B1(n14661), .B2(n13982), .C1(
        n14711), .C2(n13981), .ZN(P1_U2893) );
  AOI22_X1 U17417 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n11575), .B1(
        n11588), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13990) );
  AOI22_X1 U17418 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12262), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13989) );
  NAND2_X1 U17419 ( .A1(n11513), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n13984) );
  NAND2_X1 U17420 ( .A1(n11537), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n13983) );
  OAI211_X1 U17421 ( .C1(n14153), .C2(n13985), .A(n13984), .B(n13983), .ZN(
        n13986) );
  INV_X1 U17422 ( .A(n13986), .ZN(n13988) );
  AOI22_X1 U17423 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n14156), .B1(
        n14155), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13987) );
  NAND4_X1 U17424 ( .A1(n13990), .A2(n13989), .A3(n13988), .A4(n13987), .ZN(
        n13996) );
  AOI22_X1 U17425 ( .A1(n14162), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14161), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13994) );
  AOI22_X1 U17426 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9741), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13993) );
  AOI22_X1 U17427 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n11528), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13992) );
  NAND2_X1 U17428 ( .A1(n11523), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n13991) );
  NAND4_X1 U17429 ( .A1(n13994), .A2(n13993), .A3(n13992), .A4(n13991), .ZN(
        n13995) );
  NOR2_X1 U17430 ( .A1(n13996), .A2(n13995), .ZN(n16296) );
  AOI22_X1 U17431 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11528), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14002) );
  NAND2_X1 U17432 ( .A1(n13998), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n14001) );
  NAND2_X1 U17433 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n14000) );
  NAND2_X1 U17434 ( .A1(n11523), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n13999) );
  NAND4_X1 U17435 ( .A1(n14002), .A2(n14001), .A3(n14000), .A4(n13999), .ZN(
        n14005) );
  OAI22_X1 U17436 ( .A1(n14096), .A2(n14227), .B1(n14095), .B2(n14003), .ZN(
        n14004) );
  NOR2_X1 U17437 ( .A1(n14005), .A2(n14004), .ZN(n14015) );
  OAI22_X1 U17438 ( .A1(n14006), .A2(n14101), .B1(n14099), .B2(n14220), .ZN(
        n14011) );
  NAND2_X1 U17439 ( .A1(n11513), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n14008) );
  NAND2_X1 U17440 ( .A1(n11537), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n14007) );
  OAI211_X1 U17441 ( .C1(n14153), .C2(n14009), .A(n14008), .B(n14007), .ZN(
        n14010) );
  NOR2_X1 U17442 ( .A1(n14011), .A2(n14010), .ZN(n14014) );
  AOI22_X1 U17443 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n11575), .B1(
        n11588), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14013) );
  AOI22_X1 U17444 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12262), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14012) );
  NAND4_X1 U17445 ( .A1(n14015), .A2(n14014), .A3(n14013), .A4(n14012), .ZN(
        n14018) );
  INV_X1 U17446 ( .A(n14089), .ZN(n14017) );
  OAI21_X1 U17447 ( .B1(n14016), .B2(n14018), .A(n14017), .ZN(n15435) );
  OR2_X1 U17448 ( .A1(n14020), .A2(n14019), .ZN(n14022) );
  NAND2_X1 U17449 ( .A1(n14022), .A2(n14021), .ZN(n18997) );
  AOI22_X1 U17450 ( .A1(n19174), .A2(BUF2_REG_19__SCAN_IN), .B1(n19173), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n14025) );
  AOI22_X1 U17451 ( .A1(n19172), .A2(n14023), .B1(n19231), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n14024) );
  OAI211_X1 U17452 ( .C1(n19180), .C2(n18997), .A(n14025), .B(n14024), .ZN(
        n14026) );
  INV_X1 U17453 ( .A(n14026), .ZN(n14027) );
  OAI21_X1 U17454 ( .B1(n15435), .B2(n19236), .A(n14027), .ZN(P2_U2900) );
  AND3_X1 U17455 ( .A1(n18332), .A2(n17237), .A3(n14028), .ZN(n17209) );
  NAND2_X1 U17456 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17237), .ZN(n17238) );
  NOR2_X1 U17457 ( .A1(n16890), .A2(n17238), .ZN(n17212) );
  AOI21_X1 U17458 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17212), .A(
        P3_EBX_REG_15__SCAN_IN), .ZN(n14029) );
  NOR2_X1 U17459 ( .A1(n17209), .A2(n14029), .ZN(n14043) );
  AOI22_X1 U17460 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14034) );
  AOI22_X1 U17461 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14033) );
  AOI22_X1 U17462 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14032) );
  AOI22_X1 U17463 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14031) );
  NAND4_X1 U17464 ( .A1(n14034), .A2(n14033), .A3(n14032), .A4(n14031), .ZN(
        n14041) );
  AOI22_X1 U17465 ( .A1(n17256), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14039) );
  AOI22_X1 U17466 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14038) );
  AOI22_X1 U17467 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14037) );
  AOI22_X1 U17468 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14036) );
  NAND4_X1 U17469 ( .A1(n14039), .A2(n14038), .A3(n14037), .A4(n14036), .ZN(
        n14040) );
  NOR2_X1 U17470 ( .A1(n14041), .A2(n14040), .ZN(n17426) );
  INV_X1 U17471 ( .A(n17426), .ZN(n14042) );
  MUX2_X1 U17472 ( .A(n14043), .B(n14042), .S(n17338), .Z(P3_U2688) );
  OAI211_X1 U17473 ( .C1(n20949), .C2(n18736), .A(n9769), .B(n18780), .ZN(
        n18286) );
  NOR2_X1 U17474 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18286), .ZN(n14044) );
  NAND3_X1 U17475 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(P3_STATE2_REG_0__SCAN_IN), .ZN(n18885)
         );
  OAI21_X1 U17476 ( .B1(n14044), .B2(n18885), .A(n18445), .ZN(n18295) );
  INV_X1 U17477 ( .A(n18295), .ZN(n14046) );
  AOI22_X1 U17478 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .B1(n14045), .B2(n17872), .ZN(n18289) );
  NOR2_X1 U17479 ( .A1(n14046), .A2(n18289), .ZN(n14048) );
  NOR2_X1 U17480 ( .A1(n18887), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18336) );
  OR2_X1 U17481 ( .A1(n18336), .A2(n14046), .ZN(n18290) );
  OR2_X1 U17482 ( .A1(n18641), .A2(n18290), .ZN(n14047) );
  MUX2_X1 U17483 ( .A(n14048), .B(n14047), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  OR2_X1 U17484 ( .A1(n14679), .A2(n14049), .ZN(n14053) );
  NAND2_X1 U17485 ( .A1(n14661), .A2(n13061), .ZN(n14699) );
  INV_X1 U17486 ( .A(DATAI_14_), .ZN(n14051) );
  MUX2_X1 U17487 ( .A(n14051), .B(n14050), .S(n20130), .Z(n20069) );
  OAI22_X1 U17488 ( .A1(n14699), .A2(n20069), .B1(n14661), .B2(n13079), .ZN(
        n14052) );
  AOI21_X1 U17489 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n14701), .A(n14052), .ZN(
        n14055) );
  NOR2_X2 U17490 ( .A1(n14053), .A2(n20130), .ZN(n14702) );
  NAND2_X1 U17491 ( .A1(n14702), .A2(DATAI_30_), .ZN(n14054) );
  OAI211_X1 U17492 ( .C1(n10972), .C2(n14712), .A(n14055), .B(n14054), .ZN(
        P1_U2874) );
  INV_X1 U17493 ( .A(n14056), .ZN(n14057) );
  NAND2_X1 U17494 ( .A1(n14356), .A2(n14058), .ZN(n14061) );
  OR2_X1 U17495 ( .A1(n14396), .A2(n14059), .ZN(n14060) );
  NAND2_X1 U17496 ( .A1(n14061), .A2(n14060), .ZN(n14063) );
  AOI22_X1 U17497 ( .A1(n11167), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n14358), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14357) );
  INV_X1 U17498 ( .A(n14357), .ZN(n14062) );
  XNOR2_X1 U17499 ( .A(n14063), .B(n14062), .ZN(n14922) );
  INV_X1 U17500 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14064) );
  OAI222_X1 U17501 ( .A1(n14636), .A2(n14922), .B1(n14064), .B2(n16118), .C1(
        n10972), .C2(n14638), .ZN(P1_U2842) );
  INV_X1 U17502 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19339) );
  AOI22_X1 U17503 ( .A1(n14068), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n14067), .ZN(n14069) );
  AND2_X1 U17504 ( .A1(n14661), .A2(n14071), .ZN(n14072) );
  NAND2_X1 U17505 ( .A1(n14721), .A2(n14072), .ZN(n14074) );
  AOI22_X1 U17506 ( .A1(n14702), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14679), .ZN(n14073) );
  OAI211_X1 U17507 ( .C1(n14683), .C2(n19339), .A(n14074), .B(n14073), .ZN(
        P1_U2873) );
  AOI22_X1 U17508 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11588), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14082) );
  AOI22_X1 U17509 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12262), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14081) );
  NAND2_X1 U17510 ( .A1(n11513), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n14076) );
  NAND2_X1 U17511 ( .A1(n11537), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n14075) );
  OAI211_X1 U17512 ( .C1(n14153), .C2(n14077), .A(n14076), .B(n14075), .ZN(
        n14078) );
  INV_X1 U17513 ( .A(n14078), .ZN(n14080) );
  AOI22_X1 U17514 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n14156), .B1(
        n14155), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14079) );
  NAND4_X1 U17515 ( .A1(n14082), .A2(n14081), .A3(n14080), .A4(n14079), .ZN(
        n14088) );
  AOI22_X1 U17516 ( .A1(n14162), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14161), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14086) );
  AOI22_X1 U17517 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n11529), .B1(
        n9741), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14085) );
  AOI22_X1 U17518 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11528), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14084) );
  NAND2_X1 U17519 ( .A1(n11523), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14083) );
  NAND4_X1 U17520 ( .A1(n14086), .A2(n14085), .A3(n14084), .A4(n14083), .ZN(
        n14087) );
  OR2_X1 U17521 ( .A1(n14088), .A2(n14087), .ZN(n16291) );
  AOI22_X1 U17522 ( .A1(n11528), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14093) );
  NAND2_X1 U17523 ( .A1(n9741), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n14092) );
  NAND2_X1 U17524 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n14091) );
  NAND2_X1 U17525 ( .A1(n11523), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14090) );
  NAND4_X1 U17526 ( .A1(n14093), .A2(n14092), .A3(n14091), .A4(n14090), .ZN(
        n14098) );
  OAI22_X1 U17527 ( .A1(n14096), .A2(n14274), .B1(n14095), .B2(n14094), .ZN(
        n14097) );
  NOR2_X1 U17528 ( .A1(n14098), .A2(n14097), .ZN(n14110) );
  OAI22_X1 U17529 ( .A1(n14101), .A2(n14100), .B1(n14099), .B2(n14267), .ZN(
        n14106) );
  NAND2_X1 U17530 ( .A1(n11513), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n14103) );
  NAND2_X1 U17531 ( .A1(n11537), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n14102) );
  OAI211_X1 U17532 ( .C1(n14153), .C2(n14104), .A(n14103), .B(n14102), .ZN(
        n14105) );
  NOR2_X1 U17533 ( .A1(n14106), .A2(n14105), .ZN(n14109) );
  AOI22_X1 U17534 ( .A1(n11575), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11588), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14108) );
  AOI22_X1 U17535 ( .A1(n12262), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14107) );
  NAND4_X1 U17536 ( .A1(n14110), .A2(n14109), .A3(n14108), .A4(n14107), .ZN(
        n15427) );
  AOI22_X1 U17537 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n11575), .B1(
        n11588), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14118) );
  AOI22_X1 U17538 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12262), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14117) );
  NAND2_X1 U17539 ( .A1(n11513), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n14112) );
  NAND2_X1 U17540 ( .A1(n11537), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n14111) );
  OAI211_X1 U17541 ( .C1(n14153), .C2(n14113), .A(n14112), .B(n14111), .ZN(
        n14114) );
  INV_X1 U17542 ( .A(n14114), .ZN(n14116) );
  AOI22_X1 U17543 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n14156), .B1(
        n14155), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14115) );
  NAND4_X1 U17544 ( .A1(n14118), .A2(n14117), .A3(n14116), .A4(n14115), .ZN(
        n14124) );
  AOI22_X1 U17545 ( .A1(n14162), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14161), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14122) );
  AOI22_X1 U17546 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n11529), .B1(
        n9741), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14121) );
  AOI22_X1 U17547 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11528), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14120) );
  NAND2_X1 U17548 ( .A1(n11523), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n14119) );
  NAND4_X1 U17549 ( .A1(n14122), .A2(n14121), .A3(n14120), .A4(n14119), .ZN(
        n14123) );
  NOR2_X1 U17550 ( .A1(n14124), .A2(n14123), .ZN(n16288) );
  INV_X1 U17551 ( .A(n16288), .ZN(n14125) );
  NAND2_X1 U17552 ( .A1(n14126), .A2(n14125), .ZN(n14171) );
  AOI22_X1 U17553 ( .A1(n14326), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14307), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14139) );
  INV_X1 U17554 ( .A(n14127), .ZN(n14320) );
  INV_X1 U17555 ( .A(n14320), .ZN(n14312) );
  AOI22_X1 U17556 ( .A1(n14312), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14311), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14138) );
  AOI22_X1 U17557 ( .A1(n14325), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14265), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14137) );
  NAND2_X1 U17558 ( .A1(n11516), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14133) );
  INV_X1 U17559 ( .A(n14129), .ZN(n14132) );
  INV_X1 U17560 ( .A(n14130), .ZN(n14131) );
  NAND2_X1 U17561 ( .A1(n14132), .A2(n14131), .ZN(n14316) );
  OAI211_X1 U17562 ( .C1(n11499), .C2(n14134), .A(n14133), .B(n14316), .ZN(
        n14135) );
  INV_X1 U17563 ( .A(n14135), .ZN(n14136) );
  NAND4_X1 U17564 ( .A1(n14139), .A2(n14138), .A3(n14137), .A4(n14136), .ZN(
        n14150) );
  AOI22_X1 U17565 ( .A1(n14307), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11516), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14148) );
  INV_X1 U17566 ( .A(n14311), .ZN(n14275) );
  INV_X1 U17567 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14143) );
  INV_X1 U17568 ( .A(n14316), .ZN(n14293) );
  INV_X1 U17569 ( .A(n14265), .ZN(n14318) );
  OR2_X1 U17570 ( .A1(n14318), .A2(n14141), .ZN(n14142) );
  OAI211_X1 U17571 ( .C1(n14275), .C2(n14143), .A(n14293), .B(n14142), .ZN(
        n14144) );
  INV_X1 U17572 ( .A(n14144), .ZN(n14147) );
  AOI22_X1 U17573 ( .A1(n14326), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14325), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14146) );
  AOI22_X1 U17574 ( .A1(n14312), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14128), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14145) );
  NAND4_X1 U17575 ( .A1(n14148), .A2(n14147), .A3(n14146), .A4(n14145), .ZN(
        n14149) );
  AND2_X1 U17576 ( .A1(n14150), .A2(n14149), .ZN(n14189) );
  NAND2_X1 U17577 ( .A1(n19944), .A2(n14189), .ZN(n14170) );
  AOI22_X1 U17578 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n11588), .B1(
        n11575), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14160) );
  AOI22_X1 U17579 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12262), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14159) );
  INV_X1 U17580 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14319) );
  NAND2_X1 U17581 ( .A1(n11513), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n14152) );
  NAND2_X1 U17582 ( .A1(n11537), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n14151) );
  OAI211_X1 U17583 ( .C1(n14153), .C2(n14319), .A(n14152), .B(n14151), .ZN(
        n14154) );
  INV_X1 U17584 ( .A(n14154), .ZN(n14158) );
  AOI22_X1 U17585 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n14156), .B1(
        n14155), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14157) );
  NAND4_X1 U17586 ( .A1(n14160), .A2(n14159), .A3(n14158), .A4(n14157), .ZN(
        n14169) );
  AOI22_X1 U17587 ( .A1(n14162), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14161), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14167) );
  AOI22_X1 U17588 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n11529), .B1(
        n13998), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14166) );
  AOI22_X1 U17589 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n11528), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14165) );
  NAND2_X1 U17590 ( .A1(n11523), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14164) );
  NAND4_X1 U17591 ( .A1(n14167), .A2(n14166), .A3(n14165), .A4(n14164), .ZN(
        n14168) );
  OR2_X1 U17592 ( .A1(n14169), .A2(n14168), .ZN(n14190) );
  XNOR2_X1 U17593 ( .A(n14170), .B(n14190), .ZN(n14195) );
  INV_X1 U17594 ( .A(n14189), .ZN(n14193) );
  NOR2_X1 U17595 ( .A1(n19944), .A2(n14193), .ZN(n15464) );
  INV_X1 U17596 ( .A(n14171), .ZN(n16287) );
  AOI22_X1 U17597 ( .A1(n14326), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14307), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14179) );
  AOI22_X1 U17598 ( .A1(n14325), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n14265), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14178) );
  AOI22_X1 U17599 ( .A1(n14312), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14128), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14177) );
  NAND2_X1 U17600 ( .A1(n11516), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14173) );
  OAI211_X1 U17601 ( .C1(n14275), .C2(n14174), .A(n14316), .B(n14173), .ZN(
        n14175) );
  INV_X1 U17602 ( .A(n14175), .ZN(n14176) );
  NAND4_X1 U17603 ( .A1(n14179), .A2(n14178), .A3(n14177), .A4(n14176), .ZN(
        n14188) );
  AOI22_X1 U17604 ( .A1(n14326), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14307), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14186) );
  AOI22_X1 U17605 ( .A1(n14325), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14265), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14185) );
  AOI22_X1 U17606 ( .A1(n14312), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14128), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14184) );
  NAND2_X1 U17607 ( .A1(n11516), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n14180) );
  OAI211_X1 U17608 ( .C1(n14275), .C2(n14181), .A(n14293), .B(n14180), .ZN(
        n14182) );
  INV_X1 U17609 ( .A(n14182), .ZN(n14183) );
  NAND4_X1 U17610 ( .A1(n14186), .A2(n14185), .A3(n14184), .A4(n14183), .ZN(
        n14187) );
  AND2_X1 U17611 ( .A1(n14188), .A2(n14187), .ZN(n14192) );
  AND2_X1 U17612 ( .A1(n14190), .A2(n14189), .ZN(n14191) );
  NAND2_X1 U17613 ( .A1(n14191), .A2(n14192), .ZN(n14212) );
  OAI211_X1 U17614 ( .C1(n14192), .C2(n14191), .A(n14258), .B(n14212), .ZN(
        n15419) );
  NAND2_X1 U17615 ( .A1(n14263), .A2(n14192), .ZN(n15421) );
  NOR2_X1 U17616 ( .A1(n15421), .A2(n14193), .ZN(n14194) );
  AOI22_X1 U17617 ( .A1(n14326), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14307), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14202) );
  AOI22_X1 U17618 ( .A1(n14312), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14311), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14201) );
  AOI22_X1 U17619 ( .A1(n14325), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14265), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14200) );
  INV_X1 U17620 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14197) );
  NAND2_X1 U17621 ( .A1(n11516), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n14196) );
  OAI211_X1 U17622 ( .C1(n14197), .C2(n11499), .A(n14196), .B(n14293), .ZN(
        n14198) );
  INV_X1 U17623 ( .A(n14198), .ZN(n14199) );
  NAND4_X1 U17624 ( .A1(n14202), .A2(n14201), .A3(n14200), .A4(n14199), .ZN(
        n14211) );
  AOI22_X1 U17625 ( .A1(n14326), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14312), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14209) );
  AOI22_X1 U17626 ( .A1(n14325), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14265), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14208) );
  AOI22_X1 U17627 ( .A1(n14311), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14128), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14207) );
  INV_X1 U17628 ( .A(n14307), .ZN(n14322) );
  INV_X1 U17629 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14204) );
  NAND2_X1 U17630 ( .A1(n11516), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14203) );
  OAI211_X1 U17631 ( .C1(n14322), .C2(n14204), .A(n14316), .B(n14203), .ZN(
        n14205) );
  INV_X1 U17632 ( .A(n14205), .ZN(n14206) );
  NAND4_X1 U17633 ( .A1(n14209), .A2(n14208), .A3(n14207), .A4(n14206), .ZN(
        n14210) );
  NAND2_X1 U17634 ( .A1(n14211), .A2(n14210), .ZN(n14215) );
  NAND2_X1 U17635 ( .A1(n14212), .A2(n14215), .ZN(n14213) );
  NAND3_X1 U17636 ( .A1(n14238), .A2(n14258), .A3(n14213), .ZN(n14216) );
  NOR2_X1 U17637 ( .A1(n19944), .A2(n14215), .ZN(n15415) );
  INV_X1 U17638 ( .A(n14238), .ZN(n14235) );
  AOI22_X1 U17639 ( .A1(n14326), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14307), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14225) );
  AOI22_X1 U17640 ( .A1(n14325), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14265), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14224) );
  AOI22_X1 U17641 ( .A1(n14312), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14128), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14223) );
  NAND2_X1 U17642 ( .A1(n11516), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14219) );
  OAI211_X1 U17643 ( .C1(n14275), .C2(n14220), .A(n14316), .B(n14219), .ZN(
        n14221) );
  INV_X1 U17644 ( .A(n14221), .ZN(n14222) );
  NAND4_X1 U17645 ( .A1(n14225), .A2(n14224), .A3(n14223), .A4(n14222), .ZN(
        n14234) );
  AOI22_X1 U17646 ( .A1(n14326), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14307), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14232) );
  AOI22_X1 U17647 ( .A1(n14325), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14265), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14231) );
  AOI22_X1 U17648 ( .A1(n14312), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14128), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14230) );
  NAND2_X1 U17649 ( .A1(n11516), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n14226) );
  OAI211_X1 U17650 ( .C1(n14275), .C2(n14227), .A(n14293), .B(n14226), .ZN(
        n14228) );
  INV_X1 U17651 ( .A(n14228), .ZN(n14229) );
  NAND4_X1 U17652 ( .A1(n14232), .A2(n14231), .A3(n14230), .A4(n14229), .ZN(
        n14233) );
  AND2_X1 U17653 ( .A1(n14234), .A2(n14233), .ZN(n14240) );
  NAND2_X1 U17654 ( .A1(n14235), .A2(n14240), .ZN(n14242) );
  INV_X1 U17655 ( .A(n14240), .ZN(n14237) );
  AOI21_X1 U17656 ( .B1(n14238), .B2(n14237), .A(n14236), .ZN(n14239) );
  NAND2_X1 U17657 ( .A1(n14263), .A2(n14240), .ZN(n15410) );
  INV_X1 U17658 ( .A(n14242), .ZN(n14259) );
  AOI22_X1 U17659 ( .A1(n14326), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14312), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14248) );
  AOI22_X1 U17660 ( .A1(n14325), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14265), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14247) );
  AOI22_X1 U17661 ( .A1(n14311), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14128), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14246) );
  NAND2_X1 U17662 ( .A1(n11516), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14243) );
  OAI211_X1 U17663 ( .C1(n14322), .C2(n20934), .A(n14316), .B(n14243), .ZN(
        n14244) );
  INV_X1 U17664 ( .A(n14244), .ZN(n14245) );
  NAND4_X1 U17665 ( .A1(n14248), .A2(n14247), .A3(n14246), .A4(n14245), .ZN(
        n14257) );
  INV_X1 U17666 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n19554) );
  AOI22_X1 U17667 ( .A1(n14307), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11516), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14255) );
  INV_X1 U17668 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14250) );
  INV_X1 U17669 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n19669) );
  OR2_X1 U17670 ( .A1(n14318), .A2(n19669), .ZN(n14249) );
  OAI211_X1 U17671 ( .C1(n14275), .C2(n14250), .A(n14293), .B(n14249), .ZN(
        n14251) );
  INV_X1 U17672 ( .A(n14251), .ZN(n14254) );
  AOI22_X1 U17673 ( .A1(n14326), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14325), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14253) );
  AOI22_X1 U17674 ( .A1(n14312), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14128), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14252) );
  NAND4_X1 U17675 ( .A1(n14255), .A2(n14254), .A3(n14253), .A4(n14252), .ZN(
        n14256) );
  AND2_X1 U17676 ( .A1(n14257), .A2(n14256), .ZN(n14262) );
  NAND2_X1 U17677 ( .A1(n14259), .A2(n14262), .ZN(n15395) );
  OAI211_X1 U17678 ( .C1(n14259), .C2(n14262), .A(n15395), .B(n14258), .ZN(
        n14260) );
  INV_X1 U17679 ( .A(n14260), .ZN(n14261) );
  NAND2_X1 U17680 ( .A1(n14263), .A2(n14262), .ZN(n15402) );
  INV_X1 U17681 ( .A(n14264), .ZN(n14283) );
  AOI22_X1 U17682 ( .A1(n14326), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14307), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14272) );
  AOI22_X1 U17683 ( .A1(n14325), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14265), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14271) );
  AOI22_X1 U17684 ( .A1(n14312), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14128), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14270) );
  NAND2_X1 U17685 ( .A1(n11516), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n14266) );
  OAI211_X1 U17686 ( .C1(n14275), .C2(n14267), .A(n14316), .B(n14266), .ZN(
        n14268) );
  INV_X1 U17687 ( .A(n14268), .ZN(n14269) );
  NAND4_X1 U17688 ( .A1(n14272), .A2(n14271), .A3(n14270), .A4(n14269), .ZN(
        n14282) );
  AOI22_X1 U17689 ( .A1(n14326), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14307), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14280) );
  AOI22_X1 U17690 ( .A1(n14325), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14265), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14279) );
  AOI22_X1 U17691 ( .A1(n14312), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14128), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14278) );
  NAND2_X1 U17692 ( .A1(n11516), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n14273) );
  OAI211_X1 U17693 ( .C1(n14275), .C2(n14274), .A(n14293), .B(n14273), .ZN(
        n14276) );
  INV_X1 U17694 ( .A(n14276), .ZN(n14277) );
  NAND4_X1 U17695 ( .A1(n14280), .A2(n14279), .A3(n14278), .A4(n14277), .ZN(
        n14281) );
  AND2_X1 U17696 ( .A1(n14282), .A2(n14281), .ZN(n15396) );
  NAND2_X1 U17697 ( .A1(n19944), .A2(n15396), .ZN(n14284) );
  NOR2_X1 U17698 ( .A1(n15395), .A2(n14284), .ZN(n14304) );
  AOI22_X1 U17699 ( .A1(n14326), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14311), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14291) );
  AOI22_X1 U17700 ( .A1(n14325), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11516), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14290) );
  AOI22_X1 U17701 ( .A1(n14307), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14128), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14289) );
  OR2_X1 U17702 ( .A1(n14318), .A2(n14285), .ZN(n14286) );
  OAI211_X1 U17703 ( .C1(n14320), .C2(n14113), .A(n14316), .B(n14286), .ZN(
        n14287) );
  INV_X1 U17704 ( .A(n14287), .ZN(n14288) );
  NAND4_X1 U17705 ( .A1(n14291), .A2(n14290), .A3(n14289), .A4(n14288), .ZN(
        n14302) );
  AOI22_X1 U17706 ( .A1(n14326), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14307), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14300) );
  AOI22_X1 U17707 ( .A1(n14311), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14292), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14299) );
  AOI22_X1 U17708 ( .A1(n14312), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14325), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14298) );
  NAND2_X1 U17709 ( .A1(n11516), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n14294) );
  OAI211_X1 U17710 ( .C1(n11499), .C2(n14295), .A(n14294), .B(n14293), .ZN(
        n14296) );
  INV_X1 U17711 ( .A(n14296), .ZN(n14297) );
  NAND4_X1 U17712 ( .A1(n14300), .A2(n14299), .A3(n14298), .A4(n14297), .ZN(
        n14301) );
  AND2_X1 U17713 ( .A1(n14302), .A2(n14301), .ZN(n14303) );
  NAND2_X1 U17714 ( .A1(n14304), .A2(n14303), .ZN(n14305) );
  OAI21_X1 U17715 ( .B1(n14304), .B2(n14303), .A(n14305), .ZN(n14345) );
  INV_X1 U17716 ( .A(n14305), .ZN(n14306) );
  NOR2_X1 U17717 ( .A1(n14343), .A2(n14306), .ZN(n14334) );
  AOI22_X1 U17718 ( .A1(n14326), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14128), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14309) );
  NAND2_X1 U17719 ( .A1(n14307), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n14308) );
  OAI211_X1 U17720 ( .C1(n14310), .C2(n19564), .A(n14309), .B(n14308), .ZN(
        n14332) );
  INV_X1 U17721 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14315) );
  AOI22_X1 U17722 ( .A1(n14312), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14311), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14314) );
  AOI21_X1 U17723 ( .B1(n14265), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n14316), .ZN(n14313) );
  OAI211_X1 U17724 ( .C1(n13266), .C2(n14315), .A(n14314), .B(n14313), .ZN(
        n14331) );
  INV_X1 U17725 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14317) );
  OAI21_X1 U17726 ( .B1(n14318), .B2(n14317), .A(n14316), .ZN(n14324) );
  INV_X1 U17727 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14321) );
  OAI22_X1 U17728 ( .A1(n14322), .A2(n14321), .B1(n14320), .B2(n14319), .ZN(
        n14323) );
  AOI211_X1 U17729 ( .C1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .C2(n14311), .A(
        n14324), .B(n14323), .ZN(n14329) );
  AOI22_X1 U17730 ( .A1(n14325), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11516), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14328) );
  AOI22_X1 U17731 ( .A1(n14326), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14128), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14327) );
  NAND3_X1 U17732 ( .A1(n14329), .A2(n14328), .A3(n14327), .ZN(n14330) );
  OAI21_X1 U17733 ( .B1(n14332), .B2(n14331), .A(n14330), .ZN(n14333) );
  XNOR2_X1 U17734 ( .A(n14334), .B(n14333), .ZN(n14342) );
  AOI22_X1 U17735 ( .A1(n19174), .A2(BUF2_REG_30__SCAN_IN), .B1(n19173), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n14336) );
  AOI22_X1 U17736 ( .A1(n19172), .A2(n19184), .B1(n19231), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n14335) );
  OAI211_X1 U17737 ( .C1(n14337), .C2(n19180), .A(n14336), .B(n14335), .ZN(
        n14338) );
  INV_X1 U17738 ( .A(n14338), .ZN(n14339) );
  OAI21_X1 U17739 ( .B1(n14342), .B2(n19236), .A(n14339), .ZN(P2_U2889) );
  NOR2_X1 U17740 ( .A1(n15497), .A2(n19161), .ZN(n14340) );
  AOI21_X1 U17741 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n19161), .A(n14340), .ZN(
        n14341) );
  OAI21_X1 U17742 ( .B1(n14342), .B2(n19165), .A(n14341), .ZN(P2_U2857) );
  NAND2_X1 U17743 ( .A1(n14344), .A2(n14345), .ZN(n15391) );
  NAND2_X1 U17744 ( .A1(n15391), .A2(n19219), .ZN(n14352) );
  INV_X1 U17745 ( .A(n9778), .ZN(n14347) );
  INV_X1 U17746 ( .A(n16280), .ZN(n15647) );
  INV_X1 U17747 ( .A(n19172), .ZN(n15458) );
  OAI22_X1 U17748 ( .A1(n15458), .A2(n19187), .B1(n19205), .B2(n14348), .ZN(
        n14349) );
  AOI21_X1 U17749 ( .B1(n19232), .B2(n15647), .A(n14349), .ZN(n14351) );
  AOI22_X1 U17750 ( .A1(n19174), .A2(BUF2_REG_29__SCAN_IN), .B1(n19173), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14350) );
  OAI211_X1 U17751 ( .C1(n14343), .C2(n14352), .A(n14351), .B(n14350), .ZN(
        P2_U2890) );
  NAND2_X1 U17752 ( .A1(n14353), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n14355)
         );
  NAND3_X1 U17753 ( .A1(n14355), .A2(n14354), .A3(n19967), .ZN(P1_U2801) );
  MUX2_X1 U17754 ( .A(n14357), .B(n11224), .S(n14356), .Z(n14360) );
  AOI22_X1 U17755 ( .A1(n11167), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n14358), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14359) );
  NAND2_X1 U17756 ( .A1(n14721), .A2(n20018), .ZN(n14375) );
  INV_X1 U17757 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20776) );
  INV_X1 U17758 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20753) );
  NAND3_X1 U17759 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(P1_REIP_REG_9__SCAN_IN), .ZN(n14561) );
  NOR2_X1 U17760 ( .A1(n20753), .A2(n14561), .ZN(n16094) );
  NAND3_X1 U17761 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(n16094), .ZN(n14500) );
  NAND3_X1 U17762 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14513) );
  NOR4_X1 U17763 ( .A1(n14362), .A2(n14500), .A3(n14361), .A4(n14513), .ZN(
        n14364) );
  AND3_X1 U17764 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(P1_REIP_REG_20__SCAN_IN), .ZN(n14363) );
  AND2_X1 U17765 ( .A1(n14364), .A2(n14363), .ZN(n14466) );
  NAND2_X1 U17766 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n14467) );
  INV_X1 U17767 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14785) );
  NOR2_X1 U17768 ( .A1(n14467), .A2(n14785), .ZN(n14365) );
  AND2_X1 U17769 ( .A1(n14466), .A2(n14365), .ZN(n14452) );
  NAND3_X1 U17770 ( .A1(n14452), .A2(P1_REIP_REG_25__SCAN_IN), .A3(
        P1_REIP_REG_24__SCAN_IN), .ZN(n14423) );
  NOR2_X1 U17771 ( .A1(n20776), .A2(n14423), .ZN(n14411) );
  NAND3_X1 U17772 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .A3(n14411), .ZN(n14370) );
  INV_X1 U17773 ( .A(n14370), .ZN(n14366) );
  AND2_X1 U17774 ( .A1(n14585), .A2(n14366), .ZN(n14386) );
  NAND2_X1 U17775 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14371) );
  INV_X1 U17776 ( .A(n14371), .ZN(n14367) );
  NAND2_X1 U17777 ( .A1(n14386), .A2(n14367), .ZN(n14368) );
  AND2_X1 U17778 ( .A1(n19996), .A2(n14368), .ZN(n14378) );
  INV_X1 U17779 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14596) );
  OAI22_X1 U17780 ( .A1(n20000), .A2(n14596), .B1(n14369), .B2(n19999), .ZN(
        n14373) );
  OR2_X1 U17781 ( .A1(n14590), .A2(n14370), .ZN(n14388) );
  NOR3_X1 U17782 ( .A1(n14388), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14371), 
        .ZN(n14372) );
  AOI211_X1 U17783 ( .C1(n14378), .C2(P1_REIP_REG_31__SCAN_IN), .A(n14373), 
        .B(n14372), .ZN(n14374) );
  OAI211_X1 U17784 ( .C1(n14883), .C2(n20053), .A(n14375), .B(n14374), .ZN(
        P1_U2809) );
  NAND2_X1 U17785 ( .A1(n14376), .A2(n20018), .ZN(n14385) );
  INV_X1 U17786 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20783) );
  INV_X1 U17787 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14377) );
  OAI21_X1 U17788 ( .B1(n14388), .B2(n20783), .A(n14377), .ZN(n14379) );
  NAND2_X1 U17789 ( .A1(n14379), .A2(n14378), .ZN(n14381) );
  AOI22_X1 U17790 ( .A1(n20041), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20042), .ZN(n14380) );
  NAND2_X1 U17791 ( .A1(n14381), .A2(n14380), .ZN(n14382) );
  AOI21_X1 U17792 ( .B1(n20039), .B2(n14383), .A(n14382), .ZN(n14384) );
  OAI211_X1 U17793 ( .C1(n14922), .C2(n20053), .A(n14385), .B(n14384), .ZN(
        P1_U2810) );
  NAND2_X1 U17794 ( .A1(n14729), .A2(n20018), .ZN(n14392) );
  NOR2_X1 U17795 ( .A1(n16095), .A2(n14386), .ZN(n14399) );
  AOI22_X1 U17796 ( .A1(n20041), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20042), .ZN(n14387) );
  OAI21_X1 U17797 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(n14388), .A(n14387), 
        .ZN(n14390) );
  NOR2_X1 U17798 ( .A1(n20030), .A2(n14727), .ZN(n14389) );
  AOI211_X1 U17799 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(n14399), .A(n14390), 
        .B(n14389), .ZN(n14391) );
  OAI211_X1 U17800 ( .C1(n20053), .C2(n14932), .A(n14392), .B(n14391), .ZN(
        P1_U2811) );
  OAI21_X1 U17801 ( .B1(n14393), .B2(n14394), .A(n11135), .ZN(n14744) );
  OR2_X1 U17802 ( .A1(n14408), .A2(n14395), .ZN(n14397) );
  INV_X1 U17803 ( .A(n14733), .ZN(n14403) );
  AOI22_X1 U17804 ( .A1(n20041), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20042), .ZN(n14402) );
  NAND2_X1 U17805 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n14411), .ZN(n14398) );
  NOR2_X1 U17806 ( .A1(n14590), .A2(n14398), .ZN(n14400) );
  OAI21_X1 U17807 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n14400), .A(n14399), 
        .ZN(n14401) );
  OAI211_X1 U17808 ( .C1(n20030), .C2(n14403), .A(n14402), .B(n14401), .ZN(
        n14404) );
  AOI21_X1 U17809 ( .B1(n14941), .B2(n20024), .A(n14404), .ZN(n14405) );
  OAI21_X1 U17810 ( .B1(n14744), .B2(n14571), .A(n14405), .ZN(P1_U2812) );
  AOI21_X1 U17811 ( .B1(n14434), .B2(n14422), .A(n14406), .ZN(n14407) );
  OR2_X1 U17812 ( .A1(n14408), .A2(n14407), .ZN(n14956) );
  AOI21_X1 U17813 ( .B1(n14410), .B2(n14420), .A(n14393), .ZN(n14750) );
  NAND2_X1 U17814 ( .A1(n14750), .A2(n20018), .ZN(n14418) );
  AOI21_X1 U17815 ( .B1(n14411), .B2(n14585), .A(n16095), .ZN(n14426) );
  INV_X1 U17816 ( .A(n14411), .ZN(n14412) );
  NOR3_X1 U17817 ( .A1(n14590), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14412), 
        .ZN(n14413) );
  AOI21_X1 U17818 ( .B1(n20042), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14413), .ZN(n14414) );
  OAI21_X1 U17819 ( .B1(n20000), .B2(n14598), .A(n14414), .ZN(n14416) );
  NOR2_X1 U17820 ( .A1(n20030), .A2(n14748), .ZN(n14415) );
  AOI211_X1 U17821 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14426), .A(n14416), 
        .B(n14415), .ZN(n14417) );
  OAI211_X1 U17822 ( .C1(n20053), .C2(n14956), .A(n14418), .B(n14417), .ZN(
        P1_U2813) );
  XOR2_X1 U17823 ( .A(n14422), .B(n14434), .Z(n14973) );
  INV_X1 U17824 ( .A(n14760), .ZN(n14429) );
  NOR2_X1 U17825 ( .A1(n19999), .A2(n14756), .ZN(n14425) );
  NOR3_X1 U17826 ( .A1(n14590), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n14423), 
        .ZN(n14424) );
  AOI211_X1 U17827 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n20041), .A(n14425), .B(
        n14424), .ZN(n14428) );
  NAND2_X1 U17828 ( .A1(n14426), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14427) );
  OAI211_X1 U17829 ( .C1(n20030), .C2(n14429), .A(n14428), .B(n14427), .ZN(
        n14430) );
  AOI21_X1 U17830 ( .B1(n14973), .B2(n20024), .A(n14430), .ZN(n14431) );
  OAI21_X1 U17831 ( .B1(n14757), .B2(n14571), .A(n14431), .ZN(P1_U2814) );
  NOR2_X1 U17832 ( .A1(n14450), .A2(n14432), .ZN(n14433) );
  OR2_X1 U17833 ( .A1(n14434), .A2(n14433), .ZN(n14980) );
  AOI21_X1 U17834 ( .B1(n14437), .B2(n14436), .A(n14419), .ZN(n14771) );
  NAND2_X1 U17835 ( .A1(n14771), .A2(n20018), .ZN(n14447) );
  INV_X1 U17836 ( .A(n14769), .ZN(n14445) );
  INV_X1 U17837 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20775) );
  NAND2_X1 U17838 ( .A1(n14452), .A2(n20775), .ZN(n14438) );
  NAND2_X1 U17839 ( .A1(n14438), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14439) );
  OAI21_X1 U17840 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(P1_REIP_REG_24__SCAN_IN), 
        .A(n14439), .ZN(n14443) );
  OR2_X1 U17841 ( .A1(n14590), .A2(n14452), .ZN(n14440) );
  NAND2_X1 U17842 ( .A1(n14440), .A2(n14585), .ZN(n14468) );
  NAND2_X1 U17843 ( .A1(n14468), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14442) );
  AOI22_X1 U17844 ( .A1(n20041), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20042), .ZN(n14441) );
  OAI211_X1 U17845 ( .C1(n14590), .C2(n14443), .A(n14442), .B(n14441), .ZN(
        n14444) );
  AOI21_X1 U17846 ( .B1(n20039), .B2(n14445), .A(n14444), .ZN(n14446) );
  OAI211_X1 U17847 ( .C1(n14980), .C2(n20053), .A(n14447), .B(n14446), .ZN(
        P1_U2815) );
  OAI21_X1 U17848 ( .B1(n14448), .B2(n14449), .A(n14436), .ZN(n14782) );
  AOI21_X1 U17849 ( .B1(n14451), .B2(n14463), .A(n14450), .ZN(n14992) );
  INV_X1 U17850 ( .A(n14992), .ZN(n14457) );
  INV_X1 U17851 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20773) );
  NAND3_X1 U17852 ( .A1(n14578), .A2(n14452), .A3(n20773), .ZN(n14454) );
  NAND2_X1 U17853 ( .A1(n20041), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n14453) );
  OAI211_X1 U17854 ( .C1(n19999), .C2(n14773), .A(n14454), .B(n14453), .ZN(
        n14455) );
  AOI21_X1 U17855 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n14468), .A(n14455), 
        .ZN(n14456) );
  OAI21_X1 U17856 ( .B1(n14457), .B2(n20053), .A(n14456), .ZN(n14458) );
  AOI21_X1 U17857 ( .B1(n14775), .B2(n20039), .A(n14458), .ZN(n14459) );
  OAI21_X1 U17858 ( .B1(n14782), .B2(n14571), .A(n14459), .ZN(P1_U2816) );
  AOI21_X1 U17859 ( .B1(n14462), .B2(n14461), .A(n14448), .ZN(n14789) );
  INV_X1 U17860 ( .A(n14789), .ZN(n14668) );
  INV_X1 U17861 ( .A(n14787), .ZN(n14473) );
  INV_X1 U17862 ( .A(n14463), .ZN(n14464) );
  AOI21_X1 U17863 ( .B1(n14465), .B2(n9770), .A(n14464), .ZN(n14602) );
  INV_X1 U17864 ( .A(n14602), .ZN(n15000) );
  AOI22_X1 U17865 ( .A1(n20041), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20042), .ZN(n14471) );
  INV_X1 U17866 ( .A(n14466), .ZN(n14480) );
  OR2_X1 U17867 ( .A1(n14590), .A2(n14480), .ZN(n14491) );
  NOR2_X1 U17868 ( .A1(n14491), .A2(n14467), .ZN(n14469) );
  OAI21_X1 U17869 ( .B1(n14469), .B2(P1_REIP_REG_23__SCAN_IN), .A(n14468), 
        .ZN(n14470) );
  OAI211_X1 U17870 ( .C1(n15000), .C2(n20053), .A(n14471), .B(n14470), .ZN(
        n14472) );
  AOI21_X1 U17871 ( .B1(n14473), .B2(n20039), .A(n14472), .ZN(n14474) );
  OAI21_X1 U17872 ( .B1(n14668), .B2(n14571), .A(n14474), .ZN(P1_U2817) );
  OAI21_X1 U17873 ( .B1(n14475), .B2(n14476), .A(n14461), .ZN(n14799) );
  INV_X1 U17874 ( .A(n14477), .ZN(n14478) );
  OAI21_X1 U17875 ( .B1(n9758), .B2(n14478), .A(n9770), .ZN(n16158) );
  AOI21_X1 U17876 ( .B1(n14578), .B2(n14480), .A(n14479), .ZN(n14503) );
  OAI21_X1 U17877 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n14590), .A(n14503), 
        .ZN(n14483) );
  INV_X1 U17878 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14604) );
  OAI22_X1 U17879 ( .A1(n20000), .A2(n14604), .B1(n14791), .B2(n19999), .ZN(
        n14482) );
  INV_X1 U17880 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20768) );
  NOR3_X1 U17881 ( .A1(n14491), .A2(P1_REIP_REG_22__SCAN_IN), .A3(n20768), 
        .ZN(n14481) );
  AOI211_X1 U17882 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(n14483), .A(n14482), 
        .B(n14481), .ZN(n14484) );
  OAI21_X1 U17883 ( .B1(n16158), .B2(n20053), .A(n14484), .ZN(n14485) );
  AOI21_X1 U17884 ( .B1(n14793), .B2(n20039), .A(n14485), .ZN(n14486) );
  OAI21_X1 U17885 ( .B1(n14799), .B2(n14571), .A(n14486), .ZN(P1_U2818) );
  AOI21_X1 U17886 ( .B1(n14488), .B2(n14487), .A(n14475), .ZN(n14807) );
  NAND2_X1 U17887 ( .A1(n14807), .A2(n20018), .ZN(n14495) );
  AOI21_X1 U17888 ( .B1(n14489), .B2(n9792), .A(n9758), .ZN(n15016) );
  NOR2_X1 U17889 ( .A1(n14503), .A2(n20768), .ZN(n14493) );
  AOI22_X1 U17890 ( .A1(n20041), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20042), .ZN(n14490) );
  OAI21_X1 U17891 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n14491), .A(n14490), 
        .ZN(n14492) );
  AOI211_X1 U17892 ( .C1(n15016), .C2(n20024), .A(n14493), .B(n14492), .ZN(
        n14494) );
  OAI211_X1 U17893 ( .C1(n20030), .C2(n14805), .A(n14495), .B(n14494), .ZN(
        P1_U2819) );
  XOR2_X1 U17894 ( .A(n14497), .B(n14496), .Z(n14816) );
  INV_X1 U17895 ( .A(n14816), .ZN(n14686) );
  OAI21_X1 U17896 ( .B1(n14519), .B2(n14498), .A(n9792), .ZN(n15019) );
  AOI22_X1 U17897 ( .A1(n20041), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20042), .ZN(n14499) );
  OAI21_X1 U17898 ( .B1(n15019), .B2(n20053), .A(n14499), .ZN(n14506) );
  INV_X1 U17899 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20763) );
  NAND2_X1 U17900 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n14502) );
  INV_X1 U17901 ( .A(n14500), .ZN(n14512) );
  NAND2_X1 U17902 ( .A1(n14512), .A2(n14501), .ZN(n14539) );
  NOR2_X1 U17903 ( .A1(n14502), .A2(n14539), .ZN(n16084) );
  NAND2_X1 U17904 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n16084), .ZN(n14511) );
  NOR2_X1 U17905 ( .A1(n20763), .A2(n14511), .ZN(n14510) );
  AOI21_X1 U17906 ( .B1(n14510), .B2(P1_REIP_REG_19__SCAN_IN), .A(
        P1_REIP_REG_20__SCAN_IN), .ZN(n14504) );
  NOR2_X1 U17907 ( .A1(n14504), .A2(n14503), .ZN(n14505) );
  AOI211_X1 U17908 ( .C1(n20039), .C2(n14813), .A(n14506), .B(n14505), .ZN(
        n14507) );
  OAI21_X1 U17909 ( .B1(n14686), .B2(n14571), .A(n14507), .ZN(P1_U2820) );
  AOI21_X1 U17910 ( .B1(n14509), .B2(n14508), .A(n14496), .ZN(n16123) );
  INV_X1 U17911 ( .A(n16123), .ZN(n14691) );
  INV_X1 U17912 ( .A(n14510), .ZN(n14516) );
  NOR2_X1 U17913 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n14511), .ZN(n14532) );
  OAI21_X1 U17914 ( .B1(n14512), .B2(n16095), .A(n19995), .ZN(n14567) );
  AOI21_X1 U17915 ( .B1(n14513), .B2(n19996), .A(n14567), .ZN(n14514) );
  INV_X1 U17916 ( .A(n14514), .ZN(n16083) );
  NOR2_X1 U17917 ( .A1(n14532), .A2(n16083), .ZN(n14515) );
  MUX2_X1 U17918 ( .A(n14516), .B(n14515), .S(P1_REIP_REG_19__SCAN_IN), .Z(
        n14523) );
  AND2_X1 U17919 ( .A1(n14528), .A2(n14517), .ZN(n14518) );
  NOR2_X1 U17920 ( .A1(n14519), .A2(n14518), .ZN(n16166) );
  AOI22_X1 U17921 ( .A1(P1_EBX_REG_19__SCAN_IN), .A2(n20041), .B1(n20024), 
        .B2(n16166), .ZN(n14520) );
  OAI21_X1 U17922 ( .B1(n16126), .B2(n20030), .A(n14520), .ZN(n14521) );
  AOI211_X1 U17923 ( .C1(n20042), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n19987), .B(n14521), .ZN(n14522) );
  OAI211_X1 U17924 ( .C1(n14691), .C2(n14571), .A(n14523), .B(n14522), .ZN(
        P1_U2821) );
  OAI21_X1 U17925 ( .B1(n14524), .B2(n14525), .A(n14508), .ZN(n14824) );
  NAND2_X1 U17926 ( .A1(n14619), .A2(n14526), .ZN(n14527) );
  NAND2_X1 U17927 ( .A1(n14528), .A2(n14527), .ZN(n15046) );
  AOI21_X1 U17928 ( .B1(n20042), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n19987), .ZN(n14530) );
  AOI22_X1 U17929 ( .A1(n14820), .A2(n20039), .B1(P1_EBX_REG_18__SCAN_IN), 
        .B2(n20041), .ZN(n14529) );
  OAI211_X1 U17930 ( .C1(n20053), .C2(n15046), .A(n14530), .B(n14529), .ZN(
        n14531) );
  AOI211_X1 U17931 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n16083), .A(n14532), 
        .B(n14531), .ZN(n14533) );
  OAI21_X1 U17932 ( .B1(n14824), .B2(n14571), .A(n14533), .ZN(P1_U2822) );
  OR2_X1 U17933 ( .A1(n14534), .A2(n14546), .ZN(n14544) );
  AOI21_X1 U17934 ( .B1(n14536), .B2(n14544), .A(n14535), .ZN(n14833) );
  INV_X1 U17935 ( .A(n14833), .ZN(n14705) );
  NOR2_X1 U17936 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n14539), .ZN(n14552) );
  OAI21_X1 U17937 ( .B1(n14552), .B2(n14567), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n14543) );
  XNOR2_X1 U17938 ( .A(n14616), .B(n14614), .ZN(n16178) );
  AOI22_X1 U17939 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(n20041), .B1(n20024), 
        .B2(n16178), .ZN(n14537) );
  OAI211_X1 U17940 ( .C1(n19999), .C2(n14538), .A(n14537), .B(n20043), .ZN(
        n14541) );
  INV_X1 U17941 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20759) );
  NOR3_X1 U17942 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n20759), .A3(n14539), 
        .ZN(n14540) );
  AOI211_X1 U17943 ( .C1(n20039), .C2(n14828), .A(n14541), .B(n14540), .ZN(
        n14542) );
  OAI211_X1 U17944 ( .C1(n14705), .C2(n14571), .A(n14543), .B(n14542), .ZN(
        P1_U2824) );
  INV_X1 U17945 ( .A(n14544), .ZN(n14545) );
  AOI21_X1 U17946 ( .B1(n14546), .B2(n14534), .A(n14545), .ZN(n14847) );
  NAND2_X1 U17947 ( .A1(n14847), .A2(n20018), .ZN(n14556) );
  NAND2_X1 U17948 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n14567), .ZN(n14555) );
  INV_X1 U17949 ( .A(n14563), .ZN(n14547) );
  AOI21_X1 U17950 ( .B1(n14548), .B2(n14547), .A(n14616), .ZN(n16186) );
  AOI22_X1 U17951 ( .A1(P1_EBX_REG_15__SCAN_IN), .A2(n20041), .B1(n20024), 
        .B2(n16186), .ZN(n14549) );
  OAI211_X1 U17952 ( .C1(n19999), .C2(n14550), .A(n14549), .B(n20043), .ZN(
        n14551) );
  AOI21_X1 U17953 ( .B1(n14846), .B2(n20039), .A(n14551), .ZN(n14554) );
  INV_X1 U17954 ( .A(n14552), .ZN(n14553) );
  NAND4_X1 U17955 ( .A1(n14556), .A2(n14555), .A3(n14554), .A4(n14553), .ZN(
        P1_U2825) );
  INV_X1 U17956 ( .A(n14534), .ZN(n14558) );
  AOI21_X1 U17957 ( .B1(n14559), .B2(n14557), .A(n14558), .ZN(n14859) );
  INV_X1 U17958 ( .A(n14859), .ZN(n14708) );
  INV_X1 U17959 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20755) );
  NOR2_X1 U17960 ( .A1(n14561), .A2(n14560), .ZN(n16104) );
  NAND2_X1 U17961 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n16104), .ZN(n16099) );
  INV_X1 U17962 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20756) );
  OAI21_X1 U17963 ( .B1(n20755), .B2(n16099), .A(n20756), .ZN(n14566) );
  AND2_X1 U17964 ( .A1(n14633), .A2(n14562), .ZN(n14564) );
  OR2_X1 U17965 ( .A1(n14564), .A2(n14563), .ZN(n16193) );
  OAI22_X1 U17966 ( .A1(n20875), .A2(n19999), .B1(n20053), .B2(n16193), .ZN(
        n14565) );
  AOI211_X1 U17967 ( .C1(n14567), .C2(n14566), .A(n19987), .B(n14565), .ZN(
        n14570) );
  INV_X1 U17968 ( .A(n14857), .ZN(n14568) );
  AOI22_X1 U17969 ( .A1(n20039), .A2(n14568), .B1(n20041), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n14569) );
  OAI211_X1 U17970 ( .C1(n14708), .C2(n14571), .A(n14570), .B(n14569), .ZN(
        P1_U2826) );
  NAND2_X1 U17971 ( .A1(n20406), .A2(n20037), .ZN(n14576) );
  OAI22_X1 U17972 ( .A1(n14573), .A2(n19999), .B1(n14572), .B2(n20030), .ZN(
        n14574) );
  AOI21_X1 U17973 ( .B1(n20041), .B2(P1_EBX_REG_3__SCAN_IN), .A(n14574), .ZN(
        n14575) );
  OAI211_X1 U17974 ( .C1(n14577), .C2(n20053), .A(n14576), .B(n14575), .ZN(
        n14581) );
  NAND3_X1 U17975 ( .A1(n14578), .A2(P1_REIP_REG_1__SCAN_IN), .A3(
        P1_REIP_REG_2__SCAN_IN), .ZN(n14579) );
  AOI211_X1 U17976 ( .C1(n20739), .C2(n14579), .A(n20040), .B(n16095), .ZN(
        n14580) );
  AOI211_X1 U17977 ( .C1(n14582), .C2(n20048), .A(n14581), .B(n14580), .ZN(
        n14583) );
  INV_X1 U17978 ( .A(n14583), .ZN(P1_U2837) );
  INV_X1 U17979 ( .A(n13182), .ZN(n20139) );
  AOI22_X1 U17980 ( .A1(n20737), .A2(P1_REIP_REG_1__SCAN_IN), .B1(n20734), 
        .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n14591) );
  OAI22_X1 U17981 ( .A1(n14584), .A2(n20030), .B1(n20053), .B2(n20106), .ZN(
        n14587) );
  NOR2_X1 U17982 ( .A1(n14585), .A2(n20737), .ZN(n14586) );
  AOI211_X1 U17983 ( .C1(n20042), .C2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n14587), .B(n14586), .ZN(n14589) );
  NAND2_X1 U17984 ( .A1(n20041), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n14588) );
  OAI211_X1 U17985 ( .C1(n14591), .C2(n14590), .A(n14589), .B(n14588), .ZN(
        n14592) );
  AOI21_X1 U17986 ( .B1(n20139), .B2(n20037), .A(n14592), .ZN(n14593) );
  OAI21_X1 U17987 ( .B1(n14595), .B2(n14594), .A(n14593), .ZN(P1_U2838) );
  OAI22_X1 U17988 ( .A1(n14883), .A2(n14636), .B1(n16118), .B2(n14596), .ZN(
        P1_U2841) );
  AOI22_X1 U17989 ( .A1(n14941), .A2(n16115), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n14623), .ZN(n14597) );
  OAI21_X1 U17990 ( .B1(n14744), .B2(n14628), .A(n14597), .ZN(P1_U2844) );
  INV_X1 U17991 ( .A(n14750), .ZN(n14653) );
  OAI222_X1 U17992 ( .A1(n14638), .A2(n14653), .B1(n14598), .B2(n16118), .C1(
        n14956), .C2(n14636), .ZN(P1_U2845) );
  AOI22_X1 U17993 ( .A1(n14973), .A2(n16115), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n14623), .ZN(n14599) );
  OAI21_X1 U17994 ( .B1(n14757), .B2(n14628), .A(n14599), .ZN(P1_U2846) );
  INV_X1 U17995 ( .A(n14771), .ZN(n14660) );
  INV_X1 U17996 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14600) );
  OAI222_X1 U17997 ( .A1(n14660), .A2(n14638), .B1(n14600), .B2(n16118), .C1(
        n14980), .C2(n14636), .ZN(P1_U2847) );
  AOI22_X1 U17998 ( .A1(n14992), .A2(n16115), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n14623), .ZN(n14601) );
  OAI21_X1 U17999 ( .B1(n14782), .B2(n14628), .A(n14601), .ZN(P1_U2848) );
  AOI22_X1 U18000 ( .A1(n14602), .A2(n16115), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n14623), .ZN(n14603) );
  OAI21_X1 U18001 ( .B1(n14668), .B2(n14628), .A(n14603), .ZN(P1_U2849) );
  OAI222_X1 U18002 ( .A1(n16158), .A2(n14636), .B1(n14604), .B2(n16118), .C1(
        n14799), .C2(n14638), .ZN(P1_U2850) );
  INV_X1 U18003 ( .A(n14807), .ZN(n14678) );
  AOI22_X1 U18004 ( .A1(n15016), .A2(n16115), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n14623), .ZN(n14605) );
  OAI21_X1 U18005 ( .B1(n14678), .B2(n14638), .A(n14605), .ZN(P1_U2851) );
  INV_X1 U18006 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14606) );
  OAI222_X1 U18007 ( .A1(n14686), .A2(n14638), .B1(n14606), .B2(n16118), .C1(
        n15019), .C2(n14636), .ZN(P1_U2852) );
  AOI22_X1 U18008 ( .A1(n16166), .A2(n16115), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14623), .ZN(n14607) );
  OAI21_X1 U18009 ( .B1(n14691), .B2(n14638), .A(n14607), .ZN(P1_U2853) );
  OAI22_X1 U18010 ( .A1(n15046), .A2(n14636), .B1(n14608), .B2(n16118), .ZN(
        n14609) );
  INV_X1 U18011 ( .A(n14609), .ZN(n14610) );
  OAI21_X1 U18012 ( .B1(n14824), .B2(n14628), .A(n14610), .ZN(P1_U2854) );
  INV_X1 U18013 ( .A(n14611), .ZN(n14613) );
  INV_X1 U18014 ( .A(n14535), .ZN(n14612) );
  AOI21_X1 U18015 ( .B1(n14613), .B2(n14612), .A(n14524), .ZN(n16137) );
  INV_X1 U18016 ( .A(n16137), .ZN(n14698) );
  INV_X1 U18017 ( .A(n14614), .ZN(n14615) );
  NAND2_X1 U18018 ( .A1(n14616), .A2(n14615), .ZN(n14618) );
  NAND2_X1 U18019 ( .A1(n14618), .A2(n14617), .ZN(n14620) );
  AND2_X1 U18020 ( .A1(n14620), .A2(n14619), .ZN(n16172) );
  AOI22_X1 U18021 ( .A1(n16172), .A2(n16115), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14623), .ZN(n14621) );
  OAI21_X1 U18022 ( .B1(n14698), .B2(n14638), .A(n14621), .ZN(P1_U2855) );
  AOI22_X1 U18023 ( .A1(n16178), .A2(n16115), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n14623), .ZN(n14622) );
  OAI21_X1 U18024 ( .B1(n14705), .B2(n14638), .A(n14622), .ZN(P1_U2856) );
  INV_X1 U18025 ( .A(n14847), .ZN(n14707) );
  AOI22_X1 U18026 ( .A1(n16186), .A2(n16115), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n14623), .ZN(n14624) );
  OAI21_X1 U18027 ( .B1(n14707), .B2(n14628), .A(n14624), .ZN(P1_U2857) );
  OAI22_X1 U18028 ( .A1(n16193), .A2(n14636), .B1(n14625), .B2(n16118), .ZN(
        n14626) );
  INV_X1 U18029 ( .A(n14626), .ZN(n14627) );
  OAI21_X1 U18030 ( .B1(n14708), .B2(n14628), .A(n14627), .ZN(P1_U2858) );
  AOI21_X1 U18031 ( .B1(n9738), .B2(n14710), .A(n14630), .ZN(n14631) );
  INV_X1 U18032 ( .A(n16096), .ZN(n14709) );
  INV_X1 U18033 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14637) );
  AOI21_X1 U18034 ( .B1(n9951), .B2(n16100), .A(n14632), .ZN(n14635) );
  INV_X1 U18035 ( .A(n14633), .ZN(n14634) );
  NOR2_X1 U18036 ( .A1(n14635), .A2(n14634), .ZN(n16093) );
  INV_X1 U18037 ( .A(n16093), .ZN(n15054) );
  OAI222_X1 U18038 ( .A1(n14709), .A2(n14638), .B1(n14637), .B2(n16118), .C1(
        n14636), .C2(n15054), .ZN(P1_U2859) );
  INV_X1 U18039 ( .A(DATAI_13_), .ZN(n14640) );
  MUX2_X1 U18040 ( .A(n14640), .B(n14639), .S(n20130), .Z(n20066) );
  OAI22_X1 U18041 ( .A1(n14699), .A2(n20066), .B1(n14661), .B2(n13076), .ZN(
        n14641) );
  AOI21_X1 U18042 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n14701), .A(n14641), .ZN(
        n14643) );
  NAND2_X1 U18043 ( .A1(n14702), .A2(DATAI_29_), .ZN(n14642) );
  OAI211_X1 U18044 ( .C1(n14644), .C2(n14712), .A(n14643), .B(n14642), .ZN(
        P1_U2875) );
  INV_X1 U18045 ( .A(DATAI_12_), .ZN(n14645) );
  INV_X1 U18046 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16605) );
  MUX2_X1 U18047 ( .A(n14645), .B(n16605), .S(n20130), .Z(n20063) );
  OAI22_X1 U18048 ( .A1(n14699), .A2(n20063), .B1(n14661), .B2(n13094), .ZN(
        n14646) );
  AOI21_X1 U18049 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n14701), .A(n14646), .ZN(
        n14648) );
  NAND2_X1 U18050 ( .A1(n14702), .A2(DATAI_28_), .ZN(n14647) );
  OAI211_X1 U18051 ( .C1(n14744), .C2(n14712), .A(n14648), .B(n14647), .ZN(
        P1_U2876) );
  INV_X1 U18052 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n19318) );
  INV_X1 U18053 ( .A(n14699), .ZN(n14681) );
  AOI22_X1 U18054 ( .A1(n14681), .A2(n14649), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n14679), .ZN(n14650) );
  OAI21_X1 U18055 ( .B1(n19318), .B2(n14683), .A(n14650), .ZN(n14651) );
  AOI21_X1 U18056 ( .B1(n14702), .B2(DATAI_27_), .A(n14651), .ZN(n14652) );
  OAI21_X1 U18057 ( .B1(n14653), .B2(n14712), .A(n14652), .ZN(P1_U2877) );
  OAI22_X1 U18058 ( .A1(n14699), .A2(n20060), .B1(n14661), .B2(n13085), .ZN(
        n14654) );
  AOI21_X1 U18059 ( .B1(BUF1_REG_26__SCAN_IN), .B2(n14701), .A(n14654), .ZN(
        n14656) );
  NAND2_X1 U18060 ( .A1(n14702), .A2(DATAI_26_), .ZN(n14655) );
  OAI211_X1 U18061 ( .C1(n14757), .C2(n14712), .A(n14656), .B(n14655), .ZN(
        P1_U2878) );
  OAI22_X1 U18062 ( .A1(n14699), .A2(n20057), .B1(n14661), .B2(n13088), .ZN(
        n14657) );
  AOI21_X1 U18063 ( .B1(n14701), .B2(BUF1_REG_25__SCAN_IN), .A(n14657), .ZN(
        n14659) );
  NAND2_X1 U18064 ( .A1(n14702), .A2(DATAI_25_), .ZN(n14658) );
  OAI211_X1 U18065 ( .C1(n14660), .C2(n14712), .A(n14659), .B(n14658), .ZN(
        P1_U2879) );
  OAI22_X1 U18066 ( .A1(n14699), .A2(n20054), .B1(n14661), .B2(n13091), .ZN(
        n14662) );
  AOI21_X1 U18067 ( .B1(n14701), .B2(BUF1_REG_24__SCAN_IN), .A(n14662), .ZN(
        n14664) );
  NAND2_X1 U18068 ( .A1(n14702), .A2(DATAI_24_), .ZN(n14663) );
  OAI211_X1 U18069 ( .C1(n14782), .C2(n14712), .A(n14664), .B(n14663), .ZN(
        P1_U2880) );
  OAI22_X1 U18070 ( .A1(n14699), .A2(n20174), .B1(n14661), .B2(n13391), .ZN(
        n14665) );
  AOI21_X1 U18071 ( .B1(n14701), .B2(BUF1_REG_23__SCAN_IN), .A(n14665), .ZN(
        n14667) );
  NAND2_X1 U18072 ( .A1(n14702), .A2(DATAI_23_), .ZN(n14666) );
  OAI211_X1 U18073 ( .C1(n14668), .C2(n14712), .A(n14667), .B(n14666), .ZN(
        P1_U2881) );
  INV_X1 U18074 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n14671) );
  AOI22_X1 U18075 ( .A1(n14681), .A2(n14669), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n14679), .ZN(n14670) );
  OAI21_X1 U18076 ( .B1(n14683), .B2(n14671), .A(n14670), .ZN(n14672) );
  AOI21_X1 U18077 ( .B1(n14702), .B2(DATAI_22_), .A(n14672), .ZN(n14673) );
  OAI21_X1 U18078 ( .B1(n14799), .B2(n14712), .A(n14673), .ZN(P1_U2882) );
  OAI22_X1 U18079 ( .A1(n14699), .A2(n20165), .B1(n14661), .B2(n14674), .ZN(
        n14675) );
  AOI21_X1 U18080 ( .B1(n14701), .B2(BUF1_REG_21__SCAN_IN), .A(n14675), .ZN(
        n14677) );
  NAND2_X1 U18081 ( .A1(n14702), .A2(DATAI_21_), .ZN(n14676) );
  OAI211_X1 U18082 ( .C1(n14678), .C2(n14712), .A(n14677), .B(n14676), .ZN(
        P1_U2883) );
  INV_X1 U18083 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16593) );
  AOI22_X1 U18084 ( .A1(n14681), .A2(n14680), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n14679), .ZN(n14682) );
  OAI21_X1 U18085 ( .B1(n14683), .B2(n16593), .A(n14682), .ZN(n14684) );
  AOI21_X1 U18086 ( .B1(n14702), .B2(DATAI_20_), .A(n14684), .ZN(n14685) );
  OAI21_X1 U18087 ( .B1(n14686), .B2(n14712), .A(n14685), .ZN(P1_U2884) );
  OAI22_X1 U18088 ( .A1(n14699), .A2(n20158), .B1(n14661), .B2(n14687), .ZN(
        n14688) );
  AOI21_X1 U18089 ( .B1(n14701), .B2(BUF1_REG_19__SCAN_IN), .A(n14688), .ZN(
        n14690) );
  NAND2_X1 U18090 ( .A1(n14702), .A2(DATAI_19_), .ZN(n14689) );
  OAI211_X1 U18091 ( .C1(n14691), .C2(n14712), .A(n14690), .B(n14689), .ZN(
        P1_U2885) );
  OAI22_X1 U18092 ( .A1(n14699), .A2(n20154), .B1(n14661), .B2(n13405), .ZN(
        n14692) );
  AOI21_X1 U18093 ( .B1(n14701), .B2(BUF1_REG_18__SCAN_IN), .A(n14692), .ZN(
        n14694) );
  NAND2_X1 U18094 ( .A1(n14702), .A2(DATAI_18_), .ZN(n14693) );
  OAI211_X1 U18095 ( .C1(n14824), .C2(n14712), .A(n14694), .B(n14693), .ZN(
        P1_U2886) );
  OAI22_X1 U18096 ( .A1(n14699), .A2(n20151), .B1(n14661), .B2(n13408), .ZN(
        n14695) );
  AOI21_X1 U18097 ( .B1(n14701), .B2(BUF1_REG_17__SCAN_IN), .A(n14695), .ZN(
        n14697) );
  NAND2_X1 U18098 ( .A1(n14702), .A2(DATAI_17_), .ZN(n14696) );
  OAI211_X1 U18099 ( .C1(n14698), .C2(n14712), .A(n14697), .B(n14696), .ZN(
        P1_U2887) );
  OAI22_X1 U18100 ( .A1(n14699), .A2(n20142), .B1(n14661), .B2(n13399), .ZN(
        n14700) );
  AOI21_X1 U18101 ( .B1(n14701), .B2(BUF1_REG_16__SCAN_IN), .A(n14700), .ZN(
        n14704) );
  NAND2_X1 U18102 ( .A1(n14702), .A2(DATAI_16_), .ZN(n14703) );
  OAI211_X1 U18103 ( .C1(n14705), .C2(n14712), .A(n14704), .B(n14703), .ZN(
        P1_U2888) );
  OAI222_X1 U18104 ( .A1(n14707), .A2(n14712), .B1(n14661), .B2(n13180), .C1(
        n14711), .C2(n14706), .ZN(P1_U2889) );
  OAI222_X1 U18105 ( .A1(n14708), .A2(n14712), .B1(n13422), .B2(n14661), .C1(
        n14711), .C2(n20069), .ZN(P1_U2890) );
  OAI222_X1 U18106 ( .A1(n14709), .A2(n14712), .B1(n13430), .B2(n14661), .C1(
        n14711), .C2(n20066), .ZN(P1_U2891) );
  XOR2_X1 U18107 ( .A(n14710), .B(n9738), .Z(n16145) );
  INV_X1 U18108 ( .A(n16145), .ZN(n14713) );
  OAI222_X1 U18109 ( .A1(n14713), .A2(n14712), .B1(n13419), .B2(n14661), .C1(
        n14711), .C2(n20063), .ZN(P1_U2892) );
  AOI21_X1 U18110 ( .B1(n14716), .B2(n14734), .A(n14715), .ZN(n14717) );
  XNOR2_X1 U18111 ( .A(n14717), .B(n13195), .ZN(n14921) );
  INV_X1 U18112 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21075) );
  NOR2_X1 U18113 ( .A1(n16200), .A2(n21075), .ZN(n14898) );
  AOI21_X1 U18114 ( .B1(n16135), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14898), .ZN(n14718) );
  OAI21_X1 U18115 ( .B1(n14719), .B2(n16127), .A(n14718), .ZN(n14720) );
  OAI21_X1 U18116 ( .B1(n14921), .B2(n19970), .A(n14722), .ZN(P1_U2968) );
  MUX2_X1 U18117 ( .A(n14724), .B(n14723), .S(n14734), .Z(n14725) );
  XNOR2_X1 U18118 ( .A(n14725), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14940) );
  NOR2_X1 U18119 ( .A1(n16200), .A2(n20783), .ZN(n14934) );
  AOI21_X1 U18120 ( .B1(n16135), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14934), .ZN(n14726) );
  OAI21_X1 U18121 ( .B1(n14727), .B2(n16127), .A(n14726), .ZN(n14728) );
  AOI21_X1 U18122 ( .B1(n14729), .B2(n16152), .A(n14728), .ZN(n14730) );
  OAI21_X1 U18123 ( .B1(n19970), .B2(n14940), .A(n14730), .ZN(P1_U2970) );
  INV_X1 U18124 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20781) );
  NOR2_X1 U18125 ( .A1(n16200), .A2(n20781), .ZN(n14949) );
  NOR2_X1 U18126 ( .A1(n14818), .A2(n14731), .ZN(n14732) );
  AOI211_X1 U18127 ( .C1(n14733), .C2(n16151), .A(n14949), .B(n14732), .ZN(
        n14743) );
  INV_X1 U18128 ( .A(n14897), .ZN(n14968) );
  NAND2_X1 U18129 ( .A1(n14765), .A2(n14968), .ZN(n14735) );
  NAND2_X1 U18130 ( .A1(n14762), .A2(n14735), .ZN(n14737) );
  NAND3_X1 U18131 ( .A1(n14753), .A2(n14967), .A3(n14958), .ZN(n14736) );
  NOR2_X1 U18132 ( .A1(n14737), .A2(n14736), .ZN(n14739) );
  AND3_X1 U18133 ( .A1(n14737), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14738) );
  MUX2_X1 U18134 ( .A(n14739), .B(n14738), .S(n9721), .Z(n14741) );
  NAND2_X1 U18135 ( .A1(n14942), .A2(n11125), .ZN(n14742) );
  OAI211_X1 U18136 ( .C1(n14744), .C2(n20129), .A(n14743), .B(n14742), .ZN(
        P1_U2971) );
  XNOR2_X1 U18137 ( .A(n14746), .B(n14958), .ZN(n14961) );
  INV_X1 U18138 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20779) );
  NOR2_X1 U18139 ( .A1(n16200), .A2(n20779), .ZN(n14953) );
  AOI21_X1 U18140 ( .B1(n16135), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14953), .ZN(n14747) );
  OAI21_X1 U18141 ( .B1(n14748), .B2(n16127), .A(n14747), .ZN(n14749) );
  AOI21_X1 U18142 ( .B1(n14750), .B2(n16152), .A(n14749), .ZN(n14751) );
  OAI21_X1 U18143 ( .B1(n19970), .B2(n14961), .A(n14751), .ZN(P1_U2972) );
  MUX2_X1 U18144 ( .A(n14753), .B(n14968), .S(n9721), .Z(n14754) );
  NAND3_X1 U18145 ( .A1(n14762), .A2(n14752), .A3(n14754), .ZN(n14755) );
  XNOR2_X1 U18146 ( .A(n14755), .B(n14967), .ZN(n14975) );
  NAND2_X1 U18147 ( .A1(n16171), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14969) );
  OAI21_X1 U18148 ( .B1(n14818), .B2(n14756), .A(n14969), .ZN(n14759) );
  NOR2_X1 U18149 ( .A1(n14757), .A2(n20129), .ZN(n14758) );
  OAI21_X1 U18150 ( .B1(n19970), .B2(n14975), .A(n14761), .ZN(P1_U2973) );
  NAND2_X1 U18151 ( .A1(n14734), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14763) );
  NAND2_X1 U18152 ( .A1(n14762), .A2(n14763), .ZN(n14778) );
  NAND2_X1 U18153 ( .A1(n9721), .A2(n15002), .ZN(n14776) );
  NAND2_X1 U18154 ( .A1(n14763), .A2(n14776), .ZN(n14783) );
  NOR2_X1 U18155 ( .A1(n14783), .A2(n14993), .ZN(n14764) );
  NAND2_X1 U18156 ( .A1(n15002), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14989) );
  AOI22_X1 U18157 ( .A1(n14765), .A2(n14764), .B1(n14734), .B2(n14989), .ZN(
        n14766) );
  OR2_X1 U18158 ( .A1(n14778), .A2(n14766), .ZN(n14767) );
  XNOR2_X1 U18159 ( .A(n14767), .B(n14962), .ZN(n14983) );
  NOR2_X1 U18160 ( .A1(n16200), .A2(n20775), .ZN(n14976) );
  AOI21_X1 U18161 ( .B1(n16135), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14976), .ZN(n14768) );
  OAI21_X1 U18162 ( .B1(n14769), .B2(n16127), .A(n14768), .ZN(n14770) );
  AOI21_X1 U18163 ( .B1(n14771), .B2(n16152), .A(n14770), .ZN(n14772) );
  OAI21_X1 U18164 ( .B1(n19970), .B2(n14983), .A(n14772), .ZN(P1_U2974) );
  NOR2_X1 U18165 ( .A1(n16200), .A2(n20773), .ZN(n14986) );
  NOR2_X1 U18166 ( .A1(n14818), .A2(n14773), .ZN(n14774) );
  AOI211_X1 U18167 ( .C1(n14775), .C2(n16151), .A(n14986), .B(n14774), .ZN(
        n14781) );
  NAND2_X1 U18168 ( .A1(n14752), .A2(n14776), .ZN(n14777) );
  XNOR2_X1 U18169 ( .A(n14779), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14984) );
  NAND2_X1 U18170 ( .A1(n14984), .A2(n11125), .ZN(n14780) );
  OAI211_X1 U18171 ( .C1(n14782), .C2(n20129), .A(n14781), .B(n14780), .ZN(
        P1_U2975) );
  XNOR2_X1 U18172 ( .A(n14784), .B(n14783), .ZN(n15005) );
  NOR2_X1 U18173 ( .A1(n16200), .A2(n14785), .ZN(n14997) );
  AOI21_X1 U18174 ( .B1(n16135), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n14997), .ZN(n14786) );
  OAI21_X1 U18175 ( .B1(n14787), .B2(n16127), .A(n14786), .ZN(n14788) );
  AOI21_X1 U18176 ( .B1(n14789), .B2(n16152), .A(n14788), .ZN(n14790) );
  OAI21_X1 U18177 ( .B1(n19970), .B2(n15005), .A(n14790), .ZN(P1_U2976) );
  INV_X1 U18178 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20770) );
  OAI22_X1 U18179 ( .A1(n14818), .A2(n14791), .B1(n16200), .B2(n20770), .ZN(
        n14792) );
  AOI21_X1 U18180 ( .B1(n14793), .B2(n16151), .A(n14792), .ZN(n14798) );
  OAI21_X1 U18181 ( .B1(n14795), .B2(n9721), .A(n14794), .ZN(n14796) );
  XNOR2_X1 U18182 ( .A(n14796), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16160) );
  NAND2_X1 U18183 ( .A1(n16160), .A2(n11125), .ZN(n14797) );
  OAI211_X1 U18184 ( .C1(n14799), .C2(n20129), .A(n14798), .B(n14797), .ZN(
        P1_U2977) );
  OAI21_X1 U18185 ( .B1(n9721), .B2(n14894), .A(n14800), .ZN(n16121) );
  NAND2_X1 U18186 ( .A1(n14734), .A2(n15020), .ZN(n16120) );
  NAND2_X1 U18187 ( .A1(n9721), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16119) );
  OAI22_X1 U18188 ( .A1(n16121), .A2(n16120), .B1(n14800), .B2(n16119), .ZN(
        n14809) );
  NAND2_X1 U18189 ( .A1(n14809), .A2(n15024), .ZN(n14810) );
  INV_X1 U18190 ( .A(n16119), .ZN(n14801) );
  NAND2_X1 U18191 ( .A1(n14801), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14802) );
  OAI22_X1 U18192 ( .A1(n14810), .A2(n9721), .B1(n14800), .B2(n14802), .ZN(
        n14803) );
  XNOR2_X1 U18193 ( .A(n14803), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15018) );
  NAND2_X1 U18194 ( .A1(n16171), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15012) );
  NAND2_X1 U18195 ( .A1(n16135), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14804) );
  OAI211_X1 U18196 ( .C1(n14805), .C2(n16127), .A(n15012), .B(n14804), .ZN(
        n14806) );
  AOI21_X1 U18197 ( .B1(n14807), .B2(n16152), .A(n14806), .ZN(n14808) );
  OAI21_X1 U18198 ( .B1(n15018), .B2(n19970), .A(n14808), .ZN(P1_U2978) );
  INV_X1 U18199 ( .A(n14809), .ZN(n14812) );
  INV_X1 U18200 ( .A(n14810), .ZN(n14811) );
  AOI21_X1 U18201 ( .B1(n14812), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14811), .ZN(n15031) );
  NAND2_X1 U18202 ( .A1(n14813), .A2(n16151), .ZN(n14814) );
  NAND2_X1 U18203 ( .A1(n16171), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15025) );
  OAI211_X1 U18204 ( .C1(n14818), .C2(n21040), .A(n14814), .B(n15025), .ZN(
        n14815) );
  AOI21_X1 U18205 ( .B1(n14816), .B2(n16152), .A(n14815), .ZN(n14817) );
  OAI21_X1 U18206 ( .B1(n15031), .B2(n19970), .A(n14817), .ZN(P1_U2979) );
  NAND2_X1 U18207 ( .A1(n16171), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15045) );
  OAI21_X1 U18208 ( .B1(n14818), .B2(n10167), .A(n15045), .ZN(n14819) );
  AOI21_X1 U18209 ( .B1(n14820), .B2(n16151), .A(n14819), .ZN(n14823) );
  OR2_X1 U18210 ( .A1(n11064), .A2(n14821), .ZN(n15032) );
  NAND3_X1 U18211 ( .A1(n15032), .A2(n11125), .A3(n14800), .ZN(n14822) );
  OAI211_X1 U18212 ( .C1(n14824), .C2(n20129), .A(n14823), .B(n14822), .ZN(
        P1_U2981) );
  NOR2_X1 U18213 ( .A1(n16148), .A2(n14825), .ZN(n14842) );
  OAI21_X1 U18214 ( .B1(n14842), .B2(n14840), .A(n14839), .ZN(n14827) );
  XNOR2_X1 U18215 ( .A(n14827), .B(n14826), .ZN(n16179) );
  INV_X1 U18216 ( .A(n16179), .ZN(n14835) );
  INV_X1 U18217 ( .A(n14828), .ZN(n14831) );
  INV_X1 U18218 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14829) );
  NOR2_X1 U18219 ( .A1(n16200), .A2(n14829), .ZN(n16177) );
  AOI21_X1 U18220 ( .B1(n16135), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16177), .ZN(n14830) );
  OAI21_X1 U18221 ( .B1(n16127), .B2(n14831), .A(n14830), .ZN(n14832) );
  AOI21_X1 U18222 ( .B1(n14833), .B2(n16152), .A(n14832), .ZN(n14834) );
  OAI21_X1 U18223 ( .B1(n19970), .B2(n14835), .A(n14834), .ZN(P1_U2983) );
  INV_X1 U18224 ( .A(n14842), .ZN(n14838) );
  AOI22_X1 U18225 ( .A1(n14838), .A2(n14837), .B1(n14836), .B2(n14839), .ZN(
        n14844) );
  INV_X1 U18226 ( .A(n14839), .ZN(n14841) );
  NOR3_X1 U18227 ( .A1(n14842), .A2(n14841), .A3(n14840), .ZN(n14843) );
  NOR2_X1 U18228 ( .A1(n14844), .A2(n14843), .ZN(n16187) );
  NOR2_X1 U18229 ( .A1(n16200), .A2(n20759), .ZN(n16185) );
  AND2_X1 U18230 ( .A1(n16135), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14845) );
  AOI211_X1 U18231 ( .C1(n14846), .C2(n16151), .A(n16185), .B(n14845), .ZN(
        n14849) );
  NAND2_X1 U18232 ( .A1(n14847), .A2(n16152), .ZN(n14848) );
  OAI211_X1 U18233 ( .C1(n16187), .C2(n19970), .A(n14849), .B(n14848), .ZN(
        P1_U2984) );
  NOR2_X1 U18234 ( .A1(n9721), .A2(n16214), .ZN(n14865) );
  NOR2_X1 U18235 ( .A1(n9721), .A2(n14850), .ZN(n14862) );
  NOR3_X1 U18236 ( .A1(n9776), .A2(n14865), .A3(n14862), .ZN(n16131) );
  INV_X1 U18237 ( .A(n14851), .ZN(n14853) );
  OAI21_X1 U18238 ( .B1(n16131), .B2(n14853), .A(n14852), .ZN(n14855) );
  XNOR2_X1 U18239 ( .A(n9721), .B(n16198), .ZN(n14854) );
  XNOR2_X1 U18240 ( .A(n14855), .B(n14854), .ZN(n16195) );
  INV_X1 U18241 ( .A(n16195), .ZN(n14861) );
  AOI22_X1 U18242 ( .A1(n16135), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16171), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n14856) );
  OAI21_X1 U18243 ( .B1(n16127), .B2(n14857), .A(n14856), .ZN(n14858) );
  AOI21_X1 U18244 ( .B1(n14859), .B2(n16152), .A(n14858), .ZN(n14860) );
  OAI21_X1 U18245 ( .B1(n14861), .B2(n19970), .A(n14860), .ZN(P1_U2985) );
  AOI21_X1 U18246 ( .B1(n9776), .B2(n14863), .A(n14862), .ZN(n16142) );
  INV_X1 U18247 ( .A(n14866), .ZN(n14864) );
  NOR2_X1 U18248 ( .A1(n14865), .A2(n14864), .ZN(n16141) );
  NAND2_X1 U18249 ( .A1(n16142), .A2(n16141), .ZN(n16140) );
  NAND2_X1 U18250 ( .A1(n16140), .A2(n14866), .ZN(n14868) );
  XNOR2_X1 U18251 ( .A(n14868), .B(n14867), .ZN(n15062) );
  INV_X1 U18252 ( .A(n16089), .ZN(n14870) );
  NAND2_X1 U18253 ( .A1(n16171), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15053) );
  NAND2_X1 U18254 ( .A1(n16135), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14869) );
  OAI211_X1 U18255 ( .C1(n16127), .C2(n14870), .A(n15053), .B(n14869), .ZN(
        n14871) );
  AOI21_X1 U18256 ( .B1(n16096), .B2(n16152), .A(n14871), .ZN(n14872) );
  OAI21_X1 U18257 ( .B1(n15062), .B2(n19970), .A(n14872), .ZN(P1_U2986) );
  INV_X1 U18258 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16234) );
  NOR2_X1 U18259 ( .A1(n16148), .A2(n16234), .ZN(n14875) );
  NOR2_X1 U18260 ( .A1(n14873), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14874) );
  MUX2_X1 U18261 ( .A(n14875), .B(n14874), .S(n14734), .Z(n14876) );
  INV_X1 U18262 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16225) );
  XNOR2_X1 U18263 ( .A(n14876), .B(n16225), .ZN(n16222) );
  NAND2_X1 U18264 ( .A1(n16222), .A2(n11125), .ZN(n14881) );
  INV_X1 U18265 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n14877) );
  NOR2_X1 U18266 ( .A1(n16200), .A2(n14877), .ZN(n16219) );
  NOR2_X1 U18267 ( .A1(n16127), .A2(n14878), .ZN(n14879) );
  AOI211_X1 U18268 ( .C1(n16135), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16219), .B(n14879), .ZN(n14880) );
  OAI211_X1 U18269 ( .C1(n20129), .C2(n14882), .A(n14881), .B(n14880), .ZN(
        P1_U2988) );
  INV_X1 U18270 ( .A(n14883), .ZN(n14919) );
  NAND2_X1 U18271 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14884), .ZN(
        n14885) );
  NOR3_X1 U18272 ( .A1(n10996), .A2(n11153), .A3(n14885), .ZN(n16203) );
  NOR3_X1 U18273 ( .A1(n14887), .A2(n11040), .A3(n14886), .ZN(n16232) );
  NAND3_X1 U18274 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n16232), .ZN(n16208) );
  NOR2_X1 U18275 ( .A1(n16225), .A2(n16208), .ZN(n16215) );
  INV_X1 U18276 ( .A(n16215), .ZN(n16206) );
  NOR2_X1 U18277 ( .A1(n16214), .A2(n16206), .ZN(n14890) );
  NAND2_X1 U18278 ( .A1(n16203), .A2(n14890), .ZN(n15007) );
  NOR2_X1 U18279 ( .A1(n15055), .A2(n15007), .ZN(n15052) );
  NAND2_X1 U18280 ( .A1(n14888), .A2(n15052), .ZN(n14990) );
  AND2_X1 U18281 ( .A1(n14890), .A2(n14889), .ZN(n15008) );
  NAND2_X1 U18282 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15008), .ZN(
        n15033) );
  INV_X1 U18283 ( .A(n15033), .ZN(n14899) );
  NAND2_X1 U18284 ( .A1(n16207), .A2(n14899), .ZN(n14891) );
  INV_X1 U18285 ( .A(n16199), .ZN(n14896) );
  NOR2_X1 U18286 ( .A1(n14893), .A2(n14892), .ZN(n16183) );
  NAND3_X1 U18287 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n16183), .ZN(n15044) );
  NOR2_X1 U18288 ( .A1(n14894), .A2(n15044), .ZN(n14900) );
  NAND2_X1 U18289 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16161) );
  INV_X1 U18290 ( .A(n16161), .ZN(n14906) );
  AND3_X1 U18291 ( .A1(n14900), .A2(n14904), .A3(n14906), .ZN(n14895) );
  NAND2_X1 U18292 ( .A1(n14896), .A2(n14895), .ZN(n14966) );
  NOR3_X1 U18293 ( .A1(n14966), .A2(n14897), .A3(n14967), .ZN(n14959) );
  NAND2_X1 U18294 ( .A1(n14959), .A2(n14912), .ZN(n14937) );
  NAND3_X1 U18295 ( .A1(n13195), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14917) );
  INV_X1 U18296 ( .A(n14898), .ZN(n14916) );
  AND2_X1 U18297 ( .A1(n14900), .A2(n14899), .ZN(n14903) );
  INV_X1 U18298 ( .A(n15007), .ZN(n15059) );
  NAND2_X1 U18299 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14900), .ZN(
        n15009) );
  INV_X1 U18300 ( .A(n15009), .ZN(n14901) );
  NAND2_X1 U18301 ( .A1(n15059), .A2(n14901), .ZN(n15006) );
  NAND2_X1 U18302 ( .A1(n20099), .A2(n15006), .ZN(n14902) );
  OAI211_X1 U18303 ( .C1(n14903), .C2(n20104), .A(n14902), .B(n20097), .ZN(
        n16165) );
  INV_X1 U18304 ( .A(n14904), .ZN(n15011) );
  NOR2_X1 U18305 ( .A1(n16165), .A2(n15011), .ZN(n14905) );
  AND2_X1 U18306 ( .A1(n15043), .A2(n20097), .ZN(n16229) );
  OR2_X1 U18307 ( .A1(n14905), .A2(n16229), .ZN(n16156) );
  OR2_X1 U18308 ( .A1(n15043), .A2(n14906), .ZN(n14907) );
  NAND2_X1 U18309 ( .A1(n16156), .A2(n14907), .ZN(n14998) );
  AND2_X1 U18310 ( .A1(n16207), .A2(n15002), .ZN(n14908) );
  NOR2_X1 U18311 ( .A1(n14998), .A2(n14908), .ZN(n14985) );
  OAI22_X1 U18312 ( .A1(n20119), .A2(n14963), .B1(n14968), .B2(n15051), .ZN(
        n14909) );
  INV_X1 U18313 ( .A(n14909), .ZN(n14910) );
  NAND2_X1 U18314 ( .A1(n14985), .A2(n14910), .ZN(n14977) );
  INV_X1 U18315 ( .A(n15043), .ZN(n14911) );
  OR2_X1 U18316 ( .A1(n14977), .A2(n14911), .ZN(n14945) );
  INV_X1 U18317 ( .A(n14912), .ZN(n14913) );
  NAND2_X1 U18318 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14943) );
  OR3_X1 U18319 ( .A1(n14977), .A2(n14913), .A3(n14943), .ZN(n14914) );
  NAND2_X1 U18320 ( .A1(n14945), .A2(n14914), .ZN(n14933) );
  OAI211_X1 U18321 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15043), .A(
        n14933), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14924) );
  NAND3_X1 U18322 ( .A1(n14924), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14945), .ZN(n14915) );
  OAI211_X1 U18323 ( .C1(n14937), .C2(n14917), .A(n14916), .B(n14915), .ZN(
        n14918) );
  AOI21_X1 U18324 ( .B1(n14919), .B2(n20116), .A(n14918), .ZN(n14920) );
  OAI21_X1 U18325 ( .B1(n14921), .B2(n20091), .A(n14920), .ZN(P1_U3000) );
  INV_X1 U18326 ( .A(n14922), .ZN(n14929) );
  INV_X1 U18327 ( .A(n14937), .ZN(n14923) );
  AOI21_X1 U18328 ( .B1(n14923), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14927) );
  INV_X1 U18329 ( .A(n14924), .ZN(n14926) );
  OAI21_X1 U18330 ( .B1(n14927), .B2(n14926), .A(n14925), .ZN(n14928) );
  AOI21_X1 U18331 ( .B1(n14929), .B2(n20116), .A(n14928), .ZN(n14930) );
  OAI21_X1 U18332 ( .B1(n14931), .B2(n20091), .A(n14930), .ZN(P1_U3001) );
  INV_X1 U18333 ( .A(n14933), .ZN(n14935) );
  AOI21_X1 U18334 ( .B1(n14935), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14934), .ZN(n14936) );
  OAI21_X1 U18335 ( .B1(n14937), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14936), .ZN(n14938) );
  AOI21_X1 U18336 ( .B1(n11254), .B2(n20116), .A(n14938), .ZN(n14939) );
  OAI21_X1 U18337 ( .B1(n14940), .B2(n20091), .A(n14939), .ZN(P1_U3002) );
  INV_X1 U18338 ( .A(n14941), .ZN(n14952) );
  NAND2_X1 U18339 ( .A1(n14942), .A2(n20117), .ZN(n14951) );
  OR2_X1 U18340 ( .A1(n14977), .A2(n14943), .ZN(n14944) );
  AND2_X1 U18341 ( .A1(n14945), .A2(n14944), .ZN(n14954) );
  INV_X1 U18342 ( .A(n14959), .ZN(n14947) );
  XNOR2_X1 U18343 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14946) );
  NOR2_X1 U18344 ( .A1(n14947), .A2(n14946), .ZN(n14948) );
  AOI211_X1 U18345 ( .C1(n14954), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14949), .B(n14948), .ZN(n14950) );
  OAI211_X1 U18346 ( .C1(n20107), .C2(n14952), .A(n14951), .B(n14950), .ZN(
        P1_U3003) );
  AOI21_X1 U18347 ( .B1(n14954), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14953), .ZN(n14955) );
  OAI21_X1 U18348 ( .B1(n14956), .B2(n20107), .A(n14955), .ZN(n14957) );
  AOI21_X1 U18349 ( .B1(n14959), .B2(n14958), .A(n14957), .ZN(n14960) );
  OAI21_X1 U18350 ( .B1(n14961), .B2(n20091), .A(n14960), .ZN(P1_U3004) );
  NAND2_X1 U18351 ( .A1(n14963), .A2(n14962), .ZN(n14964) );
  OR2_X1 U18352 ( .A1(n14966), .A2(n14964), .ZN(n14978) );
  INV_X1 U18353 ( .A(n14977), .ZN(n14965) );
  AOI21_X1 U18354 ( .B1(n14978), .B2(n14965), .A(n14967), .ZN(n14972) );
  INV_X1 U18355 ( .A(n14966), .ZN(n15003) );
  NAND3_X1 U18356 ( .A1(n15003), .A2(n14968), .A3(n14967), .ZN(n14970) );
  NAND2_X1 U18357 ( .A1(n14970), .A2(n14969), .ZN(n14971) );
  AOI211_X1 U18358 ( .C1(n14973), .C2(n20116), .A(n14972), .B(n14971), .ZN(
        n14974) );
  OAI21_X1 U18359 ( .B1(n14975), .B2(n20091), .A(n14974), .ZN(P1_U3005) );
  AOI21_X1 U18360 ( .B1(n14977), .B2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n14976), .ZN(n14979) );
  OAI211_X1 U18361 ( .C1(n14980), .C2(n20107), .A(n14979), .B(n14978), .ZN(
        n14981) );
  INV_X1 U18362 ( .A(n14981), .ZN(n14982) );
  OAI21_X1 U18363 ( .B1(n14983), .B2(n20091), .A(n14982), .ZN(P1_U3006) );
  INV_X1 U18364 ( .A(n14984), .ZN(n14996) );
  INV_X1 U18365 ( .A(n14985), .ZN(n14987) );
  AOI21_X1 U18366 ( .B1(n14987), .B2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n14986), .ZN(n14988) );
  OAI21_X1 U18367 ( .B1(n14990), .B2(n14989), .A(n14988), .ZN(n14991) );
  AOI21_X1 U18368 ( .B1(n14992), .B2(n20116), .A(n14991), .ZN(n14995) );
  NAND3_X1 U18369 ( .A1(n15003), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n14993), .ZN(n14994) );
  OAI211_X1 U18370 ( .C1(n14996), .C2(n20091), .A(n14995), .B(n14994), .ZN(
        P1_U3007) );
  AOI21_X1 U18371 ( .B1(n14998), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n14997), .ZN(n14999) );
  OAI21_X1 U18372 ( .B1(n15000), .B2(n20107), .A(n14999), .ZN(n15001) );
  AOI21_X1 U18373 ( .B1(n15003), .B2(n15002), .A(n15001), .ZN(n15004) );
  OAI21_X1 U18374 ( .B1(n15005), .B2(n20091), .A(n15004), .ZN(P1_U3008) );
  INV_X1 U18375 ( .A(n15006), .ZN(n15010) );
  NOR2_X1 U18376 ( .A1(n20100), .A2(n15007), .ZN(n15034) );
  AOI22_X1 U18377 ( .A1(n16207), .A2(n15008), .B1(n15035), .B2(n15034), .ZN(
        n15056) );
  NOR2_X1 U18378 ( .A1(n15056), .A2(n15009), .ZN(n15021) );
  AOI21_X1 U18379 ( .B1(n15010), .B2(n20122), .A(n15021), .ZN(n16170) );
  NOR2_X1 U18380 ( .A1(n16170), .A2(n15011), .ZN(n16162) );
  NAND2_X1 U18381 ( .A1(n16162), .A2(n15014), .ZN(n15013) );
  OAI211_X1 U18382 ( .C1(n16156), .C2(n15014), .A(n15013), .B(n15012), .ZN(
        n15015) );
  AOI21_X1 U18383 ( .B1(n15016), .B2(n20116), .A(n15015), .ZN(n15017) );
  OAI21_X1 U18384 ( .B1(n15018), .B2(n20091), .A(n15017), .ZN(P1_U3010) );
  INV_X1 U18385 ( .A(n15019), .ZN(n15029) );
  OAI21_X1 U18386 ( .B1(n15021), .B2(n20122), .A(n15020), .ZN(n15023) );
  INV_X1 U18387 ( .A(n16165), .ZN(n15022) );
  AOI21_X1 U18388 ( .B1(n15023), .B2(n15022), .A(n15024), .ZN(n15028) );
  NAND2_X1 U18389 ( .A1(n15024), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15026) );
  OAI21_X1 U18390 ( .B1(n16170), .B2(n15026), .A(n15025), .ZN(n15027) );
  AOI211_X1 U18391 ( .C1(n15029), .C2(n20116), .A(n15028), .B(n15027), .ZN(
        n15030) );
  OAI21_X1 U18392 ( .B1(n15031), .B2(n20091), .A(n15030), .ZN(P1_U3011) );
  NAND3_X1 U18393 ( .A1(n15032), .A2(n20117), .A3(n14800), .ZN(n15050) );
  INV_X1 U18394 ( .A(n15044), .ZN(n15042) );
  INV_X1 U18395 ( .A(n15052), .ZN(n15041) );
  AND2_X1 U18396 ( .A1(n15033), .A2(n16207), .ZN(n15040) );
  INV_X1 U18397 ( .A(n15034), .ZN(n15036) );
  OAI21_X1 U18398 ( .B1(n15055), .B2(n15036), .A(n15035), .ZN(n15038) );
  NAND2_X1 U18399 ( .A1(n15038), .A2(n15037), .ZN(n15039) );
  AOI211_X1 U18400 ( .C1(n20122), .C2(n15041), .A(n15040), .B(n15039), .ZN(
        n16197) );
  OAI21_X1 U18401 ( .B1(n15043), .B2(n15042), .A(n16197), .ZN(n16173) );
  NOR3_X1 U18402 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16199), .A3(
        n15044), .ZN(n15048) );
  OAI21_X1 U18403 ( .B1(n15046), .B2(n20107), .A(n15045), .ZN(n15047) );
  AOI211_X1 U18404 ( .C1(n16173), .C2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15048), .B(n15047), .ZN(n15049) );
  NAND2_X1 U18405 ( .A1(n15050), .A2(n15049), .ZN(P1_U3013) );
  NOR2_X1 U18406 ( .A1(n15052), .A2(n15051), .ZN(n15060) );
  OAI21_X1 U18407 ( .B1(n15054), .B2(n20107), .A(n15053), .ZN(n15058) );
  AOI21_X1 U18408 ( .B1(n15056), .B2(n15055), .A(n16197), .ZN(n15057) );
  AOI211_X1 U18409 ( .C1(n15060), .C2(n15059), .A(n15058), .B(n15057), .ZN(
        n15061) );
  OAI21_X1 U18410 ( .B1(n15062), .B2(n20091), .A(n15061), .ZN(P1_U3018) );
  OAI21_X1 U18411 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n20208), .A(n20658), 
        .ZN(n15063) );
  OAI21_X1 U18412 ( .B1(n15070), .B2(n20464), .A(n15063), .ZN(n15064) );
  MUX2_X1 U18413 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15064), .S(
        n20126), .Z(P1_U3477) );
  NOR2_X1 U18414 ( .A1(n13485), .A2(n15065), .ZN(n20602) );
  OAI22_X1 U18415 ( .A1(n20602), .A2(n20208), .B1(n20383), .B2(n20249), .ZN(
        n15067) );
  NAND2_X1 U18416 ( .A1(n15067), .A2(n20510), .ZN(n15068) );
  OAI211_X1 U18417 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n10999), .A(n15068), 
        .B(n20661), .ZN(n15069) );
  OAI21_X1 U18418 ( .B1(n15071), .B2(n15070), .A(n15069), .ZN(n15072) );
  MUX2_X1 U18419 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n15072), .S(
        n20126), .Z(P1_U3475) );
  OR2_X1 U18420 ( .A1(n20464), .A2(n15073), .ZN(n15080) );
  INV_X1 U18421 ( .A(n13188), .ZN(n15075) );
  INV_X1 U18422 ( .A(n13474), .ZN(n15074) );
  NAND3_X1 U18423 ( .A1(n15076), .A2(n15075), .A3(n15074), .ZN(n15077) );
  AND2_X1 U18424 ( .A1(n15078), .A2(n15077), .ZN(n15079) );
  AND2_X1 U18425 ( .A1(n15080), .A2(n15079), .ZN(n16023) );
  INV_X1 U18426 ( .A(n15081), .ZN(n15084) );
  NOR3_X1 U18427 ( .A1(n13474), .A2(n13188), .A3(n15089), .ZN(n15082) );
  AOI21_X1 U18428 ( .B1(n15084), .B2(n15083), .A(n15082), .ZN(n15085) );
  OAI21_X1 U18429 ( .B1(n16023), .B2(n15090), .A(n15085), .ZN(n15086) );
  MUX2_X1 U18430 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15086), .S(
        n16257), .Z(P1_U3473) );
  INV_X1 U18431 ( .A(n15087), .ZN(n15091) );
  OAI22_X1 U18432 ( .A1(n15091), .A2(n15090), .B1(n15089), .B2(n15088), .ZN(
        n15092) );
  MUX2_X1 U18433 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15092), .S(
        n16257), .Z(P1_U3469) );
  INV_X1 U18434 ( .A(n15093), .ZN(n15096) );
  NOR2_X1 U18435 ( .A1(n15094), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n15095) );
  MUX2_X1 U18436 ( .A(n15096), .B(n15095), .S(n19325), .Z(n15483) );
  INV_X1 U18437 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n21076) );
  NAND2_X1 U18438 ( .A1(n12076), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n15098) );
  NAND2_X1 U18439 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15097) );
  OAI211_X1 U18440 ( .C1(n15099), .C2(n21076), .A(n15098), .B(n15097), .ZN(
        n15100) );
  AOI21_X1 U18441 ( .B1(n15101), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n15100), .ZN(n15102) );
  NOR2_X1 U18442 ( .A1(n19098), .A2(n19090), .ZN(n19034) );
  XOR2_X1 U18443 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n15103), .Z(
        n15493) );
  AOI21_X1 U18444 ( .B1(n16272), .B2(n15105), .A(n15103), .ZN(n16271) );
  OR2_X1 U18445 ( .A1(n15107), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15104) );
  AND2_X1 U18446 ( .A1(n15105), .A2(n15104), .ZN(n15155) );
  INV_X1 U18447 ( .A(n15155), .ZN(n15523) );
  NOR2_X1 U18448 ( .A1(n15134), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15106) );
  OR2_X1 U18449 ( .A1(n15107), .A2(n15106), .ZN(n15179) );
  INV_X1 U18450 ( .A(n15179), .ZN(n15532) );
  AND2_X1 U18451 ( .A1(n15130), .A2(n15210), .ZN(n15108) );
  AOI21_X1 U18452 ( .B1(n15559), .B2(n15128), .A(n15131), .ZN(n15562) );
  AOI21_X1 U18453 ( .B1(n15126), .B2(n15577), .A(n15129), .ZN(n15580) );
  AOI21_X1 U18454 ( .B1(n18993), .B2(n15124), .A(n15127), .ZN(n18991) );
  AOI21_X1 U18455 ( .B1(n15109), .B2(n15122), .A(n15125), .ZN(n19005) );
  AOI21_X1 U18456 ( .B1(n15616), .B2(n15120), .A(n15123), .ZN(n19016) );
  AOI21_X1 U18457 ( .B1(n16354), .B2(n15118), .A(n15121), .ZN(n19044) );
  AOI21_X1 U18458 ( .B1(n16370), .B2(n15116), .A(n15119), .ZN(n16363) );
  AOI21_X1 U18459 ( .B1(n16392), .B2(n15114), .A(n15117), .ZN(n19069) );
  AOI21_X1 U18460 ( .B1(n16415), .B2(n15112), .A(n15110), .ZN(n19115) );
  NOR2_X1 U18461 ( .A1(n16416), .A2(n15111), .ZN(n15346) );
  OAI21_X1 U18462 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n15113), .A(
        n15112), .ZN(n19283) );
  NAND2_X1 U18463 ( .A1(n15346), .A2(n19283), .ZN(n19112) );
  NOR2_X1 U18464 ( .A1(n19115), .A2(n19112), .ZN(n19097) );
  NAND2_X1 U18465 ( .A1(n19097), .A2(n19099), .ZN(n19079) );
  NOR2_X1 U18466 ( .A1(n19080), .A2(n19079), .ZN(n15327) );
  OAI21_X1 U18467 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n15115), .A(
        n15114), .ZN(n16409) );
  NAND2_X1 U18468 ( .A1(n15327), .A2(n16409), .ZN(n19068) );
  NOR2_X1 U18469 ( .A1(n19069), .A2(n19068), .ZN(n19061) );
  OAI21_X1 U18470 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n15117), .A(
        n15116), .ZN(n19062) );
  NAND2_X1 U18471 ( .A1(n19061), .A2(n19062), .ZN(n15314) );
  NOR2_X1 U18472 ( .A1(n16363), .A2(n15314), .ZN(n15313) );
  OAI21_X1 U18473 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n15119), .A(
        n15118), .ZN(n19051) );
  NAND2_X1 U18474 ( .A1(n15313), .A2(n19051), .ZN(n19036) );
  NOR2_X1 U18475 ( .A1(n19044), .A2(n19036), .ZN(n19035) );
  OAI21_X1 U18476 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n15121), .A(
        n15120), .ZN(n19025) );
  NAND2_X1 U18477 ( .A1(n19035), .A2(n19025), .ZN(n19015) );
  NOR2_X1 U18478 ( .A1(n19016), .A2(n19015), .ZN(n15296) );
  OAI21_X1 U18479 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n15123), .A(
        n15122), .ZN(n15604) );
  NAND2_X1 U18480 ( .A1(n15296), .A2(n15604), .ZN(n19003) );
  NOR2_X1 U18481 ( .A1(n19005), .A2(n19003), .ZN(n15280) );
  OAI21_X1 U18482 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n15125), .A(
        n15124), .ZN(n16343) );
  NAND2_X1 U18483 ( .A1(n15280), .A2(n16343), .ZN(n18989) );
  NOR2_X1 U18484 ( .A1(n18991), .A2(n18989), .ZN(n18975) );
  OAI21_X1 U18485 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n15127), .A(
        n15126), .ZN(n18977) );
  NAND2_X1 U18486 ( .A1(n18975), .A2(n18977), .ZN(n15264) );
  NOR2_X1 U18487 ( .A1(n15580), .A2(n15264), .ZN(n15250) );
  OAI21_X1 U18488 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n15129), .A(
        n15128), .ZN(n16328) );
  NAND2_X1 U18489 ( .A1(n15250), .A2(n16328), .ZN(n15234) );
  NOR2_X1 U18490 ( .A1(n15562), .A2(n15234), .ZN(n15219) );
  OAI21_X1 U18491 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n15131), .A(
        n15130), .ZN(n16321) );
  NAND2_X1 U18492 ( .A1(n15219), .A2(n16321), .ZN(n15202) );
  NOR2_X1 U18493 ( .A1(n9791), .A2(n15202), .ZN(n15185) );
  NOR2_X1 U18494 ( .A1(n15132), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15133) );
  OR2_X1 U18495 ( .A1(n15134), .A2(n15133), .ZN(n15543) );
  NOR2_X1 U18496 ( .A1(n16271), .A2(n16270), .ZN(n16269) );
  NOR2_X1 U18497 ( .A1(n19098), .A2(n16269), .ZN(n15144) );
  NOR2_X1 U18498 ( .A1(n15493), .A2(n15144), .ZN(n15143) );
  NAND2_X1 U18499 ( .A1(n9719), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n15136) );
  AOI22_X1 U18500 ( .A1(n12312), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n12142), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15135) );
  NAND2_X1 U18501 ( .A1(n15136), .A2(n15135), .ZN(n15137) );
  XNOR2_X2 U18502 ( .A(n15138), .B(n15137), .ZN(n19168) );
  INV_X1 U18503 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n15139) );
  OAI22_X1 U18504 ( .A1(n19129), .A2(n21076), .B1(n15140), .B2(n15139), .ZN(
        n15141) );
  AOI21_X1 U18505 ( .B1(n19168), .B2(n19123), .A(n15141), .ZN(n15142) );
  AOI211_X1 U18506 ( .C1(n15493), .C2(n15144), .A(n15143), .B(n19090), .ZN(
        n15147) );
  INV_X1 U18507 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n15145) );
  OAI22_X1 U18508 ( .A1(n19109), .A2(n15145), .B1(n12346), .B2(n19129), .ZN(
        n15146) );
  AOI211_X1 U18509 ( .C1(n9717), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15147), .B(n15146), .ZN(n15151) );
  INV_X1 U18510 ( .A(n15497), .ZN(n15149) );
  AOI22_X1 U18511 ( .A1(n15149), .A2(n19133), .B1(n15148), .B2(n19123), .ZN(
        n15150) );
  OAI211_X1 U18512 ( .C1(n15152), .C2(n19107), .A(n15151), .B(n15150), .ZN(
        P2_U2825) );
  INV_X1 U18513 ( .A(n15153), .ZN(n15154) );
  AOI221_X1 U18514 ( .B1(n15155), .B2(n15154), .C1(n15523), .C2(n15153), .A(
        n19090), .ZN(n15167) );
  NOR2_X1 U18515 ( .A1(n15157), .A2(n15158), .ZN(n15159) );
  OR2_X1 U18516 ( .A1(n15174), .A2(n15160), .ZN(n15161) );
  AOI22_X1 U18517 ( .A1(n15656), .A2(n19123), .B1(P2_EBX_REG_28__SCAN_IN), 
        .B2(n19126), .ZN(n15165) );
  INV_X1 U18518 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15162) );
  OAI22_X1 U18519 ( .A1(n15162), .A2(n18992), .B1(n12332), .B2(n19129), .ZN(
        n15163) );
  INV_X1 U18520 ( .A(n15163), .ZN(n15164) );
  OAI211_X1 U18521 ( .C1(n15659), .C2(n19085), .A(n15165), .B(n15164), .ZN(
        n15166) );
  AOI211_X1 U18522 ( .C1(n15168), .C2(n19125), .A(n15167), .B(n15166), .ZN(
        n15169) );
  INV_X1 U18523 ( .A(n15169), .ZN(P2_U2827) );
  AOI21_X1 U18524 ( .B1(n15170), .B2(n10160), .A(n15157), .ZN(n15673) );
  INV_X1 U18525 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n15178) );
  AND2_X1 U18526 ( .A1(n15171), .A2(n15172), .ZN(n15173) );
  OR2_X1 U18527 ( .A1(n15174), .A2(n15173), .ZN(n15666) );
  INV_X1 U18528 ( .A(n15666), .ZN(n15176) );
  INV_X1 U18529 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15530) );
  OAI22_X1 U18530 ( .A1(n15530), .A2(n18992), .B1(n19871), .B2(n19129), .ZN(
        n15175) );
  AOI21_X1 U18531 ( .B1(n15176), .B2(n19123), .A(n15175), .ZN(n15177) );
  OAI21_X1 U18532 ( .B1(n19109), .B2(n15178), .A(n15177), .ZN(n15182) );
  AOI221_X1 U18533 ( .B1(n15532), .B2(n15180), .C1(n15179), .C2(n9884), .A(
        n19090), .ZN(n15181) );
  AOI211_X1 U18534 ( .C1(n19133), .C2(n15673), .A(n15182), .B(n15181), .ZN(
        n15183) );
  OAI21_X1 U18535 ( .B1(n15184), .B2(n19107), .A(n15183), .ZN(P2_U2828) );
  INV_X1 U18536 ( .A(n15543), .ZN(n15188) );
  NOR2_X1 U18537 ( .A1(n19098), .A2(n15185), .ZN(n15187) );
  OAI21_X1 U18538 ( .B1(n15188), .B2(n15187), .A(n19117), .ZN(n15186) );
  AOI21_X1 U18539 ( .B1(n15188), .B2(n15187), .A(n15186), .ZN(n15191) );
  OAI22_X1 U18540 ( .A1(n19109), .A2(n15189), .B1(n19869), .B2(n19129), .ZN(
        n15190) );
  AOI211_X1 U18541 ( .C1(n9717), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15191), .B(n15190), .ZN(n15199) );
  NAND2_X1 U18542 ( .A1(n15208), .A2(n15192), .ZN(n15193) );
  NAND2_X1 U18543 ( .A1(n10160), .A2(n15193), .ZN(n15678) );
  OR2_X1 U18544 ( .A1(n15195), .A2(n15194), .ZN(n15196) );
  NAND2_X1 U18545 ( .A1(n15171), .A2(n15196), .ZN(n15679) );
  OAI22_X1 U18546 ( .A1(n15678), .A2(n19085), .B1(n15679), .B2(n19121), .ZN(
        n15197) );
  INV_X1 U18547 ( .A(n15197), .ZN(n15198) );
  OAI211_X1 U18548 ( .C1(n15200), .C2(n19107), .A(n15199), .B(n15198), .ZN(
        P2_U2829) );
  MUX2_X1 U18549 ( .A(n10017), .B(P2_EBX_REG_25__SCAN_IN), .S(n15201), .Z(
        n15217) );
  AND2_X1 U18550 ( .A1(n9740), .A2(n15202), .ZN(n15204) );
  OAI21_X1 U18551 ( .B1(n9791), .B2(n15204), .A(n19117), .ZN(n15203) );
  AOI21_X1 U18552 ( .B1(n9791), .B2(n15204), .A(n15203), .ZN(n15205) );
  INV_X1 U18553 ( .A(n15205), .ZN(n15216) );
  OR2_X1 U18554 ( .A1(n15228), .A2(n15206), .ZN(n15207) );
  NAND2_X1 U18555 ( .A1(n15208), .A2(n15207), .ZN(n15550) );
  INV_X1 U18556 ( .A(n15550), .ZN(n15694) );
  XNOR2_X1 U18557 ( .A(n9773), .B(n15209), .ZN(n15692) );
  INV_X1 U18558 ( .A(n15692), .ZN(n15212) );
  OAI22_X1 U18559 ( .A1(n15210), .A2(n18992), .B1(n19867), .B2(n19129), .ZN(
        n15211) );
  AOI21_X1 U18560 ( .B1(n19123), .B2(n15212), .A(n15211), .ZN(n15213) );
  OAI21_X1 U18561 ( .B1(n19109), .B2(n10017), .A(n15213), .ZN(n15214) );
  AOI21_X1 U18562 ( .B1(n15694), .B2(n19133), .A(n15214), .ZN(n15215) );
  OAI211_X1 U18563 ( .C1(n15217), .C2(n19107), .A(n15216), .B(n15215), .ZN(
        P2_U2830) );
  MUX2_X1 U18564 ( .A(P2_EBX_REG_24__SCAN_IN), .B(n15223), .S(n15218), .Z(
        n15233) );
  INV_X1 U18565 ( .A(n16321), .ZN(n15222) );
  NOR2_X1 U18566 ( .A1(n19098), .A2(n15219), .ZN(n15221) );
  OAI21_X1 U18567 ( .B1(n15222), .B2(n15221), .A(n19117), .ZN(n15220) );
  AOI21_X1 U18568 ( .B1(n15222), .B2(n15221), .A(n15220), .ZN(n15225) );
  OAI22_X1 U18569 ( .A1(n19109), .A2(n15223), .B1(n9888), .B2(n18992), .ZN(
        n15224) );
  AOI211_X1 U18570 ( .C1(n19060), .C2(P2_REIP_REG_24__SCAN_IN), .A(n15225), 
        .B(n15224), .ZN(n15232) );
  AND2_X1 U18571 ( .A1(n15239), .A2(n15226), .ZN(n15227) );
  NOR2_X1 U18572 ( .A1(n15228), .A2(n15227), .ZN(n16317) );
  AND2_X1 U18573 ( .A1(n15243), .A2(n15229), .ZN(n15230) );
  NOR2_X1 U18574 ( .A1(n9773), .A2(n15230), .ZN(n15711) );
  AOI22_X1 U18575 ( .A1(n16317), .A2(n19133), .B1(n15711), .B2(n19123), .ZN(
        n15231) );
  OAI211_X1 U18576 ( .C1(n15233), .C2(n19107), .A(n15232), .B(n15231), .ZN(
        P2_U2831) );
  NAND2_X1 U18577 ( .A1(n9740), .A2(n15234), .ZN(n15235) );
  XNOR2_X1 U18578 ( .A(n15562), .B(n15235), .ZN(n15236) );
  AOI22_X1 U18579 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n9717), .B1(
        n19117), .B2(n15236), .ZN(n15248) );
  NAND2_X1 U18580 ( .A1(n15257), .A2(n15237), .ZN(n15238) );
  NAND2_X1 U18581 ( .A1(n15239), .A2(n15238), .ZN(n16282) );
  INV_X1 U18582 ( .A(n16282), .ZN(n15246) );
  NAND2_X1 U18583 ( .A1(n15240), .A2(n15241), .ZN(n15242) );
  AND2_X1 U18584 ( .A1(n15243), .A2(n15242), .ZN(n15719) );
  INV_X1 U18585 ( .A(n15719), .ZN(n15470) );
  AOI22_X1 U18586 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(n19126), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19060), .ZN(n15244) );
  OAI21_X1 U18587 ( .B1(n19121), .B2(n15470), .A(n15244), .ZN(n15245) );
  AOI21_X1 U18588 ( .B1(n15246), .B2(n19133), .A(n15245), .ZN(n15247) );
  OAI211_X1 U18589 ( .C1(n15249), .C2(n19107), .A(n15248), .B(n15247), .ZN(
        P2_U2832) );
  NOR2_X1 U18590 ( .A1(n19098), .A2(n15250), .ZN(n15251) );
  XOR2_X1 U18591 ( .A(n16328), .B(n15251), .Z(n15253) );
  AOI22_X1 U18592 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n19126), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19060), .ZN(n15252) );
  OAI21_X1 U18593 ( .B1(n19090), .B2(n15253), .A(n15252), .ZN(n15254) );
  AOI21_X1 U18594 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n9717), .A(
        n15254), .ZN(n15262) );
  INV_X1 U18595 ( .A(n15255), .ZN(n15258) );
  OAI21_X1 U18596 ( .B1(n15258), .B2(n10131), .A(n15257), .ZN(n16290) );
  INV_X1 U18597 ( .A(n16290), .ZN(n16324) );
  OAI21_X1 U18598 ( .B1(n15260), .B2(n15259), .A(n15240), .ZN(n15737) );
  INV_X1 U18599 ( .A(n15737), .ZN(n16299) );
  AOI22_X1 U18600 ( .A1(n16324), .A2(n19133), .B1(n16299), .B2(n19123), .ZN(
        n15261) );
  OAI211_X1 U18601 ( .C1(n15263), .C2(n19107), .A(n15262), .B(n15261), .ZN(
        P2_U2833) );
  AND2_X1 U18602 ( .A1(n9740), .A2(n15264), .ZN(n15266) );
  OAI21_X1 U18603 ( .B1(n15580), .B2(n15266), .A(n19117), .ZN(n15265) );
  AOI21_X1 U18604 ( .B1(n15580), .B2(n15266), .A(n15265), .ZN(n15269) );
  AOI22_X1 U18605 ( .A1(n19126), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n19060), .ZN(n15267) );
  INV_X1 U18606 ( .A(n15267), .ZN(n15268) );
  AOI211_X1 U18607 ( .C1(n9717), .C2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15269), .B(n15268), .ZN(n15277) );
  OR2_X1 U18608 ( .A1(n15764), .A2(n15270), .ZN(n15271) );
  NAND2_X1 U18609 ( .A1(n15255), .A2(n15271), .ZN(n15745) );
  OR2_X1 U18610 ( .A1(n15272), .A2(n15765), .ZN(n15274) );
  INV_X1 U18611 ( .A(n15259), .ZN(n15273) );
  AND2_X1 U18612 ( .A1(n15274), .A2(n15273), .ZN(n15742) );
  INV_X1 U18613 ( .A(n15742), .ZN(n15475) );
  OAI22_X1 U18614 ( .A1(n15745), .A2(n19085), .B1(n15475), .B2(n19121), .ZN(
        n15275) );
  INV_X1 U18615 ( .A(n15275), .ZN(n15276) );
  OAI211_X1 U18616 ( .C1(n15278), .C2(n19107), .A(n15277), .B(n15276), .ZN(
        P2_U2834) );
  INV_X1 U18617 ( .A(n15279), .ZN(n15295) );
  NOR2_X1 U18618 ( .A1(n19098), .A2(n15280), .ZN(n15281) );
  XNOR2_X1 U18619 ( .A(n15281), .B(n16343), .ZN(n15282) );
  NAND2_X1 U18620 ( .A1(n15282), .A2(n19117), .ZN(n15294) );
  AOI21_X1 U18621 ( .B1(n13958), .B2(n15283), .A(n14019), .ZN(n16433) );
  NAND2_X1 U18622 ( .A1(n19123), .A2(n16433), .ZN(n15286) );
  AOI21_X1 U18623 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n9717), .A(
        n19276), .ZN(n15285) );
  OAI211_X1 U18624 ( .C1(n19129), .C2(n15287), .A(n15286), .B(n15285), .ZN(
        n15292) );
  NAND2_X1 U18625 ( .A1(n13726), .A2(n15289), .ZN(n15290) );
  NAND2_X1 U18626 ( .A1(n15431), .A2(n15290), .ZN(n16341) );
  NOR2_X1 U18627 ( .A1(n16341), .A2(n19085), .ZN(n15291) );
  AOI211_X1 U18628 ( .C1(P2_EBX_REG_18__SCAN_IN), .C2(n19126), .A(n15292), .B(
        n15291), .ZN(n15293) );
  OAI211_X1 U18629 ( .C1(n19107), .C2(n15295), .A(n15294), .B(n15293), .ZN(
        P2_U2837) );
  NOR2_X1 U18630 ( .A1(n19098), .A2(n15296), .ZN(n15297) );
  XNOR2_X1 U18631 ( .A(n15297), .B(n15604), .ZN(n15298) );
  NAND2_X1 U18632 ( .A1(n15298), .A2(n19117), .ZN(n15311) );
  AND2_X1 U18633 ( .A1(n16443), .A2(n15299), .ZN(n15300) );
  NOR2_X1 U18634 ( .A1(n9808), .A2(n15300), .ZN(n19175) );
  NAND2_X1 U18635 ( .A1(n19123), .A2(n19175), .ZN(n15302) );
  AOI21_X1 U18636 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n9717), .A(
        n19276), .ZN(n15301) );
  OAI211_X1 U18637 ( .C1(n19129), .C2(n19856), .A(n15302), .B(n15301), .ZN(
        n15309) );
  INV_X1 U18638 ( .A(n15303), .ZN(n15307) );
  NAND2_X1 U18639 ( .A1(n15305), .A2(n15304), .ZN(n15306) );
  NAND2_X1 U18640 ( .A1(n15307), .A2(n15306), .ZN(n19142) );
  NOR2_X1 U18641 ( .A1(n19142), .A2(n19085), .ZN(n15308) );
  AOI211_X1 U18642 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n19126), .A(n15309), .B(
        n15308), .ZN(n15310) );
  OAI211_X1 U18643 ( .C1(n19107), .C2(n15312), .A(n15311), .B(n15310), .ZN(
        P2_U2839) );
  NOR2_X1 U18644 ( .A1(n9740), .A2(n19090), .ZN(n19134) );
  NOR2_X1 U18645 ( .A1(n19098), .A2(n15313), .ZN(n19052) );
  AOI21_X1 U18646 ( .B1(n16363), .B2(n15314), .A(n19090), .ZN(n15315) );
  AOI22_X1 U18647 ( .A1(n16363), .A2(n19134), .B1(n19052), .B2(n15315), .ZN(
        n15326) );
  OAI22_X1 U18648 ( .A1(n19109), .A2(n11781), .B1(n16370), .B2(n18992), .ZN(
        n15316) );
  AOI211_X1 U18649 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n19060), .A(n19276), 
        .B(n15316), .ZN(n15325) );
  OR2_X1 U18650 ( .A1(n15318), .A2(n15317), .ZN(n15320) );
  NAND2_X1 U18651 ( .A1(n15320), .A2(n15319), .ZN(n19193) );
  OAI22_X1 U18652 ( .A1(n15321), .A2(n19085), .B1(n19193), .B2(n19121), .ZN(
        n15322) );
  AOI21_X1 U18653 ( .B1(n15323), .B2(n19125), .A(n15322), .ZN(n15324) );
  NAND3_X1 U18654 ( .A1(n15326), .A2(n15325), .A3(n15324), .ZN(P2_U2844) );
  NOR2_X1 U18655 ( .A1(n19098), .A2(n15327), .ZN(n15328) );
  XNOR2_X1 U18656 ( .A(n15328), .B(n16409), .ZN(n15329) );
  NAND2_X1 U18657 ( .A1(n15329), .A2(n19117), .ZN(n15344) );
  OR2_X1 U18658 ( .A1(n15330), .A2(n12994), .ZN(n15332) );
  NAND2_X1 U18659 ( .A1(n15332), .A2(n15331), .ZN(n19162) );
  NAND2_X1 U18660 ( .A1(n19126), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n15333) );
  OAI21_X1 U18661 ( .B1(n19085), .B2(n19162), .A(n15333), .ZN(n15342) );
  AOI21_X1 U18662 ( .B1(n15336), .B2(n15334), .A(n15335), .ZN(n19202) );
  NAND2_X1 U18663 ( .A1(n19123), .A2(n19202), .ZN(n15339) );
  AND2_X1 U18664 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n9717), .ZN(
        n15337) );
  NOR2_X1 U18665 ( .A1(n19276), .A2(n15337), .ZN(n15338) );
  OAI211_X1 U18666 ( .C1(n19129), .C2(n15340), .A(n15339), .B(n15338), .ZN(
        n15341) );
  NOR2_X1 U18667 ( .A1(n15342), .A2(n15341), .ZN(n15343) );
  OAI211_X1 U18668 ( .C1(n19107), .C2(n15345), .A(n15344), .B(n15343), .ZN(
        P2_U2847) );
  NOR2_X1 U18669 ( .A1(n19098), .A2(n15346), .ZN(n15347) );
  XNOR2_X1 U18670 ( .A(n15347), .B(n19283), .ZN(n15365) );
  NAND2_X1 U18671 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15348), .ZN(
        n15349) );
  AND2_X1 U18672 ( .A1(n15350), .A2(n15349), .ZN(n15354) );
  INV_X1 U18673 ( .A(n15351), .ZN(n15352) );
  NAND3_X1 U18674 ( .A1(n15354), .A2(n15353), .A3(n15352), .ZN(n15355) );
  NAND2_X1 U18675 ( .A1(n15356), .A2(n15355), .ZN(n19218) );
  NOR2_X1 U18676 ( .A1(n19218), .A2(n19130), .ZN(n15364) );
  AOI21_X1 U18677 ( .B1(P2_REIP_REG_4__SCAN_IN), .B2(n19060), .A(n19276), .ZN(
        n15359) );
  AOI22_X1 U18678 ( .A1(n19126), .A2(P2_EBX_REG_4__SCAN_IN), .B1(n19125), .B2(
        n15357), .ZN(n15358) );
  OAI211_X1 U18679 ( .C1(n19121), .C2(n15360), .A(n15359), .B(n15358), .ZN(
        n15361) );
  AOI21_X1 U18680 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n9717), .A(
        n15361), .ZN(n15362) );
  OAI21_X1 U18681 ( .B1(n19085), .B2(n19277), .A(n15362), .ZN(n15363) );
  AOI211_X1 U18682 ( .C1(n15365), .C2(n19117), .A(n15364), .B(n15363), .ZN(
        n15366) );
  INV_X1 U18683 ( .A(n15366), .ZN(P2_U2851) );
  NOR2_X1 U18684 ( .A1(n19098), .A2(n15376), .ZN(n15367) );
  XNOR2_X1 U18685 ( .A(n15367), .B(n19292), .ZN(n15368) );
  NAND2_X1 U18686 ( .A1(n15368), .A2(n19117), .ZN(n15375) );
  AOI22_X1 U18687 ( .A1(n19060), .A2(P2_REIP_REG_2__SCAN_IN), .B1(n19126), 
        .B2(P2_EBX_REG_2__SCAN_IN), .ZN(n15369) );
  OAI21_X1 U18688 ( .B1(n15370), .B2(n19107), .A(n15369), .ZN(n15373) );
  INV_X1 U18689 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n15371) );
  OAI22_X1 U18690 ( .A1(n19905), .A2(n19121), .B1(n15371), .B2(n18992), .ZN(
        n15372) );
  AOI211_X1 U18691 ( .C1(n19133), .C2(n19295), .A(n15373), .B(n15372), .ZN(
        n15374) );
  OAI211_X1 U18692 ( .C1(n19210), .C2(n19130), .A(n15375), .B(n15374), .ZN(
        P2_U2853) );
  AOI211_X1 U18693 ( .C1(n15378), .C2(n15377), .A(n19098), .B(n15376), .ZN(
        n15933) );
  NAND2_X1 U18694 ( .A1(n15933), .A2(n19117), .ZN(n15387) );
  AOI22_X1 U18695 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(n19126), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n9717), .ZN(n15380) );
  NAND2_X1 U18696 ( .A1(n15623), .A2(n19134), .ZN(n15379) );
  OAI211_X1 U18697 ( .C1(n19107), .C2(n15381), .A(n15380), .B(n15379), .ZN(
        n15382) );
  AOI21_X1 U18698 ( .B1(P2_REIP_REG_1__SCAN_IN), .B2(n19060), .A(n15382), .ZN(
        n15383) );
  OAI21_X1 U18699 ( .B1(n19121), .B2(n15384), .A(n15383), .ZN(n15385) );
  AOI21_X1 U18700 ( .B1(n15917), .B2(n19133), .A(n15385), .ZN(n15386) );
  OAI211_X1 U18701 ( .C1(n19915), .C2(n19130), .A(n15387), .B(n15386), .ZN(
        P2_U2854) );
  NAND2_X1 U18702 ( .A1(n15390), .A2(n15389), .ZN(n16275) );
  INV_X1 U18703 ( .A(n14343), .ZN(n15392) );
  NAND3_X1 U18704 ( .A1(n15392), .A2(n19151), .A3(n15391), .ZN(n15394) );
  NAND2_X1 U18705 ( .A1(n19161), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15393) );
  NAND2_X1 U18706 ( .A1(n14264), .A2(n15395), .ZN(n15397) );
  XNOR2_X1 U18707 ( .A(n15397), .B(n15396), .ZN(n15440) );
  NOR2_X1 U18708 ( .A1(n15659), .A2(n19161), .ZN(n15398) );
  AOI21_X1 U18709 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n19161), .A(n15398), .ZN(
        n15399) );
  OAI21_X1 U18710 ( .B1(n15440), .B2(n19165), .A(n15399), .ZN(P2_U2859) );
  INV_X1 U18711 ( .A(n15673), .ZN(n15405) );
  AOI21_X1 U18712 ( .B1(n15400), .B2(n15402), .A(n15401), .ZN(n15445) );
  NAND2_X1 U18713 ( .A1(n15445), .A2(n19151), .ZN(n15404) );
  NAND2_X1 U18714 ( .A1(n19161), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15403) );
  OAI211_X1 U18715 ( .C1(n15405), .C2(n19161), .A(n15404), .B(n15403), .ZN(
        P2_U2860) );
  AOI21_X1 U18716 ( .B1(n15407), .B2(n15410), .A(n15409), .ZN(n15450) );
  NAND2_X1 U18717 ( .A1(n15450), .A2(n19151), .ZN(n15412) );
  NAND2_X1 U18718 ( .A1(n19161), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15411) );
  OAI211_X1 U18719 ( .C1(n15678), .C2(n19161), .A(n15412), .B(n15411), .ZN(
        P2_U2861) );
  OAI21_X1 U18720 ( .B1(n15413), .B2(n15415), .A(n15414), .ZN(n15456) );
  NOR2_X1 U18721 ( .A1(n15550), .A2(n19161), .ZN(n15416) );
  AOI21_X1 U18722 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n19161), .A(n15416), .ZN(
        n15417) );
  OAI21_X1 U18723 ( .B1(n15456), .B2(n19165), .A(n15417), .ZN(P2_U2862) );
  AOI21_X1 U18724 ( .B1(n15418), .B2(n15419), .A(n9757), .ZN(n15420) );
  XOR2_X1 U18725 ( .A(n15421), .B(n15420), .Z(n15462) );
  NAND2_X1 U18726 ( .A1(n19161), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n15423) );
  NAND2_X1 U18727 ( .A1(n16317), .A2(n19164), .ZN(n15422) );
  OAI211_X1 U18728 ( .C1(n15462), .C2(n19165), .A(n15423), .B(n15422), .ZN(
        P2_U2863) );
  OAI21_X1 U18729 ( .B1(n15424), .B2(n15427), .A(n15426), .ZN(n15478) );
  NOR2_X1 U18730 ( .A1(n15745), .A2(n19161), .ZN(n15428) );
  AOI21_X1 U18731 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n19161), .A(n15428), .ZN(
        n15429) );
  OAI21_X1 U18732 ( .B1(n15478), .B2(n19165), .A(n15429), .ZN(P2_U2866) );
  AND2_X1 U18733 ( .A1(n15431), .A2(n15430), .ZN(n15432) );
  OR2_X1 U18734 ( .A1(n15432), .A2(n9751), .ZN(n18998) );
  NOR2_X1 U18735 ( .A1(n18998), .A2(n19161), .ZN(n15433) );
  AOI21_X1 U18736 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19161), .A(n15433), .ZN(
        n15434) );
  OAI21_X1 U18737 ( .B1(n15435), .B2(n19165), .A(n15434), .ZN(P2_U2868) );
  INV_X1 U18738 ( .A(n19189), .ZN(n15436) );
  OAI22_X1 U18739 ( .A1(n15458), .A2(n15436), .B1(n19205), .B2(n20977), .ZN(
        n15437) );
  AOI21_X1 U18740 ( .B1(n19232), .B2(n15656), .A(n15437), .ZN(n15439) );
  AOI22_X1 U18741 ( .A1(n19174), .A2(BUF2_REG_28__SCAN_IN), .B1(n19173), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15438) );
  OAI211_X1 U18742 ( .C1(n15440), .C2(n19236), .A(n15439), .B(n15438), .ZN(
        P2_U2891) );
  AOI22_X1 U18743 ( .A1(n19174), .A2(BUF2_REG_27__SCAN_IN), .B1(n19173), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15443) );
  AOI22_X1 U18744 ( .A1(n19172), .A2(n15441), .B1(n19231), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n15442) );
  OAI211_X1 U18745 ( .C1(n19180), .C2(n15666), .A(n15443), .B(n15442), .ZN(
        n15444) );
  AOI21_X1 U18746 ( .B1(n15445), .B2(n19219), .A(n15444), .ZN(n15446) );
  INV_X1 U18747 ( .A(n15446), .ZN(P2_U2892) );
  AOI22_X1 U18748 ( .A1(n19174), .A2(BUF2_REG_26__SCAN_IN), .B1(n19173), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15448) );
  AOI22_X1 U18749 ( .A1(n19172), .A2(n19194), .B1(n19231), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15447) );
  OAI211_X1 U18750 ( .C1(n19180), .C2(n15679), .A(n15448), .B(n15447), .ZN(
        n15449) );
  AOI21_X1 U18751 ( .B1(n15450), .B2(n19219), .A(n15449), .ZN(n15451) );
  INV_X1 U18752 ( .A(n15451), .ZN(P2_U2893) );
  AOI22_X1 U18753 ( .A1(n19174), .A2(BUF2_REG_25__SCAN_IN), .B1(n19173), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15453) );
  AOI22_X1 U18754 ( .A1(n19172), .A2(n19197), .B1(n19231), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n15452) );
  OAI211_X1 U18755 ( .C1(n15692), .C2(n19180), .A(n15453), .B(n15452), .ZN(
        n15454) );
  INV_X1 U18756 ( .A(n15454), .ZN(n15455) );
  OAI21_X1 U18757 ( .B1(n15456), .B2(n19236), .A(n15455), .ZN(P2_U2894) );
  INV_X1 U18758 ( .A(n19200), .ZN(n15457) );
  OAI22_X1 U18759 ( .A1(n15458), .A2(n15457), .B1(n19205), .B2(n12850), .ZN(
        n15459) );
  AOI21_X1 U18760 ( .B1(n19232), .B2(n15711), .A(n15459), .ZN(n15461) );
  AOI22_X1 U18761 ( .A1(n19174), .A2(BUF2_REG_24__SCAN_IN), .B1(n19173), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15460) );
  OAI211_X1 U18762 ( .C1(n15462), .C2(n19236), .A(n15461), .B(n15460), .ZN(
        P2_U2895) );
  NOR2_X1 U18763 ( .A1(n15463), .A2(n15464), .ZN(n15466) );
  NOR2_X1 U18764 ( .A1(n15466), .A2(n15465), .ZN(n16284) );
  AOI22_X1 U18765 ( .A1(n19174), .A2(BUF2_REG_23__SCAN_IN), .B1(n19173), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n15469) );
  AOI22_X1 U18766 ( .A1(n19172), .A2(n15467), .B1(n19231), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n15468) );
  OAI211_X1 U18767 ( .C1(n19180), .C2(n15470), .A(n15469), .B(n15468), .ZN(
        n15471) );
  AOI21_X1 U18768 ( .B1(n16284), .B2(n19219), .A(n15471), .ZN(n15472) );
  INV_X1 U18769 ( .A(n15472), .ZN(P2_U2896) );
  AOI22_X1 U18770 ( .A1(n19174), .A2(BUF2_REG_21__SCAN_IN), .B1(n19173), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n15474) );
  AOI22_X1 U18771 ( .A1(n19172), .A2(n19208), .B1(n19231), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15473) );
  OAI211_X1 U18772 ( .C1(n19180), .C2(n15475), .A(n15474), .B(n15473), .ZN(
        n15476) );
  INV_X1 U18773 ( .A(n15476), .ZN(n15477) );
  OAI21_X1 U18774 ( .B1(n15478), .B2(n19236), .A(n15477), .ZN(P2_U2898) );
  INV_X1 U18775 ( .A(n15502), .ZN(n15479) );
  NAND2_X1 U18776 ( .A1(n15483), .A2(n11763), .ZN(n15484) );
  XNOR2_X1 U18777 ( .A(n15484), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15485) );
  XNOR2_X1 U18778 ( .A(n15486), .B(n15485), .ZN(n15640) );
  NAND2_X1 U18779 ( .A1(n15508), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15487) );
  XNOR2_X1 U18780 ( .A(n15487), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15638) );
  NOR2_X1 U18781 ( .A1(n15488), .A2(n19291), .ZN(n15491) );
  NAND2_X1 U18782 ( .A1(n19276), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n15632) );
  NAND2_X1 U18783 ( .A1(n19284), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15489) );
  OAI211_X1 U18784 ( .C1(n16281), .C2(n13674), .A(n15632), .B(n15489), .ZN(
        n15490) );
  AOI211_X1 U18785 ( .C1(n15638), .C2(n19288), .A(n15491), .B(n15490), .ZN(
        n15492) );
  OAI21_X1 U18786 ( .B1(n15640), .B2(n16421), .A(n15492), .ZN(P2_U2983) );
  NAND2_X1 U18787 ( .A1(n15493), .A2(n16417), .ZN(n15496) );
  AOI21_X1 U18788 ( .B1(n19284), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15494), .ZN(n15495) );
  OAI211_X1 U18789 ( .C1(n13674), .C2(n15497), .A(n15496), .B(n15495), .ZN(
        n15498) );
  AOI21_X1 U18790 ( .B1(n15499), .B2(n19288), .A(n15498), .ZN(n15500) );
  OAI21_X1 U18791 ( .B1(n15501), .B2(n16421), .A(n15500), .ZN(P2_U2984) );
  NAND2_X1 U18792 ( .A1(n15503), .A2(n15502), .ZN(n15505) );
  XOR2_X1 U18793 ( .A(n15505), .B(n15504), .Z(n15653) );
  INV_X1 U18794 ( .A(n15506), .ZN(n15507) );
  AOI21_X1 U18795 ( .B1(n15507), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15509) );
  NOR2_X1 U18796 ( .A1(n15509), .A2(n15508), .ZN(n15651) );
  NAND2_X1 U18797 ( .A1(n16271), .A2(n16417), .ZN(n15511) );
  NOR2_X1 U18798 ( .A1(n9725), .A2(n19873), .ZN(n15645) );
  AOI21_X1 U18799 ( .B1(n19284), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15645), .ZN(n15510) );
  OAI211_X1 U18800 ( .C1(n13674), .C2(n16275), .A(n15511), .B(n15510), .ZN(
        n15512) );
  AOI21_X1 U18801 ( .B1(n15651), .B2(n19288), .A(n15512), .ZN(n15513) );
  OAI21_X1 U18802 ( .B1(n15653), .B2(n16421), .A(n15513), .ZN(P2_U2985) );
  XNOR2_X1 U18803 ( .A(n15516), .B(n15518), .ZN(n15528) );
  INV_X1 U18804 ( .A(n15516), .ZN(n15517) );
  AOI22_X1 U18805 ( .A1(n15528), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n15518), .B2(n15517), .ZN(n15522) );
  XNOR2_X1 U18806 ( .A(n15520), .B(n15519), .ZN(n15521) );
  XNOR2_X1 U18807 ( .A(n15522), .B(n15521), .ZN(n15664) );
  XNOR2_X1 U18808 ( .A(n15506), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15662) );
  NOR2_X1 U18809 ( .A1(n15523), .A2(n19291), .ZN(n15526) );
  NAND2_X1 U18810 ( .A1(n19276), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15654) );
  NAND2_X1 U18811 ( .A1(n19284), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15524) );
  OAI211_X1 U18812 ( .C1(n15659), .C2(n13674), .A(n15654), .B(n15524), .ZN(
        n15525) );
  AOI211_X1 U18813 ( .C1(n15662), .C2(n19288), .A(n15526), .B(n15525), .ZN(
        n15527) );
  OAI21_X1 U18814 ( .B1(n15664), .B2(n16421), .A(n15527), .ZN(P2_U2986) );
  XNOR2_X1 U18815 ( .A(n15528), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15677) );
  NAND2_X1 U18816 ( .A1(n15673), .A2(n19294), .ZN(n15529) );
  NAND2_X1 U18817 ( .A1(n19276), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15665) );
  OAI211_X1 U18818 ( .C1(n16428), .C2(n15530), .A(n15529), .B(n15665), .ZN(
        n15531) );
  AOI21_X1 U18819 ( .B1(n16417), .B2(n15532), .A(n15531), .ZN(n15534) );
  OR2_X1 U18820 ( .A1(n15540), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15674) );
  NAND3_X1 U18821 ( .A1(n15674), .A2(n19288), .A3(n15506), .ZN(n15533) );
  OAI211_X1 U18822 ( .C1(n15677), .C2(n16421), .A(n15534), .B(n15533), .ZN(
        P2_U2987) );
  AOI21_X1 U18823 ( .B1(n15535), .B2(n15547), .A(n15546), .ZN(n15536) );
  XOR2_X1 U18824 ( .A(n15537), .B(n15536), .Z(n15689) );
  AND2_X1 U18825 ( .A1(n15551), .A2(n15538), .ZN(n15539) );
  NOR2_X1 U18826 ( .A1(n15540), .A2(n15539), .ZN(n15687) );
  NOR2_X1 U18827 ( .A1(n9725), .A2(n19869), .ZN(n15681) );
  NOR2_X1 U18828 ( .A1(n15678), .A2(n13674), .ZN(n15541) );
  AOI211_X1 U18829 ( .C1(n19284), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15681), .B(n15541), .ZN(n15542) );
  OAI21_X1 U18830 ( .B1(n19291), .B2(n15543), .A(n15542), .ZN(n15544) );
  AOI21_X1 U18831 ( .B1(n15687), .B2(n19288), .A(n15544), .ZN(n15545) );
  OAI21_X1 U18832 ( .B1(n15689), .B2(n16421), .A(n15545), .ZN(P2_U2988) );
  NAND2_X1 U18833 ( .A1(n10143), .A2(n15547), .ZN(n15548) );
  XNOR2_X1 U18834 ( .A(n15535), .B(n15548), .ZN(n15702) );
  NAND2_X1 U18835 ( .A1(n19276), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15691) );
  NAND2_X1 U18836 ( .A1(n19284), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15549) );
  OAI211_X1 U18837 ( .C1(n15550), .C2(n13674), .A(n15691), .B(n15549), .ZN(
        n15554) );
  INV_X1 U18838 ( .A(n15708), .ZN(n15552) );
  OAI21_X1 U18839 ( .B1(n15552), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15551), .ZN(n15690) );
  NOR2_X1 U18840 ( .A1(n15690), .A2(n16418), .ZN(n15553) );
  AOI211_X1 U18841 ( .C1(n16417), .C2(n9791), .A(n15554), .B(n15553), .ZN(
        n15555) );
  OAI21_X1 U18842 ( .B1(n15702), .B2(n16421), .A(n15555), .ZN(P2_U2989) );
  NOR2_X1 U18843 ( .A1(n15556), .A2(n15735), .ZN(n15732) );
  OAI21_X1 U18844 ( .B1(n15732), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15706), .ZN(n15727) );
  XOR2_X1 U18845 ( .A(n15558), .B(n15557), .Z(n15718) );
  NAND2_X1 U18846 ( .A1(n15718), .A2(n19285), .ZN(n15564) );
  OAI22_X1 U18847 ( .A1(n16428), .A2(n15559), .B1(n12060), .B2(n9725), .ZN(
        n15561) );
  NOR2_X1 U18848 ( .A1(n16282), .A2(n13674), .ZN(n15560) );
  AOI211_X1 U18849 ( .C1(n15562), .C2(n16417), .A(n15561), .B(n15560), .ZN(
        n15563) );
  OAI211_X1 U18850 ( .C1(n16418), .C2(n15727), .A(n15564), .B(n15563), .ZN(
        P2_U2991) );
  OAI21_X1 U18851 ( .B1(n15565), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15556), .ZN(n15752) );
  NAND2_X1 U18852 ( .A1(n15567), .A2(n15566), .ZN(n15576) );
  INV_X1 U18853 ( .A(n15813), .ZN(n15569) );
  INV_X1 U18854 ( .A(n15612), .ZN(n15570) );
  NAND2_X1 U18855 ( .A1(n15603), .A2(n15602), .ZN(n15601) );
  INV_X1 U18856 ( .A(n15593), .ZN(n15572) );
  XOR2_X1 U18857 ( .A(n15576), .B(n15575), .Z(n15741) );
  NAND2_X1 U18858 ( .A1(n15741), .A2(n19285), .ZN(n15582) );
  NAND2_X1 U18859 ( .A1(n19276), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15744) );
  OAI21_X1 U18860 ( .B1(n16428), .B2(n15577), .A(n15744), .ZN(n15579) );
  NOR2_X1 U18861 ( .A1(n15745), .A2(n13674), .ZN(n15578) );
  AOI211_X1 U18862 ( .C1(n16417), .C2(n15580), .A(n15579), .B(n15578), .ZN(
        n15581) );
  OAI211_X1 U18863 ( .C1(n16418), .C2(n15752), .A(n15582), .B(n15581), .ZN(
        P2_U2993) );
  INV_X1 U18864 ( .A(n15583), .ZN(n15584) );
  NAND2_X1 U18865 ( .A1(n15585), .A2(n15584), .ZN(n15587) );
  AOI21_X1 U18866 ( .B1(n16338), .B2(n16337), .A(n16335), .ZN(n15586) );
  XOR2_X1 U18867 ( .A(n15587), .B(n15586), .Z(n15787) );
  OAI22_X1 U18868 ( .A1(n16428), .A2(n18993), .B1(n12047), .B2(n9725), .ZN(
        n15589) );
  NOR2_X1 U18869 ( .A1(n18998), .A2(n13674), .ZN(n15588) );
  AOI211_X1 U18870 ( .C1(n18991), .C2(n16417), .A(n15589), .B(n15588), .ZN(
        n15592) );
  XNOR2_X1 U18871 ( .A(n15590), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15785) );
  NAND2_X1 U18872 ( .A1(n15785), .A2(n19288), .ZN(n15591) );
  OAI211_X1 U18873 ( .C1(n15787), .C2(n16421), .A(n15592), .B(n15591), .ZN(
        P2_U2995) );
  NAND2_X1 U18874 ( .A1(n15594), .A2(n15593), .ZN(n15596) );
  XOR2_X1 U18875 ( .A(n15596), .B(n15595), .Z(n15805) );
  NAND2_X1 U18876 ( .A1(n19276), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15788) );
  NAND2_X1 U18877 ( .A1(n19284), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15597) );
  OAI211_X1 U18878 ( .C1(n19009), .C2(n13674), .A(n15788), .B(n15597), .ZN(
        n15600) );
  INV_X1 U18879 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15889) );
  OAI21_X1 U18880 ( .B1(n15603), .B2(n15602), .A(n15601), .ZN(n15812) );
  NOR2_X1 U18881 ( .A1(n19142), .A2(n13674), .ZN(n15606) );
  OAI22_X1 U18882 ( .A1(n19856), .A2(n9725), .B1(n19291), .B2(n15604), .ZN(
        n15605) );
  AOI211_X1 U18883 ( .C1(n19284), .C2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n15606), .B(n15605), .ZN(n15610) );
  NOR2_X1 U18884 ( .A1(n15789), .A2(n16446), .ZN(n15608) );
  INV_X1 U18885 ( .A(n16339), .ZN(n15607) );
  OAI211_X1 U18886 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15608), .A(
        n15607), .B(n19288), .ZN(n15609) );
  OAI211_X1 U18887 ( .C1(n15812), .C2(n16421), .A(n15610), .B(n15609), .ZN(
        P2_U2998) );
  NAND2_X1 U18888 ( .A1(n15612), .A2(n15611), .ZN(n15613) );
  XNOR2_X1 U18889 ( .A(n15614), .B(n15613), .ZN(n16452) );
  XNOR2_X1 U18890 ( .A(n15789), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16449) );
  INV_X1 U18891 ( .A(n19016), .ZN(n15615) );
  OAI22_X1 U18892 ( .A1(n16428), .A2(n15616), .B1(n19291), .B2(n15615), .ZN(
        n15619) );
  OAI22_X1 U18893 ( .A1(n13674), .A2(n19020), .B1(n15617), .B2(n9725), .ZN(
        n15618) );
  AOI211_X1 U18894 ( .C1(n16449), .C2(n19288), .A(n15619), .B(n15618), .ZN(
        n15620) );
  OAI21_X1 U18895 ( .B1(n16452), .B2(n16421), .A(n15620), .ZN(P2_U2999) );
  AOI21_X1 U18896 ( .B1(n15914), .B2(n15622), .A(n15621), .ZN(n15916) );
  INV_X1 U18897 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15623) );
  AOI22_X1 U18898 ( .A1(n15916), .A2(n19285), .B1(n16417), .B2(n15623), .ZN(
        n15630) );
  AOI21_X1 U18899 ( .B1(n15914), .B2(n15625), .A(n15624), .ZN(n15911) );
  NAND2_X1 U18900 ( .A1(n19276), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n15912) );
  INV_X1 U18901 ( .A(n15912), .ZN(n15626) );
  AOI21_X1 U18902 ( .B1(n19288), .B2(n15911), .A(n15626), .ZN(n15629) );
  NAND2_X1 U18903 ( .A1(n15917), .A2(n19294), .ZN(n15628) );
  NAND2_X1 U18904 ( .A1(n19284), .A2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15627) );
  NAND4_X1 U18905 ( .A1(n15630), .A2(n15629), .A3(n15628), .A4(n15627), .ZN(
        P2_U3013) );
  NOR4_X1 U18906 ( .A1(n15644), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15642), .A4(n20856), .ZN(n15637) );
  OAI211_X1 U18907 ( .C1(n15631), .C2(n20856), .A(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n15695), .ZN(n15633) );
  AND2_X1 U18908 ( .A1(n15633), .A2(n15632), .ZN(n15634) );
  OAI211_X1 U18909 ( .C1(n16281), .C2(n16466), .A(n15635), .B(n15634), .ZN(
        n15636) );
  OAI21_X1 U18910 ( .B1(n15640), .B2(n16498), .A(n15639), .ZN(P2_U3015) );
  INV_X1 U18911 ( .A(n15641), .ZN(n15670) );
  NOR3_X1 U18912 ( .A1(n15670), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n15669), .ZN(n15661) );
  AOI21_X1 U18913 ( .B1(n15695), .B2(n15667), .A(n15661), .ZN(n15643) );
  NOR2_X1 U18914 ( .A1(n15643), .A2(n15642), .ZN(n15650) );
  NAND2_X1 U18915 ( .A1(n10152), .A2(n15648), .ZN(n15649) );
  OAI21_X1 U18916 ( .B1(n15653), .B2(n16498), .A(n15652), .ZN(P2_U3017) );
  INV_X1 U18917 ( .A(n15654), .ZN(n15655) );
  AOI21_X1 U18918 ( .B1(n16493), .B2(n15656), .A(n15655), .ZN(n15658) );
  NAND3_X1 U18919 ( .A1(n15667), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n15695), .ZN(n15657) );
  OAI211_X1 U18920 ( .C1(n15659), .C2(n16466), .A(n15658), .B(n15657), .ZN(
        n15660) );
  AOI211_X1 U18921 ( .C1(n15662), .C2(n16460), .A(n15661), .B(n15660), .ZN(
        n15663) );
  OAI21_X1 U18922 ( .B1(n15664), .B2(n16498), .A(n15663), .ZN(P2_U3018) );
  OAI21_X1 U18923 ( .B1(n16479), .B2(n15666), .A(n15665), .ZN(n15672) );
  INV_X1 U18924 ( .A(n15667), .ZN(n15668) );
  AOI21_X1 U18925 ( .B1(n15670), .B2(n15669), .A(n15668), .ZN(n15671) );
  AOI211_X1 U18926 ( .C1(n16494), .C2(n15673), .A(n15672), .B(n15671), .ZN(
        n15676) );
  NAND3_X1 U18927 ( .A1(n15674), .A2(n16460), .A3(n15506), .ZN(n15675) );
  OAI211_X1 U18928 ( .C1(n15677), .C2(n16498), .A(n15676), .B(n15675), .ZN(
        P2_U3019) );
  XNOR2_X1 U18929 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15685) );
  INV_X1 U18930 ( .A(n15678), .ZN(n15682) );
  NOR2_X1 U18931 ( .A1(n16479), .A2(n15679), .ZN(n15680) );
  AOI211_X1 U18932 ( .C1(n15682), .C2(n16494), .A(n15681), .B(n15680), .ZN(
        n15684) );
  NAND3_X1 U18933 ( .A1(n15709), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15695), .ZN(n15683) );
  OAI211_X1 U18934 ( .C1(n15698), .C2(n15685), .A(n15684), .B(n15683), .ZN(
        n15686) );
  AOI21_X1 U18935 ( .B1(n15687), .B2(n16460), .A(n15686), .ZN(n15688) );
  OAI21_X1 U18936 ( .B1(n15689), .B2(n16498), .A(n15688), .ZN(P2_U3020) );
  INV_X1 U18937 ( .A(n15690), .ZN(n15700) );
  OAI21_X1 U18938 ( .B1(n16479), .B2(n15692), .A(n15691), .ZN(n15693) );
  AOI21_X1 U18939 ( .B1(n15694), .B2(n16494), .A(n15693), .ZN(n15697) );
  NAND3_X1 U18940 ( .A1(n15709), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n15695), .ZN(n15696) );
  OAI211_X1 U18941 ( .C1(n15698), .C2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15697), .B(n15696), .ZN(n15699) );
  AOI21_X1 U18942 ( .B1(n15700), .B2(n16460), .A(n15699), .ZN(n15701) );
  OAI21_X1 U18943 ( .B1(n15702), .B2(n16498), .A(n15701), .ZN(P2_U3021) );
  XOR2_X1 U18944 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n10158), .Z(
        n15703) );
  XNOR2_X1 U18945 ( .A(n15704), .B(n15703), .ZN(n16318) );
  INV_X1 U18946 ( .A(n16318), .ZN(n15717) );
  NAND2_X1 U18947 ( .A1(n15706), .A2(n15705), .ZN(n15707) );
  AND2_X1 U18948 ( .A1(n15708), .A2(n15707), .ZN(n16316) );
  OAI21_X1 U18949 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15710), .A(
        n15709), .ZN(n15714) );
  AOI22_X1 U18950 ( .A1(n16493), .A2(n15711), .B1(P2_REIP_REG_24__SCAN_IN), 
        .B2(n19276), .ZN(n15713) );
  NAND2_X1 U18951 ( .A1(n16317), .A2(n16494), .ZN(n15712) );
  NAND3_X1 U18952 ( .A1(n15714), .A2(n15713), .A3(n15712), .ZN(n15715) );
  AOI21_X1 U18953 ( .B1(n16316), .B2(n16460), .A(n15715), .ZN(n15716) );
  OAI21_X1 U18954 ( .B1(n15717), .B2(n16498), .A(n15716), .ZN(P2_U3022) );
  NAND2_X1 U18955 ( .A1(n15718), .A2(n16485), .ZN(n15726) );
  INV_X1 U18956 ( .A(n15734), .ZN(n15749) );
  AOI22_X1 U18957 ( .A1(n16493), .A2(n15719), .B1(P2_REIP_REG_23__SCAN_IN), 
        .B2(n19276), .ZN(n15720) );
  OAI21_X1 U18958 ( .B1(n16282), .B2(n16466), .A(n15720), .ZN(n15724) );
  INV_X1 U18959 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15735) );
  AOI211_X1 U18960 ( .C1(n15722), .C2(n15735), .A(n15721), .B(n15736), .ZN(
        n15723) );
  AOI211_X1 U18961 ( .C1(n15749), .C2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15724), .B(n15723), .ZN(n15725) );
  OAI211_X1 U18962 ( .C1(n15727), .C2(n16503), .A(n15726), .B(n15725), .ZN(
        P2_U3023) );
  NAND2_X1 U18963 ( .A1(n15729), .A2(n15728), .ZN(n15731) );
  XOR2_X1 U18964 ( .A(n15731), .B(n15730), .Z(n16322) );
  AOI21_X1 U18965 ( .B1(n15735), .B2(n15556), .A(n15732), .ZN(n16323) );
  NAND2_X1 U18966 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19276), .ZN(n15733) );
  OAI221_X1 U18967 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15736), 
        .C1(n15735), .C2(n15734), .A(n15733), .ZN(n15739) );
  OAI22_X1 U18968 ( .A1(n16290), .A2(n16466), .B1(n16479), .B2(n15737), .ZN(
        n15738) );
  AOI211_X1 U18969 ( .C1(n16323), .C2(n16460), .A(n15739), .B(n15738), .ZN(
        n15740) );
  OAI21_X1 U18970 ( .B1(n16322), .B2(n16498), .A(n15740), .ZN(P2_U3024) );
  NAND2_X1 U18971 ( .A1(n15741), .A2(n16485), .ZN(n15751) );
  NAND2_X1 U18972 ( .A1(n16493), .A2(n15742), .ZN(n15743) );
  OAI211_X1 U18973 ( .C1(n15745), .C2(n16466), .A(n15744), .B(n15743), .ZN(
        n15748) );
  INV_X1 U18974 ( .A(n15767), .ZN(n15777) );
  NOR4_X1 U18975 ( .A1(n15907), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15746), .A4(n15777), .ZN(n15747) );
  AOI211_X1 U18976 ( .C1(n15749), .C2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15748), .B(n15747), .ZN(n15750) );
  OAI211_X1 U18977 ( .C1(n15752), .C2(n16503), .A(n15751), .B(n15750), .ZN(
        P2_U3025) );
  NAND2_X1 U18978 ( .A1(n15754), .A2(n15753), .ZN(n15758) );
  NAND2_X1 U18979 ( .A1(n15756), .A2(n15755), .ZN(n15757) );
  XOR2_X1 U18980 ( .A(n15758), .B(n15757), .Z(n16332) );
  INV_X1 U18981 ( .A(n16332), .ZN(n15775) );
  INV_X1 U18982 ( .A(n15590), .ZN(n16340) );
  AOI21_X1 U18983 ( .B1(n16340), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15759) );
  NOR2_X1 U18984 ( .A1(n15759), .A2(n15565), .ZN(n16331) );
  INV_X1 U18985 ( .A(n15887), .ZN(n16430) );
  AND2_X1 U18986 ( .A1(n15818), .A2(n15796), .ZN(n16447) );
  INV_X1 U18987 ( .A(n16447), .ZN(n15760) );
  NOR4_X1 U18988 ( .A1(n15760), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n21013), .A4(n15790), .ZN(n16434) );
  AOI211_X1 U18989 ( .C1(n16432), .C2(n16431), .A(n16430), .B(n16434), .ZN(
        n15776) );
  NOR2_X1 U18990 ( .A1(n15776), .A2(n15761), .ZN(n15773) );
  NOR2_X1 U18991 ( .A1(n9751), .A2(n15762), .ZN(n15763) );
  OR2_X1 U18992 ( .A1(n15764), .A2(n15763), .ZN(n18984) );
  AOI21_X1 U18993 ( .B1(n15766), .B2(n14021), .A(n15765), .ZN(n18986) );
  NOR2_X1 U18994 ( .A1(n9725), .A2(n18980), .ZN(n16330) );
  OAI211_X1 U18995 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n15767), .B(n15818), .ZN(
        n15768) );
  NOR2_X1 U18996 ( .A1(n15769), .A2(n15768), .ZN(n15770) );
  AOI211_X1 U18997 ( .C1(n16493), .C2(n18986), .A(n16330), .B(n15770), .ZN(
        n15771) );
  OAI21_X1 U18998 ( .B1(n18984), .B2(n16466), .A(n15771), .ZN(n15772) );
  AOI211_X1 U18999 ( .C1(n16331), .C2(n16460), .A(n15773), .B(n15772), .ZN(
        n15774) );
  OAI21_X1 U19000 ( .B1(n15775), .B2(n16498), .A(n15774), .ZN(P2_U3026) );
  INV_X1 U19001 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15781) );
  NOR2_X1 U19002 ( .A1(n15776), .A2(n15781), .ZN(n15784) );
  NOR2_X1 U19003 ( .A1(n15777), .A2(n15907), .ZN(n15780) );
  NOR2_X1 U19004 ( .A1(n12047), .A2(n9725), .ZN(n15779) );
  NOR2_X1 U19005 ( .A1(n18998), .A2(n16466), .ZN(n15778) );
  AOI211_X1 U19006 ( .C1(n15781), .C2(n15780), .A(n15779), .B(n15778), .ZN(
        n15782) );
  OAI21_X1 U19007 ( .B1(n16479), .B2(n18997), .A(n15782), .ZN(n15783) );
  AOI211_X1 U19008 ( .C1(n15785), .C2(n16460), .A(n15784), .B(n15783), .ZN(
        n15786) );
  OAI21_X1 U19009 ( .B1(n15787), .B2(n16498), .A(n15786), .ZN(P2_U3027) );
  OAI21_X1 U19010 ( .B1(n16466), .B2(n19009), .A(n15788), .ZN(n15792) );
  INV_X1 U19011 ( .A(n15789), .ZN(n15817) );
  AOI21_X1 U19012 ( .B1(n15817), .B2(n16460), .A(n16447), .ZN(n15806) );
  NOR3_X1 U19013 ( .A1(n15806), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15790), .ZN(n15791) );
  AOI211_X1 U19014 ( .C1(n16493), .C2(n19010), .A(n15792), .B(n15791), .ZN(
        n15804) );
  INV_X1 U19015 ( .A(n15793), .ZN(n15794) );
  NOR2_X1 U19016 ( .A1(n15794), .A2(n16460), .ZN(n15795) );
  OR2_X1 U19017 ( .A1(n16339), .A2(n15795), .ZN(n15801) );
  OR2_X1 U19018 ( .A1(n16491), .A2(n15796), .ZN(n15797) );
  NAND2_X1 U19019 ( .A1(n15887), .A2(n15797), .ZN(n16445) );
  NOR2_X1 U19020 ( .A1(n15798), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15799) );
  NOR2_X1 U19021 ( .A1(n16445), .A2(n15799), .ZN(n15800) );
  NAND2_X1 U19022 ( .A1(n15801), .A2(n15800), .ZN(n15809) );
  NOR2_X1 U19023 ( .A1(n16491), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15802) );
  OAI21_X1 U19024 ( .B1(n15809), .B2(n15802), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15803) );
  OAI211_X1 U19025 ( .C1(n15805), .C2(n16498), .A(n15804), .B(n15803), .ZN(
        P2_U3029) );
  OAI22_X1 U19026 ( .A1(n16466), .A2(n19142), .B1(n19856), .B2(n9725), .ZN(
        n15808) );
  NOR3_X1 U19027 ( .A1(n15806), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n16446), .ZN(n15807) );
  AOI211_X1 U19028 ( .C1(n16493), .C2(n19175), .A(n15808), .B(n15807), .ZN(
        n15811) );
  NAND2_X1 U19029 ( .A1(n15809), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15810) );
  OAI211_X1 U19030 ( .C1(n15812), .C2(n16498), .A(n15811), .B(n15810), .ZN(
        P2_U3030) );
  NAND2_X1 U19031 ( .A1(n15814), .A2(n15813), .ZN(n15815) );
  XNOR2_X1 U19032 ( .A(n15816), .B(n15815), .ZN(n16345) );
  INV_X1 U19033 ( .A(n16345), .ZN(n15837) );
  AOI21_X1 U19034 ( .B1(n15834), .B2(n15844), .A(n15817), .ZN(n16344) );
  INV_X1 U19035 ( .A(n15888), .ZN(n15819) );
  NAND2_X1 U19036 ( .A1(n15818), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16455) );
  NOR2_X1 U19037 ( .A1(n15819), .A2(n16455), .ZN(n15863) );
  NAND2_X1 U19038 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15822) );
  NOR2_X1 U19039 ( .A1(n15820), .A2(n15819), .ZN(n15821) );
  OAI21_X1 U19040 ( .B1(n15821), .B2(n16491), .A(n15887), .ZN(n15862) );
  AOI21_X1 U19041 ( .B1(n15863), .B2(n15822), .A(n15862), .ZN(n15858) );
  INV_X1 U19042 ( .A(n15823), .ZN(n15825) );
  AOI21_X1 U19043 ( .B1(n15825), .B2(n15852), .A(n9793), .ZN(n19183) );
  OR2_X1 U19044 ( .A1(n15827), .A2(n15826), .ZN(n15828) );
  NAND2_X1 U19045 ( .A1(n15829), .A2(n15828), .ZN(n19146) );
  OAI22_X1 U19046 ( .A1(n16466), .A2(n19146), .B1(n12030), .B2(n9725), .ZN(
        n15832) );
  NOR3_X1 U19047 ( .A1(n16455), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n15830), .ZN(n15831) );
  AOI211_X1 U19048 ( .C1(n16493), .C2(n19183), .A(n15832), .B(n15831), .ZN(
        n15833) );
  OAI21_X1 U19049 ( .B1(n15858), .B2(n15834), .A(n15833), .ZN(n15835) );
  AOI21_X1 U19050 ( .B1(n16344), .B2(n16460), .A(n15835), .ZN(n15836) );
  OAI21_X1 U19051 ( .B1(n15837), .B2(n16498), .A(n15836), .ZN(P2_U3032) );
  INV_X1 U19052 ( .A(n15838), .ZN(n15840) );
  NOR2_X1 U19053 ( .A1(n15840), .A2(n15839), .ZN(n15843) );
  XOR2_X1 U19054 ( .A(n15843), .B(n15842), .Z(n16349) );
  INV_X1 U19055 ( .A(n15844), .ZN(n15845) );
  AOI21_X1 U19056 ( .B1(n15846), .B2(n16356), .A(n15845), .ZN(n16348) );
  AOI21_X1 U19057 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15863), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15857) );
  INV_X1 U19058 ( .A(n19045), .ZN(n15848) );
  OAI22_X1 U19059 ( .A1(n16466), .A2(n15848), .B1(n9725), .B2(n15847), .ZN(
        n15849) );
  INV_X1 U19060 ( .A(n15849), .ZN(n15856) );
  OR2_X1 U19061 ( .A1(n15851), .A2(n15850), .ZN(n15853) );
  NAND2_X1 U19062 ( .A1(n15853), .A2(n15852), .ZN(n19188) );
  INV_X1 U19063 ( .A(n19188), .ZN(n15854) );
  NAND2_X1 U19064 ( .A1(n16493), .A2(n15854), .ZN(n15855) );
  OAI211_X1 U19065 ( .C1(n15858), .C2(n15857), .A(n15856), .B(n15855), .ZN(
        n15859) );
  AOI21_X1 U19066 ( .B1(n16348), .B2(n16460), .A(n15859), .ZN(n15860) );
  OAI21_X1 U19067 ( .B1(n16498), .B2(n16349), .A(n15860), .ZN(P2_U3033) );
  NAND3_X1 U19068 ( .A1(n16355), .A2(n16356), .A3(n16460), .ZN(n15879) );
  NOR2_X1 U19069 ( .A1(n12024), .A2(n9725), .ZN(n15861) );
  AOI221_X1 U19070 ( .B1(n15863), .B2(n11794), .C1(n15862), .C2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n15861), .ZN(n15878) );
  OR2_X1 U19071 ( .A1(n15865), .A2(n15864), .ZN(n15867) );
  NAND2_X1 U19072 ( .A1(n15867), .A2(n15866), .ZN(n19149) );
  INV_X1 U19073 ( .A(n19149), .ZN(n19053) );
  XNOR2_X1 U19074 ( .A(n15319), .B(n15868), .ZN(n19191) );
  INV_X1 U19075 ( .A(n19191), .ZN(n15869) );
  AOI22_X1 U19076 ( .A1(n16494), .A2(n19053), .B1(n16493), .B2(n15869), .ZN(
        n15877) );
  INV_X1 U19077 ( .A(n15871), .ZN(n15872) );
  OR2_X1 U19078 ( .A1(n15873), .A2(n15872), .ZN(n15874) );
  XNOR2_X1 U19079 ( .A(n15875), .B(n15874), .ZN(n16357) );
  NAND2_X1 U19080 ( .A1(n16357), .A2(n16485), .ZN(n15876) );
  NAND4_X1 U19081 ( .A1(n15879), .A2(n15878), .A3(n15877), .A4(n15876), .ZN(
        P2_U3034) );
  NAND3_X1 U19082 ( .A1(n15880), .A2(n15897), .A3(n16373), .ZN(n15885) );
  INV_X1 U19083 ( .A(n15881), .ZN(n15882) );
  NOR2_X1 U19084 ( .A1(n15883), .A2(n15882), .ZN(n15884) );
  XNOR2_X1 U19085 ( .A(n15885), .B(n15884), .ZN(n16364) );
  OAI21_X1 U19086 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n9977), .A(
        n15886), .ZN(n16365) );
  OAI21_X1 U19087 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16491), .A(
        n15887), .ZN(n16458) );
  NOR2_X1 U19088 ( .A1(n12021), .A2(n9725), .ZN(n15891) );
  AOI211_X1 U19089 ( .C1(n16380), .C2(n15889), .A(n15888), .B(n16455), .ZN(
        n15890) );
  AOI211_X1 U19090 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16458), .A(
        n15891), .B(n15890), .ZN(n15894) );
  INV_X1 U19091 ( .A(n19193), .ZN(n15892) );
  AOI22_X1 U19092 ( .A1(n16494), .A2(n16367), .B1(n16493), .B2(n15892), .ZN(
        n15893) );
  OAI211_X1 U19093 ( .C1(n16365), .C2(n16503), .A(n15894), .B(n15893), .ZN(
        n15895) );
  INV_X1 U19094 ( .A(n15895), .ZN(n15896) );
  OAI21_X1 U19095 ( .B1(n16364), .B2(n16498), .A(n15896), .ZN(P2_U3035) );
  INV_X1 U19096 ( .A(n15897), .ZN(n16371) );
  OR2_X1 U19097 ( .A1(n16371), .A2(n15898), .ZN(n15899) );
  XNOR2_X1 U19098 ( .A(n15900), .B(n15899), .ZN(n16387) );
  NOR2_X1 U19099 ( .A1(n12010), .A2(n9725), .ZN(n15905) );
  OR2_X1 U19100 ( .A1(n15901), .A2(n15335), .ZN(n15903) );
  NAND2_X1 U19101 ( .A1(n15903), .A2(n16454), .ZN(n19199) );
  NOR2_X1 U19102 ( .A1(n16479), .A2(n19199), .ZN(n15904) );
  AOI211_X1 U19103 ( .C1(n16494), .C2(n19073), .A(n15905), .B(n15904), .ZN(
        n15906) );
  OAI21_X1 U19104 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15907), .A(
        n15906), .ZN(n15909) );
  NOR2_X1 U19105 ( .A1(n16388), .A2(n16503), .ZN(n15908) );
  AOI211_X1 U19106 ( .C1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n16430), .A(
        n15909), .B(n15908), .ZN(n15910) );
  OAI21_X1 U19107 ( .B1(n16498), .B2(n16387), .A(n15910), .ZN(P2_U3037) );
  AOI22_X1 U19108 ( .A1(n16460), .A2(n15911), .B1(n16493), .B2(n19920), .ZN(
        n15913) );
  OAI211_X1 U19109 ( .C1(n16490), .C2(n15914), .A(n15913), .B(n15912), .ZN(
        n15915) );
  INV_X1 U19110 ( .A(n15915), .ZN(n15922) );
  AOI22_X1 U19111 ( .A1(n15917), .A2(n16494), .B1(n16485), .B2(n15916), .ZN(
        n15921) );
  INV_X1 U19112 ( .A(n15918), .ZN(n15919) );
  OAI211_X1 U19113 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n16431), .B(n15919), .ZN(n15920) );
  NAND3_X1 U19114 ( .A1(n15922), .A2(n15921), .A3(n15920), .ZN(P2_U3045) );
  INV_X1 U19115 ( .A(n15935), .ZN(n16508) );
  AOI22_X1 U19116 ( .A1(n19098), .A2(n15923), .B1(n19138), .B2(n9740), .ZN(
        n15934) );
  OAI222_X1 U19117 ( .A1(n16508), .A2(n12829), .B1(n19889), .B2(n15924), .C1(
        n12874), .C2(n15934), .ZN(n15931) );
  AOI22_X1 U19118 ( .A1(n15926), .A2(n15925), .B1(P2_FLUSH_REG_SCAN_IN), .B2(
        n16506), .ZN(n15927) );
  OAI21_X1 U19119 ( .B1(n19757), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n15927), 
        .ZN(n15981) );
  INV_X1 U19120 ( .A(n15928), .ZN(n15929) );
  OAI21_X1 U19121 ( .B1(n15929), .B2(n19889), .A(n15981), .ZN(n15930) );
  AOI22_X1 U19122 ( .A1(n15931), .A2(n15981), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15930), .ZN(n15932) );
  INV_X1 U19123 ( .A(n15932), .ZN(P2_U3601) );
  AOI21_X1 U19124 ( .B1(n19098), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n15933), .ZN(n15944) );
  NAND2_X1 U19125 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15934), .ZN(n15945) );
  INV_X1 U19126 ( .A(n15945), .ZN(n15936) );
  AOI222_X1 U19127 ( .A1(n15938), .A2(n15937), .B1(n15944), .B2(n15936), .C1(
        n19917), .C2(n15935), .ZN(n15941) );
  INV_X1 U19128 ( .A(n15981), .ZN(n15940) );
  NAND2_X1 U19129 ( .A1(n15940), .A2(n21077), .ZN(n15939) );
  OAI21_X1 U19130 ( .B1(n15941), .B2(n15940), .A(n15939), .ZN(P2_U3600) );
  INV_X1 U19131 ( .A(n15942), .ZN(n15943) );
  OAI222_X1 U19132 ( .A1(n19210), .A2(n16508), .B1(n15945), .B2(n15944), .C1(
        n19889), .C2(n15943), .ZN(n15946) );
  MUX2_X1 U19133 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n15946), .S(
        n15981), .Z(P2_U3599) );
  OAI22_X1 U19134 ( .A1(n19567), .A2(n16508), .B1(n15947), .B2(n19889), .ZN(
        n15948) );
  MUX2_X1 U19135 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15948), .S(
        n15981), .Z(P2_U3596) );
  AOI22_X1 U19136 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15949), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15956) );
  AOI22_X1 U19137 ( .A1(n15950), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15955) );
  AOI22_X1 U19138 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15951), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15954) );
  AOI22_X1 U19139 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15952), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15953) );
  NAND4_X1 U19140 ( .A1(n15956), .A2(n15955), .A3(n15954), .A4(n15953), .ZN(
        n15962) );
  AOI22_X1 U19141 ( .A1(n17256), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15960) );
  AOI22_X1 U19142 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15959) );
  AOI22_X1 U19143 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15958) );
  AOI22_X1 U19144 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15957) );
  NAND4_X1 U19145 ( .A1(n15960), .A2(n15959), .A3(n15958), .A4(n15957), .ZN(
        n15961) );
  NOR2_X1 U19146 ( .A1(n15962), .A2(n15961), .ZN(n17435) );
  INV_X1 U19147 ( .A(n17238), .ZN(n15963) );
  NOR2_X1 U19148 ( .A1(n17338), .A2(n17212), .ZN(n17224) );
  OAI21_X1 U19149 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n15963), .A(n17224), .ZN(
        n15964) );
  OAI21_X1 U19150 ( .B1(n17435), .B2(n17332), .A(n15964), .ZN(P3_U2690) );
  NOR2_X1 U19151 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18887), .ZN(n18301) );
  NAND2_X1 U19152 ( .A1(n18772), .A2(n18927), .ZN(n15970) );
  NAND2_X1 U19153 ( .A1(n18931), .A2(n15966), .ZN(n17492) );
  AOI21_X1 U19154 ( .B1(n15969), .B2(n15968), .A(n15967), .ZN(n15994) );
  OAI21_X1 U19155 ( .B1(n15970), .B2(n17492), .A(n15994), .ZN(n15971) );
  NOR3_X1 U19156 ( .A1(n16079), .A2(n15972), .A3(n15971), .ZN(n18757) );
  INV_X1 U19157 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18287) );
  OAI22_X1 U19158 ( .A1(n18757), .A2(n18792), .B1(n18287), .B2(n18885), .ZN(
        n15973) );
  INV_X1 U19159 ( .A(n18736), .ZN(n18738) );
  AOI21_X1 U19160 ( .B1(n18738), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15975) );
  NOR3_X1 U19161 ( .A1(n15975), .A2(n18733), .A3(n15974), .ZN(n18775) );
  NAND3_X1 U19162 ( .A1(n18912), .A2(n18946), .A3(n18775), .ZN(n15976) );
  OAI21_X1 U19163 ( .B1(n18912), .B2(n18780), .A(n15976), .ZN(P3_U3284) );
  INV_X1 U19164 ( .A(n15977), .ZN(n15978) );
  NOR4_X1 U19165 ( .A1(n11913), .A2(n15978), .A3(n19944), .A4(n19889), .ZN(
        n15979) );
  NAND2_X1 U19166 ( .A1(n15981), .A2(n15979), .ZN(n15980) );
  OAI21_X1 U19167 ( .B1(n15981), .B2(n20966), .A(n15980), .ZN(P2_U3595) );
  INV_X1 U19168 ( .A(n15982), .ZN(n15992) );
  OAI21_X1 U19169 ( .B1(n18309), .B2(n17554), .A(n15983), .ZN(n15984) );
  OAI21_X1 U19170 ( .B1(n15985), .B2(n15984), .A(n18927), .ZN(n16667) );
  NOR3_X1 U19171 ( .A1(n15987), .A2(n15986), .A3(n16667), .ZN(n15991) );
  AOI21_X1 U19172 ( .B1(n18318), .B2(n15989), .A(n15988), .ZN(n15990) );
  AOI211_X1 U19173 ( .C1(n15992), .C2(n18773), .A(n15991), .B(n15990), .ZN(
        n15993) );
  NAND2_X1 U19174 ( .A1(n18766), .A2(n16006), .ZN(n18106) );
  NOR2_X2 U19175 ( .A1(n18281), .A2(n18106), .ZN(n18181) );
  INV_X1 U19176 ( .A(n18181), .ZN(n18194) );
  OAI21_X1 U19177 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n9788), .A(
        n15995), .ZN(n16546) );
  INV_X1 U19178 ( .A(n18229), .ZN(n16063) );
  INV_X1 U19179 ( .A(n16518), .ZN(n18030) );
  NAND3_X1 U19180 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18077) );
  NOR3_X1 U19181 ( .A1(n18222), .A2(n18217), .A3(n18245), .ZN(n18076) );
  NAND3_X1 U19182 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n18076), .ZN(n18185) );
  NOR2_X1 U19183 ( .A1(n18077), .A2(n18185), .ZN(n18157) );
  NAND2_X1 U19184 ( .A1(n15997), .A2(n18157), .ZN(n18070) );
  NOR2_X1 U19185 ( .A1(n18030), .A2(n18070), .ZN(n16000) );
  NAND2_X1 U19186 ( .A1(n9745), .A2(n18911), .ZN(n18187) );
  NAND2_X1 U19187 ( .A1(n16000), .A2(n18187), .ZN(n18026) );
  NOR2_X1 U19188 ( .A1(n18012), .A2(n18018), .ZN(n17973) );
  NAND2_X1 U19189 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17973), .ZN(
        n17975) );
  NOR2_X1 U19190 ( .A1(n15999), .A2(n17975), .ZN(n16519) );
  NAND2_X1 U19191 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n16519), .ZN(
        n17611) );
  OAI21_X1 U19192 ( .B1(n18026), .B2(n17611), .A(n9745), .ZN(n16004) );
  OAI21_X1 U19193 ( .B1(n18911), .B2(n10060), .A(n18254), .ZN(n18250) );
  NAND2_X1 U19194 ( .A1(n18076), .A2(n18250), .ZN(n18186) );
  NOR2_X1 U19195 ( .A1(n18186), .A2(n18077), .ZN(n18152) );
  INV_X1 U19196 ( .A(n18152), .ZN(n15998) );
  INV_X1 U19197 ( .A(n18071), .ZN(n15996) );
  NAND2_X1 U19198 ( .A1(n15997), .A2(n15996), .ZN(n16569) );
  NOR2_X1 U19199 ( .A1(n15998), .A2(n16569), .ZN(n18027) );
  INV_X1 U19200 ( .A(n18027), .ZN(n18072) );
  NOR3_X1 U19201 ( .A1(n20842), .A2(n18030), .A3(n18072), .ZN(n18011) );
  NAND2_X1 U19202 ( .A1(n17973), .A2(n18011), .ZN(n17977) );
  OAI21_X1 U19203 ( .B1(n15999), .B2(n17977), .A(n18768), .ZN(n16003) );
  INV_X1 U19204 ( .A(n18282), .ZN(n18749) );
  AOI21_X1 U19205 ( .B1(n16000), .B2(n16519), .A(n18749), .ZN(n16001) );
  INV_X1 U19206 ( .A(n16001), .ZN(n16002) );
  AND4_X1 U19207 ( .A1(n18265), .A2(n16004), .A3(n16003), .A4(n16002), .ZN(
        n16064) );
  OAI21_X1 U19208 ( .B1(n18162), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16064), .ZN(n16564) );
  AOI21_X1 U19209 ( .B1(n16063), .B2(n17613), .A(n16564), .ZN(n16009) );
  NAND2_X1 U19210 ( .A1(n18767), .A2(n18265), .ZN(n18257) );
  AOI21_X1 U19211 ( .B1(n17978), .B2(n16527), .A(n18257), .ZN(n16008) );
  INV_X1 U19212 ( .A(n16005), .ZN(n16528) );
  NAND2_X1 U19213 ( .A1(n18766), .A2(n18265), .ZN(n18274) );
  NOR3_X1 U19214 ( .A1(n16528), .A2(n16006), .A3(n18274), .ZN(n16007) );
  NOR2_X1 U19215 ( .A1(n16008), .A2(n16007), .ZN(n16067) );
  OAI21_X1 U19216 ( .B1(n18125), .B2(n16009), .A(n16067), .ZN(n16017) );
  INV_X1 U19217 ( .A(n18257), .ZN(n18277) );
  NAND2_X1 U19218 ( .A1(n18766), .A2(n17458), .ZN(n18153) );
  NOR2_X1 U19219 ( .A1(n16011), .A2(n16010), .ZN(n18734) );
  OAI21_X1 U19220 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18282), .A(
        n18735), .ZN(n18246) );
  NOR2_X1 U19221 ( .A1(n16569), .A2(n18246), .ZN(n16012) );
  AOI22_X1 U19222 ( .A1(n18768), .A2(n18027), .B1(n18157), .B2(n16012), .ZN(
        n16568) );
  NOR3_X1 U19223 ( .A1(n16568), .A2(n16013), .A3(n17975), .ZN(n17996) );
  NAND2_X1 U19224 ( .A1(n17974), .A2(n17996), .ZN(n16551) );
  OAI21_X1 U19225 ( .B1(n18153), .B2(n17981), .A(n16551), .ZN(n16014) );
  AOI22_X1 U19226 ( .A1(n17978), .A2(n18277), .B1(n18265), .B2(n16014), .ZN(
        n16070) );
  NOR2_X1 U19227 ( .A1(n16070), .A2(n16533), .ZN(n16016) );
  AOI22_X1 U19228 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16017), .B1(
        n16016), .B2(n16015), .ZN(n16018) );
  NAND2_X1 U19229 ( .A1(n18198), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16542) );
  OAI211_X1 U19230 ( .C1(n18194), .C2(n16546), .A(n16018), .B(n16542), .ZN(
        P3_U2833) );
  AOI21_X1 U19231 ( .B1(n16019), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n20573), .ZN(n16020) );
  AND2_X1 U19232 ( .A1(n16021), .A2(n16020), .ZN(n16024) );
  OAI22_X1 U19233 ( .A1(n16023), .A2(n16022), .B1(n16024), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n16027) );
  INV_X1 U19234 ( .A(n16024), .ZN(n16025) );
  OR2_X1 U19235 ( .A1(n16025), .A2(n20541), .ZN(n16026) );
  AND2_X1 U19236 ( .A1(n16027), .A2(n16026), .ZN(n16029) );
  INV_X1 U19237 ( .A(n16029), .ZN(n16031) );
  OAI21_X1 U19238 ( .B1(n16029), .B2(n20459), .A(n16028), .ZN(n16030) );
  OAI21_X1 U19239 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16031), .A(
        n16030), .ZN(n16032) );
  AOI222_X1 U19240 ( .A1(n21022), .A2(n16033), .B1(n21022), .B2(n16032), .C1(
        n16033), .C2(n16032), .ZN(n16036) );
  OAI211_X1 U19241 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n16036), .A(
        n16035), .B(n16034), .ZN(n16043) );
  INV_X1 U19242 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19971) );
  NAND2_X1 U19243 ( .A1(n20868), .A2(n19971), .ZN(n16038) );
  AOI21_X1 U19244 ( .B1(n16039), .B2(n16038), .A(n16037), .ZN(n16040) );
  NAND2_X1 U19245 ( .A1(n16041), .A2(n16040), .ZN(n16042) );
  NAND2_X1 U19246 ( .A1(n16044), .A2(n20812), .ZN(n16047) );
  OAI21_X1 U19247 ( .B1(n16045), .B2(n20819), .A(n16052), .ZN(n16046) );
  OAI21_X1 U19248 ( .B1(n16048), .B2(n16047), .A(n16046), .ZN(n16262) );
  AOI221_X1 U19249 ( .B1(n20815), .B2(n20714), .C1(n16049), .C2(n20714), .A(
        n16262), .ZN(n16266) );
  INV_X1 U19250 ( .A(n16049), .ZN(n16053) );
  AOI21_X1 U19251 ( .B1(n20724), .B2(n20811), .A(n16056), .ZN(n16051) );
  OAI211_X1 U19252 ( .C1(n16053), .C2(n16052), .A(n16051), .B(n16050), .ZN(
        n16054) );
  NOR2_X1 U19253 ( .A1(n16266), .A2(n16054), .ZN(n16059) );
  NAND2_X1 U19254 ( .A1(n16056), .A2(n16055), .ZN(n16057) );
  NAND2_X1 U19255 ( .A1(n20815), .A2(n16057), .ZN(n16058) );
  OAI22_X1 U19256 ( .A1(n16059), .A2(n20815), .B1(n16266), .B2(n16058), .ZN(
        P1_U3161) );
  NAND2_X1 U19257 ( .A1(n16527), .A2(n16066), .ZN(n16531) );
  NOR2_X1 U19258 ( .A1(n16061), .A2(n16060), .ZN(n16062) );
  XNOR2_X1 U19259 ( .A(n16062), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16526) );
  NAND2_X1 U19260 ( .A1(n18265), .A2(n16063), .ZN(n18267) );
  OAI22_X1 U19261 ( .A1(n18267), .A2(n16527), .B1(n18198), .B2(n16064), .ZN(
        n16065) );
  INV_X1 U19262 ( .A(n16065), .ZN(n16547) );
  AOI21_X1 U19263 ( .B1(n16547), .B2(n16067), .A(n16066), .ZN(n16068) );
  AOI21_X1 U19264 ( .B1(n18181), .B2(n16526), .A(n16068), .ZN(n16069) );
  NAND2_X1 U19265 ( .A1(n18198), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16521) );
  OAI211_X1 U19266 ( .C1(n16070), .C2(n16531), .A(n16069), .B(n16521), .ZN(
        P3_U2832) );
  INV_X1 U19267 ( .A(HOLD), .ZN(n20719) );
  INV_X1 U19268 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20733) );
  NAND2_X1 U19269 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20733), .ZN(n20723) );
  INV_X1 U19270 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20725) );
  NOR2_X1 U19271 ( .A1(n12916), .A2(n20725), .ZN(n20726) );
  NAND2_X1 U19272 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n16071) );
  AOI22_X1 U19273 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20724), .B1(n20726), 
        .B2(n16071), .ZN(n16073) );
  OAI211_X1 U19274 ( .C1(n20719), .C2(n20723), .A(n16073), .B(n16072), .ZN(
        P1_U3195) );
  AND2_X1 U19275 ( .A1(n16074), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR3_X1 U19276 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n16510), .A3(n16075), 
        .ZN(n16505) );
  AOI221_X1 U19277 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .C1(P2_STATE2_REG_0__SCAN_IN), .C2(
        P2_STATE2_REG_1__SCAN_IN), .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n16076)
         );
  NOR3_X1 U19278 ( .A1(n16505), .A2(n16506), .A3(n16076), .ZN(P2_U3178) );
  INV_X1 U19279 ( .A(n16507), .ZN(n19936) );
  AOI221_X1 U19280 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16506), .C1(n19936), .C2(
        n16506), .A(n19765), .ZN(n19932) );
  AND2_X1 U19281 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n19932), .ZN(
        P2_U3047) );
  INV_X1 U19282 ( .A(n16080), .ZN(n18748) );
  NAND2_X1 U19283 ( .A1(n17478), .A2(n16080), .ZN(n17475) );
  AOI22_X1 U19284 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17485), .B1(
        P3_EAX_REG_0__SCAN_IN), .B2(n17486), .ZN(n16082) );
  NAND2_X1 U19285 ( .A1(n18332), .A2(n9929), .ZN(n17427) );
  NOR2_X1 U19286 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17427), .ZN(n17487) );
  INV_X1 U19287 ( .A(n17487), .ZN(n16081) );
  OAI211_X1 U19288 ( .C1(n17967), .C2(n17490), .A(n16082), .B(n16081), .ZN(
        P3_U2735) );
  AOI22_X1 U19289 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n20042), .B1(
        P1_EBX_REG_17__SCAN_IN), .B2(n20041), .ZN(n16088) );
  AOI21_X1 U19290 ( .B1(n20039), .B2(n16136), .A(n19987), .ZN(n16087) );
  AOI22_X1 U19291 ( .A1(n16137), .A2(n20018), .B1(n20024), .B2(n16172), .ZN(
        n16086) );
  OAI21_X1 U19292 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n16084), .A(n16083), 
        .ZN(n16085) );
  NAND4_X1 U19293 ( .A1(n16088), .A2(n16087), .A3(n16086), .A4(n16085), .ZN(
        P1_U2823) );
  AOI22_X1 U19294 ( .A1(n16089), .A2(n20039), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n20041), .ZN(n16090) );
  OAI211_X1 U19295 ( .C1(n19999), .C2(n16091), .A(n16090), .B(n20043), .ZN(
        n16092) );
  AOI21_X1 U19296 ( .B1(n20024), .B2(n16093), .A(n16092), .ZN(n16098) );
  OAI21_X1 U19297 ( .B1(n16095), .B2(n16094), .A(n19995), .ZN(n16103) );
  AOI22_X1 U19298 ( .A1(n16096), .A2(n20018), .B1(P1_REIP_REG_13__SCAN_IN), 
        .B2(n16103), .ZN(n16097) );
  OAI211_X1 U19299 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n16099), .A(n16098), 
        .B(n16097), .ZN(P1_U2827) );
  AOI22_X1 U19300 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20042), .B1(
        P1_EBX_REG_12__SCAN_IN), .B2(n20041), .ZN(n16108) );
  XNOR2_X1 U19301 ( .A(n16101), .B(n16100), .ZN(n16213) );
  AOI21_X1 U19302 ( .B1(n20024), .B2(n16213), .A(n19987), .ZN(n16107) );
  INV_X1 U19303 ( .A(n16102), .ZN(n16144) );
  AOI22_X1 U19304 ( .A1(n16145), .A2(n20018), .B1(n16144), .B2(n20039), .ZN(
        n16106) );
  OAI21_X1 U19305 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(n16104), .A(n16103), 
        .ZN(n16105) );
  NAND4_X1 U19306 ( .A1(n16108), .A2(n16107), .A3(n16106), .A4(n16105), .ZN(
        P1_U2828) );
  AOI21_X1 U19307 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n19995), .A(
        P1_REIP_REG_10__SCAN_IN), .ZN(n16113) );
  OAI22_X1 U19308 ( .A1(n16109), .A2(n20000), .B1(n20053), .B2(n16235), .ZN(
        n16110) );
  AOI211_X1 U19309 ( .C1(n20042), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n19987), .B(n16110), .ZN(n16112) );
  AOI22_X1 U19310 ( .A1(n16153), .A2(n20018), .B1(n20039), .B2(n16150), .ZN(
        n16111) );
  OAI211_X1 U19311 ( .C1(n16114), .C2(n16113), .A(n16112), .B(n16111), .ZN(
        P1_U2830) );
  INV_X1 U19312 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n20833) );
  AOI22_X1 U19313 ( .A1(n16145), .A2(n16116), .B1(n16115), .B2(n16213), .ZN(
        n16117) );
  OAI21_X1 U19314 ( .B1(n16118), .B2(n20833), .A(n16117), .ZN(P1_U2860) );
  AOI22_X1 U19315 ( .A1(n16135), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n16171), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16125) );
  NAND2_X1 U19316 ( .A1(n16120), .A2(n16119), .ZN(n16122) );
  XOR2_X1 U19317 ( .A(n16122), .B(n16121), .Z(n16167) );
  AOI22_X1 U19318 ( .A1(n16123), .A2(n16152), .B1(n11125), .B2(n16167), .ZN(
        n16124) );
  OAI211_X1 U19319 ( .C1(n16127), .C2(n16126), .A(n16125), .B(n16124), .ZN(
        P1_U2980) );
  INV_X1 U19320 ( .A(n16128), .ZN(n16129) );
  AOI21_X1 U19321 ( .B1(n16131), .B2(n16130), .A(n16129), .ZN(n16133) );
  NOR2_X1 U19322 ( .A1(n16133), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16132) );
  MUX2_X1 U19323 ( .A(n16133), .B(n16132), .S(n14734), .Z(n16134) );
  XNOR2_X1 U19324 ( .A(n16134), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16176) );
  AOI22_X1 U19325 ( .A1(n16135), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n16171), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16139) );
  AOI22_X1 U19326 ( .A1(n16137), .A2(n16152), .B1(n16136), .B2(n16151), .ZN(
        n16138) );
  OAI211_X1 U19327 ( .C1(n19970), .C2(n16176), .A(n16139), .B(n16138), .ZN(
        P1_U2982) );
  OAI21_X1 U19328 ( .B1(n16142), .B2(n16141), .A(n16140), .ZN(n16143) );
  INV_X1 U19329 ( .A(n16143), .ZN(n16218) );
  AOI22_X1 U19330 ( .A1(n16135), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n16171), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16147) );
  AOI22_X1 U19331 ( .A1(n16145), .A2(n16152), .B1(n16144), .B2(n16151), .ZN(
        n16146) );
  OAI211_X1 U19332 ( .C1(n16218), .C2(n19970), .A(n16147), .B(n16146), .ZN(
        P1_U2987) );
  MUX2_X1 U19333 ( .A(n16148), .B(n14873), .S(n14734), .Z(n16149) );
  XNOR2_X1 U19334 ( .A(n16149), .B(n16234), .ZN(n16239) );
  AOI22_X1 U19335 ( .A1(n16135), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n16171), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n16155) );
  AOI22_X1 U19336 ( .A1(n16153), .A2(n16152), .B1(n16151), .B2(n16150), .ZN(
        n16154) );
  OAI211_X1 U19337 ( .C1(n19970), .C2(n16239), .A(n16155), .B(n16154), .ZN(
        P1_U2989) );
  INV_X1 U19338 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16157) );
  OAI22_X1 U19339 ( .A1(n16158), .A2(n20107), .B1(n16157), .B2(n16156), .ZN(
        n16159) );
  AOI21_X1 U19340 ( .B1(n20117), .B2(n16160), .A(n16159), .ZN(n16164) );
  OAI211_X1 U19341 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16162), .B(n16161), .ZN(
        n16163) );
  OAI211_X1 U19342 ( .C1(n20770), .C2(n16200), .A(n16164), .B(n16163), .ZN(
        P1_U3009) );
  AOI22_X1 U19343 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16165), .B1(
        n16171), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16169) );
  AOI22_X1 U19344 ( .A1(n16167), .A2(n20117), .B1(n20116), .B2(n16166), .ZN(
        n16168) );
  OAI211_X1 U19345 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n16170), .A(
        n16169), .B(n16168), .ZN(P1_U3012) );
  AOI22_X1 U19346 ( .A1(n16172), .A2(n20116), .B1(n16171), .B2(
        P1_REIP_REG_17__SCAN_IN), .ZN(n16175) );
  NOR2_X1 U19347 ( .A1(n16199), .A2(n16198), .ZN(n16184) );
  OAI221_X1 U19348 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n16183), 
        .C1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n16184), .A(n16173), .ZN(
        n16174) );
  OAI211_X1 U19349 ( .C1(n16176), .C2(n20091), .A(n16175), .B(n16174), .ZN(
        P1_U3014) );
  OAI21_X1 U19350 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n16184), .ZN(n16182) );
  AOI21_X1 U19351 ( .B1(n16178), .B2(n20116), .A(n16177), .ZN(n16181) );
  OAI21_X1 U19352 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16199), .A(
        n16197), .ZN(n16188) );
  AOI22_X1 U19353 ( .A1(n16179), .A2(n20117), .B1(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n16188), .ZN(n16180) );
  OAI211_X1 U19354 ( .C1(n16183), .C2(n16182), .A(n16181), .B(n16180), .ZN(
        P1_U3015) );
  INV_X1 U19355 ( .A(n16184), .ZN(n16192) );
  AOI21_X1 U19356 ( .B1(n16186), .B2(n20116), .A(n16185), .ZN(n16191) );
  INV_X1 U19357 ( .A(n16187), .ZN(n16189) );
  AOI22_X1 U19358 ( .A1(n16189), .A2(n20117), .B1(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16188), .ZN(n16190) );
  OAI211_X1 U19359 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16192), .A(
        n16191), .B(n16190), .ZN(P1_U3016) );
  OAI22_X1 U19360 ( .A1(n16193), .A2(n20107), .B1(n20756), .B2(n16200), .ZN(
        n16194) );
  AOI21_X1 U19361 ( .B1(n20117), .B2(n16195), .A(n16194), .ZN(n16196) );
  OAI221_X1 U19362 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16199), 
        .C1(n16198), .C2(n16197), .A(n16196), .ZN(P1_U3017) );
  NOR2_X1 U19363 ( .A1(n16200), .A2(n20753), .ZN(n16212) );
  INV_X1 U19364 ( .A(n16208), .ZN(n16202) );
  AOI21_X1 U19365 ( .B1(n16203), .B2(n16202), .A(n16201), .ZN(n16205) );
  AOI211_X1 U19366 ( .C1(n16207), .C2(n16206), .A(n16205), .B(n16204), .ZN(
        n16226) );
  NOR2_X1 U19367 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16208), .ZN(
        n16221) );
  NAND2_X1 U19368 ( .A1(n16221), .A2(n16209), .ZN(n16210) );
  AOI21_X1 U19369 ( .B1(n16226), .B2(n16210), .A(n16214), .ZN(n16211) );
  AOI211_X1 U19370 ( .C1(n20116), .C2(n16213), .A(n16212), .B(n16211), .ZN(
        n16217) );
  NAND3_X1 U19371 ( .A1(n16215), .A2(n16231), .A3(n16214), .ZN(n16216) );
  OAI211_X1 U19372 ( .C1(n16218), .C2(n20091), .A(n16217), .B(n16216), .ZN(
        P1_U3019) );
  AOI21_X1 U19373 ( .B1(n16220), .B2(n20116), .A(n16219), .ZN(n16224) );
  AOI22_X1 U19374 ( .A1(n20117), .A2(n16222), .B1(n16231), .B2(n16221), .ZN(
        n16223) );
  OAI211_X1 U19375 ( .C1(n16226), .C2(n16225), .A(n16224), .B(n16223), .ZN(
        P1_U3020) );
  NOR2_X1 U19376 ( .A1(n16228), .A2(n16227), .ZN(n16230) );
  AOI21_X1 U19377 ( .B1(n16230), .B2(n16232), .A(n16229), .ZN(n16242) );
  NAND2_X1 U19378 ( .A1(n16232), .A2(n16231), .ZN(n16246) );
  AOI221_X1 U19379 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n16234), .C2(n16233), .A(
        n16246), .ZN(n16237) );
  INV_X1 U19380 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20750) );
  OAI22_X1 U19381 ( .A1(n16235), .A2(n20107), .B1(n20750), .B2(n16200), .ZN(
        n16236) );
  AOI211_X1 U19382 ( .C1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n16242), .A(
        n16237), .B(n16236), .ZN(n16238) );
  OAI21_X1 U19383 ( .B1(n20091), .B2(n16239), .A(n16238), .ZN(P1_U3021) );
  AOI21_X1 U19384 ( .B1(n16241), .B2(n20116), .A(n16240), .ZN(n16245) );
  AOI22_X1 U19385 ( .A1(n16243), .A2(n20117), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16242), .ZN(n16244) );
  OAI211_X1 U19386 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n16246), .A(
        n16245), .B(n16244), .ZN(P1_U3022) );
  INV_X1 U19387 ( .A(n16247), .ZN(n16254) );
  NAND2_X1 U19388 ( .A1(n20005), .A2(n20116), .ZN(n16249) );
  OAI211_X1 U19389 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16250), .A(
        n16249), .B(n16248), .ZN(n16251) );
  AOI21_X1 U19390 ( .B1(n16252), .B2(n20117), .A(n16251), .ZN(n16253) );
  OAI21_X1 U19391 ( .B1(n16254), .B2(n11040), .A(n16253), .ZN(P1_U3024) );
  NAND3_X1 U19392 ( .A1(n20036), .A2(n16256), .A3(n16255), .ZN(n16258) );
  OAI22_X1 U19393 ( .A1(n16259), .A2(n16258), .B1(n10603), .B2(n16257), .ZN(
        P1_U3468) );
  NAND4_X1 U19394 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20811), .A4(n20819), .ZN(n16260) );
  NAND2_X1 U19395 ( .A1(n16261), .A2(n16260), .ZN(n20715) );
  OAI21_X1 U19396 ( .B1(n16263), .B2(n20715), .A(n16262), .ZN(n16264) );
  OAI221_X1 U19397 ( .B1(n20814), .B2(n20547), .C1(n20814), .C2(n20819), .A(
        n16264), .ZN(n16265) );
  AOI221_X1 U19398 ( .B1(n16266), .B2(n20714), .C1(n20815), .C2(n20714), .A(
        n16265), .ZN(P1_U3162) );
  NOR2_X1 U19399 ( .A1(n16266), .A2(n20815), .ZN(n16268) );
  OAI21_X1 U19400 ( .B1(n16268), .B2(n20547), .A(n16267), .ZN(P1_U3466) );
  AOI211_X1 U19401 ( .C1(n16271), .C2(n16270), .A(n16269), .B(n19090), .ZN(
        n16274) );
  OAI22_X1 U19402 ( .A1(n16272), .A2(n18992), .B1(n19873), .B2(n19129), .ZN(
        n16273) );
  AOI211_X1 U19403 ( .C1(P2_EBX_REG_29__SCAN_IN), .C2(n19126), .A(n16274), .B(
        n16273), .ZN(n16279) );
  INV_X1 U19404 ( .A(n16275), .ZN(n16276) );
  AOI22_X1 U19405 ( .A1(n16277), .A2(n19125), .B1(n16276), .B2(n19133), .ZN(
        n16278) );
  OAI211_X1 U19406 ( .C1(n16280), .C2(n19121), .A(n16279), .B(n16278), .ZN(
        P2_U2826) );
  AOI22_X1 U19407 ( .A1(n19164), .A2(n16281), .B1(n15139), .B2(n19161), .ZN(
        P2_U2856) );
  INV_X1 U19408 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n16286) );
  NOR2_X1 U19409 ( .A1(n16282), .A2(n19161), .ZN(n16283) );
  AOI21_X1 U19410 ( .B1(n16284), .B2(n19151), .A(n16283), .ZN(n16285) );
  OAI21_X1 U19411 ( .B1(n19164), .B2(n16286), .A(n16285), .ZN(P2_U2864) );
  AOI21_X1 U19412 ( .B1(n16288), .B2(n15426), .A(n16287), .ZN(n16300) );
  AOI22_X1 U19413 ( .A1(n16300), .A2(n19151), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n19161), .ZN(n16289) );
  OAI21_X1 U19414 ( .B1(n19161), .B2(n16290), .A(n16289), .ZN(P2_U2865) );
  NOR2_X1 U19415 ( .A1(n14089), .A2(n16291), .ZN(n16292) );
  OR2_X1 U19416 ( .A1(n15424), .A2(n16292), .ZN(n16306) );
  OAI22_X1 U19417 ( .A1(n16306), .A2(n19165), .B1(n19164), .B2(n16293), .ZN(
        n16294) );
  INV_X1 U19418 ( .A(n16294), .ZN(n16295) );
  OAI21_X1 U19419 ( .B1(n19161), .B2(n18984), .A(n16295), .ZN(P2_U2867) );
  AOI21_X1 U19420 ( .B1(n16296), .B2(n13760), .A(n14016), .ZN(n16312) );
  AOI22_X1 U19421 ( .A1(n16312), .A2(n19151), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n19161), .ZN(n16297) );
  OAI21_X1 U19422 ( .B1(n19161), .B2(n16341), .A(n16297), .ZN(P2_U2869) );
  AOI22_X1 U19423 ( .A1(n19172), .A2(n16298), .B1(n19231), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16303) );
  AOI22_X1 U19424 ( .A1(n19174), .A2(BUF2_REG_22__SCAN_IN), .B1(n19173), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n16302) );
  AOI22_X1 U19425 ( .A1(n16300), .A2(n19219), .B1(n19232), .B2(n16299), .ZN(
        n16301) );
  NAND3_X1 U19426 ( .A1(n16303), .A2(n16302), .A3(n16301), .ZN(P2_U2897) );
  AOI22_X1 U19427 ( .A1(n19172), .A2(n16304), .B1(n19231), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16310) );
  AOI22_X1 U19428 ( .A1(n19174), .A2(BUF2_REG_20__SCAN_IN), .B1(n19173), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16309) );
  INV_X1 U19429 ( .A(n18986), .ZN(n16305) );
  OAI22_X1 U19430 ( .A1(n16306), .A2(n19236), .B1(n19180), .B2(n16305), .ZN(
        n16307) );
  INV_X1 U19431 ( .A(n16307), .ZN(n16308) );
  NAND3_X1 U19432 ( .A1(n16310), .A2(n16309), .A3(n16308), .ZN(P2_U2899) );
  AOI22_X1 U19433 ( .A1(n19172), .A2(n16311), .B1(n19231), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16315) );
  AOI22_X1 U19434 ( .A1(n19174), .A2(BUF2_REG_18__SCAN_IN), .B1(n19173), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16314) );
  AOI22_X1 U19435 ( .A1(n16312), .A2(n19219), .B1(n19232), .B2(n16433), .ZN(
        n16313) );
  NAND3_X1 U19436 ( .A1(n16315), .A2(n16314), .A3(n16313), .ZN(P2_U2901) );
  AOI22_X1 U19437 ( .A1(n19284), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19276), .ZN(n16320) );
  AOI222_X1 U19438 ( .A1(n16318), .A2(n19285), .B1(n19294), .B2(n16317), .C1(
        n19288), .C2(n16316), .ZN(n16319) );
  OAI211_X1 U19439 ( .C1(n19291), .C2(n16321), .A(n16320), .B(n16319), .ZN(
        P2_U2990) );
  AOI22_X1 U19440 ( .A1(n19284), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19276), .ZN(n16327) );
  INV_X1 U19441 ( .A(n16322), .ZN(n16325) );
  AOI222_X1 U19442 ( .A1(n16325), .A2(n19285), .B1(n19294), .B2(n16324), .C1(
        n19288), .C2(n16323), .ZN(n16326) );
  OAI211_X1 U19443 ( .C1(n19291), .C2(n16328), .A(n16327), .B(n16326), .ZN(
        P2_U2992) );
  NOR2_X1 U19444 ( .A1(n19291), .A2(n18977), .ZN(n16329) );
  AOI211_X1 U19445 ( .C1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n19284), .A(
        n16330), .B(n16329), .ZN(n16334) );
  OAI211_X1 U19446 ( .C1(n13674), .C2(n18984), .A(n16334), .B(n16333), .ZN(
        P2_U2994) );
  AOI22_X1 U19447 ( .A1(n19284), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19276), .ZN(n16342) );
  INV_X1 U19448 ( .A(n16335), .ZN(n16336) );
  INV_X1 U19449 ( .A(n16341), .ZN(n16436) );
  AOI22_X1 U19450 ( .A1(n19284), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19276), .ZN(n16347) );
  INV_X1 U19451 ( .A(n19146), .ZN(n19030) );
  AOI222_X1 U19452 ( .A1(n16345), .A2(n19285), .B1(n19294), .B2(n19030), .C1(
        n19288), .C2(n16344), .ZN(n16346) );
  OAI211_X1 U19453 ( .C1(n19291), .C2(n19025), .A(n16347), .B(n16346), .ZN(
        P2_U3000) );
  AOI22_X1 U19454 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19276), .B1(n16417), 
        .B2(n19044), .ZN(n16353) );
  INV_X1 U19455 ( .A(n16348), .ZN(n16350) );
  OAI22_X1 U19456 ( .A1(n16350), .A2(n16418), .B1(n16421), .B2(n16349), .ZN(
        n16351) );
  AOI21_X1 U19457 ( .B1(n19294), .B2(n19045), .A(n16351), .ZN(n16352) );
  OAI211_X1 U19458 ( .C1(n16428), .C2(n16354), .A(n16353), .B(n16352), .ZN(
        P2_U3001) );
  AOI22_X1 U19459 ( .A1(n19284), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19276), .ZN(n16362) );
  NAND3_X1 U19460 ( .A1(n16356), .A2(n16355), .A3(n19288), .ZN(n16359) );
  NAND2_X1 U19461 ( .A1(n16357), .A2(n19285), .ZN(n16358) );
  OAI211_X1 U19462 ( .C1(n13674), .C2(n19149), .A(n16359), .B(n16358), .ZN(
        n16360) );
  INV_X1 U19463 ( .A(n16360), .ZN(n16361) );
  OAI211_X1 U19464 ( .C1(n19291), .C2(n19051), .A(n16362), .B(n16361), .ZN(
        P2_U3002) );
  AOI22_X1 U19465 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19276), .B1(n16417), 
        .B2(n16363), .ZN(n16369) );
  OAI22_X1 U19466 ( .A1(n16365), .A2(n16418), .B1(n16364), .B2(n16421), .ZN(
        n16366) );
  AOI21_X1 U19467 ( .B1(n19294), .B2(n16367), .A(n16366), .ZN(n16368) );
  OAI211_X1 U19468 ( .C1(n16428), .C2(n16370), .A(n16369), .B(n16368), .ZN(
        P2_U3003) );
  AOI22_X1 U19469 ( .A1(n19284), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19276), .ZN(n16386) );
  NOR2_X1 U19470 ( .A1(n16372), .A2(n16371), .ZN(n16376) );
  NAND2_X1 U19471 ( .A1(n16374), .A2(n16373), .ZN(n16375) );
  XNOR2_X1 U19472 ( .A(n16376), .B(n16375), .ZN(n16464) );
  INV_X1 U19473 ( .A(n16464), .ZN(n16384) );
  NOR2_X1 U19474 ( .A1(n16377), .A2(n13027), .ZN(n16378) );
  OR2_X1 U19475 ( .A1(n16379), .A2(n16378), .ZN(n19154) );
  INV_X1 U19476 ( .A(n19154), .ZN(n19064) );
  NAND2_X1 U19477 ( .A1(n16381), .A2(n16380), .ZN(n16382) );
  AND2_X1 U19478 ( .A1(n16383), .A2(n16382), .ZN(n16461) );
  AOI222_X1 U19479 ( .A1(n16384), .A2(n19285), .B1(n19294), .B2(n19064), .C1(
        n19288), .C2(n16461), .ZN(n16385) );
  OAI211_X1 U19480 ( .C1(n19291), .C2(n19062), .A(n16386), .B(n16385), .ZN(
        P2_U3004) );
  AOI22_X1 U19481 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19276), .B1(n16417), 
        .B2(n19069), .ZN(n16391) );
  OAI22_X1 U19482 ( .A1(n16388), .A2(n16418), .B1(n16421), .B2(n16387), .ZN(
        n16389) );
  AOI21_X1 U19483 ( .B1(n19294), .B2(n19073), .A(n16389), .ZN(n16390) );
  OAI211_X1 U19484 ( .C1(n16428), .C2(n16392), .A(n16391), .B(n16390), .ZN(
        P2_U3005) );
  AOI22_X1 U19485 ( .A1(n19284), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19276), .ZN(n16408) );
  INV_X1 U19486 ( .A(n16393), .ZN(n16394) );
  XNOR2_X1 U19487 ( .A(n16395), .B(n16394), .ZN(n16465) );
  NAND2_X1 U19488 ( .A1(n16465), .A2(n19288), .ZN(n16405) );
  NAND2_X1 U19489 ( .A1(n13909), .A2(n16396), .ZN(n16398) );
  NAND2_X1 U19490 ( .A1(n16398), .A2(n16397), .ZN(n16403) );
  INV_X1 U19491 ( .A(n16399), .ZN(n16401) );
  NAND2_X1 U19492 ( .A1(n16401), .A2(n16400), .ZN(n16402) );
  XNOR2_X1 U19493 ( .A(n16403), .B(n16402), .ZN(n16469) );
  NAND2_X1 U19494 ( .A1(n16469), .A2(n19285), .ZN(n16404) );
  OAI211_X1 U19495 ( .C1(n13674), .C2(n19162), .A(n16405), .B(n16404), .ZN(
        n16406) );
  INV_X1 U19496 ( .A(n16406), .ZN(n16407) );
  OAI211_X1 U19497 ( .C1(n19291), .C2(n16409), .A(n16408), .B(n16407), .ZN(
        P2_U3006) );
  AOI22_X1 U19498 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19276), .B1(n16417), 
        .B2(n19115), .ZN(n16414) );
  OAI22_X1 U19499 ( .A1(n16411), .A2(n16421), .B1(n16418), .B2(n16410), .ZN(
        n16412) );
  AOI21_X1 U19500 ( .B1(n19294), .B2(n19116), .A(n16412), .ZN(n16413) );
  OAI211_X1 U19501 ( .C1(n16428), .C2(n16415), .A(n16414), .B(n16413), .ZN(
        P2_U3009) );
  AOI22_X1 U19502 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19276), .B1(n16417), 
        .B2(n16416), .ZN(n16427) );
  NOR3_X1 U19503 ( .A1(n16420), .A2(n16419), .A3(n16418), .ZN(n16424) );
  NOR2_X1 U19504 ( .A1(n16422), .A2(n16421), .ZN(n16423) );
  AOI211_X1 U19505 ( .C1(n19294), .C2(n16425), .A(n16424), .B(n16423), .ZN(
        n16426) );
  OAI211_X1 U19506 ( .C1(n16429), .C2(n16428), .A(n16427), .B(n16426), .ZN(
        P2_U3011) );
  AOI21_X1 U19507 ( .B1(n16432), .B2(n16431), .A(n16430), .ZN(n16442) );
  AND2_X1 U19508 ( .A1(n16493), .A2(n16433), .ZN(n16435) );
  AOI211_X1 U19509 ( .C1(n19276), .C2(P2_REIP_REG_18__SCAN_IN), .A(n16435), 
        .B(n16434), .ZN(n16440) );
  AOI222_X1 U19510 ( .A1(n16438), .A2(n16485), .B1(n16460), .B2(n16437), .C1(
        n16494), .C2(n16436), .ZN(n16439) );
  OAI211_X1 U19511 ( .C1(n16442), .C2(n16441), .A(n16440), .B(n16439), .ZN(
        P2_U3028) );
  OAI21_X1 U19512 ( .B1(n9793), .B2(n9829), .A(n16443), .ZN(n19182) );
  OAI22_X1 U19513 ( .A1(n16479), .A2(n19182), .B1(n15617), .B2(n9725), .ZN(
        n16444) );
  AOI221_X1 U19514 ( .B1(n16447), .B2(n16446), .C1(n16445), .C2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(n16444), .ZN(n16451) );
  AOI22_X1 U19515 ( .A1(n16449), .A2(n16460), .B1(n16494), .B2(n16448), .ZN(
        n16450) );
  OAI211_X1 U19516 ( .C1(n16452), .C2(n16498), .A(n16451), .B(n16450), .ZN(
        P2_U3031) );
  NOR2_X1 U19517 ( .A1(n12015), .A2(n9725), .ZN(n16457) );
  XNOR2_X1 U19518 ( .A(n16454), .B(n16453), .ZN(n19196) );
  OAI22_X1 U19519 ( .A1(n16455), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n19196), .B2(n16479), .ZN(n16456) );
  AOI211_X1 U19520 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n16458), .A(
        n16457), .B(n16456), .ZN(n16463) );
  NOR2_X1 U19521 ( .A1(n16466), .A2(n19154), .ZN(n16459) );
  AOI21_X1 U19522 ( .B1(n16461), .B2(n16460), .A(n16459), .ZN(n16462) );
  OAI211_X1 U19523 ( .C1(n16464), .C2(n16498), .A(n16463), .B(n16462), .ZN(
        P2_U3036) );
  AOI22_X1 U19524 ( .A1(n16481), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16493), .B2(n19202), .ZN(n16476) );
  INV_X1 U19525 ( .A(n16465), .ZN(n16467) );
  OAI22_X1 U19526 ( .A1(n16467), .A2(n16503), .B1(n16466), .B2(n19162), .ZN(
        n16468) );
  AOI21_X1 U19527 ( .B1(n16485), .B2(n16469), .A(n16468), .ZN(n16475) );
  NAND2_X1 U19528 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19276), .ZN(n16474) );
  NOR3_X1 U19529 ( .A1(n20980), .A2(n16471), .A3(n16470), .ZN(n16483) );
  OAI221_X1 U19530 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16472), .C2(n16482), .A(
        n16483), .ZN(n16473) );
  NAND4_X1 U19531 ( .A1(n16476), .A2(n16475), .A3(n16474), .A4(n16473), .ZN(
        P2_U3038) );
  OAI21_X1 U19532 ( .B1(n16478), .B2(n16477), .A(n15334), .ZN(n19204) );
  OAI22_X1 U19533 ( .A1(n16479), .A2(n19204), .B1(n12005), .B2(n9725), .ZN(
        n16480) );
  AOI221_X1 U19534 ( .B1(n16483), .B2(n16482), .C1(n16481), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16480), .ZN(n16488) );
  AOI22_X1 U19535 ( .A1(n16486), .A2(n16485), .B1(n16494), .B2(n16484), .ZN(
        n16487) );
  OAI211_X1 U19536 ( .C1(n16503), .C2(n16489), .A(n16488), .B(n16487), .ZN(
        P2_U3039) );
  MUX2_X1 U19537 ( .A(n16491), .B(n16490), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n16496) );
  INV_X1 U19538 ( .A(n16492), .ZN(n19122) );
  AOI22_X1 U19539 ( .A1(n16494), .A2(n12816), .B1(n16493), .B2(n19122), .ZN(
        n16495) );
  OAI211_X1 U19540 ( .C1(n16498), .C2(n16497), .A(n16496), .B(n16495), .ZN(
        n16499) );
  INV_X1 U19541 ( .A(n16499), .ZN(n16501) );
  OAI211_X1 U19542 ( .C1(n16503), .C2(n16502), .A(n16501), .B(n16500), .ZN(
        P2_U3046) );
  AOI211_X1 U19543 ( .C1(n16507), .C2(n16506), .A(n16505), .B(n16504), .ZN(
        n16515) );
  MUX2_X1 U19544 ( .A(n16508), .B(n16509), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n16513) );
  INV_X1 U19545 ( .A(n16509), .ZN(n16512) );
  NAND2_X1 U19546 ( .A1(n16510), .A2(n19952), .ZN(n16511) );
  OAI22_X1 U19547 ( .A1(n16513), .A2(n19947), .B1(n16512), .B2(n16511), .ZN(
        n16514) );
  OAI211_X1 U19548 ( .C1(n16517), .C2(n16516), .A(n16515), .B(n16514), .ZN(
        P2_U3176) );
  OAI22_X1 U19549 ( .A1(n18156), .A2(n17972), .B1(n17808), .B2(n17833), .ZN(
        n17847) );
  NAND2_X1 U19550 ( .A1(n16518), .A2(n17769), .ZN(n17701) );
  INV_X1 U19551 ( .A(n17701), .ZN(n17619) );
  NAND2_X1 U19552 ( .A1(n16519), .A2(n17619), .ZN(n17629) );
  OAI21_X1 U19553 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16535), .A(
        n16520), .ZN(n16697) );
  NOR2_X1 U19554 ( .A1(n17817), .A2(n16697), .ZN(n16525) );
  INV_X1 U19555 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16700) );
  OAI221_X1 U19556 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16523), .C1(
        n16700), .C2(n16522), .A(n16521), .ZN(n16524) );
  AOI211_X1 U19557 ( .C1(n17861), .C2(n16526), .A(n16525), .B(n16524), .ZN(
        n16530) );
  AOI21_X1 U19558 ( .B1(n17978), .B2(n16527), .A(n17972), .ZN(n16544) );
  NOR2_X1 U19559 ( .A1(n16528), .A2(n17808), .ZN(n16534) );
  OAI21_X1 U19560 ( .B1(n16544), .B2(n16534), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16529) );
  OAI211_X1 U19561 ( .C1(n17629), .C2(n16531), .A(n16530), .B(n16529), .ZN(
        P3_U2800) );
  INV_X1 U19562 ( .A(n17978), .ZN(n16532) );
  NOR2_X1 U19563 ( .A1(n16532), .A2(n16533), .ZN(n16562) );
  NOR2_X1 U19564 ( .A1(n16533), .A2(n17981), .ZN(n16561) );
  OAI21_X1 U19565 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16561), .A(
        n16534), .ZN(n16541) );
  AOI21_X1 U19566 ( .B1(n16719), .B2(n16536), .A(n16535), .ZN(n16713) );
  OAI21_X1 U19567 ( .B1(n16537), .B2(n17730), .A(n16713), .ZN(n16540) );
  OAI221_X1 U19568 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n9828), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n18678), .A(n16538), .ZN(
        n16539) );
  NAND4_X1 U19569 ( .A1(n16542), .A2(n16541), .A3(n16540), .A4(n16539), .ZN(
        n16543) );
  AOI221_X1 U19570 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16544), 
        .C1(n16562), .C2(n16544), .A(n16543), .ZN(n16545) );
  OAI21_X1 U19571 ( .B1(n17879), .B2(n16546), .A(n16545), .ZN(P3_U2801) );
  OAI21_X1 U19572 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18267), .A(
        n16547), .ZN(n16549) );
  AOI21_X1 U19573 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16549), .A(
        n16548), .ZN(n16557) );
  INV_X1 U19574 ( .A(n16550), .ZN(n16553) );
  OAI22_X1 U19575 ( .A1(n16553), .A2(n18153), .B1(n16552), .B2(n16551), .ZN(
        n16554) );
  AOI22_X1 U19576 ( .A1(n16555), .A2(n18181), .B1(n18265), .B2(n16554), .ZN(
        n16556) );
  OAI211_X1 U19577 ( .C1(n16558), .C2(n18257), .A(n16557), .B(n16556), .ZN(
        P3_U2831) );
  INV_X1 U19578 ( .A(n17625), .ZN(n16559) );
  AOI21_X1 U19579 ( .B1(n17795), .B2(n16559), .A(n17626), .ZN(n17616) );
  NAND2_X1 U19580 ( .A1(n16560), .A2(n17616), .ZN(n16575) );
  AOI21_X1 U19581 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17868), .A(
        n16560), .ZN(n17615) );
  NOR2_X1 U19582 ( .A1(n17616), .A2(n17615), .ZN(n17614) );
  NOR2_X1 U19583 ( .A1(n17614), .A2(n18106), .ZN(n16566) );
  OAI22_X1 U19584 ( .A1(n16562), .A2(n18029), .B1(n16561), .B2(n18153), .ZN(
        n16563) );
  AOI211_X1 U19585 ( .C1(n16566), .C2(n16565), .A(n16564), .B(n16563), .ZN(
        n16567) );
  NOR2_X1 U19586 ( .A1(n16567), .A2(n17613), .ZN(n16572) );
  INV_X1 U19587 ( .A(n17833), .ZN(n18154) );
  INV_X1 U19588 ( .A(n18153), .ZN(n18192) );
  AOI22_X1 U19589 ( .A1(n18767), .A2(n17777), .B1(n18154), .B2(n18192), .ZN(
        n18078) );
  OAI21_X1 U19590 ( .B1(n18078), .B2(n16569), .A(n16568), .ZN(n18043) );
  NAND2_X1 U19591 ( .A1(n16570), .A2(n18043), .ZN(n18037) );
  NOR4_X1 U19592 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18281), .A3(
        n17611), .A4(n18037), .ZN(n16571) );
  AOI221_X1 U19593 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(n18125), .C1(n16572), 
        .C2(n18280), .A(n16571), .ZN(n16574) );
  NAND3_X1 U19594 ( .A1(n17626), .A2(n18181), .A3(n17615), .ZN(n16573) );
  OAI211_X1 U19595 ( .C1(n16575), .C2(n18274), .A(n16574), .B(n16573), .ZN(
        P3_U2834) );
  NOR3_X1 U19596 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16577) );
  NOR4_X1 U19597 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16576) );
  NAND4_X1 U19598 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16577), .A3(n16576), .A4(
        U215), .ZN(U213) );
  INV_X1 U19599 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19241) );
  INV_X2 U19600 ( .A(U214), .ZN(n16622) );
  NOR2_X1 U19601 ( .A1(n16622), .A2(n16578), .ZN(n16619) );
  INV_X1 U19602 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16657) );
  OAI222_X1 U19603 ( .A1(U212), .A2(n19241), .B1(n16624), .B2(n19339), .C1(
        U214), .C2(n16657), .ZN(U216) );
  INV_X1 U19604 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n19329) );
  AOI22_X1 U19605 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16621), .ZN(n16579) );
  OAI21_X1 U19606 ( .B1(n19329), .B2(n16624), .A(n16579), .ZN(U217) );
  INV_X1 U19607 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16581) );
  AOI22_X1 U19608 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16621), .ZN(n16580) );
  OAI21_X1 U19609 ( .B1(n16581), .B2(n16624), .A(n16580), .ZN(U218) );
  AOI22_X1 U19610 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16621), .ZN(n16582) );
  OAI21_X1 U19611 ( .B1(n16583), .B2(n16624), .A(n16582), .ZN(U219) );
  AOI22_X1 U19612 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16621), .ZN(n16584) );
  OAI21_X1 U19613 ( .B1(n19318), .B2(n16624), .A(n16584), .ZN(U220) );
  AOI22_X1 U19614 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16621), .ZN(n16585) );
  OAI21_X1 U19615 ( .B1(n20859), .B2(n16624), .A(n16585), .ZN(U221) );
  INV_X1 U19616 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n19311) );
  AOI22_X1 U19617 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16621), .ZN(n16586) );
  OAI21_X1 U19618 ( .B1(n19311), .B2(n16624), .A(n16586), .ZN(U222) );
  INV_X1 U19619 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n16648) );
  OAI222_X1 U19620 ( .A1(U212), .A2(n16648), .B1(n16624), .B2(n16587), .C1(
        U214), .C2(n13090), .ZN(U223) );
  INV_X1 U19621 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16589) );
  AOI22_X1 U19622 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16621), .ZN(n16588) );
  OAI21_X1 U19623 ( .B1(n16589), .B2(n16624), .A(n16588), .ZN(U224) );
  AOI22_X1 U19624 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16621), .ZN(n16590) );
  OAI21_X1 U19625 ( .B1(n14671), .B2(n16624), .A(n16590), .ZN(U225) );
  INV_X1 U19626 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20887) );
  AOI22_X1 U19627 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16621), .ZN(n16591) );
  OAI21_X1 U19628 ( .B1(n20887), .B2(n16624), .A(n16591), .ZN(U226) );
  AOI22_X1 U19629 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16621), .ZN(n16592) );
  OAI21_X1 U19630 ( .B1(n16593), .B2(n16624), .A(n16592), .ZN(U227) );
  INV_X1 U19631 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16595) );
  AOI22_X1 U19632 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16621), .ZN(n16594) );
  OAI21_X1 U19633 ( .B1(n16595), .B2(n16624), .A(n16594), .ZN(U228) );
  INV_X1 U19634 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16597) );
  AOI22_X1 U19635 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16621), .ZN(n16596) );
  OAI21_X1 U19636 ( .B1(n16597), .B2(n16624), .A(n16596), .ZN(U229) );
  INV_X1 U19637 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16599) );
  AOI22_X1 U19638 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16621), .ZN(n16598) );
  OAI21_X1 U19639 ( .B1(n16599), .B2(n16624), .A(n16598), .ZN(U230) );
  INV_X1 U19640 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16601) );
  AOI22_X1 U19641 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16621), .ZN(n16600) );
  OAI21_X1 U19642 ( .B1(n16601), .B2(n16624), .A(n16600), .ZN(U231) );
  AOI22_X1 U19643 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n16619), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16621), .ZN(n16602) );
  OAI21_X1 U19644 ( .B1(n13441), .B2(U214), .A(n16602), .ZN(U232) );
  INV_X1 U19645 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16638) );
  AOI22_X1 U19646 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16619), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16622), .ZN(n16603) );
  OAI21_X1 U19647 ( .B1(n16638), .B2(U212), .A(n16603), .ZN(U233) );
  INV_X1 U19648 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16636) );
  AOI22_X1 U19649 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n16619), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16622), .ZN(n16604) );
  OAI21_X1 U19650 ( .B1(n16636), .B2(U212), .A(n16604), .ZN(U234) );
  INV_X1 U19651 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n20891) );
  OAI222_X1 U19652 ( .A1(U212), .A2(n20891), .B1(n16624), .B2(n16605), .C1(
        U214), .C2(n13418), .ZN(U235) );
  INV_X1 U19653 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16635) );
  AOI22_X1 U19654 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16619), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16622), .ZN(n16606) );
  OAI21_X1 U19655 ( .B1(n16635), .B2(U212), .A(n16606), .ZN(U236) );
  AOI22_X1 U19656 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16621), .ZN(n16607) );
  OAI21_X1 U19657 ( .B1(n16608), .B2(n16624), .A(n16607), .ZN(U237) );
  AOI22_X1 U19658 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16621), .ZN(n16609) );
  OAI21_X1 U19659 ( .B1(n21045), .B2(n16624), .A(n16609), .ZN(U238) );
  AOI22_X1 U19660 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16621), .ZN(n16610) );
  OAI21_X1 U19661 ( .B1(n16611), .B2(n16624), .A(n16610), .ZN(U239) );
  AOI22_X1 U19662 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16619), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16621), .ZN(n16612) );
  OAI21_X1 U19663 ( .B1(n13427), .B2(U214), .A(n16612), .ZN(U240) );
  INV_X1 U19664 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16614) );
  AOI22_X1 U19665 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16621), .ZN(n16613) );
  OAI21_X1 U19666 ( .B1(n16614), .B2(n16624), .A(n16613), .ZN(U241) );
  INV_X1 U19667 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n20946) );
  AOI22_X1 U19668 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16619), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16622), .ZN(n16615) );
  OAI21_X1 U19669 ( .B1(n20946), .B2(U212), .A(n16615), .ZN(U242) );
  AOI222_X1 U19670 ( .A1(n16621), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n16619), 
        .B2(BUF1_REG_4__SCAN_IN), .C1(n16622), .C2(P1_DATAO_REG_4__SCAN_IN), 
        .ZN(n16616) );
  INV_X1 U19671 ( .A(n16616), .ZN(U243) );
  INV_X1 U19672 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16629) );
  AOI22_X1 U19673 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16619), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16622), .ZN(n16617) );
  OAI21_X1 U19674 ( .B1(n16629), .B2(U212), .A(n16617), .ZN(U244) );
  INV_X1 U19675 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16628) );
  OAI222_X1 U19676 ( .A1(U212), .A2(n16628), .B1(n16624), .B2(n16618), .C1(
        U214), .C2(n13106), .ZN(U245) );
  INV_X1 U19677 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16627) );
  AOI22_X1 U19678 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16619), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16622), .ZN(n16620) );
  OAI21_X1 U19679 ( .B1(n16627), .B2(U212), .A(n16620), .ZN(U246) );
  AOI22_X1 U19680 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16622), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16621), .ZN(n16623) );
  OAI21_X1 U19681 ( .B1(n16625), .B2(n16624), .A(n16623), .ZN(U247) );
  INV_X1 U19682 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16626) );
  AOI22_X1 U19683 ( .A1(n16656), .A2(n16626), .B1(n18296), .B2(U215), .ZN(U251) );
  INV_X1 U19684 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18304) );
  AOI22_X1 U19685 ( .A1(n16656), .A2(n16627), .B1(n18304), .B2(U215), .ZN(U252) );
  AOI22_X1 U19686 ( .A1(n16656), .A2(n16628), .B1(n18308), .B2(U215), .ZN(U253) );
  INV_X1 U19687 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18312) );
  AOI22_X1 U19688 ( .A1(n16656), .A2(n16629), .B1(n18312), .B2(U215), .ZN(U254) );
  INV_X1 U19689 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n20998) );
  INV_X1 U19690 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18317) );
  AOI22_X1 U19691 ( .A1(n16651), .A2(n20998), .B1(n18317), .B2(U215), .ZN(U255) );
  INV_X1 U19692 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18321) );
  AOI22_X1 U19693 ( .A1(n16656), .A2(n20946), .B1(n18321), .B2(U215), .ZN(U256) );
  INV_X1 U19694 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16630) );
  INV_X1 U19695 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18325) );
  AOI22_X1 U19696 ( .A1(n16656), .A2(n16630), .B1(n18325), .B2(U215), .ZN(U257) );
  INV_X1 U19697 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16631) );
  INV_X1 U19698 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18329) );
  AOI22_X1 U19699 ( .A1(n16656), .A2(n16631), .B1(n18329), .B2(U215), .ZN(U258) );
  INV_X1 U19700 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16632) );
  INV_X1 U19701 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17583) );
  AOI22_X1 U19702 ( .A1(n16656), .A2(n16632), .B1(n17583), .B2(U215), .ZN(U259) );
  INV_X1 U19703 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16633) );
  INV_X1 U19704 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17585) );
  AOI22_X1 U19705 ( .A1(n16651), .A2(n16633), .B1(n17585), .B2(U215), .ZN(U260) );
  INV_X1 U19706 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16634) );
  INV_X1 U19707 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17587) );
  AOI22_X1 U19708 ( .A1(n16656), .A2(n16634), .B1(n17587), .B2(U215), .ZN(U261) );
  INV_X1 U19709 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17589) );
  AOI22_X1 U19710 ( .A1(n16656), .A2(n16635), .B1(n17589), .B2(U215), .ZN(U262) );
  INV_X1 U19711 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17593) );
  AOI22_X1 U19712 ( .A1(n16656), .A2(n20891), .B1(n17593), .B2(U215), .ZN(U263) );
  INV_X1 U19713 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17596) );
  AOI22_X1 U19714 ( .A1(n16651), .A2(n16636), .B1(n17596), .B2(U215), .ZN(U264) );
  INV_X1 U19715 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n16637) );
  AOI22_X1 U19716 ( .A1(n16656), .A2(n16638), .B1(n16637), .B2(U215), .ZN(U265) );
  OAI22_X1 U19717 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16651), .ZN(n16639) );
  INV_X1 U19718 ( .A(n16639), .ZN(U266) );
  OAI22_X1 U19719 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16656), .ZN(n16640) );
  INV_X1 U19720 ( .A(n16640), .ZN(U267) );
  OAI22_X1 U19721 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16656), .ZN(n16641) );
  INV_X1 U19722 ( .A(n16641), .ZN(U268) );
  OAI22_X1 U19723 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16651), .ZN(n16642) );
  INV_X1 U19724 ( .A(n16642), .ZN(U269) );
  INV_X1 U19725 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n16643) );
  INV_X1 U19726 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n20937) );
  AOI22_X1 U19727 ( .A1(n16651), .A2(n16643), .B1(n20937), .B2(U215), .ZN(U270) );
  OAI22_X1 U19728 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16651), .ZN(n16644) );
  INV_X1 U19729 ( .A(n16644), .ZN(U271) );
  OAI22_X1 U19730 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16651), .ZN(n16645) );
  INV_X1 U19731 ( .A(n16645), .ZN(U272) );
  OAI22_X1 U19732 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16656), .ZN(n16646) );
  INV_X1 U19733 ( .A(n16646), .ZN(U273) );
  OAI22_X1 U19734 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16656), .ZN(n16647) );
  INV_X1 U19735 ( .A(n16647), .ZN(U274) );
  AOI22_X1 U19736 ( .A1(n16656), .A2(n16648), .B1(n17382), .B2(U215), .ZN(U275) );
  INV_X1 U19737 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n16649) );
  INV_X1 U19738 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n19310) );
  AOI22_X1 U19739 ( .A1(n16651), .A2(n16649), .B1(n19310), .B2(U215), .ZN(U276) );
  INV_X1 U19740 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n16650) );
  AOI22_X1 U19741 ( .A1(n16651), .A2(n16650), .B1(n17370), .B2(U215), .ZN(U277) );
  INV_X1 U19742 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n16652) );
  INV_X1 U19743 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n20947) );
  AOI22_X1 U19744 ( .A1(n16656), .A2(n16652), .B1(n20947), .B2(U215), .ZN(U278) );
  INV_X1 U19745 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16653) );
  AOI22_X1 U19746 ( .A1(n16656), .A2(n16653), .B1(n17361), .B2(U215), .ZN(U279) );
  OAI22_X1 U19747 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16656), .ZN(n16654) );
  INV_X1 U19748 ( .A(n16654), .ZN(U280) );
  INV_X1 U19749 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n16655) );
  INV_X1 U19750 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19330) );
  AOI22_X1 U19751 ( .A1(n16656), .A2(n16655), .B1(n19330), .B2(U215), .ZN(U281) );
  INV_X1 U19752 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19337) );
  AOI22_X1 U19753 ( .A1(n16656), .A2(n19241), .B1(n19337), .B2(U215), .ZN(U282) );
  INV_X1 U19754 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17493) );
  AOI222_X1 U19755 ( .A1(n16657), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19241), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n17493), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16658) );
  INV_X2 U19756 ( .A(n16660), .ZN(n16659) );
  INV_X1 U19757 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18839) );
  INV_X1 U19758 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19850) );
  AOI22_X1 U19759 ( .A1(n16659), .A2(n18839), .B1(n19850), .B2(n16660), .ZN(
        U347) );
  INV_X1 U19760 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18837) );
  INV_X1 U19761 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19849) );
  AOI22_X1 U19762 ( .A1(n16659), .A2(n18837), .B1(n19849), .B2(n16660), .ZN(
        U348) );
  INV_X1 U19763 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18834) );
  INV_X1 U19764 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19848) );
  AOI22_X1 U19765 ( .A1(n16659), .A2(n18834), .B1(n19848), .B2(n16660), .ZN(
        U349) );
  INV_X1 U19766 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18833) );
  INV_X1 U19767 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19847) );
  AOI22_X1 U19768 ( .A1(n16659), .A2(n18833), .B1(n19847), .B2(n16660), .ZN(
        U350) );
  INV_X1 U19769 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18831) );
  INV_X1 U19770 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19846) );
  AOI22_X1 U19771 ( .A1(n16659), .A2(n18831), .B1(n19846), .B2(n16660), .ZN(
        U351) );
  INV_X1 U19772 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18830) );
  INV_X1 U19773 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19844) );
  AOI22_X1 U19774 ( .A1(n16659), .A2(n18830), .B1(n19844), .B2(n16660), .ZN(
        U352) );
  INV_X1 U19775 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18828) );
  INV_X1 U19776 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19843) );
  AOI22_X1 U19777 ( .A1(n16659), .A2(n18828), .B1(n19843), .B2(n16660), .ZN(
        U353) );
  INV_X1 U19778 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18826) );
  AOI22_X1 U19779 ( .A1(n16659), .A2(n18826), .B1(n19842), .B2(n16660), .ZN(
        U354) );
  INV_X1 U19780 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n21036) );
  INV_X1 U19781 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20965) );
  AOI22_X1 U19782 ( .A1(n16659), .A2(n21036), .B1(n20965), .B2(n16660), .ZN(
        U355) );
  INV_X1 U19783 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18872) );
  INV_X1 U19784 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19874) );
  AOI22_X1 U19785 ( .A1(n16659), .A2(n18872), .B1(n19874), .B2(n16660), .ZN(
        U356) );
  INV_X1 U19786 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n20933) );
  INV_X1 U19787 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19872) );
  AOI22_X1 U19788 ( .A1(n16659), .A2(n20933), .B1(n19872), .B2(n16660), .ZN(
        U357) );
  INV_X1 U19789 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n20902) );
  INV_X1 U19790 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19870) );
  AOI22_X1 U19791 ( .A1(n16659), .A2(n20902), .B1(n19870), .B2(n16660), .ZN(
        U358) );
  INV_X1 U19792 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18868) );
  INV_X1 U19793 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20936) );
  AOI22_X1 U19794 ( .A1(n16659), .A2(n18868), .B1(n20936), .B2(n16660), .ZN(
        U359) );
  INV_X1 U19795 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18866) );
  INV_X1 U19796 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19868) );
  AOI22_X1 U19797 ( .A1(n16659), .A2(n18866), .B1(n19868), .B2(n16660), .ZN(
        U360) );
  INV_X1 U19798 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18863) );
  INV_X1 U19799 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19866) );
  AOI22_X1 U19800 ( .A1(n16659), .A2(n18863), .B1(n19866), .B2(n16660), .ZN(
        U361) );
  INV_X1 U19801 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18861) );
  INV_X1 U19802 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19865) );
  AOI22_X1 U19803 ( .A1(n16659), .A2(n18861), .B1(n19865), .B2(n16660), .ZN(
        U362) );
  INV_X1 U19804 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18859) );
  INV_X1 U19805 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19864) );
  AOI22_X1 U19806 ( .A1(n16659), .A2(n18859), .B1(n19864), .B2(n16660), .ZN(
        U363) );
  INV_X1 U19807 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18858) );
  INV_X1 U19808 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19863) );
  AOI22_X1 U19809 ( .A1(n16659), .A2(n18858), .B1(n19863), .B2(n16660), .ZN(
        U364) );
  INV_X1 U19810 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18824) );
  INV_X1 U19811 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19841) );
  AOI22_X1 U19812 ( .A1(n16659), .A2(n18824), .B1(n19841), .B2(n16660), .ZN(
        U365) );
  INV_X1 U19813 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18857) );
  INV_X1 U19814 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19862) );
  AOI22_X1 U19815 ( .A1(n16659), .A2(n18857), .B1(n19862), .B2(n16660), .ZN(
        U366) );
  INV_X1 U19816 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18855) );
  INV_X1 U19817 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19861) );
  AOI22_X1 U19818 ( .A1(n16659), .A2(n18855), .B1(n19861), .B2(n16660), .ZN(
        U367) );
  INV_X1 U19819 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n20829) );
  INV_X1 U19820 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19860) );
  AOI22_X1 U19821 ( .A1(n16659), .A2(n20829), .B1(n19860), .B2(n16660), .ZN(
        U368) );
  INV_X1 U19822 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18853) );
  INV_X1 U19823 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19859) );
  AOI22_X1 U19824 ( .A1(n16659), .A2(n18853), .B1(n19859), .B2(n16660), .ZN(
        U369) );
  INV_X1 U19825 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18851) );
  INV_X1 U19826 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19857) );
  AOI22_X1 U19827 ( .A1(n16659), .A2(n18851), .B1(n19857), .B2(n16660), .ZN(
        U370) );
  INV_X1 U19828 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18849) );
  INV_X1 U19829 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19855) );
  AOI22_X1 U19830 ( .A1(n16659), .A2(n18849), .B1(n19855), .B2(n16660), .ZN(
        U371) );
  INV_X1 U19831 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18846) );
  INV_X1 U19832 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19854) );
  AOI22_X1 U19833 ( .A1(n16659), .A2(n18846), .B1(n19854), .B2(n16660), .ZN(
        U372) );
  INV_X1 U19834 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18845) );
  INV_X1 U19835 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19853) );
  AOI22_X1 U19836 ( .A1(n16659), .A2(n18845), .B1(n19853), .B2(n16660), .ZN(
        U373) );
  INV_X1 U19837 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18843) );
  INV_X1 U19838 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19852) );
  AOI22_X1 U19839 ( .A1(n16659), .A2(n18843), .B1(n19852), .B2(n16660), .ZN(
        U374) );
  INV_X1 U19840 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18841) );
  INV_X1 U19841 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19851) );
  AOI22_X1 U19842 ( .A1(n16659), .A2(n18841), .B1(n19851), .B2(n16660), .ZN(
        U375) );
  INV_X1 U19843 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18821) );
  INV_X1 U19844 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19840) );
  AOI22_X1 U19845 ( .A1(n16659), .A2(n18821), .B1(n19840), .B2(n16660), .ZN(
        U376) );
  INV_X1 U19846 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16661) );
  INV_X1 U19847 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18820) );
  NAND2_X1 U19848 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18820), .ZN(n18808) );
  AOI22_X1 U19849 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18808), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18818), .ZN(n18884) );
  OAI21_X1 U19850 ( .B1(n18818), .B2(n16661), .A(n18882), .ZN(P3_U2633) );
  OAI21_X1 U19851 ( .B1(n16662), .B2(n17551), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16663) );
  OAI21_X1 U19852 ( .B1(n16664), .B2(n18796), .A(n16663), .ZN(P3_U2634) );
  AOI21_X1 U19853 ( .B1(n18818), .B2(n18820), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16665) );
  AOI22_X1 U19854 ( .A1(n18942), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16665), 
        .B2(n18943), .ZN(P3_U2635) );
  NOR2_X1 U19855 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18805) );
  OAI21_X1 U19856 ( .B1(n18805), .B2(BS16), .A(n18884), .ZN(n18883) );
  OAI21_X1 U19857 ( .B1(n18884), .B2(n16666), .A(n18883), .ZN(P3_U2636) );
  AND3_X1 U19858 ( .A1(n16668), .A2(n16667), .A3(n18772), .ZN(n18776) );
  NOR2_X1 U19859 ( .A1(n18776), .A2(n18792), .ZN(n18925) );
  OAI21_X1 U19860 ( .B1(n18925), .B2(n18287), .A(n16669), .ZN(P3_U2637) );
  NOR4_X1 U19861 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A3(P3_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n16679) );
  NOR4_X1 U19862 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_6__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n16678) );
  NOR4_X1 U19863 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(n16670) );
  INV_X1 U19864 ( .A(P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20978) );
  INV_X1 U19865 ( .A(P3_DATAWIDTH_REG_8__SCAN_IN), .ZN(n20919) );
  NAND3_X1 U19866 ( .A1(n16670), .A2(n20978), .A3(n20919), .ZN(n16676) );
  NOR4_X1 U19867 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_19__SCAN_IN), .A3(P3_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_21__SCAN_IN), .ZN(n16674) );
  NOR4_X1 U19868 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_15__SCAN_IN), .A3(P3_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(n16673) );
  NOR4_X1 U19869 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16672) );
  NOR4_X1 U19870 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16671) );
  NAND4_X1 U19871 ( .A1(n16674), .A2(n16673), .A3(n16672), .A4(n16671), .ZN(
        n16675) );
  AOI211_X1 U19872 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(n16676), .B(n16675), .ZN(n16677) );
  NAND3_X1 U19873 ( .A1(n16679), .A2(n16678), .A3(n16677), .ZN(n18921) );
  NOR2_X1 U19874 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18921), .ZN(n18923) );
  OR4_X1 U19875 ( .A1(n18921), .A2(P3_REIP_REG_0__SCAN_IN), .A3(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A4(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16680) );
  INV_X1 U19876 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18879) );
  AOI22_X1 U19877 ( .A1(n18923), .A2(n16680), .B1(n18921), .B2(n18879), .ZN(
        P3_U2638) );
  INV_X1 U19878 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20995) );
  AOI22_X1 U19879 ( .A1(P3_BYTEENABLE_REG_3__SCAN_IN), .A2(n18921), .B1(n18923), .B2(n20995), .ZN(n16681) );
  NAND2_X1 U19880 ( .A1(n16681), .A2(n16680), .ZN(P3_U2639) );
  NAND2_X1 U19881 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16682), .ZN(
        n16685) );
  OAI21_X1 U19882 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16682), .A(
        n16685), .ZN(n17634) );
  INV_X1 U19883 ( .A(n17634), .ZN(n16733) );
  NOR2_X1 U19884 ( .A1(n16683), .A2(n16933), .ZN(n16732) );
  NOR2_X1 U19885 ( .A1(n16733), .A2(n16732), .ZN(n16731) );
  NOR2_X1 U19886 ( .A1(n16731), .A2(n16933), .ZN(n16722) );
  AOI21_X1 U19887 ( .B1(n16726), .B2(n16685), .A(n16684), .ZN(n17610) );
  NAND2_X1 U19888 ( .A1(n16697), .A2(n16699), .ZN(n16695) );
  NAND2_X1 U19889 ( .A1(n9959), .A2(n16974), .ZN(n17036) );
  INV_X1 U19890 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16738) );
  NAND2_X1 U19891 ( .A1(n16739), .A2(n16738), .ZN(n16737) );
  NOR2_X1 U19892 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16737), .ZN(n16720) );
  INV_X1 U19893 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17092) );
  NAND2_X1 U19894 ( .A1(n16720), .A2(n17092), .ZN(n16696) );
  NOR2_X1 U19895 ( .A1(n17049), .A2(n16696), .ZN(n16705) );
  INV_X1 U19896 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17061) );
  INV_X1 U19897 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18875) );
  NOR2_X1 U19898 ( .A1(n18867), .A2(n16686), .ZN(n16730) );
  NAND4_X1 U19899 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(P3_REIP_REG_28__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16730), .ZN(n16691) );
  NOR3_X1 U19900 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18875), .A3(n16691), 
        .ZN(n16690) );
  INV_X1 U19901 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n16687) );
  OAI22_X1 U19902 ( .A1(n16688), .A2(n17035), .B1(n16687), .B2(n17050), .ZN(
        n16689) );
  AOI211_X1 U19903 ( .C1(n16705), .C2(n17061), .A(n16690), .B(n16689), .ZN(
        n16694) );
  NOR2_X1 U19904 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16691), .ZN(n16703) );
  NAND3_X1 U19905 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(P3_REIP_REG_28__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16692) );
  NAND2_X1 U19906 ( .A1(n17041), .A2(n17053), .ZN(n17051) );
  AOI21_X1 U19907 ( .B1(n16692), .B2(n17051), .A(n16736), .ZN(n16701) );
  INV_X1 U19908 ( .A(n16701), .ZN(n16716) );
  OAI21_X1 U19909 ( .B1(n16703), .B2(n16716), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n16693) );
  OAI211_X1 U19910 ( .C1(n16695), .C2(n17036), .A(n16694), .B(n16693), .ZN(
        P3_U2640) );
  NAND2_X1 U19911 ( .A1(n17015), .A2(n16696), .ZN(n16709) );
  INV_X1 U19912 ( .A(n16697), .ZN(n16698) );
  XNOR2_X1 U19913 ( .A(n16699), .B(n16698), .ZN(n16704) );
  OAI22_X1 U19914 ( .A1(n16701), .A2(n18875), .B1(n16700), .B2(n17035), .ZN(
        n16702) );
  AOI211_X1 U19915 ( .C1(n16704), .C2(n16974), .A(n16703), .B(n16702), .ZN(
        n16707) );
  OAI21_X1 U19916 ( .B1(n17019), .B2(n16705), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16706) );
  OAI211_X1 U19917 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16709), .A(n16707), .B(
        n16706), .ZN(P3_U2641) );
  NAND2_X1 U19918 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16723) );
  NOR2_X1 U19919 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16723), .ZN(n16708) );
  AOI22_X1 U19920 ( .A1(n17019), .A2(P3_EBX_REG_29__SCAN_IN), .B1(n16730), 
        .B2(n16708), .ZN(n16718) );
  INV_X1 U19921 ( .A(n16720), .ZN(n16710) );
  AOI21_X1 U19922 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16710), .A(n16709), .ZN(
        n16715) );
  AOI211_X1 U19923 ( .C1(n16713), .C2(n16712), .A(n16711), .B(n18799), .ZN(
        n16714) );
  OAI211_X1 U19924 ( .C1(n16719), .C2(n17035), .A(n16718), .B(n16717), .ZN(
        P3_U2642) );
  AOI211_X1 U19925 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16737), .A(n16720), .B(
        n17049), .ZN(n16729) );
  AOI211_X1 U19926 ( .C1(n17610), .C2(n16722), .A(n16721), .B(n18799), .ZN(
        n16728) );
  AOI22_X1 U19927 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n16736), .B1(n17019), 
        .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16725) );
  OAI211_X1 U19928 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16730), .B(n16723), .ZN(n16724) );
  OAI211_X1 U19929 ( .C1(n17035), .C2(n16726), .A(n16725), .B(n16724), .ZN(
        n16727) );
  OR3_X1 U19930 ( .A1(n16729), .A2(n16728), .A3(n16727), .ZN(P3_U2643) );
  INV_X1 U19931 ( .A(n16730), .ZN(n16742) );
  AOI211_X1 U19932 ( .C1(n16733), .C2(n16732), .A(n16731), .B(n18799), .ZN(
        n16735) );
  OAI22_X1 U19933 ( .A1(n17607), .A2(n17035), .B1(n17050), .B2(n16738), .ZN(
        n16734) );
  AOI211_X1 U19934 ( .C1(n16736), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16735), 
        .B(n16734), .ZN(n16741) );
  OAI211_X1 U19935 ( .C1(n16739), .C2(n16738), .A(n17015), .B(n16737), .ZN(
        n16740) );
  OAI211_X1 U19936 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n16742), .A(n16741), 
        .B(n16740), .ZN(P3_U2644) );
  AOI21_X1 U19937 ( .B1(n17015), .B2(n16743), .A(n17019), .ZN(n16753) );
  NOR2_X1 U19938 ( .A1(n16743), .A2(n17049), .ZN(n16757) );
  AOI211_X1 U19939 ( .C1(n17648), .C2(n16745), .A(n16744), .B(n18799), .ZN(
        n16750) );
  NAND2_X1 U19940 ( .A1(n17031), .A2(n18865), .ZN(n16746) );
  OAI22_X1 U19941 ( .A1(n16748), .A2(n17035), .B1(n16747), .B2(n16746), .ZN(
        n16749) );
  AOI211_X1 U19942 ( .C1(n16757), .C2(n16754), .A(n16750), .B(n16749), .ZN(
        n16752) );
  NOR2_X1 U19943 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17041), .ZN(n16762) );
  OAI21_X1 U19944 ( .B1(n16761), .B2(n17041), .A(n17053), .ZN(n16771) );
  OAI21_X1 U19945 ( .B1(n16762), .B2(n16771), .A(P3_REIP_REG_25__SCAN_IN), 
        .ZN(n16751) );
  OAI211_X1 U19946 ( .C1(n16754), .C2(n16753), .A(n16752), .B(n16751), .ZN(
        P3_U2646) );
  INV_X1 U19947 ( .A(n16771), .ZN(n16765) );
  INV_X1 U19948 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18862) );
  AOI22_X1 U19949 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16992), .B1(
        n17019), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n16764) );
  AOI211_X1 U19950 ( .C1(n17660), .C2(n16756), .A(n16755), .B(n18799), .ZN(
        n16760) );
  INV_X1 U19951 ( .A(n16757), .ZN(n16758) );
  AOI21_X1 U19952 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16772), .A(n16758), .ZN(
        n16759) );
  AOI211_X1 U19953 ( .C1(n16762), .C2(n16761), .A(n16760), .B(n16759), .ZN(
        n16763) );
  OAI211_X1 U19954 ( .C1(n16765), .C2(n18862), .A(n16764), .B(n16763), .ZN(
        P3_U2647) );
  NAND2_X1 U19955 ( .A1(n17031), .A2(n18860), .ZN(n16776) );
  AOI211_X1 U19956 ( .C1(n17677), .C2(n16767), .A(n16766), .B(n18799), .ZN(
        n16770) );
  OAI22_X1 U19957 ( .A1(n16768), .A2(n17035), .B1(n17050), .B2(n16773), .ZN(
        n16769) );
  AOI211_X1 U19958 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n16771), .A(n16770), 
        .B(n16769), .ZN(n16775) );
  OAI211_X1 U19959 ( .C1(n16782), .C2(n16773), .A(n17015), .B(n16772), .ZN(
        n16774) );
  OAI211_X1 U19960 ( .C1(n16777), .C2(n16776), .A(n16775), .B(n16774), .ZN(
        P3_U2648) );
  NAND2_X1 U19961 ( .A1(n17031), .A2(n16785), .ZN(n16867) );
  NOR2_X1 U19962 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16867), .ZN(n16778) );
  AOI22_X1 U19963 ( .A1(n17019), .A2(P3_EBX_REG_22__SCAN_IN), .B1(n16779), 
        .B2(n16778), .ZN(n16789) );
  AOI211_X1 U19964 ( .C1(n17693), .C2(n16781), .A(n16780), .B(n18799), .ZN(
        n16784) );
  AOI211_X1 U19965 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16797), .A(n16782), .B(
        n17049), .ZN(n16783) );
  AOI211_X1 U19966 ( .C1(n16992), .C2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16784), .B(n16783), .ZN(n16788) );
  NAND2_X1 U19967 ( .A1(n17053), .A2(n16785), .ZN(n16869) );
  OAI21_X1 U19968 ( .B1(n16786), .B2(n16869), .A(n17051), .ZN(n16809) );
  INV_X1 U19969 ( .A(n16809), .ZN(n16796) );
  NOR3_X1 U19970 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16786), .A3(n16867), 
        .ZN(n16792) );
  OAI21_X1 U19971 ( .B1(n16796), .B2(n16792), .A(P3_REIP_REG_22__SCAN_IN), 
        .ZN(n16787) );
  NAND3_X1 U19972 ( .A1(n16789), .A2(n16788), .A3(n16787), .ZN(P3_U2649) );
  AOI211_X1 U19973 ( .C1(n17712), .C2(n16791), .A(n16790), .B(n18799), .ZN(
        n16795) );
  INV_X1 U19974 ( .A(n16792), .ZN(n16793) );
  OAI21_X1 U19975 ( .B1(n17141), .B2(n17050), .A(n16793), .ZN(n16794) );
  AOI211_X1 U19976 ( .C1(n16796), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16795), 
        .B(n16794), .ZN(n16799) );
  OAI211_X1 U19977 ( .C1(n16804), .C2(n17141), .A(n17015), .B(n16797), .ZN(
        n16798) );
  OAI211_X1 U19978 ( .C1(n17035), .C2(n17704), .A(n16799), .B(n16798), .ZN(
        P3_U2650) );
  INV_X1 U19979 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18856) );
  NOR2_X1 U19980 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16867), .ZN(n16800) );
  AOI22_X1 U19981 ( .A1(n17019), .A2(P3_EBX_REG_20__SCAN_IN), .B1(n16801), 
        .B2(n16800), .ZN(n16808) );
  AOI211_X1 U19982 ( .C1(n17721), .C2(n16803), .A(n16802), .B(n18799), .ZN(
        n16806) );
  AOI211_X1 U19983 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16820), .A(n16804), .B(
        n17049), .ZN(n16805) );
  AOI211_X1 U19984 ( .C1(n16992), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16806), .B(n16805), .ZN(n16807) );
  OAI211_X1 U19985 ( .C1(n18856), .C2(n16809), .A(n16808), .B(n16807), .ZN(
        P3_U2651) );
  INV_X1 U19986 ( .A(n16811), .ZN(n16810) );
  OAI21_X1 U19987 ( .B1(n16810), .B2(n16869), .A(n17051), .ZN(n16846) );
  INV_X1 U19988 ( .A(n16867), .ZN(n16847) );
  INV_X1 U19989 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18854) );
  NAND3_X1 U19990 ( .A1(n16811), .A2(n16847), .A3(n18854), .ZN(n16832) );
  AOI21_X1 U19991 ( .B1(n16846), .B2(n16832), .A(n20997), .ZN(n16819) );
  NOR3_X1 U19992 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16812), .A3(n16867), 
        .ZN(n16818) );
  AOI211_X1 U19993 ( .C1(n17729), .C2(n16814), .A(n16813), .B(n18799), .ZN(
        n16817) );
  INV_X1 U19994 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16815) );
  OAI21_X1 U19995 ( .B1(n16815), .B2(n17035), .A(n18280), .ZN(n16816) );
  NOR4_X1 U19996 ( .A1(n16819), .A2(n16818), .A3(n16817), .A4(n16816), .ZN(
        n16822) );
  OAI211_X1 U19997 ( .C1(n16824), .C2(n16823), .A(n17015), .B(n16820), .ZN(
        n16821) );
  OAI211_X1 U19998 ( .C1(n16823), .C2(n17050), .A(n16822), .B(n16821), .ZN(
        P3_U2652) );
  AOI211_X1 U19999 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16839), .A(n16824), .B(
        n17049), .ZN(n16831) );
  INV_X1 U20000 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17181) );
  OAI21_X1 U20001 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17728), .A(
        n16825), .ZN(n17739) );
  INV_X1 U20002 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17037) );
  NAND2_X1 U20003 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17037), .ZN(
        n17023) );
  OAI21_X1 U20004 ( .B1(n16826), .B2(n17023), .A(n9959), .ZN(n16828) );
  AOI21_X1 U20005 ( .B1(n17739), .B2(n16828), .A(n18799), .ZN(n16827) );
  OAI21_X1 U20006 ( .B1(n17739), .B2(n16828), .A(n16827), .ZN(n16829) );
  OAI211_X1 U20007 ( .C1(n17050), .C2(n17181), .A(n18280), .B(n16829), .ZN(
        n16830) );
  AOI211_X1 U20008 ( .C1(n16992), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16831), .B(n16830), .ZN(n16833) );
  OAI211_X1 U20009 ( .C1(n16846), .C2(n18854), .A(n16833), .B(n16832), .ZN(
        P3_U2653) );
  INV_X1 U20010 ( .A(n16858), .ZN(n16834) );
  OAI21_X1 U20011 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16834), .A(
        n16835), .ZN(n17767) );
  AOI21_X1 U20012 ( .B1(n16857), .B2(n17767), .A(n16933), .ZN(n16836) );
  AOI21_X1 U20013 ( .B1(n9958), .B2(n16835), .A(n17728), .ZN(n17755) );
  XOR2_X1 U20014 ( .A(n16836), .B(n17755), .Z(n16844) );
  NOR3_X1 U20015 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16837), .A3(n16867), 
        .ZN(n16838) );
  AOI211_X1 U20016 ( .C1(n17019), .C2(P3_EBX_REG_17__SCAN_IN), .A(n18125), .B(
        n16838), .ZN(n16842) );
  OAI211_X1 U20017 ( .C1(n16848), .C2(n16840), .A(n17015), .B(n16839), .ZN(
        n16841) );
  OAI211_X1 U20018 ( .C1(n17035), .C2(n9958), .A(n16842), .B(n16841), .ZN(
        n16843) );
  AOI21_X1 U20019 ( .B1(n16844), .B2(n16974), .A(n16843), .ZN(n16845) );
  OAI21_X1 U20020 ( .B1(n18852), .B2(n16846), .A(n16845), .ZN(P3_U2654) );
  NAND2_X1 U20021 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16847), .ZN(n16856) );
  INV_X1 U20022 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18850) );
  INV_X1 U20023 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18848) );
  OAI21_X1 U20024 ( .B1(n18848), .B2(n16869), .A(n17051), .ZN(n16868) );
  AOI211_X1 U20025 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16861), .A(n16848), .B(
        n17049), .ZN(n16854) );
  INV_X1 U20026 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16852) );
  OR2_X1 U20027 ( .A1(n16933), .A2(n16857), .ZN(n16850) );
  OAI21_X1 U20028 ( .B1(n16857), .B2(n16933), .A(n17767), .ZN(n16849) );
  OAI211_X1 U20029 ( .C1(n17767), .C2(n16850), .A(n16974), .B(n16849), .ZN(
        n16851) );
  OAI211_X1 U20030 ( .C1(n16852), .C2(n17035), .A(n18280), .B(n16851), .ZN(
        n16853) );
  AOI211_X1 U20031 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17019), .A(n16854), .B(
        n16853), .ZN(n16855) );
  OAI221_X1 U20032 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n16856), .C1(n18850), 
        .C2(n16868), .A(n16855), .ZN(P3_U2655) );
  INV_X1 U20033 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17775) );
  NOR2_X1 U20034 ( .A1(n16857), .A2(n17036), .ZN(n16860) );
  OAI21_X1 U20035 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17764), .A(
        n16858), .ZN(n17787) );
  OAI21_X1 U20036 ( .B1(n16933), .B2(n17037), .A(n16974), .ZN(n17048) );
  AOI211_X1 U20037 ( .C1(n9959), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n17048), .B(n17787), .ZN(n16859) );
  AOI211_X1 U20038 ( .C1(n16860), .C2(n17787), .A(n18198), .B(n16859), .ZN(
        n16864) );
  OAI211_X1 U20039 ( .C1(n16871), .C2(n16862), .A(n17015), .B(n16861), .ZN(
        n16863) );
  OAI211_X1 U20040 ( .C1(n17035), .C2(n17775), .A(n16864), .B(n16863), .ZN(
        n16865) );
  AOI21_X1 U20041 ( .B1(n17019), .B2(P3_EBX_REG_15__SCAN_IN), .A(n16865), .ZN(
        n16866) );
  OAI221_X1 U20042 ( .B1(n16868), .B2(n18848), .C1(n16868), .C2(n16867), .A(
        n16866), .ZN(P3_U2656) );
  INV_X1 U20043 ( .A(n16869), .ZN(n16880) );
  NOR2_X1 U20044 ( .A1(n17041), .A2(n16870), .ZN(n16886) );
  AOI22_X1 U20045 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n17051), .B1(
        P3_REIP_REG_13__SCAN_IN), .B2(n16886), .ZN(n16879) );
  AOI211_X1 U20046 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16889), .A(n16871), .B(
        n17049), .ZN(n16877) );
  INV_X1 U20047 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16875) );
  INV_X1 U20048 ( .A(n17829), .ZN(n16898) );
  NOR2_X1 U20049 ( .A1(n17961), .A2(n17901), .ZN(n16981) );
  NAND2_X1 U20050 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16981), .ZN(
        n16970) );
  NOR2_X1 U20051 ( .A1(n16898), .A2(n16970), .ZN(n17800) );
  INV_X1 U20052 ( .A(n17800), .ZN(n16897) );
  OR2_X1 U20053 ( .A1(n17803), .A2(n16897), .ZN(n16882) );
  AOI21_X1 U20054 ( .B1(n16875), .B2(n16882), .A(n17764), .ZN(n17793) );
  OR2_X1 U20055 ( .A1(n16970), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16958) );
  NOR3_X1 U20056 ( .A1(n16898), .A2(n17803), .A3(n16958), .ZN(n16881) );
  NOR2_X1 U20057 ( .A1(n16933), .A2(n16881), .ZN(n16873) );
  AOI21_X1 U20058 ( .B1(n17793), .B2(n16873), .A(n18799), .ZN(n16872) );
  OAI21_X1 U20059 ( .B1(n17793), .B2(n16873), .A(n16872), .ZN(n16874) );
  OAI211_X1 U20060 ( .C1(n16875), .C2(n17035), .A(n16874), .B(n18280), .ZN(
        n16876) );
  AOI211_X1 U20061 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17019), .A(n16877), .B(
        n16876), .ZN(n16878) );
  OAI21_X1 U20062 ( .B1(n16880), .B2(n16879), .A(n16878), .ZN(P3_U2657) );
  AOI22_X1 U20063 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n16992), .B1(
        n17019), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n16894) );
  NOR2_X1 U20064 ( .A1(n16881), .A2(n17036), .ZN(n16885) );
  INV_X1 U20065 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17820) );
  NOR2_X1 U20066 ( .A1(n17820), .A2(n16897), .ZN(n16883) );
  OAI21_X1 U20067 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16883), .A(
        n16882), .ZN(n17806) );
  AOI211_X1 U20068 ( .C1(n9959), .C2(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n17048), .B(n17806), .ZN(n16884) );
  AOI211_X1 U20069 ( .C1(n16885), .C2(n17806), .A(n18125), .B(n16884), .ZN(
        n16893) );
  INV_X1 U20070 ( .A(n16886), .ZN(n16888) );
  OAI21_X1 U20071 ( .B1(n16902), .B2(n17041), .A(n17053), .ZN(n16909) );
  NOR2_X1 U20072 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17041), .ZN(n16901) );
  NOR2_X1 U20073 ( .A1(n16909), .A2(n16901), .ZN(n16887) );
  MUX2_X1 U20074 ( .A(n16888), .B(n16887), .S(P3_REIP_REG_13__SCAN_IN), .Z(
        n16892) );
  OAI211_X1 U20075 ( .C1(n16895), .C2(n16890), .A(n17015), .B(n16889), .ZN(
        n16891) );
  NAND4_X1 U20076 ( .A1(n16894), .A2(n16893), .A3(n16892), .A4(n16891), .ZN(
        P3_U2658) );
  AOI211_X1 U20077 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16914), .A(n16895), .B(
        n17049), .ZN(n16896) );
  AOI21_X1 U20078 ( .B1(n16992), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16896), .ZN(n16905) );
  AOI22_X1 U20079 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16897), .B1(
        n17800), .B2(n17820), .ZN(n17816) );
  OAI21_X1 U20080 ( .B1(n16898), .B2(n16958), .A(n9959), .ZN(n16899) );
  XOR2_X1 U20081 ( .A(n17816), .B(n16899), .Z(n16900) );
  AOI22_X1 U20082 ( .A1(n17019), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n16974), 
        .B2(n16900), .ZN(n16904) );
  AOI22_X1 U20083 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16909), .B1(n16902), 
        .B2(n16901), .ZN(n16903) );
  NAND4_X1 U20084 ( .A1(n16905), .A2(n16904), .A3(n16903), .A4(n18280), .ZN(
        P3_U2659) );
  NAND2_X1 U20085 ( .A1(n17871), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17870) );
  NOR2_X1 U20086 ( .A1(n17961), .A2(n17870), .ZN(n16957) );
  NAND2_X1 U20087 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16957), .ZN(
        n16944) );
  INV_X1 U20088 ( .A(n16944), .ZN(n16932) );
  NAND2_X1 U20089 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16932), .ZN(
        n16931) );
  INV_X1 U20090 ( .A(n16931), .ZN(n16919) );
  NAND2_X1 U20091 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16919), .ZN(
        n16918) );
  AOI21_X1 U20092 ( .B1(n16917), .B2(n16918), .A(n17800), .ZN(n17832) );
  OAI21_X1 U20093 ( .B1(n16906), .B2(n16958), .A(n9959), .ZN(n16907) );
  XNOR2_X1 U20094 ( .A(n17832), .B(n16907), .ZN(n16913) );
  NOR2_X1 U20095 ( .A1(n17041), .A2(n16921), .ZN(n16925) );
  AOI21_X1 U20096 ( .B1(n16908), .B2(n16925), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16911) );
  INV_X1 U20097 ( .A(n16909), .ZN(n16910) );
  OAI22_X1 U20098 ( .A1(n16911), .A2(n16910), .B1(n17050), .B2(n20906), .ZN(
        n16912) );
  AOI211_X1 U20099 ( .C1(n16974), .C2(n16913), .A(n18125), .B(n16912), .ZN(
        n16916) );
  OAI211_X1 U20100 ( .C1(n16922), .C2(n20906), .A(n17015), .B(n16914), .ZN(
        n16915) );
  OAI211_X1 U20101 ( .C1(n17035), .C2(n16917), .A(n16916), .B(n16915), .ZN(
        P3_U2660) );
  OAI21_X1 U20102 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16919), .A(
        n16918), .ZN(n17845) );
  OAI21_X1 U20103 ( .B1(n17827), .B2(n16958), .A(n9959), .ZN(n16934) );
  XOR2_X1 U20104 ( .A(n17845), .B(n16934), .Z(n16920) );
  AOI22_X1 U20105 ( .A1(n17019), .A2(P3_EBX_REG_10__SCAN_IN), .B1(n16974), 
        .B2(n16920), .ZN(n16928) );
  AOI21_X1 U20106 ( .B1(n17031), .B2(n16921), .A(n17045), .ZN(n16947) );
  NAND2_X1 U20107 ( .A1(n16925), .A2(n18836), .ZN(n16940) );
  AOI21_X1 U20108 ( .B1(n16947), .B2(n16940), .A(n18838), .ZN(n16924) );
  AOI211_X1 U20109 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16929), .A(n16922), .B(
        n17049), .ZN(n16923) );
  AOI211_X1 U20110 ( .C1(n16992), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16924), .B(n16923), .ZN(n16927) );
  NAND3_X1 U20111 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16925), .A3(n18838), 
        .ZN(n16926) );
  NAND4_X1 U20112 ( .A1(n16928), .A2(n16927), .A3(n18280), .A4(n16926), .ZN(
        P3_U2661) );
  OAI211_X1 U20113 ( .C1(n16942), .C2(n16930), .A(n17015), .B(n16929), .ZN(
        n16938) );
  OAI21_X1 U20114 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16932), .A(
        n16931), .ZN(n17856) );
  OAI221_X1 U20115 ( .B1(n17856), .B2(n16932), .C1(n17856), .C2(n17037), .A(
        n16974), .ZN(n16935) );
  NAND2_X1 U20116 ( .A1(n16974), .A2(n16933), .ZN(n17025) );
  AOI22_X1 U20117 ( .A1(n16935), .A2(n17025), .B1(n17856), .B2(n16934), .ZN(
        n16936) );
  AOI211_X1 U20118 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n16992), .A(
        n18125), .B(n16936), .ZN(n16937) );
  NAND2_X1 U20119 ( .A1(n16938), .A2(n16937), .ZN(n16939) );
  AOI21_X1 U20120 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17019), .A(n16939), .ZN(
        n16941) );
  OAI211_X1 U20121 ( .C1(n16947), .C2(n18836), .A(n16941), .B(n16940), .ZN(
        P3_U2662) );
  AOI211_X1 U20122 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16964), .A(n16942), .B(
        n17049), .ZN(n16943) );
  AOI21_X1 U20123 ( .B1(n16992), .B2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16943), .ZN(n16954) );
  OAI21_X1 U20124 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16957), .A(
        n16944), .ZN(n17875) );
  OAI21_X1 U20125 ( .B1(n17886), .B2(n16958), .A(n9959), .ZN(n16945) );
  XOR2_X1 U20126 ( .A(n17875), .B(n16945), .Z(n16946) );
  AOI22_X1 U20127 ( .A1(n17019), .A2(P3_EBX_REG_8__SCAN_IN), .B1(n16974), .B2(
        n16946), .ZN(n16953) );
  INV_X1 U20128 ( .A(n16947), .ZN(n16951) );
  NOR2_X1 U20129 ( .A1(n16948), .A2(n17041), .ZN(n16949) );
  AOI22_X1 U20130 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16951), .B1(n16950), 
        .B2(n16949), .ZN(n16952) );
  NAND4_X1 U20131 ( .A1(n16954), .A2(n16953), .A3(n16952), .A4(n18280), .ZN(
        P3_U2663) );
  NAND2_X1 U20132 ( .A1(n17031), .A2(n18832), .ZN(n16968) );
  INV_X1 U20133 ( .A(n16956), .ZN(n16955) );
  AOI21_X1 U20134 ( .B1(n17031), .B2(n16955), .A(n17045), .ZN(n16984) );
  INV_X1 U20135 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20920) );
  NAND3_X1 U20136 ( .A1(n17031), .A2(n16956), .A3(n20920), .ZN(n16972) );
  AOI21_X1 U20137 ( .B1(n16984), .B2(n16972), .A(n18832), .ZN(n16963) );
  AOI21_X1 U20138 ( .B1(n17886), .B2(n16970), .A(n16957), .ZN(n16960) );
  NAND2_X1 U20139 ( .A1(n16958), .A2(n9959), .ZN(n16959) );
  INV_X1 U20140 ( .A(n16959), .ZN(n16973) );
  INV_X1 U20141 ( .A(n16960), .ZN(n17892) );
  AOI221_X1 U20142 ( .B1(n16960), .B2(n16973), .C1(n17892), .C2(n16959), .A(
        n18799), .ZN(n16962) );
  OAI22_X1 U20143 ( .A1(n17886), .A2(n17035), .B1(n17050), .B2(n17310), .ZN(
        n16961) );
  NOR4_X1 U20144 ( .A1(n18125), .A2(n16963), .A3(n16962), .A4(n16961), .ZN(
        n16966) );
  OAI211_X1 U20145 ( .C1(n16969), .C2(n17310), .A(n17015), .B(n16964), .ZN(
        n16965) );
  OAI211_X1 U20146 ( .C1(n16968), .C2(n16967), .A(n16966), .B(n16965), .ZN(
        P3_U2664) );
  AOI211_X1 U20147 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16988), .A(n16969), .B(
        n17049), .ZN(n16979) );
  INV_X1 U20148 ( .A(n16981), .ZN(n16971) );
  OAI21_X1 U20149 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16981), .A(
        n16970), .ZN(n17902) );
  AOI211_X1 U20150 ( .C1(n9959), .C2(n16971), .A(n17048), .B(n17902), .ZN(
        n16978) );
  OAI21_X1 U20151 ( .B1(n17035), .B2(n17905), .A(n16972), .ZN(n16977) );
  NAND3_X1 U20152 ( .A1(n16974), .A2(n16973), .A3(n17902), .ZN(n16975) );
  OAI211_X1 U20153 ( .C1(n17050), .C2(n17311), .A(n18280), .B(n16975), .ZN(
        n16976) );
  NOR4_X1 U20154 ( .A1(n16979), .A2(n16978), .A3(n16977), .A4(n16976), .ZN(
        n16980) );
  OAI21_X1 U20155 ( .B1(n16984), .B2(n20920), .A(n16980), .ZN(P3_U2665) );
  NAND2_X1 U20156 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17911), .ZN(
        n16995) );
  OAI21_X1 U20157 ( .B1(n16995), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n9959), .ZN(n16994) );
  INV_X1 U20158 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16982) );
  AOI21_X1 U20159 ( .B1(n16982), .B2(n16995), .A(n16981), .ZN(n17917) );
  XOR2_X1 U20160 ( .A(n16994), .B(n17917), .Z(n16983) );
  OAI21_X1 U20161 ( .B1(n16983), .B2(n18799), .A(n18280), .ZN(n16987) );
  AOI221_X1 U20162 ( .B1(n17041), .B2(n18829), .C1(n16985), .C2(n18829), .A(
        n16984), .ZN(n16986) );
  AOI211_X1 U20163 ( .C1(n16992), .C2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n16987), .B(n16986), .ZN(n16990) );
  OAI211_X1 U20164 ( .C1(n16993), .C2(n17307), .A(n17015), .B(n16988), .ZN(
        n16989) );
  OAI211_X1 U20165 ( .C1(n17307), .C2(n17050), .A(n16990), .B(n16989), .ZN(
        P3_U2666) );
  NOR2_X1 U20166 ( .A1(n17002), .A2(n17041), .ZN(n17009) );
  NOR2_X1 U20167 ( .A1(n17045), .A2(n17009), .ZN(n17011) );
  INV_X1 U20168 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18827) );
  NAND2_X1 U20169 ( .A1(n18932), .A2(n18948), .ZN(n18951) );
  AOI21_X1 U20170 ( .B1(n17006), .B2(n18780), .A(n18951), .ZN(n16991) );
  AOI211_X1 U20171 ( .C1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n16992), .A(
        n18125), .B(n16991), .ZN(n17004) );
  NOR2_X1 U20172 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17041), .ZN(n17001) );
  AOI211_X1 U20173 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17014), .A(n16993), .B(
        n17049), .ZN(n17000) );
  INV_X1 U20174 ( .A(n16994), .ZN(n16997) );
  NOR2_X1 U20175 ( .A1(n17961), .A2(n17926), .ZN(n17005) );
  OAI21_X1 U20176 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17005), .A(
        n16995), .ZN(n17929) );
  OR2_X1 U20177 ( .A1(n17926), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17925) );
  OAI22_X1 U20178 ( .A1(n9959), .A2(n17929), .B1(n17023), .B2(n17925), .ZN(
        n16996) );
  AOI21_X1 U20179 ( .B1(n16997), .B2(n17929), .A(n16996), .ZN(n16998) );
  OAI22_X1 U20180 ( .A1(n16998), .A2(n18799), .B1(n17050), .B2(n20981), .ZN(
        n16999) );
  AOI211_X1 U20181 ( .C1(n17002), .C2(n17001), .A(n17000), .B(n16999), .ZN(
        n17003) );
  OAI211_X1 U20182 ( .C1(n17011), .C2(n18827), .A(n17004), .B(n17003), .ZN(
        P3_U2667) );
  INV_X1 U20183 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17018) );
  NAND2_X1 U20184 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17021) );
  AOI21_X1 U20185 ( .B1(n17018), .B2(n17021), .A(n17005), .ZN(n17943) );
  INV_X1 U20186 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17955) );
  OAI21_X1 U20187 ( .B1(n17955), .B2(n17023), .A(n9959), .ZN(n17022) );
  XOR2_X1 U20188 ( .A(n17943), .B(n17022), .Z(n17008) );
  NOR2_X1 U20189 ( .A1(n18914), .A2(n18736), .ZN(n17007) );
  OAI21_X1 U20190 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n17007), .A(
        n17006), .ZN(n18888) );
  OAI22_X1 U20191 ( .A1(n18799), .A2(n17008), .B1(n18951), .B2(n18888), .ZN(
        n17013) );
  INV_X1 U20192 ( .A(n17009), .ZN(n17010) );
  OAI22_X1 U20193 ( .A1(n17011), .A2(n18825), .B1(n17030), .B2(n17010), .ZN(
        n17012) );
  AOI211_X1 U20194 ( .C1(n17019), .C2(P3_EBX_REG_3__SCAN_IN), .A(n17013), .B(
        n17012), .ZN(n17017) );
  OAI211_X1 U20195 ( .C1(n17020), .C2(n17319), .A(n17015), .B(n17014), .ZN(
        n17016) );
  OAI211_X1 U20196 ( .C1(n17035), .C2(n17018), .A(n17017), .B(n17016), .ZN(
        P3_U2668) );
  AOI22_X1 U20197 ( .A1(n17019), .A2(P3_EBX_REG_2__SCAN_IN), .B1(
        P3_REIP_REG_2__SCAN_IN), .B2(n17045), .ZN(n17034) );
  NOR2_X1 U20198 ( .A1(n17955), .A2(n17035), .ZN(n17029) );
  OR2_X1 U20199 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), .ZN(
        n17038) );
  AOI211_X1 U20200 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17038), .A(n17020), .B(
        n17049), .ZN(n17028) );
  OAI21_X1 U20201 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17021), .ZN(n17951) );
  INV_X1 U20202 ( .A(n17951), .ZN(n17024) );
  AOI211_X1 U20203 ( .C1(n17024), .C2(n17023), .A(n18799), .B(n17022), .ZN(
        n17027) );
  NAND2_X1 U20204 ( .A1(n17040), .A2(n18900), .ZN(n18740) );
  OAI21_X1 U20205 ( .B1(n18736), .B2(n18914), .A(n18740), .ZN(n18894) );
  OAI22_X1 U20206 ( .A1(n18894), .A2(n18951), .B1(n17951), .B2(n17025), .ZN(
        n17026) );
  NOR4_X1 U20207 ( .A1(n17029), .A2(n17028), .A3(n17027), .A4(n17026), .ZN(
        n17033) );
  OAI211_X1 U20208 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17031), .B(n17030), .ZN(n17032) );
  NAND3_X1 U20209 ( .A1(n17034), .A2(n17033), .A3(n17032), .ZN(P3_U2669) );
  OAI21_X1 U20210 ( .B1(n17037), .B2(n17036), .A(n17035), .ZN(n17044) );
  NAND2_X1 U20211 ( .A1(n17038), .A2(n17327), .ZN(n17336) );
  NAND2_X1 U20212 ( .A1(n17040), .A2(n17039), .ZN(n18901) );
  OAI22_X1 U20213 ( .A1(n17049), .A2(n17336), .B1(n18901), .B2(n18951), .ZN(
        n17043) );
  INV_X1 U20214 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17335) );
  OAI22_X1 U20215 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17041), .B1(n17050), 
        .B2(n17335), .ZN(n17042) );
  AOI211_X1 U20216 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n17044), .A(
        n17043), .B(n17042), .ZN(n17047) );
  NAND2_X1 U20217 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17045), .ZN(n17046) );
  OAI211_X1 U20218 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n17048), .A(
        n17047), .B(n17046), .ZN(P3_U2670) );
  NAND2_X1 U20219 ( .A1(n17050), .A2(n17049), .ZN(n17052) );
  AOI22_X1 U20220 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17052), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n17051), .ZN(n17055) );
  NAND3_X1 U20221 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18896), .A3(
        n17053), .ZN(n17054) );
  OAI211_X1 U20222 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18951), .A(
        n17055), .B(n17054), .ZN(P3_U2671) );
  NAND4_X1 U20223 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(P3_EBX_REG_25__SCAN_IN), .A4(P3_EBX_REG_24__SCAN_IN), .ZN(n17056)
         );
  NOR3_X1 U20224 ( .A1(n17141), .A2(n17154), .A3(n17056), .ZN(n17057) );
  NAND4_X1 U20225 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n17093), .A4(n17057), .ZN(n17060) );
  NOR2_X1 U20226 ( .A1(n17061), .A2(n17060), .ZN(n17087) );
  NAND2_X1 U20227 ( .A1(n17332), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17059) );
  NAND2_X1 U20228 ( .A1(n17087), .A2(n18332), .ZN(n17058) );
  OAI22_X1 U20229 ( .A1(n17087), .A2(n17059), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17058), .ZN(P3_U2672) );
  NAND2_X1 U20230 ( .A1(n17061), .A2(n17060), .ZN(n17062) );
  NAND2_X1 U20231 ( .A1(n17062), .A2(n17332), .ZN(n17086) );
  AOI22_X1 U20232 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17067) );
  AOI22_X1 U20233 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17066) );
  AOI22_X1 U20234 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17065) );
  AOI22_X1 U20235 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17064) );
  NAND4_X1 U20236 ( .A1(n17067), .A2(n17066), .A3(n17065), .A4(n17064), .ZN(
        n17073) );
  AOI22_X1 U20237 ( .A1(n17256), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17071) );
  AOI22_X1 U20238 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17070) );
  AOI22_X1 U20239 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17069) );
  AOI22_X1 U20240 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17068) );
  NAND4_X1 U20241 ( .A1(n17071), .A2(n17070), .A3(n17069), .A4(n17068), .ZN(
        n17072) );
  NOR2_X1 U20242 ( .A1(n17073), .A2(n17072), .ZN(n17085) );
  AOI22_X1 U20243 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U20244 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17220), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17083) );
  AOI22_X1 U20245 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17074) );
  OAI21_X1 U20246 ( .B1(n17075), .B2(n17312), .A(n17074), .ZN(n17081) );
  AOI22_X1 U20247 ( .A1(n15951), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17079) );
  AOI22_X1 U20248 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17078) );
  AOI22_X1 U20249 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17077) );
  AOI22_X1 U20250 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17076) );
  NAND4_X1 U20251 ( .A1(n17079), .A2(n17078), .A3(n17077), .A4(n17076), .ZN(
        n17080) );
  AOI211_X1 U20252 ( .C1(n17288), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n17081), .B(n17080), .ZN(n17082) );
  NAND3_X1 U20253 ( .A1(n17084), .A2(n17083), .A3(n17082), .ZN(n17089) );
  NAND2_X1 U20254 ( .A1(n17090), .A2(n17089), .ZN(n17088) );
  XNOR2_X1 U20255 ( .A(n17085), .B(n17088), .ZN(n17348) );
  OAI22_X1 U20256 ( .A1(n17087), .A2(n17086), .B1(n17348), .B2(n17332), .ZN(
        P3_U2673) );
  OAI21_X1 U20257 ( .B1(n17090), .B2(n17089), .A(n17088), .ZN(n17356) );
  OAI222_X1 U20258 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17103), .B1(
        P3_EBX_REG_29__SCAN_IN), .B2(n17093), .C1(n17092), .C2(n17091), .ZN(
        n17094) );
  OAI21_X1 U20259 ( .B1(n17356), .B2(n17332), .A(n17094), .ZN(P3_U2674) );
  OAI21_X1 U20260 ( .B1(n17099), .B2(n17096), .A(n17095), .ZN(n17365) );
  NAND3_X1 U20261 ( .A1(n17098), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17332), 
        .ZN(n17097) );
  OAI221_X1 U20262 ( .B1(n17098), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17332), 
        .C2(n17365), .A(n17097), .ZN(P3_U2676) );
  AOI21_X1 U20263 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17332), .A(n17107), .ZN(
        n17102) );
  AOI21_X1 U20264 ( .B1(n17100), .B2(n17104), .A(n17099), .ZN(n17366) );
  INV_X1 U20265 ( .A(n17366), .ZN(n17101) );
  OAI22_X1 U20266 ( .A1(n17103), .A2(n17102), .B1(n17101), .B2(n17332), .ZN(
        P3_U2677) );
  AOI21_X1 U20267 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17332), .A(n17112), .ZN(
        n17106) );
  OAI21_X1 U20268 ( .B1(n17108), .B2(n17105), .A(n17104), .ZN(n17375) );
  OAI22_X1 U20269 ( .A1(n17107), .A2(n17106), .B1(n17332), .B2(n17375), .ZN(
        P3_U2678) );
  AOI21_X1 U20270 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17332), .A(n17118), .ZN(
        n17111) );
  AOI21_X1 U20271 ( .B1(n17109), .B2(n17114), .A(n17108), .ZN(n17376) );
  INV_X1 U20272 ( .A(n17376), .ZN(n17110) );
  OAI22_X1 U20273 ( .A1(n17112), .A2(n17111), .B1(n17332), .B2(n17110), .ZN(
        P3_U2679) );
  AOI21_X1 U20274 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17332), .A(n17113), .ZN(
        n17117) );
  OAI21_X1 U20275 ( .B1(n17116), .B2(n17115), .A(n17114), .ZN(n17387) );
  OAI22_X1 U20276 ( .A1(n17118), .A2(n17117), .B1(n17332), .B2(n17387), .ZN(
        P3_U2680) );
  AOI22_X1 U20277 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17122) );
  AOI22_X1 U20278 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17121) );
  AOI22_X1 U20279 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17220), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17120) );
  AOI22_X1 U20280 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17119) );
  NAND4_X1 U20281 ( .A1(n17122), .A2(n17121), .A3(n17120), .A4(n17119), .ZN(
        n17128) );
  AOI22_X1 U20282 ( .A1(n15951), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17126) );
  AOI22_X1 U20283 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17125) );
  AOI22_X1 U20284 ( .A1(n17256), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17124) );
  AOI22_X1 U20285 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17123) );
  NAND4_X1 U20286 ( .A1(n17126), .A2(n17125), .A3(n17124), .A4(n17123), .ZN(
        n17127) );
  NOR2_X1 U20287 ( .A1(n17128), .A2(n17127), .ZN(n17391) );
  NAND3_X1 U20288 ( .A1(n17130), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17332), 
        .ZN(n17129) );
  OAI221_X1 U20289 ( .B1(n17130), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17332), 
        .C2(n17391), .A(n17129), .ZN(P3_U2681) );
  AOI22_X1 U20290 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17134) );
  AOI22_X1 U20291 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17133) );
  AOI22_X1 U20292 ( .A1(n12439), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17132) );
  AOI22_X1 U20293 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17131) );
  NAND4_X1 U20294 ( .A1(n17134), .A2(n17133), .A3(n17132), .A4(n17131), .ZN(
        n17140) );
  AOI22_X1 U20295 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17138) );
  AOI22_X1 U20296 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17137) );
  AOI22_X1 U20297 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17136) );
  AOI22_X1 U20298 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17135) );
  NAND4_X1 U20299 ( .A1(n17138), .A2(n17137), .A3(n17136), .A4(n17135), .ZN(
        n17139) );
  NOR2_X1 U20300 ( .A1(n17140), .A2(n17139), .ZN(n17397) );
  AOI22_X1 U20301 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17154), .B1(n17142), 
        .B2(n17141), .ZN(n17143) );
  AOI22_X1 U20302 ( .A1(n17338), .A2(n17397), .B1(n17143), .B2(n17332), .ZN(
        P3_U2682) );
  AOI22_X1 U20303 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17147) );
  AOI22_X1 U20304 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17146) );
  AOI22_X1 U20305 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17145) );
  AOI22_X1 U20306 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17144) );
  NAND4_X1 U20307 ( .A1(n17147), .A2(n17146), .A3(n17145), .A4(n17144), .ZN(
        n17153) );
  AOI22_X1 U20308 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17151) );
  AOI22_X1 U20309 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17150) );
  AOI22_X1 U20310 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17149) );
  AOI22_X1 U20311 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17148) );
  NAND4_X1 U20312 ( .A1(n17151), .A2(n17150), .A3(n17149), .A4(n17148), .ZN(
        n17152) );
  NOR2_X1 U20313 ( .A1(n17153), .A2(n17152), .ZN(n17402) );
  OAI21_X1 U20314 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17169), .A(n17154), .ZN(
        n17155) );
  AOI22_X1 U20315 ( .A1(n17338), .A2(n17402), .B1(n17155), .B2(n17332), .ZN(
        P3_U2683) );
  INV_X1 U20316 ( .A(n17170), .ZN(n17156) );
  OAI21_X1 U20317 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17156), .A(n17332), .ZN(
        n17168) );
  AOI22_X1 U20318 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17161) );
  AOI22_X1 U20319 ( .A1(n17190), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17160) );
  AOI22_X1 U20320 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17159) );
  AOI22_X1 U20321 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17158) );
  NAND4_X1 U20322 ( .A1(n17161), .A2(n17160), .A3(n17159), .A4(n17158), .ZN(
        n17167) );
  AOI22_X1 U20323 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17165) );
  AOI22_X1 U20324 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17164) );
  AOI22_X1 U20325 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17163) );
  AOI22_X1 U20326 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17162) );
  NAND4_X1 U20327 ( .A1(n17165), .A2(n17164), .A3(n17163), .A4(n17162), .ZN(
        n17166) );
  NOR2_X1 U20328 ( .A1(n17167), .A2(n17166), .ZN(n17406) );
  OAI22_X1 U20329 ( .A1(n17169), .A2(n17168), .B1(n17406), .B2(n17332), .ZN(
        P3_U2684) );
  NAND2_X1 U20330 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17170), .ZN(n17185) );
  AOI22_X1 U20331 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U20332 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U20333 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17171) );
  OAI21_X1 U20334 ( .B1(n9769), .B2(n17329), .A(n17171), .ZN(n17177) );
  AOI22_X1 U20335 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17175) );
  AOI22_X1 U20336 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17174) );
  AOI22_X1 U20337 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17173) );
  AOI22_X1 U20338 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17172) );
  NAND4_X1 U20339 ( .A1(n17175), .A2(n17174), .A3(n17173), .A4(n17172), .ZN(
        n17176) );
  AOI211_X1 U20340 ( .C1(n17220), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n17177), .B(n17176), .ZN(n17178) );
  NAND3_X1 U20341 ( .A1(n17180), .A2(n17179), .A3(n17178), .ZN(n17407) );
  INV_X1 U20342 ( .A(n17407), .ZN(n17184) );
  NAND3_X1 U20343 ( .A1(n17182), .A2(n17209), .A3(n17181), .ZN(n17183) );
  OAI221_X1 U20344 ( .B1(n17338), .B2(n17185), .C1(n17332), .C2(n17184), .A(
        n17183), .ZN(P3_U2685) );
  NAND2_X1 U20345 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17209), .ZN(n17208) );
  AOI22_X1 U20346 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17286), .ZN(n17189) );
  AOI22_X1 U20347 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17274), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n9726), .ZN(n17188) );
  AOI22_X1 U20348 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17187) );
  AOI22_X1 U20349 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17220), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17269), .ZN(n17186) );
  NAND4_X1 U20350 ( .A1(n17189), .A2(n17188), .A3(n17187), .A4(n17186), .ZN(
        n17196) );
  AOI22_X1 U20351 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n15949), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17254), .ZN(n17194) );
  AOI22_X1 U20352 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17190), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17193) );
  AOI22_X1 U20353 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17192) );
  AOI22_X1 U20354 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17287), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17191) );
  NAND4_X1 U20355 ( .A1(n17194), .A2(n17193), .A3(n17192), .A4(n17191), .ZN(
        n17195) );
  NOR2_X1 U20356 ( .A1(n17196), .A2(n17195), .ZN(n17416) );
  NAND3_X1 U20357 ( .A1(n17208), .A2(P3_EBX_REG_17__SCAN_IN), .A3(n17332), 
        .ZN(n17197) );
  OAI221_X1 U20358 ( .B1(n17208), .B2(P3_EBX_REG_17__SCAN_IN), .C1(n17332), 
        .C2(n17416), .A(n17197), .ZN(P3_U2686) );
  AOI22_X1 U20359 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17201) );
  AOI22_X1 U20360 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12439), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17200) );
  AOI22_X1 U20361 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17199) );
  AOI22_X1 U20362 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17198) );
  NAND4_X1 U20363 ( .A1(n17201), .A2(n17200), .A3(n17199), .A4(n17198), .ZN(
        n17207) );
  AOI22_X1 U20364 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17205) );
  AOI22_X1 U20365 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17204) );
  AOI22_X1 U20366 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17203) );
  AOI22_X1 U20367 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17202) );
  NAND4_X1 U20368 ( .A1(n17205), .A2(n17204), .A3(n17203), .A4(n17202), .ZN(
        n17206) );
  NOR2_X1 U20369 ( .A1(n17207), .A2(n17206), .ZN(n17422) );
  INV_X1 U20370 ( .A(n17208), .ZN(n17211) );
  AOI21_X1 U20371 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17332), .A(n17209), .ZN(
        n17210) );
  OAI22_X1 U20372 ( .A1(n17422), .A2(n17332), .B1(n17211), .B2(n17210), .ZN(
        P3_U2687) );
  NAND2_X1 U20373 ( .A1(n18332), .A2(n17212), .ZN(n17226) );
  AOI22_X1 U20374 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17223) );
  AOI22_X1 U20375 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U20376 ( .A1(n17287), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17213) );
  OAI21_X1 U20377 ( .B1(n9771), .B2(n17312), .A(n17213), .ZN(n17219) );
  AOI22_X1 U20378 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17217) );
  AOI22_X1 U20379 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17216) );
  AOI22_X1 U20380 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17215) );
  AOI22_X1 U20381 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17291), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17214) );
  NAND4_X1 U20382 ( .A1(n17217), .A2(n17216), .A3(n17215), .A4(n17214), .ZN(
        n17218) );
  AOI211_X1 U20383 ( .C1(n17220), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n17219), .B(n17218), .ZN(n17221) );
  NAND3_X1 U20384 ( .A1(n17223), .A2(n17222), .A3(n17221), .ZN(n17430) );
  AOI22_X1 U20385 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17224), .B1(n17338), 
        .B2(n17430), .ZN(n17225) );
  OAI21_X1 U20386 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17226), .A(n17225), .ZN(
        P3_U2689) );
  AOI22_X1 U20387 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17230) );
  AOI22_X1 U20388 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17229) );
  AOI22_X1 U20389 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U20390 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17227) );
  NAND4_X1 U20391 ( .A1(n17230), .A2(n17229), .A3(n17228), .A4(n17227), .ZN(
        n17236) );
  AOI22_X1 U20392 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17234) );
  AOI22_X1 U20393 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17233) );
  AOI22_X1 U20394 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17232) );
  AOI22_X1 U20395 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15949), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17231) );
  NAND4_X1 U20396 ( .A1(n17234), .A2(n17233), .A3(n17232), .A4(n17231), .ZN(
        n17235) );
  NOR2_X1 U20397 ( .A1(n17236), .A2(n17235), .ZN(n17438) );
  AND2_X1 U20398 ( .A1(n18332), .A2(n17237), .ZN(n17251) );
  OAI21_X1 U20399 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17251), .A(n17238), .ZN(
        n17239) );
  AOI22_X1 U20400 ( .A1(n17338), .A2(n17438), .B1(n17239), .B2(n17332), .ZN(
        P3_U2691) );
  AOI22_X1 U20401 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17243) );
  AOI22_X1 U20402 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17242) );
  AOI22_X1 U20403 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n9726), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17241) );
  AOI22_X1 U20404 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17240) );
  NAND4_X1 U20405 ( .A1(n17243), .A2(n17242), .A3(n17241), .A4(n17240), .ZN(
        n17249) );
  AOI22_X1 U20406 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U20407 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17246) );
  AOI22_X1 U20408 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17245) );
  AOI22_X1 U20409 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15949), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17244) );
  NAND4_X1 U20410 ( .A1(n17247), .A2(n17246), .A3(n17245), .A4(n17244), .ZN(
        n17248) );
  NOR2_X1 U20411 ( .A1(n17249), .A2(n17248), .ZN(n17441) );
  AND2_X1 U20412 ( .A1(n20906), .A2(n17250), .ZN(n17252) );
  AOI221_X1 U20413 ( .B1(n17441), .B2(n17338), .C1(n17252), .C2(n17332), .A(
        n17251), .ZN(P3_U2692) );
  NAND2_X1 U20414 ( .A1(n18332), .A2(n17253), .ZN(n17267) );
  NOR2_X1 U20415 ( .A1(n17338), .A2(n17253), .ZN(n17282) );
  AOI22_X1 U20416 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17265) );
  AOI22_X1 U20417 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17264) );
  AOI22_X1 U20418 ( .A1(n15951), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17255) );
  OAI21_X1 U20419 ( .B1(n9771), .B2(n17329), .A(n17255), .ZN(n17262) );
  AOI22_X1 U20420 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17260) );
  AOI22_X1 U20421 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17259) );
  AOI22_X1 U20422 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17258) );
  AOI22_X1 U20423 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17257) );
  NAND4_X1 U20424 ( .A1(n17260), .A2(n17259), .A3(n17258), .A4(n17257), .ZN(
        n17261) );
  AOI211_X1 U20425 ( .C1(n17274), .C2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        n17262), .B(n17261), .ZN(n17263) );
  NAND3_X1 U20426 ( .A1(n17265), .A2(n17264), .A3(n17263), .ZN(n17446) );
  AOI22_X1 U20427 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17282), .B1(n17338), 
        .B2(n17446), .ZN(n17266) );
  OAI21_X1 U20428 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17267), .A(n17266), .ZN(
        P3_U2693) );
  AOI22_X1 U20429 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n9726), .ZN(n17273) );
  AOI22_X1 U20430 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17292), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17254), .ZN(n17272) );
  AOI22_X1 U20431 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17256), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17271) );
  AOI22_X1 U20432 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17269), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17270) );
  NAND4_X1 U20433 ( .A1(n17273), .A2(n17272), .A3(n17271), .A4(n17270), .ZN(
        n17280) );
  AOI22_X1 U20434 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n12577), .ZN(n17278) );
  AOI22_X1 U20435 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17289), .ZN(n17277) );
  AOI22_X1 U20436 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17286), .ZN(n17276) );
  AOI22_X1 U20437 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17288), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17275) );
  NAND4_X1 U20438 ( .A1(n17278), .A2(n17277), .A3(n17276), .A4(n17275), .ZN(
        n17279) );
  NOR2_X1 U20439 ( .A1(n17280), .A2(n17279), .ZN(n17450) );
  INV_X1 U20440 ( .A(n17281), .ZN(n17306) );
  OAI21_X1 U20441 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17306), .A(n17282), .ZN(
        n17283) );
  OAI21_X1 U20442 ( .B1(n17450), .B2(n17332), .A(n17283), .ZN(P3_U2694) );
  NOR2_X1 U20443 ( .A1(n17284), .A2(n17340), .ZN(n17322) );
  AOI22_X1 U20444 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17332), .B1(n17285), .B2(
        n17322), .ZN(n17305) );
  AOI22_X1 U20445 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17303) );
  AOI22_X1 U20446 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17287), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17302) );
  AOI22_X1 U20447 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17290) );
  OAI21_X1 U20448 ( .B1(n10163), .B2(n21100), .A(n17290), .ZN(n17299) );
  AOI22_X1 U20449 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17256), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17297) );
  AOI22_X1 U20450 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17296) );
  AOI22_X1 U20451 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17295) );
  AOI22_X1 U20452 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17294) );
  NAND4_X1 U20453 ( .A1(n17297), .A2(n17296), .A3(n17295), .A4(n17294), .ZN(
        n17298) );
  AOI211_X1 U20454 ( .C1(n17300), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n17299), .B(n17298), .ZN(n17301) );
  NAND3_X1 U20455 ( .A1(n17303), .A2(n17302), .A3(n17301), .ZN(n17454) );
  INV_X1 U20456 ( .A(n17454), .ZN(n17304) );
  OAI22_X1 U20457 ( .A1(n17306), .A2(n17305), .B1(n17304), .B2(n17332), .ZN(
        P3_U2695) );
  NAND2_X1 U20458 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17316), .ZN(n17315) );
  OAI21_X1 U20459 ( .B1(n17311), .B2(n17315), .A(n17332), .ZN(n17313) );
  NOR3_X1 U20460 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17311), .A3(n17307), .ZN(
        n17308) );
  AOI22_X1 U20461 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17338), .B1(
        n17322), .B2(n17308), .ZN(n17309) );
  OAI21_X1 U20462 ( .B1(n17310), .B2(n17313), .A(n17309), .ZN(P3_U2696) );
  AND2_X1 U20463 ( .A1(n17311), .A2(n17315), .ZN(n17314) );
  OAI22_X1 U20464 ( .A1(n17314), .A2(n17313), .B1(n17312), .B2(n17332), .ZN(
        P3_U2697) );
  INV_X1 U20465 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17318) );
  OAI21_X1 U20466 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17316), .A(n17315), .ZN(
        n17317) );
  AOI22_X1 U20467 ( .A1(n17338), .A2(n17318), .B1(n17317), .B2(n17332), .ZN(
        P3_U2698) );
  NOR4_X1 U20468 ( .A1(n17319), .A2(n17323), .A3(n17327), .A4(n17340), .ZN(
        n17326) );
  AOI21_X1 U20469 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17332), .A(n17326), .ZN(
        n17321) );
  OAI22_X1 U20470 ( .A1(n17322), .A2(n17321), .B1(n17320), .B2(n17332), .ZN(
        P3_U2699) );
  NOR3_X1 U20471 ( .A1(n17323), .A2(n17327), .A3(n17340), .ZN(n17331) );
  AOI21_X1 U20472 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17332), .A(n17331), .ZN(
        n17325) );
  INV_X1 U20473 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17324) );
  OAI22_X1 U20474 ( .A1(n17326), .A2(n17325), .B1(n17324), .B2(n17332), .ZN(
        P3_U2700) );
  NOR2_X1 U20475 ( .A1(n17327), .A2(n17340), .ZN(n17328) );
  AOI21_X1 U20476 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n17332), .A(n17328), .ZN(
        n17330) );
  OAI22_X1 U20477 ( .A1(n17331), .A2(n17330), .B1(n17329), .B2(n17332), .ZN(
        P3_U2701) );
  INV_X1 U20478 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17333) );
  OAI222_X1 U20479 ( .A1(n17336), .A2(n17340), .B1(n17335), .B2(n17334), .C1(
        n17333), .C2(n17332), .ZN(P3_U2702) );
  AOI22_X1 U20480 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17338), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17337), .ZN(n17339) );
  OAI21_X1 U20481 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17340), .A(n17339), .ZN(
        P3_U2703) );
  NAND2_X1 U20482 ( .A1(n17478), .A2(n17341), .ZN(n17383) );
  INV_X1 U20483 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17501) );
  INV_X1 U20484 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17505) );
  INV_X1 U20485 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17507) );
  INV_X1 U20486 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17509) );
  INV_X1 U20487 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17514) );
  INV_X1 U20488 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17516) );
  INV_X1 U20489 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17603) );
  NAND3_X1 U20490 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_4__SCAN_IN), .ZN(n17428) );
  INV_X1 U20491 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17545) );
  INV_X1 U20492 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17574) );
  NAND4_X1 U20493 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n17429)
         );
  NAND3_X1 U20494 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_14__SCAN_IN), .ZN(n17342) );
  NAND2_X1 U20495 ( .A1(n18332), .A2(n17345), .ZN(n17377) );
  NAND2_X1 U20496 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17353), .ZN(n17352) );
  NOR2_X1 U20497 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n17352), .ZN(n17346) );
  INV_X1 U20498 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17571) );
  NOR2_X2 U20499 ( .A1(n17347), .A2(n17471), .ZN(n17418) );
  OAI22_X1 U20500 ( .A1(n17348), .A2(n17490), .B1(n19330), .B2(n17383), .ZN(
        n17349) );
  AOI21_X1 U20501 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17418), .A(n17349), .ZN(
        n17350) );
  OAI221_X1 U20502 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17352), .C1(n17571), 
        .C2(n17351), .A(n17350), .ZN(P3_U2705) );
  AOI22_X1 U20503 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17418), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17417), .ZN(n17355) );
  OAI211_X1 U20504 ( .C1(n17353), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17471), .B(
        n17352), .ZN(n17354) );
  OAI211_X1 U20505 ( .C1(n17356), .C2(n17490), .A(n17355), .B(n17354), .ZN(
        P3_U2706) );
  AOI22_X1 U20506 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17418), .B1(n17480), .B2(
        n17357), .ZN(n17360) );
  OAI211_X1 U20507 ( .C1(n9795), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17471), .B(
        n17358), .ZN(n17359) );
  OAI211_X1 U20508 ( .C1(n17383), .C2(n17361), .A(n17360), .B(n17359), .ZN(
        P3_U2707) );
  AOI22_X1 U20509 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17418), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17417), .ZN(n17364) );
  AOI211_X1 U20510 ( .C1(n17501), .C2(n17367), .A(n9795), .B(n17478), .ZN(
        n17362) );
  INV_X1 U20511 ( .A(n17362), .ZN(n17363) );
  OAI211_X1 U20512 ( .C1(n17365), .C2(n17490), .A(n17364), .B(n17363), .ZN(
        P3_U2708) );
  AOI22_X1 U20513 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17418), .B1(n17480), .B2(
        n17366), .ZN(n17369) );
  OAI211_X1 U20514 ( .C1(n17371), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17471), .B(
        n17367), .ZN(n17368) );
  OAI211_X1 U20515 ( .C1(n17383), .C2(n17370), .A(n17369), .B(n17368), .ZN(
        P3_U2709) );
  AOI22_X1 U20516 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17418), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17417), .ZN(n17374) );
  AOI211_X1 U20517 ( .C1(n17505), .C2(n17378), .A(n17371), .B(n17478), .ZN(
        n17372) );
  INV_X1 U20518 ( .A(n17372), .ZN(n17373) );
  OAI211_X1 U20519 ( .C1(n17375), .C2(n17490), .A(n17374), .B(n17373), .ZN(
        P3_U2710) );
  AOI22_X1 U20520 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17418), .B1(n17480), .B2(
        n17376), .ZN(n17381) );
  OAI21_X1 U20521 ( .B1(n17507), .B2(n17478), .A(n17377), .ZN(n17379) );
  NAND2_X1 U20522 ( .A1(n17379), .A2(n17378), .ZN(n17380) );
  OAI211_X1 U20523 ( .C1(n17383), .C2(n17382), .A(n17381), .B(n17380), .ZN(
        P3_U2711) );
  AOI22_X1 U20524 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17418), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17417), .ZN(n17386) );
  INV_X1 U20525 ( .A(n17388), .ZN(n17384) );
  OAI221_X1 U20526 ( .B1(P3_EAX_REG_23__SCAN_IN), .B2(n17384), .C1(n17509), 
        .C2(n17388), .A(n17471), .ZN(n17385) );
  OAI211_X1 U20527 ( .C1(n17387), .C2(n17490), .A(n17386), .B(n17385), .ZN(
        P3_U2712) );
  AOI22_X1 U20528 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17418), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n17417), .ZN(n17390) );
  OAI211_X1 U20529 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17393), .A(n17471), .B(
        n17388), .ZN(n17389) );
  OAI211_X1 U20530 ( .C1(n17391), .C2(n17490), .A(n17390), .B(n17389), .ZN(
        P3_U2713) );
  AOI22_X1 U20531 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17418), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17417), .ZN(n17396) );
  NOR2_X1 U20532 ( .A1(n17392), .A2(n17419), .ZN(n17413) );
  NAND2_X1 U20533 ( .A1(n9835), .A2(n17413), .ZN(n17403) );
  INV_X1 U20534 ( .A(n17403), .ZN(n17399) );
  NAND2_X1 U20535 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17399), .ZN(n17398) );
  AOI211_X1 U20536 ( .C1(n17514), .C2(n17398), .A(n17393), .B(n17478), .ZN(
        n17394) );
  INV_X1 U20537 ( .A(n17394), .ZN(n17395) );
  OAI211_X1 U20538 ( .C1(n17397), .C2(n17490), .A(n17396), .B(n17395), .ZN(
        P3_U2714) );
  AOI22_X1 U20539 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17418), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17417), .ZN(n17401) );
  OAI211_X1 U20540 ( .C1(n17399), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17471), .B(
        n17398), .ZN(n17400) );
  OAI211_X1 U20541 ( .C1(n17402), .C2(n17490), .A(n17401), .B(n17400), .ZN(
        P3_U2715) );
  AOI22_X1 U20542 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17418), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17417), .ZN(n17405) );
  AND3_X1 U20543 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .A3(n17413), .ZN(n17411) );
  OAI211_X1 U20544 ( .C1(n17411), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17471), .B(
        n17403), .ZN(n17404) );
  OAI211_X1 U20545 ( .C1(n17406), .C2(n17490), .A(n17405), .B(n17404), .ZN(
        P3_U2716) );
  AOI22_X1 U20546 ( .A1(n17413), .A2(P3_EAX_REG_17__SCAN_IN), .B1(
        P3_EAX_REG_18__SCAN_IN), .B2(n17471), .ZN(n17410) );
  AOI22_X1 U20547 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17417), .B1(n17480), .B2(
        n17407), .ZN(n17409) );
  NAND2_X1 U20548 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17418), .ZN(n17408) );
  OAI211_X1 U20549 ( .C1(n17411), .C2(n17410), .A(n17409), .B(n17408), .ZN(
        P3_U2717) );
  AOI22_X1 U20550 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17418), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17417), .ZN(n17415) );
  NAND2_X1 U20551 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17413), .ZN(n17412) );
  OAI211_X1 U20552 ( .C1(n17413), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17471), .B(
        n17412), .ZN(n17414) );
  OAI211_X1 U20553 ( .C1(n17416), .C2(n17490), .A(n17415), .B(n17414), .ZN(
        P3_U2718) );
  AOI22_X1 U20554 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17418), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17417), .ZN(n17421) );
  OAI211_X1 U20555 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17423), .A(n17471), .B(
        n17419), .ZN(n17420) );
  OAI211_X1 U20556 ( .C1(n17422), .C2(n17490), .A(n17421), .B(n17420), .ZN(
        P3_U2719) );
  AOI211_X1 U20557 ( .C1(n17603), .C2(n17431), .A(n17478), .B(n17423), .ZN(
        n17424) );
  AOI21_X1 U20558 ( .B1(n17485), .B2(BUF2_REG_15__SCAN_IN), .A(n17424), .ZN(
        n17425) );
  OAI21_X1 U20559 ( .B1(n17426), .B2(n17490), .A(n17425), .ZN(P3_U2720) );
  INV_X1 U20560 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17550) );
  NOR2_X1 U20561 ( .A1(n17550), .A2(n17427), .ZN(n17484) );
  NAND2_X1 U20562 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17484), .ZN(n17477) );
  NAND2_X1 U20563 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17476), .ZN(n17467) );
  NAND2_X1 U20564 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17463), .ZN(n17457) );
  NAND3_X1 U20565 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(n17443), .ZN(n17434) );
  AOI22_X1 U20566 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17485), .B1(n17480), .B2(
        n17430), .ZN(n17433) );
  NAND3_X1 U20567 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17471), .A3(n17431), 
        .ZN(n17432) );
  OAI211_X1 U20568 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17434), .A(n17433), .B(
        n17432), .ZN(P3_U2721) );
  INV_X1 U20569 ( .A(n17434), .ZN(n17437) );
  AOI22_X1 U20570 ( .A1(n17443), .A2(P3_EAX_REG_12__SCAN_IN), .B1(
        P3_EAX_REG_13__SCAN_IN), .B2(n17471), .ZN(n17436) );
  OAI222_X1 U20571 ( .A1(n17475), .A2(n17596), .B1(n17437), .B2(n17436), .C1(
        n17490), .C2(n17435), .ZN(P3_U2722) );
  AND2_X1 U20572 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17443), .ZN(n17440) );
  AOI21_X1 U20573 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17471), .A(n17443), .ZN(
        n17439) );
  OAI222_X1 U20574 ( .A1(n17475), .A2(n17593), .B1(n17440), .B2(n17439), .C1(
        n17490), .C2(n17438), .ZN(P3_U2723) );
  INV_X1 U20575 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17532) );
  INV_X1 U20576 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n20872) );
  NOR2_X1 U20577 ( .A1(n20872), .A2(n17457), .ZN(n17449) );
  NAND2_X1 U20578 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17449), .ZN(n17448) );
  NOR2_X1 U20579 ( .A1(n17532), .A2(n17448), .ZN(n17444) );
  AOI21_X1 U20580 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17471), .A(n17444), .ZN(
        n17442) );
  OAI222_X1 U20581 ( .A1(n17475), .A2(n17589), .B1(n17443), .B2(n17442), .C1(
        n17490), .C2(n17441), .ZN(P3_U2724) );
  AOI211_X1 U20582 ( .C1(n17532), .C2(n17448), .A(n17478), .B(n17444), .ZN(
        n17445) );
  AOI21_X1 U20583 ( .B1(n17480), .B2(n17446), .A(n17445), .ZN(n17447) );
  OAI21_X1 U20584 ( .B1(n17587), .B2(n17475), .A(n17447), .ZN(P3_U2725) );
  INV_X1 U20585 ( .A(n17448), .ZN(n17452) );
  AOI21_X1 U20586 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17471), .A(n17449), .ZN(
        n17451) );
  OAI222_X1 U20587 ( .A1(n17475), .A2(n17585), .B1(n17452), .B2(n17451), .C1(
        n17490), .C2(n17450), .ZN(P3_U2726) );
  NAND2_X1 U20588 ( .A1(n17471), .A2(n17453), .ZN(n17456) );
  AOI22_X1 U20589 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17485), .B1(n17480), .B2(
        n17454), .ZN(n17455) );
  OAI221_X1 U20590 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n17457), .C1(n20872), 
        .C2(n17456), .A(n17455), .ZN(P3_U2727) );
  INV_X1 U20591 ( .A(n17457), .ZN(n17460) );
  AOI21_X1 U20592 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17471), .A(n17463), .ZN(
        n17459) );
  OAI222_X1 U20593 ( .A1(n17475), .A2(n18329), .B1(n17460), .B2(n17459), .C1(
        n17490), .C2(n17458), .ZN(P3_U2728) );
  INV_X1 U20594 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17541) );
  NOR2_X1 U20595 ( .A1(n17541), .A2(n17467), .ZN(n17470) );
  AOI22_X1 U20596 ( .A1(n17470), .A2(P3_EAX_REG_5__SCAN_IN), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n17471), .ZN(n17462) );
  OAI222_X1 U20597 ( .A1(n18325), .A2(n17475), .B1(n17463), .B2(n17462), .C1(
        n17490), .C2(n17461), .ZN(P3_U2729) );
  AND2_X1 U20598 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17470), .ZN(n17466) );
  AOI21_X1 U20599 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17471), .A(n17470), .ZN(
        n17465) );
  OAI222_X1 U20600 ( .A1(n18321), .A2(n17475), .B1(n17466), .B2(n17465), .C1(
        n17490), .C2(n17464), .ZN(P3_U2730) );
  INV_X1 U20601 ( .A(n17467), .ZN(n17474) );
  AOI21_X1 U20602 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17471), .A(n17474), .ZN(
        n17469) );
  OAI222_X1 U20603 ( .A1(n18317), .A2(n17475), .B1(n17470), .B2(n17469), .C1(
        n17490), .C2(n17468), .ZN(P3_U2731) );
  AOI21_X1 U20604 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17471), .A(n17476), .ZN(
        n17473) );
  OAI222_X1 U20605 ( .A1(n18312), .A2(n17475), .B1(n17474), .B2(n17473), .C1(
        n17490), .C2(n17472), .ZN(P3_U2732) );
  INV_X1 U20606 ( .A(n17476), .ZN(n17482) );
  OAI21_X1 U20607 ( .B1(n17545), .B2(n17478), .A(n17477), .ZN(n17481) );
  AOI222_X1 U20608 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17485), .B1(n17482), .B2(
        n17481), .C1(n17480), .C2(n17479), .ZN(n17483) );
  INV_X1 U20609 ( .A(n17483), .ZN(P3_U2733) );
  AOI22_X1 U20610 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17485), .B1(n17484), .B2(
        n17574), .ZN(n17489) );
  OAI21_X1 U20611 ( .B1(n17487), .B2(n17486), .A(P3_EAX_REG_1__SCAN_IN), .ZN(
        n17488) );
  OAI211_X1 U20612 ( .C1(n17491), .C2(n17490), .A(n17489), .B(n17488), .ZN(
        P3_U2734) );
  NOR2_X1 U20613 ( .A1(n17526), .A2(n17493), .ZN(P3_U2736) );
  NAND2_X1 U20614 ( .A1(n20825), .A2(n17494), .ZN(n17522) );
  CLKBUF_X1 U20615 ( .A(n20824), .Z(n17547) );
  AOI22_X1 U20616 ( .A1(n17547), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17512), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17495) );
  OAI21_X1 U20617 ( .B1(n17571), .B2(n17522), .A(n17495), .ZN(P3_U2737) );
  INV_X1 U20618 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17497) );
  AOI22_X1 U20619 ( .A1(n20824), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17512), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17496) );
  OAI21_X1 U20620 ( .B1(n17497), .B2(n17522), .A(n17496), .ZN(P3_U2738) );
  INV_X1 U20621 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17499) );
  AOI22_X1 U20622 ( .A1(n20824), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17512), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17498) );
  OAI21_X1 U20623 ( .B1(n17499), .B2(n17522), .A(n17498), .ZN(P3_U2739) );
  AOI22_X1 U20624 ( .A1(n20824), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17512), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17500) );
  OAI21_X1 U20625 ( .B1(n17501), .B2(n17522), .A(n17500), .ZN(P3_U2740) );
  INV_X1 U20626 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17503) );
  AOI22_X1 U20627 ( .A1(n17547), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17512), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17502) );
  OAI21_X1 U20628 ( .B1(n17503), .B2(n17522), .A(n17502), .ZN(P3_U2741) );
  AOI22_X1 U20629 ( .A1(n17547), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17512), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17504) );
  OAI21_X1 U20630 ( .B1(n17505), .B2(n17522), .A(n17504), .ZN(P3_U2742) );
  AOI22_X1 U20631 ( .A1(n17547), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17512), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17506) );
  OAI21_X1 U20632 ( .B1(n17507), .B2(n17522), .A(n17506), .ZN(P3_U2743) );
  AOI22_X1 U20633 ( .A1(n17547), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17512), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17508) );
  OAI21_X1 U20634 ( .B1(n17509), .B2(n17522), .A(n17508), .ZN(P3_U2744) );
  INV_X1 U20635 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17511) );
  AOI22_X1 U20636 ( .A1(n17547), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17512), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17510) );
  OAI21_X1 U20637 ( .B1(n17511), .B2(n17522), .A(n17510), .ZN(P3_U2745) );
  AOI22_X1 U20638 ( .A1(n17547), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17512), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17513) );
  OAI21_X1 U20639 ( .B1(n17514), .B2(n17522), .A(n17513), .ZN(P3_U2746) );
  AOI22_X1 U20640 ( .A1(n17547), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n20823), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17515) );
  OAI21_X1 U20641 ( .B1(n17516), .B2(n17522), .A(n17515), .ZN(P3_U2747) );
  INV_X1 U20642 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n20961) );
  INV_X1 U20643 ( .A(n17522), .ZN(n17518) );
  AOI22_X1 U20644 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17518), .B1(n20824), 
        .B2(P3_UWORD_REG_3__SCAN_IN), .ZN(n17517) );
  OAI21_X1 U20645 ( .B1(n17526), .B2(n20961), .A(n17517), .ZN(P3_U2748) );
  INV_X1 U20646 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n20855) );
  AOI22_X1 U20647 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17518), .B1(n20824), 
        .B2(P3_UWORD_REG_2__SCAN_IN), .ZN(n17519) );
  OAI21_X1 U20648 ( .B1(n17526), .B2(n20855), .A(n17519), .ZN(P3_U2749) );
  INV_X1 U20649 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17557) );
  AOI22_X1 U20650 ( .A1(n17547), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n20823), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17520) );
  OAI21_X1 U20651 ( .B1(n17557), .B2(n17522), .A(n17520), .ZN(P3_U2750) );
  INV_X1 U20652 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n21031) );
  AOI22_X1 U20653 ( .A1(n17547), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n20823), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17521) );
  OAI21_X1 U20654 ( .B1(n21031), .B2(n17522), .A(n17521), .ZN(P3_U2751) );
  AOI22_X1 U20655 ( .A1(n17547), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n20823), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17523) );
  OAI21_X1 U20656 ( .B1(n17603), .B2(n17549), .A(n17523), .ZN(P3_U2752) );
  INV_X1 U20657 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17598) );
  AOI22_X1 U20658 ( .A1(n17547), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n20823), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17524) );
  OAI21_X1 U20659 ( .B1(n17598), .B2(n17549), .A(n17524), .ZN(P3_U2753) );
  INV_X1 U20660 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n20848) );
  AOI22_X1 U20661 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n20825), .B1(n20824), 
        .B2(P3_LWORD_REG_13__SCAN_IN), .ZN(n17525) );
  OAI21_X1 U20662 ( .B1(n17526), .B2(n20848), .A(n17525), .ZN(P3_U2754) );
  INV_X1 U20663 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17528) );
  AOI22_X1 U20664 ( .A1(n17547), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n20823), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17527) );
  OAI21_X1 U20665 ( .B1(n17528), .B2(n17549), .A(n17527), .ZN(P3_U2755) );
  INV_X1 U20666 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17530) );
  AOI22_X1 U20667 ( .A1(n17547), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n20823), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17529) );
  OAI21_X1 U20668 ( .B1(n17530), .B2(n17549), .A(n17529), .ZN(P3_U2756) );
  AOI22_X1 U20669 ( .A1(n17547), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n20823), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17531) );
  OAI21_X1 U20670 ( .B1(n17532), .B2(n17549), .A(n17531), .ZN(P3_U2757) );
  INV_X1 U20671 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17534) );
  AOI22_X1 U20672 ( .A1(n17547), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n20823), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17533) );
  OAI21_X1 U20673 ( .B1(n17534), .B2(n17549), .A(n17533), .ZN(P3_U2758) );
  AOI22_X1 U20674 ( .A1(n17547), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n20823), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17535) );
  OAI21_X1 U20675 ( .B1(n20872), .B2(n17549), .A(n17535), .ZN(P3_U2759) );
  INV_X1 U20676 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17537) );
  AOI22_X1 U20677 ( .A1(n17547), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n20823), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17536) );
  OAI21_X1 U20678 ( .B1(n17537), .B2(n17549), .A(n17536), .ZN(P3_U2760) );
  INV_X1 U20679 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17539) );
  AOI22_X1 U20680 ( .A1(n17547), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n20823), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17538) );
  OAI21_X1 U20681 ( .B1(n17539), .B2(n17549), .A(n17538), .ZN(P3_U2761) );
  AOI22_X1 U20682 ( .A1(n17547), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n20823), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17540) );
  OAI21_X1 U20683 ( .B1(n17541), .B2(n17549), .A(n17540), .ZN(P3_U2763) );
  INV_X1 U20684 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17543) );
  AOI22_X1 U20685 ( .A1(n17547), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n20823), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17542) );
  OAI21_X1 U20686 ( .B1(n17543), .B2(n17549), .A(n17542), .ZN(P3_U2764) );
  AOI22_X1 U20687 ( .A1(n17547), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n20823), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17544) );
  OAI21_X1 U20688 ( .B1(n17545), .B2(n17549), .A(n17544), .ZN(P3_U2765) );
  AOI22_X1 U20689 ( .A1(n17547), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n20823), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17546) );
  OAI21_X1 U20690 ( .B1(n17574), .B2(n17549), .A(n17546), .ZN(P3_U2766) );
  AOI22_X1 U20691 ( .A1(n17547), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n20823), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17548) );
  OAI21_X1 U20692 ( .B1(n17550), .B2(n17549), .A(n17548), .ZN(P3_U2767) );
  INV_X1 U20693 ( .A(n18927), .ZN(n18933) );
  NAND2_X1 U20694 ( .A1(n17553), .A2(n17554), .ZN(n17595) );
  INV_X2 U20695 ( .A(n17602), .ZN(n17590) );
  AOI22_X1 U20696 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17590), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17599), .ZN(n17555) );
  OAI21_X1 U20697 ( .B1(n18296), .B2(n17595), .A(n17555), .ZN(P3_U2768) );
  INV_X1 U20698 ( .A(n17595), .ZN(n17600) );
  AOI22_X1 U20699 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17600), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17599), .ZN(n17556) );
  OAI21_X1 U20700 ( .B1(n17557), .B2(n17602), .A(n17556), .ZN(P3_U2769) );
  AOI22_X1 U20701 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17590), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17599), .ZN(n17558) );
  OAI21_X1 U20702 ( .B1(n18308), .B2(n17595), .A(n17558), .ZN(P3_U2770) );
  AOI22_X1 U20703 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17590), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17599), .ZN(n17559) );
  OAI21_X1 U20704 ( .B1(n18312), .B2(n17595), .A(n17559), .ZN(P3_U2771) );
  AOI22_X1 U20705 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17590), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17599), .ZN(n17560) );
  OAI21_X1 U20706 ( .B1(n18317), .B2(n17595), .A(n17560), .ZN(P3_U2772) );
  AOI22_X1 U20707 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17590), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17599), .ZN(n17561) );
  OAI21_X1 U20708 ( .B1(n18321), .B2(n17595), .A(n17561), .ZN(P3_U2773) );
  AOI22_X1 U20709 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17590), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17599), .ZN(n17562) );
  OAI21_X1 U20710 ( .B1(n18325), .B2(n17595), .A(n17562), .ZN(P3_U2774) );
  AOI22_X1 U20711 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17590), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17599), .ZN(n17563) );
  OAI21_X1 U20712 ( .B1(n18329), .B2(n17595), .A(n17563), .ZN(P3_U2775) );
  AOI22_X1 U20713 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17590), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17599), .ZN(n17564) );
  OAI21_X1 U20714 ( .B1(n17583), .B2(n17595), .A(n17564), .ZN(P3_U2776) );
  AOI22_X1 U20715 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17590), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17599), .ZN(n17565) );
  OAI21_X1 U20716 ( .B1(n17585), .B2(n17595), .A(n17565), .ZN(P3_U2777) );
  AOI22_X1 U20717 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17590), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17599), .ZN(n17566) );
  OAI21_X1 U20718 ( .B1(n17587), .B2(n17595), .A(n17566), .ZN(P3_U2778) );
  AOI22_X1 U20719 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17590), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17581), .ZN(n17567) );
  OAI21_X1 U20720 ( .B1(n17589), .B2(n17592), .A(n17567), .ZN(P3_U2779) );
  AOI22_X1 U20721 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17590), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17581), .ZN(n17568) );
  OAI21_X1 U20722 ( .B1(n17593), .B2(n17592), .A(n17568), .ZN(P3_U2780) );
  AOI22_X1 U20723 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17590), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17581), .ZN(n17569) );
  OAI21_X1 U20724 ( .B1(n17596), .B2(n17592), .A(n17569), .ZN(P3_U2781) );
  AOI22_X1 U20725 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17600), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17581), .ZN(n17570) );
  OAI21_X1 U20726 ( .B1(n17571), .B2(n17602), .A(n17570), .ZN(P3_U2782) );
  AOI22_X1 U20727 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17590), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17581), .ZN(n17572) );
  OAI21_X1 U20728 ( .B1(n18296), .B2(n17592), .A(n17572), .ZN(P3_U2783) );
  AOI22_X1 U20729 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17600), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17581), .ZN(n17573) );
  OAI21_X1 U20730 ( .B1(n17574), .B2(n17602), .A(n17573), .ZN(P3_U2784) );
  AOI22_X1 U20731 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17590), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17581), .ZN(n17575) );
  OAI21_X1 U20732 ( .B1(n18308), .B2(n17592), .A(n17575), .ZN(P3_U2785) );
  AOI22_X1 U20733 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17590), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17581), .ZN(n17576) );
  OAI21_X1 U20734 ( .B1(n18312), .B2(n17592), .A(n17576), .ZN(P3_U2786) );
  AOI22_X1 U20735 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17590), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17581), .ZN(n17577) );
  OAI21_X1 U20736 ( .B1(n18317), .B2(n17592), .A(n17577), .ZN(P3_U2787) );
  AOI22_X1 U20737 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17590), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17581), .ZN(n17578) );
  OAI21_X1 U20738 ( .B1(n18321), .B2(n17592), .A(n17578), .ZN(P3_U2788) );
  AOI22_X1 U20739 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17590), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17581), .ZN(n17579) );
  OAI21_X1 U20740 ( .B1(n18325), .B2(n17592), .A(n17579), .ZN(P3_U2789) );
  AOI22_X1 U20741 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17590), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17581), .ZN(n17580) );
  OAI21_X1 U20742 ( .B1(n18329), .B2(n17592), .A(n17580), .ZN(P3_U2790) );
  AOI22_X1 U20743 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17590), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17581), .ZN(n17582) );
  OAI21_X1 U20744 ( .B1(n17583), .B2(n17592), .A(n17582), .ZN(P3_U2791) );
  AOI22_X1 U20745 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17590), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17599), .ZN(n17584) );
  OAI21_X1 U20746 ( .B1(n17585), .B2(n17592), .A(n17584), .ZN(P3_U2792) );
  AOI22_X1 U20747 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17590), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17599), .ZN(n17586) );
  OAI21_X1 U20748 ( .B1(n17587), .B2(n17592), .A(n17586), .ZN(P3_U2793) );
  AOI22_X1 U20749 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17590), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17599), .ZN(n17588) );
  OAI21_X1 U20750 ( .B1(n17589), .B2(n17592), .A(n17588), .ZN(P3_U2794) );
  AOI22_X1 U20751 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17590), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17599), .ZN(n17591) );
  OAI21_X1 U20752 ( .B1(n17593), .B2(n17592), .A(n17591), .ZN(P3_U2795) );
  AOI22_X1 U20753 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17590), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17599), .ZN(n17594) );
  OAI21_X1 U20754 ( .B1(n17596), .B2(n17595), .A(n17594), .ZN(P3_U2796) );
  AOI22_X1 U20755 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17600), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17599), .ZN(n17597) );
  OAI21_X1 U20756 ( .B1(n17598), .B2(n17602), .A(n17597), .ZN(P3_U2797) );
  AOI22_X1 U20757 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17600), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17599), .ZN(n17601) );
  OAI21_X1 U20758 ( .B1(n17603), .B2(n17602), .A(n17601), .ZN(P3_U2798) );
  INV_X1 U20759 ( .A(n17872), .ZN(n17927) );
  OAI21_X1 U20760 ( .B1(n17605), .B2(n18804), .A(n17968), .ZN(n17606) );
  AOI21_X1 U20761 ( .B1(n17927), .B2(n17604), .A(n17606), .ZN(n17635) );
  OAI21_X1 U20762 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17750), .A(
        n17635), .ZN(n17624) );
  NOR2_X1 U20763 ( .A1(n17802), .A2(n17604), .ZN(n17609) );
  XNOR2_X1 U20764 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B(n17607), .ZN(
        n17608) );
  AOI22_X1 U20765 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17624), .B1(
        n17609), .B2(n17608), .ZN(n17623) );
  AOI22_X1 U20766 ( .A1(n18198), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n17730), 
        .B2(n17610), .ZN(n17622) );
  NOR2_X1 U20767 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17611), .ZN(
        n17620) );
  OAI22_X1 U20768 ( .A1(n17978), .A2(n17972), .B1(n17612), .B2(n17808), .ZN(
        n17642) );
  NOR2_X1 U20769 ( .A1(n17988), .A2(n17642), .ZN(n17628) );
  AOI211_X1 U20770 ( .C1(n17972), .C2(n17808), .A(n17628), .B(n17613), .ZN(
        n17618) );
  AOI211_X1 U20771 ( .C1(n17616), .C2(n17615), .A(n17614), .B(n17879), .ZN(
        n17617) );
  AOI211_X1 U20772 ( .C1(n17620), .C2(n17619), .A(n17618), .B(n17617), .ZN(
        n17621) );
  NAND3_X1 U20773 ( .A1(n17623), .A2(n17622), .A3(n17621), .ZN(P3_U2802) );
  AOI22_X1 U20774 ( .A1(n18198), .A2(P3_REIP_REG_27__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17624), .ZN(n17633) );
  NOR2_X1 U20775 ( .A1(n17626), .A2(n17625), .ZN(n17627) );
  XNOR2_X1 U20776 ( .A(n17627), .B(n17795), .ZN(n17984) );
  AOI21_X1 U20777 ( .B1(n17988), .B2(n17629), .A(n17628), .ZN(n17631) );
  NOR3_X1 U20778 ( .A1(n17802), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        n17604), .ZN(n17630) );
  AOI211_X1 U20779 ( .C1(n17861), .C2(n17984), .A(n17631), .B(n17630), .ZN(
        n17632) );
  OAI211_X1 U20780 ( .C1(n17817), .C2(n17634), .A(n17633), .B(n17632), .ZN(
        P3_U2803) );
  AOI221_X1 U20781 ( .B1(n17637), .B2(n17636), .C1(n18313), .C2(n17636), .A(
        n17635), .ZN(n17638) );
  AOI221_X1 U20782 ( .B1(n17730), .B2(n17639), .C1(n17692), .C2(n17639), .A(
        n17638), .ZN(n17645) );
  OAI21_X1 U20783 ( .B1(n17641), .B2(n17995), .A(n17640), .ZN(n17992) );
  AOI22_X1 U20784 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17642), .B1(
        n17861), .B2(n17992), .ZN(n17644) );
  NOR2_X1 U20785 ( .A1(n20842), .A2(n17701), .ZN(n17683) );
  NAND4_X1 U20786 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17973), .A3(
        n17683), .A4(n17995), .ZN(n17643) );
  NAND2_X1 U20787 ( .A1(n18198), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17993) );
  NAND4_X1 U20788 ( .A1(n17645), .A2(n17644), .A3(n17643), .A4(n17993), .ZN(
        P3_U2804) );
  OAI21_X1 U20789 ( .B1(n17646), .B2(n18804), .A(n17968), .ZN(n17647) );
  AOI21_X1 U20790 ( .B1(n18678), .B2(n17655), .A(n17647), .ZN(n17680) );
  OAI21_X1 U20791 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17750), .A(
        n17680), .ZN(n17663) );
  AOI22_X1 U20792 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17663), .B1(
        n17730), .B2(n17648), .ZN(n17659) );
  XNOR2_X1 U20793 ( .A(n17649), .B(n18006), .ZN(n17997) );
  XNOR2_X1 U20794 ( .A(n17650), .B(n18006), .ZN(n18001) );
  OAI21_X1 U20795 ( .B1(n17795), .B2(n17652), .A(n17651), .ZN(n17653) );
  XNOR2_X1 U20796 ( .A(n17653), .B(n18006), .ZN(n18000) );
  OAI22_X1 U20797 ( .A1(n17972), .A2(n18001), .B1(n17879), .B2(n18000), .ZN(
        n17654) );
  AOI21_X1 U20798 ( .B1(n17881), .B2(n17997), .A(n17654), .ZN(n17658) );
  NAND2_X1 U20799 ( .A1(n18198), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18004) );
  NOR2_X1 U20800 ( .A1(n17802), .A2(n17655), .ZN(n17665) );
  OAI211_X1 U20801 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17665), .B(n17656), .ZN(n17657) );
  NAND4_X1 U20802 ( .A1(n17659), .A2(n17658), .A3(n18004), .A4(n17657), .ZN(
        P3_U2805) );
  INV_X1 U20803 ( .A(n17683), .ZN(n17672) );
  NAND2_X1 U20804 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18018), .ZN(
        n17671) );
  INV_X1 U20805 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17664) );
  AOI22_X1 U20806 ( .A1(n18198), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n17730), 
        .B2(n17660), .ZN(n17661) );
  INV_X1 U20807 ( .A(n17661), .ZN(n17662) );
  AOI221_X1 U20808 ( .B1(n17665), .B2(n17664), .C1(n17663), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17662), .ZN(n17670) );
  OAI22_X1 U20809 ( .A1(n18008), .A2(n17972), .B1(n17666), .B2(n17808), .ZN(
        n17682) );
  OAI21_X1 U20810 ( .B1(n17668), .B2(n18018), .A(n17667), .ZN(n18017) );
  AOI22_X1 U20811 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17682), .B1(
        n17861), .B2(n18017), .ZN(n17669) );
  OAI211_X1 U20812 ( .C1(n17672), .C2(n17671), .A(n17670), .B(n17669), .ZN(
        P3_U2806) );
  OAI22_X1 U20813 ( .A1(n17795), .A2(n20842), .B1(n17673), .B2(n17685), .ZN(
        n17674) );
  NOR2_X1 U20814 ( .A1(n17674), .A2(n17715), .ZN(n17675) );
  XNOR2_X1 U20815 ( .A(n17675), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18025) );
  AOI21_X1 U20816 ( .B1(n17676), .B2(n18678), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17679) );
  OAI21_X1 U20817 ( .B1(n17730), .B2(n17692), .A(n17677), .ZN(n17678) );
  NAND2_X1 U20818 ( .A1(n18198), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18024) );
  OAI211_X1 U20819 ( .C1(n17680), .C2(n17679), .A(n17678), .B(n18024), .ZN(
        n17681) );
  AOI221_X1 U20820 ( .B1(n17683), .B2(n18012), .C1(n17682), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17681), .ZN(n17684) );
  OAI21_X1 U20821 ( .B1(n17879), .B2(n18025), .A(n17684), .ZN(P3_U2807) );
  NAND2_X1 U20822 ( .A1(n17972), .A2(n17808), .ZN(n17717) );
  INV_X1 U20823 ( .A(n17972), .ZN(n17960) );
  NAND2_X1 U20824 ( .A1(n17960), .A2(n18104), .ZN(n17782) );
  OAI21_X1 U20825 ( .B1(n18036), .B2(n17808), .A(n17782), .ZN(n17770) );
  AOI21_X1 U20826 ( .B1(n18030), .B2(n17717), .A(n17770), .ZN(n17714) );
  INV_X1 U20827 ( .A(n17685), .ZN(n17687) );
  AOI21_X1 U20828 ( .B1(n17687), .B2(n17686), .A(n17715), .ZN(n17688) );
  XNOR2_X1 U20829 ( .A(n17688), .B(n20842), .ZN(n18039) );
  AOI22_X1 U20830 ( .A1(n17690), .A2(n17689), .B1(n17927), .B2(n17694), .ZN(
        n17691) );
  NAND2_X1 U20831 ( .A1(n17691), .A2(n17968), .ZN(n17719) );
  AOI21_X1 U20832 ( .B1(n17692), .B2(n20989), .A(n17719), .ZN(n17703) );
  AOI22_X1 U20833 ( .A1(n18198), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n17730), 
        .B2(n17693), .ZN(n17697) );
  NOR2_X1 U20834 ( .A1(n17802), .A2(n17694), .ZN(n17702) );
  OAI211_X1 U20835 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17702), .B(n17695), .ZN(n17696) );
  OAI211_X1 U20836 ( .C1(n17703), .C2(n17698), .A(n17697), .B(n17696), .ZN(
        n17699) );
  AOI21_X1 U20837 ( .B1(n17861), .B2(n18039), .A(n17699), .ZN(n17700) );
  OAI221_X1 U20838 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17701), 
        .C1(n20842), .C2(n17714), .A(n17700), .ZN(P3_U2808) );
  INV_X1 U20839 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18048) );
  INV_X1 U20840 ( .A(n17702), .ZN(n17705) );
  NAND2_X1 U20841 ( .A1(n18198), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18052) );
  OAI221_X1 U20842 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17705), .C1(
        n17704), .C2(n17703), .A(n18052), .ZN(n17711) );
  INV_X1 U20843 ( .A(n18033), .ZN(n18047) );
  OR3_X1 U20844 ( .A1(n17749), .A2(n17868), .A3(n17706), .ZN(n17726) );
  OAI22_X1 U20845 ( .A1(n18047), .A2(n17726), .B1(n17746), .B2(n17707), .ZN(
        n17708) );
  XOR2_X1 U20846 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17708), .Z(
        n18051) );
  INV_X1 U20847 ( .A(n18051), .ZN(n17709) );
  NAND2_X1 U20848 ( .A1(n18033), .A2(n18048), .ZN(n18054) );
  NOR2_X1 U20849 ( .A1(n18071), .A2(n17749), .ZN(n18045) );
  NAND2_X1 U20850 ( .A1(n17769), .A2(n18045), .ZN(n17738) );
  OAI22_X1 U20851 ( .A1(n17709), .A2(n17879), .B1(n18054), .B2(n17738), .ZN(
        n17710) );
  AOI211_X1 U20852 ( .C1(n17730), .C2(n17712), .A(n17711), .B(n17710), .ZN(
        n17713) );
  OAI21_X1 U20853 ( .B1(n17714), .B2(n18048), .A(n17713), .ZN(P3_U2809) );
  AOI221_X1 U20854 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17726), 
        .C1(n17737), .C2(n17744), .A(n17715), .ZN(n17716) );
  XNOR2_X1 U20855 ( .A(n17716), .B(n18031), .ZN(n18055) );
  NAND2_X1 U20856 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18045), .ZN(
        n18057) );
  AOI21_X1 U20857 ( .B1(n17717), .B2(n18057), .A(n17770), .ZN(n17736) );
  NAND2_X1 U20858 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18031), .ZN(
        n18064) );
  OAI22_X1 U20859 ( .A1(n17736), .A2(n18031), .B1(n17738), .B2(n18064), .ZN(
        n17718) );
  AOI21_X1 U20860 ( .B1(n17861), .B2(n18055), .A(n17718), .ZN(n17725) );
  NAND2_X1 U20861 ( .A1(n18198), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17724) );
  OAI221_X1 U20862 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18678), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n17720), .A(n17719), .ZN(
        n17723) );
  OAI21_X1 U20863 ( .B1(n17730), .B2(n17692), .A(n17721), .ZN(n17722) );
  NAND4_X1 U20864 ( .A1(n17725), .A2(n17724), .A3(n17723), .A4(n17722), .ZN(
        P3_U2810) );
  OAI21_X1 U20865 ( .B1(n17746), .B2(n17744), .A(n17726), .ZN(n17727) );
  XNOR2_X1 U20866 ( .A(n17727), .B(n17737), .ZN(n18065) );
  INV_X1 U20867 ( .A(n17968), .ZN(n17954) );
  AOI21_X1 U20868 ( .B1(n17927), .B2(n16826), .A(n17954), .ZN(n17753) );
  OAI21_X1 U20869 ( .B1(n17728), .B2(n18804), .A(n17753), .ZN(n17741) );
  AOI22_X1 U20870 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17741), .B1(
        n17730), .B2(n17729), .ZN(n17733) );
  NOR2_X1 U20871 ( .A1(n17802), .A2(n16826), .ZN(n17743) );
  OAI211_X1 U20872 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17743), .B(n17731), .ZN(n17732) );
  OAI211_X1 U20873 ( .C1(n20997), .C2(n18280), .A(n17733), .B(n17732), .ZN(
        n17734) );
  AOI21_X1 U20874 ( .B1(n17861), .B2(n18065), .A(n17734), .ZN(n17735) );
  OAI221_X1 U20875 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17738), 
        .C1(n17737), .C2(n17736), .A(n17735), .ZN(P3_U2811) );
  AOI21_X1 U20876 ( .B1(n17769), .B2(n18071), .A(n17770), .ZN(n17760) );
  INV_X1 U20877 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17742) );
  OAI22_X1 U20878 ( .A1(n18280), .A2(n18854), .B1(n17817), .B2(n17739), .ZN(
        n17740) );
  AOI221_X1 U20879 ( .B1(n17743), .B2(n17742), .C1(n17741), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17740), .ZN(n17748) );
  OAI21_X1 U20880 ( .B1(n17749), .B2(n17868), .A(n17744), .ZN(n17745) );
  XOR2_X1 U20881 ( .A(n17746), .B(n17745), .Z(n18082) );
  NOR2_X1 U20882 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18071), .ZN(
        n18081) );
  AOI22_X1 U20883 ( .A1(n17861), .A2(n18082), .B1(n17769), .B2(n18081), .ZN(
        n17747) );
  OAI211_X1 U20884 ( .C1(n17760), .C2(n17749), .A(n17748), .B(n17747), .ZN(
        P3_U2812) );
  AOI21_X1 U20885 ( .B1(n18678), .B2(n17751), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17752) );
  OAI22_X1 U20886 ( .A1(n17753), .A2(n17752), .B1(n18280), .B2(n18852), .ZN(
        n17754) );
  AOI21_X1 U20887 ( .B1(n17755), .B2(n17962), .A(n17754), .ZN(n17759) );
  OAI21_X1 U20888 ( .B1(n17757), .B2(n20847), .A(n17756), .ZN(n18087) );
  NOR2_X1 U20889 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18093), .ZN(
        n18086) );
  AOI22_X1 U20890 ( .A1(n17861), .A2(n18087), .B1(n17769), .B2(n18086), .ZN(
        n17758) );
  OAI211_X1 U20891 ( .C1(n17760), .C2(n20847), .A(n17759), .B(n17758), .ZN(
        P3_U2813) );
  AOI21_X1 U20892 ( .B1(n17795), .B2(n17762), .A(n17761), .ZN(n17763) );
  XNOR2_X1 U20893 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17763), .ZN(
        n18098) );
  AOI21_X1 U20894 ( .B1(n17927), .B2(n12724), .A(n17954), .ZN(n17791) );
  OAI21_X1 U20895 ( .B1(n17764), .B2(n18804), .A(n17791), .ZN(n17774) );
  NOR2_X1 U20896 ( .A1(n17802), .A2(n12724), .ZN(n17776) );
  OAI211_X1 U20897 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17776), .B(n17765), .ZN(n17766) );
  NAND2_X1 U20898 ( .A1(n18198), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n18096) );
  OAI211_X1 U20899 ( .C1(n17817), .C2(n17767), .A(n17766), .B(n18096), .ZN(
        n17768) );
  AOI21_X1 U20900 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17774), .A(
        n17768), .ZN(n17772) );
  AOI22_X1 U20901 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17770), .B1(
        n17769), .B2(n18093), .ZN(n17771) );
  OAI211_X1 U20902 ( .C1(n17879), .C2(n18098), .A(n17772), .B(n17771), .ZN(
        P3_U2814) );
  NOR2_X1 U20903 ( .A1(n18280), .A2(n18848), .ZN(n17773) );
  AOI221_X1 U20904 ( .B1(n17776), .B2(n17775), .C1(n17774), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17773), .ZN(n17786) );
  NOR2_X1 U20905 ( .A1(n18036), .A2(n17808), .ZN(n17784) );
  OAI21_X1 U20906 ( .B1(n18118), .B2(n17833), .A(n18103), .ZN(n18111) );
  NAND2_X1 U20907 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17778) );
  NAND2_X1 U20908 ( .A1(n18100), .A2(n17777), .ZN(n18135) );
  NOR2_X1 U20909 ( .A1(n17778), .A2(n18135), .ZN(n17794) );
  NOR2_X1 U20910 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17794), .ZN(
        n18108) );
  NOR2_X1 U20911 ( .A1(n18144), .A2(n17778), .ZN(n17779) );
  NAND2_X1 U20912 ( .A1(n17867), .A2(n17868), .ZN(n17853) );
  NOR3_X1 U20913 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17848), .A3(
        n17853), .ZN(n17814) );
  AOI22_X1 U20914 ( .A1(n17779), .A2(n18154), .B1(n17814), .B2(n18117), .ZN(
        n17780) );
  AOI221_X1 U20915 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18143), 
        .C1(n17868), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17780), .ZN(
        n17781) );
  XNOR2_X1 U20916 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17781), .ZN(
        n18105) );
  OAI22_X1 U20917 ( .A1(n18108), .A2(n17782), .B1(n17879), .B2(n18105), .ZN(
        n17783) );
  AOI21_X1 U20918 ( .B1(n17784), .B2(n18111), .A(n17783), .ZN(n17785) );
  OAI211_X1 U20919 ( .C1(n17817), .C2(n17787), .A(n17786), .B(n17785), .ZN(
        P3_U2815) );
  INV_X1 U20920 ( .A(n18100), .ZN(n18116) );
  NOR3_X1 U20921 ( .A1(n18116), .A2(n18117), .A3(n17833), .ZN(n17788) );
  OAI22_X1 U20922 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17788), .B1(
        n17833), .B2(n18118), .ZN(n18115) );
  AOI21_X1 U20923 ( .B1(n17789), .B2(n18678), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17790) );
  OAI22_X1 U20924 ( .A1(n17791), .A2(n17790), .B1(n18280), .B2(n18847), .ZN(
        n17792) );
  AOI21_X1 U20925 ( .B1(n17793), .B2(n17962), .A(n17792), .ZN(n17798) );
  INV_X1 U20926 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18120) );
  AOI221_X1 U20927 ( .B1(n18117), .B2(n18120), .C1(n18135), .C2(n18120), .A(
        n17794), .ZN(n18127) );
  NAND2_X1 U20928 ( .A1(n17795), .A2(n18154), .ZN(n17854) );
  NOR2_X1 U20929 ( .A1(n18116), .A2(n17854), .ZN(n17810) );
  AOI22_X1 U20930 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17810), .B1(
        n10159), .B2(n17814), .ZN(n17796) );
  XNOR2_X1 U20931 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17796), .ZN(
        n18126) );
  AOI22_X1 U20932 ( .A1(n17960), .A2(n18127), .B1(n17861), .B2(n18126), .ZN(
        n17797) );
  OAI211_X1 U20933 ( .C1(n17808), .C2(n18115), .A(n17798), .B(n17797), .ZN(
        P3_U2816) );
  NAND2_X1 U20934 ( .A1(n18100), .A2(n18117), .ZN(n18140) );
  AOI21_X1 U20935 ( .B1(n17927), .B2(n17801), .A(n17954), .ZN(n17799) );
  OAI21_X1 U20936 ( .B1(n17800), .B2(n18804), .A(n17799), .ZN(n17819) );
  NOR2_X1 U20937 ( .A1(n17802), .A2(n17801), .ZN(n17821) );
  OAI211_X1 U20938 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17821), .B(n17803), .ZN(n17805) );
  NAND2_X1 U20939 ( .A1(n18198), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17804) );
  OAI211_X1 U20940 ( .C1(n17817), .C2(n17806), .A(n17805), .B(n17804), .ZN(
        n17807) );
  AOI21_X1 U20941 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17819), .A(
        n17807), .ZN(n17813) );
  INV_X1 U20942 ( .A(n18135), .ZN(n17809) );
  NOR2_X1 U20943 ( .A1(n18116), .A2(n17833), .ZN(n18132) );
  OAI22_X1 U20944 ( .A1(n17809), .A2(n17972), .B1(n18132), .B2(n17808), .ZN(
        n17822) );
  AOI21_X1 U20945 ( .B1(n17814), .B2(n18143), .A(n17810), .ZN(n17811) );
  XNOR2_X1 U20946 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17811), .ZN(
        n18131) );
  AOI22_X1 U20947 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17822), .B1(
        n17861), .B2(n18131), .ZN(n17812) );
  OAI211_X1 U20948 ( .C1(n17864), .C2(n18140), .A(n17813), .B(n17812), .ZN(
        P3_U2817) );
  INV_X1 U20949 ( .A(n18160), .ZN(n17849) );
  NOR2_X1 U20950 ( .A1(n17849), .A2(n17854), .ZN(n17834) );
  AOI21_X1 U20951 ( .B1(n17834), .B2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n17814), .ZN(n17815) );
  XNOR2_X1 U20952 ( .A(n17815), .B(n18143), .ZN(n18149) );
  NAND2_X1 U20953 ( .A1(n18198), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18147) );
  OAI21_X1 U20954 ( .B1(n17817), .B2(n17816), .A(n18147), .ZN(n17818) );
  AOI221_X1 U20955 ( .B1(n17821), .B2(n17820), .C1(n17819), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17818), .ZN(n17825) );
  OAI21_X1 U20956 ( .B1(n18144), .B2(n17864), .A(n18143), .ZN(n17823) );
  NAND2_X1 U20957 ( .A1(n17823), .A2(n17822), .ZN(n17824) );
  OAI211_X1 U20958 ( .C1(n18149), .C2(n17879), .A(n17825), .B(n17824), .ZN(
        P3_U2818) );
  OR2_X1 U20959 ( .A1(n17849), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18166) );
  NAND2_X1 U20960 ( .A1(n18678), .A2(n17871), .ZN(n17826) );
  INV_X1 U20961 ( .A(n17826), .ZN(n17887) );
  NOR2_X1 U20962 ( .A1(n17827), .A2(n17826), .ZN(n17858) );
  NAND2_X1 U20963 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17858), .ZN(
        n17842) );
  NAND2_X1 U20964 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n17963), .ZN(
        n17828) );
  AOI22_X1 U20965 ( .A1(n17829), .A2(n17887), .B1(n17842), .B2(n17828), .ZN(
        n17831) );
  INV_X1 U20966 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18840) );
  NOR2_X1 U20967 ( .A1(n18280), .A2(n18840), .ZN(n17830) );
  AOI211_X1 U20968 ( .C1(n17832), .C2(n17962), .A(n17831), .B(n17830), .ZN(
        n17838) );
  AOI22_X1 U20969 ( .A1(n17960), .A2(n18156), .B1(n17881), .B2(n17833), .ZN(
        n17863) );
  OAI21_X1 U20970 ( .B1(n18160), .B2(n17864), .A(n17863), .ZN(n17836) );
  INV_X1 U20971 ( .A(n17834), .ZN(n17840) );
  OAI21_X1 U20972 ( .B1(n17853), .B2(n17848), .A(n17840), .ZN(n17835) );
  XOR2_X1 U20973 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17835), .Z(
        n18150) );
  AOI22_X1 U20974 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17836), .B1(
        n17861), .B2(n18150), .ZN(n17837) );
  OAI211_X1 U20975 ( .C1(n17864), .C2(n18166), .A(n17838), .B(n17837), .ZN(
        P3_U2819) );
  OAI221_X1 U20976 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17853), .C1(
        n18176), .C2(n17854), .A(n17852), .ZN(n17841) );
  NAND4_X1 U20977 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17867), .A3(
        n18176), .A4(n17868), .ZN(n17839) );
  AND3_X1 U20978 ( .A1(n17841), .A2(n17840), .A3(n17839), .ZN(n18171) );
  OAI211_X1 U20979 ( .C1(n17858), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n17963), .B(n17842), .ZN(n17844) );
  NAND2_X1 U20980 ( .A1(n18198), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n17843) );
  OAI211_X1 U20981 ( .C1(n17952), .C2(n17845), .A(n17844), .B(n17843), .ZN(
        n17846) );
  AOI21_X1 U20982 ( .B1(n17861), .B2(n18171), .A(n17846), .ZN(n17851) );
  NAND3_X1 U20983 ( .A1(n17849), .A2(n17848), .A3(n17847), .ZN(n17850) );
  OAI211_X1 U20984 ( .C1(n17863), .C2(n17852), .A(n17851), .B(n17850), .ZN(
        P3_U2820) );
  NAND2_X1 U20985 ( .A1(n17854), .A2(n17853), .ZN(n17855) );
  XNOR2_X1 U20986 ( .A(n17855), .B(n18176), .ZN(n18180) );
  NAND2_X1 U20987 ( .A1(n18198), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n18182) );
  INV_X1 U20988 ( .A(n18182), .ZN(n17860) );
  AOI22_X1 U20989 ( .A1(n17869), .A2(n17887), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17963), .ZN(n17857) );
  OAI22_X1 U20990 ( .A1(n17858), .A2(n17857), .B1(n17952), .B2(n17856), .ZN(
        n17859) );
  AOI211_X1 U20991 ( .C1(n17861), .C2(n18180), .A(n17860), .B(n17859), .ZN(
        n17862) );
  OAI221_X1 U20992 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17864), .C1(
        n18176), .C2(n17863), .A(n17862), .ZN(P3_U2821) );
  OAI21_X1 U20993 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17866), .A(
        n17865), .ZN(n18200) );
  NOR2_X1 U20994 ( .A1(n18154), .A2(n17867), .ZN(n18191) );
  XNOR2_X1 U20995 ( .A(n18191), .B(n17868), .ZN(n18195) );
  AOI211_X1 U20996 ( .C1(n17873), .C2(n17870), .A(n17869), .B(n18313), .ZN(
        n17877) );
  OAI21_X1 U20997 ( .B1(n17872), .B2(n17871), .A(n17968), .ZN(n17885) );
  INV_X1 U20998 ( .A(n17885), .ZN(n17874) );
  OAI22_X1 U20999 ( .A1(n17952), .A2(n17875), .B1(n17874), .B2(n17873), .ZN(
        n17876) );
  AOI211_X1 U21000 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n18198), .A(n17877), .B(
        n17876), .ZN(n17878) );
  OAI21_X1 U21001 ( .B1(n17879), .B2(n18195), .A(n17878), .ZN(n17880) );
  AOI21_X1 U21002 ( .B1(n18195), .B2(n17881), .A(n17880), .ZN(n17882) );
  OAI21_X1 U21003 ( .B1(n17972), .B2(n18200), .A(n17882), .ZN(P3_U2822) );
  OAI21_X1 U21004 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17884), .A(
        n17883), .ZN(n18202) );
  NOR2_X1 U21005 ( .A1(n18280), .A2(n18832), .ZN(n18206) );
  AOI221_X1 U21006 ( .B1(n17887), .B2(n17886), .C1(n17885), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18206), .ZN(n17895) );
  AOI21_X1 U21007 ( .B1(n17890), .B2(n17889), .A(n17888), .ZN(n17891) );
  XOR2_X1 U21008 ( .A(n17891), .B(n18203), .Z(n18210) );
  OAI22_X1 U21009 ( .A1(n17972), .A2(n18210), .B1(n17892), .B2(n17952), .ZN(
        n17893) );
  INV_X1 U21010 ( .A(n17893), .ZN(n17894) );
  OAI211_X1 U21011 ( .C1(n17971), .C2(n18202), .A(n17895), .B(n17894), .ZN(
        P3_U2823) );
  OAI21_X1 U21012 ( .B1(n17897), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n17896), .ZN(n18212) );
  NOR2_X1 U21013 ( .A1(n18313), .A2(n17901), .ZN(n17906) );
  OAI21_X1 U21014 ( .B1(n17900), .B2(n17899), .A(n17898), .ZN(n18211) );
  OAI22_X1 U21015 ( .A1(n17971), .A2(n18211), .B1(n18280), .B2(n20920), .ZN(
        n17904) );
  OAI21_X1 U21016 ( .B1(n17901), .B2(n18313), .A(n17963), .ZN(n17914) );
  OAI22_X1 U21017 ( .A1(n17952), .A2(n17902), .B1(n17905), .B2(n17914), .ZN(
        n17903) );
  AOI211_X1 U21018 ( .C1(n17906), .C2(n17905), .A(n17904), .B(n17903), .ZN(
        n17907) );
  OAI21_X1 U21019 ( .B1(n17972), .B2(n18212), .A(n17907), .ZN(P3_U2824) );
  OAI21_X1 U21020 ( .B1(n17910), .B2(n17909), .A(n17908), .ZN(n18219) );
  AOI21_X1 U21021 ( .B1(n17911), .B2(n17968), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17915) );
  OAI21_X1 U21022 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17913), .A(
        n17912), .ZN(n18225) );
  OAI22_X1 U21023 ( .A1(n17915), .A2(n17914), .B1(n17971), .B2(n18225), .ZN(
        n17916) );
  AOI21_X1 U21024 ( .B1(n17917), .B2(n17962), .A(n17916), .ZN(n17918) );
  NAND2_X1 U21025 ( .A1(n18198), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18218) );
  OAI211_X1 U21026 ( .C1(n17972), .C2(n18219), .A(n17918), .B(n18218), .ZN(
        P3_U2825) );
  OAI21_X1 U21027 ( .B1(n17921), .B2(n17920), .A(n17919), .ZN(n18236) );
  OAI21_X1 U21028 ( .B1(n17924), .B2(n17923), .A(n17922), .ZN(n18230) );
  OAI22_X1 U21029 ( .A1(n17972), .A2(n18230), .B1(n18313), .B2(n17925), .ZN(
        n17931) );
  AOI21_X1 U21030 ( .B1(n17927), .B2(n17926), .A(n17954), .ZN(n17940) );
  OAI22_X1 U21031 ( .A1(n17952), .A2(n17929), .B1(n17928), .B2(n17940), .ZN(
        n17930) );
  AOI211_X1 U21032 ( .C1(n18198), .C2(P3_REIP_REG_4__SCAN_IN), .A(n17931), .B(
        n17930), .ZN(n17932) );
  OAI21_X1 U21033 ( .B1(n17971), .B2(n18236), .A(n17932), .ZN(P3_U2826) );
  OAI21_X1 U21034 ( .B1(n17935), .B2(n17934), .A(n17933), .ZN(n18239) );
  AOI21_X1 U21035 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17968), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17941) );
  OAI21_X1 U21036 ( .B1(n17938), .B2(n17937), .A(n17936), .ZN(n17939) );
  XNOR2_X1 U21037 ( .A(n17939), .B(n18245), .ZN(n18238) );
  OAI22_X1 U21038 ( .A1(n17941), .A2(n17940), .B1(n17971), .B2(n18238), .ZN(
        n17942) );
  AOI21_X1 U21039 ( .B1(n17943), .B2(n17962), .A(n17942), .ZN(n17944) );
  NAND2_X1 U21040 ( .A1(n18198), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18243) );
  OAI211_X1 U21041 ( .C1(n17972), .C2(n18239), .A(n17944), .B(n18243), .ZN(
        P3_U2827) );
  OAI21_X1 U21042 ( .B1(n17947), .B2(n17946), .A(n17945), .ZN(n18256) );
  OAI21_X1 U21043 ( .B1(n17950), .B2(n17949), .A(n17948), .ZN(n18263) );
  OAI22_X1 U21044 ( .A1(n17952), .A2(n17951), .B1(n17971), .B2(n18263), .ZN(
        n17953) );
  AOI221_X1 U21045 ( .B1(n18678), .B2(n17955), .C1(n17954), .C2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17953), .ZN(n17956) );
  NAND2_X1 U21046 ( .A1(n18198), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18261) );
  OAI211_X1 U21047 ( .C1(n17972), .C2(n18256), .A(n17956), .B(n18261), .ZN(
        P3_U2828) );
  OAI21_X1 U21048 ( .B1(n17958), .B2(n17966), .A(n17957), .ZN(n18273) );
  NAND2_X1 U21049 ( .A1(n18911), .A2(n17967), .ZN(n17959) );
  XNOR2_X1 U21050 ( .A(n17959), .B(n17958), .ZN(n18270) );
  AOI22_X1 U21051 ( .A1(n17960), .A2(n18270), .B1(n18198), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17965) );
  AOI22_X1 U21052 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17963), .B1(
        n17962), .B2(n17961), .ZN(n17964) );
  OAI211_X1 U21053 ( .C1(n17971), .C2(n18273), .A(n17965), .B(n17964), .ZN(
        P3_U2829) );
  AOI21_X1 U21054 ( .B1(n17967), .B2(n18911), .A(n17966), .ZN(n18278) );
  INV_X1 U21055 ( .A(n18278), .ZN(n18276) );
  NAND3_X1 U21056 ( .A1(n18893), .A2(n18804), .A3(n17968), .ZN(n17969) );
  AOI22_X1 U21057 ( .A1(n18198), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17969), .ZN(n17970) );
  OAI221_X1 U21058 ( .B1(n18278), .B2(n17972), .C1(n18276), .C2(n17971), .A(
        n17970), .ZN(P3_U2830) );
  NAND2_X1 U21059 ( .A1(n18280), .A2(n18281), .ZN(n18266) );
  NOR2_X1 U21060 ( .A1(n20842), .A2(n18037), .ZN(n18022) );
  NAND3_X1 U21061 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17973), .A3(
        n18022), .ZN(n17990) );
  NOR2_X1 U21062 ( .A1(n17995), .A2(n17990), .ZN(n17983) );
  NOR2_X1 U21063 ( .A1(n18768), .A2(n9745), .ZN(n18060) );
  AOI21_X1 U21064 ( .B1(n18749), .B2(n18060), .A(n17974), .ZN(n17980) );
  OR2_X1 U21065 ( .A1(n17975), .A2(n18026), .ZN(n17976) );
  AOI22_X1 U21066 ( .A1(n18768), .A2(n17977), .B1(n18735), .B2(n17976), .ZN(
        n17999) );
  OAI21_X1 U21067 ( .B1(n17978), .B2(n18029), .A(n17999), .ZN(n17979) );
  AOI211_X1 U21068 ( .C1(n18192), .C2(n17981), .A(n17980), .B(n17979), .ZN(
        n17989) );
  INV_X1 U21069 ( .A(n17989), .ZN(n17982) );
  NAND2_X1 U21070 ( .A1(n18198), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17986) );
  OAI211_X1 U21071 ( .C1(n17988), .C2(n18266), .A(n17987), .B(n17986), .ZN(
        P3_U2835) );
  AOI211_X1 U21072 ( .C1(n17995), .C2(n17990), .A(n17989), .B(n18281), .ZN(
        n17991) );
  AOI21_X1 U21073 ( .B1(n18181), .B2(n17992), .A(n17991), .ZN(n17994) );
  OAI211_X1 U21074 ( .C1(n18266), .C2(n17995), .A(n17994), .B(n17993), .ZN(
        P3_U2836) );
  AOI22_X1 U21075 ( .A1(n17997), .A2(n18192), .B1(n17996), .B2(n18006), .ZN(
        n17998) );
  OAI21_X1 U21076 ( .B1(n17999), .B2(n18006), .A(n17998), .ZN(n18003) );
  OAI22_X1 U21077 ( .A1(n18257), .A2(n18001), .B1(n18194), .B2(n18000), .ZN(
        n18002) );
  AOI21_X1 U21078 ( .B1(n18265), .B2(n18003), .A(n18002), .ZN(n18005) );
  OAI211_X1 U21079 ( .C1(n18266), .C2(n18006), .A(n18005), .B(n18004), .ZN(
        P3_U2837) );
  OAI21_X1 U21080 ( .B1(n20842), .B2(n18026), .A(n18735), .ZN(n18007) );
  OAI211_X1 U21081 ( .C1(n18008), .C2(n18029), .A(n18266), .B(n18007), .ZN(
        n18009) );
  AOI21_X1 U21082 ( .B1(n18192), .B2(n18010), .A(n18009), .ZN(n18015) );
  INV_X1 U21083 ( .A(n18011), .ZN(n18013) );
  AOI21_X1 U21084 ( .B1(n18768), .B2(n18013), .A(n18012), .ZN(n18014) );
  AOI21_X1 U21085 ( .B1(n18015), .B2(n18014), .A(n18125), .ZN(n18021) );
  AOI21_X1 U21086 ( .B1(n18229), .B2(n18015), .A(n18018), .ZN(n18016) );
  AOI22_X1 U21087 ( .A1(n18181), .A2(n18017), .B1(n18021), .B2(n18016), .ZN(
        n18020) );
  NAND4_X1 U21088 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18265), .A3(
        n18022), .A4(n18018), .ZN(n18019) );
  OAI211_X1 U21089 ( .C1(n18862), .C2(n18280), .A(n18020), .B(n18019), .ZN(
        P3_U2838) );
  OAI221_X1 U21090 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18022), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n18266), .A(n18021), .ZN(
        n18023) );
  OAI211_X1 U21091 ( .C1(n18025), .C2(n18194), .A(n18024), .B(n18023), .ZN(
        P3_U2839) );
  AND2_X1 U21092 ( .A1(n9745), .A2(n18026), .ZN(n18035) );
  INV_X1 U21093 ( .A(n18768), .ZN(n18251) );
  AOI21_X1 U21094 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18027), .A(
        n18251), .ZN(n18028) );
  AOI221_X1 U21095 ( .B1(n18070), .B2(n18282), .C1(n18057), .C2(n18282), .A(
        n18028), .ZN(n18059) );
  NAND2_X1 U21096 ( .A1(n18029), .A2(n18153), .ZN(n18151) );
  AOI22_X1 U21097 ( .A1(n18282), .A2(n18031), .B1(n18030), .B2(n18151), .ZN(
        n18032) );
  NAND2_X1 U21098 ( .A1(n18059), .A2(n18032), .ZN(n18046) );
  OAI22_X1 U21099 ( .A1(n18162), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n18033), .B2(n18251), .ZN(n18034) );
  NOR4_X1 U21100 ( .A1(n18035), .A2(n20842), .A3(n18046), .A4(n18034), .ZN(
        n18038) );
  NOR2_X1 U21101 ( .A1(n18036), .A2(n18153), .ZN(n18112) );
  AOI21_X1 U21102 ( .B1(n18767), .B2(n18104), .A(n18112), .ZN(n18044) );
  AOI22_X1 U21103 ( .A1(n18038), .A2(n18044), .B1(n20842), .B2(n18037), .ZN(
        n18040) );
  AOI22_X1 U21104 ( .A1(n18265), .A2(n18040), .B1(n18181), .B2(n18039), .ZN(
        n18042) );
  NAND2_X1 U21105 ( .A1(n18198), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18041) );
  OAI211_X1 U21106 ( .C1(n18266), .C2(n20842), .A(n18042), .B(n18041), .ZN(
        P3_U2840) );
  NAND3_X1 U21107 ( .A1(n18265), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n18043), .ZN(n18069) );
  INV_X1 U21108 ( .A(n18060), .ZN(n18264) );
  NAND2_X1 U21109 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18157), .ZN(
        n18174) );
  NOR2_X1 U21110 ( .A1(n18080), .A2(n18174), .ZN(n18090) );
  OAI221_X1 U21111 ( .B1(n9746), .B2(n18045), .C1(n9746), .C2(n18090), .A(
        n18092), .ZN(n18056) );
  AOI211_X1 U21112 ( .C1(n18047), .C2(n18264), .A(n18046), .B(n18056), .ZN(
        n18049) );
  NOR3_X1 U21113 ( .A1(n18198), .A2(n18049), .A3(n18048), .ZN(n18050) );
  AOI21_X1 U21114 ( .B1(n18181), .B2(n18051), .A(n18050), .ZN(n18053) );
  OAI211_X1 U21115 ( .C1(n18054), .C2(n18069), .A(n18053), .B(n18052), .ZN(
        P3_U2841) );
  AOI22_X1 U21116 ( .A1(n18198), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18181), 
        .B2(n18055), .ZN(n18063) );
  AOI21_X1 U21117 ( .B1(n18057), .B2(n18151), .A(n18056), .ZN(n18058) );
  AOI21_X1 U21118 ( .B1(n18059), .B2(n18058), .A(n18125), .ZN(n18066) );
  NOR3_X1 U21119 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18060), .A3(
        n18945), .ZN(n18061) );
  OAI21_X1 U21120 ( .B1(n18066), .B2(n18061), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18062) );
  OAI211_X1 U21121 ( .C1(n18064), .C2(n18069), .A(n18063), .B(n18062), .ZN(
        P3_U2842) );
  AOI22_X1 U21122 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18066), .B1(
        n18181), .B2(n18065), .ZN(n18068) );
  NAND2_X1 U21123 ( .A1(n18198), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18067) );
  OAI211_X1 U21124 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18069), .A(
        n18068), .B(n18067), .ZN(P3_U2843) );
  INV_X1 U21125 ( .A(n18735), .ZN(n18744) );
  INV_X1 U21126 ( .A(n18187), .ZN(n18247) );
  NOR3_X1 U21127 ( .A1(n18247), .A2(n18093), .A3(n18070), .ZN(n18074) );
  AOI22_X1 U21128 ( .A1(n18768), .A2(n18072), .B1(n18071), .B2(n18151), .ZN(
        n18073) );
  OAI211_X1 U21129 ( .C1(n18744), .C2(n18074), .A(n18092), .B(n18073), .ZN(
        n18085) );
  OAI221_X1 U21130 ( .B1(n18085), .B2(n20847), .C1(n18085), .C2(n18735), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18084) );
  INV_X1 U21131 ( .A(n18250), .ZN(n18075) );
  NAND2_X1 U21132 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18226) );
  OAI22_X1 U21133 ( .A1(n18075), .A2(n18251), .B1(n18246), .B2(n18226), .ZN(
        n18241) );
  NAND2_X1 U21134 ( .A1(n18076), .A2(n18241), .ZN(n18214) );
  NOR2_X1 U21135 ( .A1(n18077), .A2(n18214), .ZN(n18099) );
  INV_X1 U21136 ( .A(n18099), .ZN(n18079) );
  AOI21_X1 U21137 ( .B1(n18079), .B2(n18078), .A(n18281), .ZN(n18170) );
  NOR2_X1 U21138 ( .A1(n18080), .A2(n18184), .ZN(n18094) );
  AOI22_X1 U21139 ( .A1(n18181), .A2(n18082), .B1(n18094), .B2(n18081), .ZN(
        n18083) );
  OAI221_X1 U21140 ( .B1(n18198), .B2(n18084), .C1(n18280), .C2(n18854), .A(
        n18083), .ZN(P3_U2844) );
  NAND2_X1 U21141 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18085), .ZN(
        n18089) );
  AOI22_X1 U21142 ( .A1(n18181), .A2(n18087), .B1(n18094), .B2(n18086), .ZN(
        n18088) );
  OAI221_X1 U21143 ( .B1(n18198), .B2(n18089), .C1(n18280), .C2(n18852), .A(
        n18088), .ZN(P3_U2845) );
  AOI21_X1 U21144 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n9746), .A(
        n18090), .ZN(n18091) );
  OAI22_X1 U21145 ( .A1(n18749), .A2(n18157), .B1(n18152), .B2(n18251), .ZN(
        n18134) );
  AOI211_X1 U21146 ( .C1(n18167), .C2(n18118), .A(n18091), .B(n18134), .ZN(
        n18102) );
  AOI221_X1 U21147 ( .B1(n18229), .B2(n18092), .C1(n18102), .C2(n18092), .A(
        n18198), .ZN(n18095) );
  AOI22_X1 U21148 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18095), .B1(
        n18094), .B2(n18093), .ZN(n18097) );
  OAI211_X1 U21149 ( .C1(n18098), .C2(n18194), .A(n18097), .B(n18096), .ZN(
        P3_U2846) );
  NAND3_X1 U21150 ( .A1(n18100), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n18099), .ZN(n18119) );
  AOI211_X1 U21151 ( .C1(n18103), .C2(n18119), .A(n18102), .B(n18101), .ZN(
        n18110) );
  NAND2_X1 U21152 ( .A1(n18767), .A2(n18104), .ZN(n18107) );
  OAI22_X1 U21153 ( .A1(n18108), .A2(n18107), .B1(n18106), .B2(n18105), .ZN(
        n18109) );
  AOI211_X1 U21154 ( .C1(n18112), .C2(n18111), .A(n18110), .B(n18109), .ZN(
        n18114) );
  INV_X1 U21155 ( .A(n18266), .ZN(n18260) );
  AOI22_X1 U21156 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18260), .B1(
        n18198), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n18113) );
  OAI21_X1 U21157 ( .B1(n18114), .B2(n18281), .A(n18113), .ZN(P3_U2847) );
  INV_X1 U21158 ( .A(n18115), .ZN(n18124) );
  NOR2_X1 U21159 ( .A1(n18116), .A2(n18174), .ZN(n18142) );
  NOR2_X1 U21160 ( .A1(n9746), .A2(n18142), .ZN(n18137) );
  AOI211_X1 U21161 ( .C1(n18117), .C2(n18264), .A(n18137), .B(n18134), .ZN(
        n18122) );
  OAI21_X1 U21162 ( .B1(n18120), .B2(n18167), .A(n18118), .ZN(n18121) );
  AOI22_X1 U21163 ( .A1(n18122), .A2(n18121), .B1(n18120), .B2(n18119), .ZN(
        n18123) );
  AOI21_X1 U21164 ( .B1(n18124), .B2(n18192), .A(n18123), .ZN(n18130) );
  AOI22_X1 U21165 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18260), .B1(
        n18125), .B2(P3_REIP_REG_14__SCAN_IN), .ZN(n18129) );
  AOI22_X1 U21166 ( .A1(n18277), .A2(n18127), .B1(n18181), .B2(n18126), .ZN(
        n18128) );
  OAI211_X1 U21167 ( .C1(n18130), .C2(n18281), .A(n18129), .B(n18128), .ZN(
        P3_U2848) );
  AOI22_X1 U21168 ( .A1(n18198), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18181), 
        .B2(n18131), .ZN(n18139) );
  INV_X1 U21169 ( .A(n18144), .ZN(n18161) );
  OAI22_X1 U21170 ( .A1(n18162), .A2(n18161), .B1(n18132), .B2(n18153), .ZN(
        n18133) );
  AOI211_X1 U21171 ( .C1(n18767), .C2(n18135), .A(n18134), .B(n18133), .ZN(
        n18141) );
  OAI211_X1 U21172 ( .C1(n18162), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18265), .B(n18141), .ZN(n18136) );
  OAI211_X1 U21173 ( .C1(n18137), .C2(n18136), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18280), .ZN(n18138) );
  OAI211_X1 U21174 ( .C1(n18140), .C2(n18184), .A(n18139), .B(n18138), .ZN(
        P3_U2849) );
  OAI211_X1 U21175 ( .C1(n18142), .C2(n9746), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n18141), .ZN(n18146) );
  OAI22_X1 U21176 ( .A1(n18144), .A2(n18184), .B1(n18143), .B2(n18281), .ZN(
        n18145) );
  AOI22_X1 U21177 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18260), .B1(
        n18146), .B2(n18145), .ZN(n18148) );
  OAI211_X1 U21178 ( .C1(n18149), .C2(n18194), .A(n18148), .B(n18147), .ZN(
        P3_U2850) );
  AOI22_X1 U21179 ( .A1(n18198), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18181), 
        .B2(n18150), .ZN(n18165) );
  INV_X1 U21180 ( .A(n18151), .ZN(n18159) );
  OAI22_X1 U21181 ( .A1(n18154), .A2(n18153), .B1(n18152), .B2(n18251), .ZN(
        n18155) );
  AOI211_X1 U21182 ( .C1(n18767), .C2(n18156), .A(n18281), .B(n18155), .ZN(
        n18178) );
  NOR2_X1 U21183 ( .A1(n18749), .A2(n18157), .ZN(n18175) );
  AOI221_X1 U21184 ( .B1(n18176), .B2(n9745), .C1(n18174), .C2(n9745), .A(
        n18175), .ZN(n18158) );
  OAI211_X1 U21185 ( .C1(n18160), .C2(n18159), .A(n18178), .B(n18158), .ZN(
        n18168) );
  OAI22_X1 U21186 ( .A1(n18162), .A2(n18161), .B1(n9746), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18163) );
  OAI211_X1 U21187 ( .C1(n18168), .C2(n18163), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18280), .ZN(n18164) );
  OAI211_X1 U21188 ( .C1(n18166), .C2(n18184), .A(n18165), .B(n18164), .ZN(
        P3_U2851) );
  OAI221_X1 U21189 ( .B1(n18168), .B2(n18167), .C1(n18168), .C2(n18176), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18173) );
  NOR2_X1 U21190 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18176), .ZN(
        n18169) );
  AOI22_X1 U21191 ( .A1(n18181), .A2(n18171), .B1(n18170), .B2(n18169), .ZN(
        n18172) );
  OAI221_X1 U21192 ( .B1(n18198), .B2(n18173), .C1(n18280), .C2(n18838), .A(
        n18172), .ZN(P3_U2852) );
  OAI21_X1 U21193 ( .B1(n18175), .B2(n9745), .A(n18174), .ZN(n18177) );
  AOI211_X1 U21194 ( .C1(n18178), .C2(n18177), .A(n18198), .B(n18176), .ZN(
        n18179) );
  AOI21_X1 U21195 ( .B1(n18181), .B2(n18180), .A(n18179), .ZN(n18183) );
  OAI211_X1 U21196 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18184), .A(
        n18183), .B(n18182), .ZN(P3_U2853) );
  AOI211_X1 U21197 ( .C1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n18229), .B(n18281), .ZN(n18208) );
  AOI22_X1 U21198 ( .A1(n18768), .A2(n18186), .B1(n18735), .B2(n18185), .ZN(
        n18188) );
  OAI221_X1 U21199 ( .B1(n18281), .B2(n18188), .C1(n18281), .C2(n18187), .A(
        n18266), .ZN(n18221) );
  NOR2_X1 U21200 ( .A1(n18208), .A2(n18221), .ZN(n18204) );
  INV_X1 U21201 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18189) );
  NOR2_X1 U21202 ( .A1(n18204), .A2(n18189), .ZN(n18197) );
  NOR4_X1 U21203 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18201), .A3(
        n18203), .A4(n18214), .ZN(n18190) );
  AOI21_X1 U21204 ( .B1(n18192), .B2(n18191), .A(n18190), .ZN(n18193) );
  OAI22_X1 U21205 ( .A1(n18195), .A2(n18194), .B1(n18193), .B2(n18281), .ZN(
        n18196) );
  AOI211_X1 U21206 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n18198), .A(n18197), .B(
        n18196), .ZN(n18199) );
  OAI21_X1 U21207 ( .B1(n18257), .B2(n18200), .A(n18199), .ZN(P3_U2854) );
  NOR2_X1 U21208 ( .A1(n18201), .A2(n18214), .ZN(n18207) );
  OAI22_X1 U21209 ( .A1(n18204), .A2(n18203), .B1(n18274), .B2(n18202), .ZN(
        n18205) );
  AOI211_X1 U21210 ( .C1(n18208), .C2(n18207), .A(n18206), .B(n18205), .ZN(
        n18209) );
  OAI21_X1 U21211 ( .B1(n18257), .B2(n18210), .A(n18209), .ZN(P3_U2855) );
  OAI22_X1 U21212 ( .A1(n18257), .A2(n18212), .B1(n18274), .B2(n18211), .ZN(
        n18213) );
  AOI21_X1 U21213 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18221), .A(
        n18213), .ZN(n18216) );
  OR3_X1 U21214 ( .A1(n18281), .A2(n18214), .A3(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18215) );
  OAI211_X1 U21215 ( .C1(n20920), .C2(n18280), .A(n18216), .B(n18215), .ZN(
        P3_U2856) );
  NAND3_X1 U21216 ( .A1(n18265), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18241), .ZN(n18231) );
  NOR2_X1 U21217 ( .A1(n18217), .A2(n18231), .ZN(n18223) );
  OAI21_X1 U21218 ( .B1(n18257), .B2(n18219), .A(n18218), .ZN(n18220) );
  AOI221_X1 U21219 ( .B1(n18223), .B2(n18222), .C1(n18221), .C2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n18220), .ZN(n18224) );
  OAI21_X1 U21220 ( .B1(n18274), .B2(n18225), .A(n18224), .ZN(P3_U2857) );
  OAI21_X1 U21221 ( .B1(n18247), .B2(n18226), .A(n18735), .ZN(n18227) );
  OAI211_X1 U21222 ( .C1(n18251), .C2(n18250), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n18227), .ZN(n18228) );
  NAND2_X1 U21223 ( .A1(n18265), .A2(n18228), .ZN(n18237) );
  AOI22_X1 U21224 ( .A1(n18229), .A2(n18265), .B1(n18266), .B2(n18237), .ZN(
        n18233) );
  OAI22_X1 U21225 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18231), .B1(
        n18230), .B2(n18257), .ZN(n18232) );
  AOI21_X1 U21226 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18233), .A(
        n18232), .ZN(n18235) );
  NAND2_X1 U21227 ( .A1(n18198), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n18234) );
  OAI211_X1 U21228 ( .C1(n18236), .C2(n18274), .A(n18235), .B(n18234), .ZN(
        P3_U2858) );
  INV_X1 U21229 ( .A(n18237), .ZN(n18242) );
  OAI22_X1 U21230 ( .A1(n18257), .A2(n18239), .B1(n18274), .B2(n18238), .ZN(
        n18240) );
  AOI221_X1 U21231 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18242), .C1(
        n18241), .C2(n18242), .A(n18240), .ZN(n18244) );
  OAI211_X1 U21232 ( .C1(n18266), .C2(n18245), .A(n18244), .B(n18243), .ZN(
        P3_U2859) );
  NOR2_X1 U21233 ( .A1(n10060), .A2(n18246), .ZN(n18255) );
  NAND2_X1 U21234 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18249) );
  OAI21_X1 U21235 ( .B1(n18247), .B2(n10060), .A(n18735), .ZN(n18248) );
  OAI21_X1 U21236 ( .B1(n18249), .B2(n18251), .A(n18248), .ZN(n18253) );
  NOR2_X1 U21237 ( .A1(n18251), .A2(n18250), .ZN(n18252) );
  AOI221_X1 U21238 ( .B1(n18255), .B2(n18254), .C1(n18253), .C2(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n18252), .ZN(n18258) );
  OAI22_X1 U21239 ( .A1(n18258), .A2(n18281), .B1(n18257), .B2(n18256), .ZN(
        n18259) );
  AOI21_X1 U21240 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n18260), .A(
        n18259), .ZN(n18262) );
  OAI211_X1 U21241 ( .C1(n18263), .C2(n18274), .A(n18262), .B(n18261), .ZN(
        P3_U2860) );
  NAND3_X1 U21242 ( .A1(n18265), .A2(n18911), .A3(n18264), .ZN(n18284) );
  AOI21_X1 U21243 ( .B1(n18266), .B2(n18284), .A(n10060), .ZN(n18269) );
  AOI211_X1 U21244 ( .C1(n18749), .C2(n18911), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18267), .ZN(n18268) );
  AOI211_X1 U21245 ( .C1(n18277), .C2(n18270), .A(n18269), .B(n18268), .ZN(
        n18272) );
  NAND2_X1 U21246 ( .A1(n18198), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18271) );
  OAI211_X1 U21247 ( .C1(n18273), .C2(n18274), .A(n18272), .B(n18271), .ZN(
        P3_U2861) );
  INV_X1 U21248 ( .A(n18274), .ZN(n18279) );
  INV_X1 U21249 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18922) );
  NOR2_X1 U21250 ( .A1(n18280), .A2(n18922), .ZN(n18275) );
  AOI221_X1 U21251 ( .B1(n18279), .B2(n18278), .C1(n18277), .C2(n18276), .A(
        n18275), .ZN(n18285) );
  OAI211_X1 U21252 ( .C1(n18282), .C2(n18281), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18280), .ZN(n18283) );
  NAND3_X1 U21253 ( .A1(n18285), .A2(n18284), .A3(n18283), .ZN(P3_U2862) );
  AOI211_X1 U21254 ( .C1(n18287), .C2(n18286), .A(n18893), .B(n18945), .ZN(
        n18786) );
  OAI21_X1 U21255 ( .B1(n18786), .B2(n18336), .A(n18295), .ZN(n18288) );
  OAI221_X1 U21256 ( .B1(n18752), .B2(n18929), .C1(n18752), .C2(n18295), .A(
        n18288), .ZN(P3_U2863) );
  INV_X1 U21257 ( .A(n18289), .ZN(n18291) );
  AOI21_X1 U21258 ( .B1(n18291), .B2(n18754), .A(n18290), .ZN(n18294) );
  OAI221_X1 U21259 ( .B1(n18641), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18641), .C2(n18291), .A(n18295), .ZN(n18292) );
  AOI22_X1 U21260 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18294), .B1(
        n18292), .B2(n21008), .ZN(P3_U2865) );
  INV_X1 U21261 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18761) );
  NOR2_X1 U21262 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18761), .ZN(
        n18585) );
  NOR2_X1 U21263 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n21008), .ZN(
        n18470) );
  NOR2_X1 U21264 ( .A1(n18585), .A2(n18470), .ZN(n18293) );
  OAI22_X1 U21265 ( .A1(n18294), .A2(n18761), .B1(n18293), .B2(n18292), .ZN(
        P3_U2866) );
  NOR2_X1 U21266 ( .A1(n18762), .A2(n18295), .ZN(P3_U2867) );
  NAND2_X1 U21267 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18298) );
  NOR2_X1 U21268 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18298), .ZN(
        n18677) );
  NAND2_X1 U21269 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18677), .ZN(
        n18721) );
  NAND2_X1 U21270 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18678), .ZN(n18646) );
  NOR2_X2 U21271 ( .A1(n18445), .A2(n18296), .ZN(n18673) );
  INV_X1 U21272 ( .A(n18298), .ZN(n18297) );
  NAND2_X1 U21273 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18297), .ZN(
        n18672) );
  NOR2_X2 U21274 ( .A1(n18752), .A2(n18672), .ZN(n18727) );
  NAND2_X1 U21275 ( .A1(n18754), .A2(n18752), .ZN(n18755) );
  NAND2_X1 U21276 ( .A1(n21008), .A2(n18761), .ZN(n18377) );
  NOR2_X1 U21277 ( .A1(n18727), .A2(n18396), .ZN(n18357) );
  NOR2_X1 U21278 ( .A1(n18794), .A2(n18357), .ZN(n18330) );
  AND2_X1 U21279 ( .A1(n18678), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18679) );
  NAND2_X1 U21280 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18752), .ZN(
        n18356) );
  AOI22_X1 U21281 ( .A1(n18673), .A2(n18330), .B1(n18679), .B2(n18664), .ZN(
        n18303) );
  INV_X1 U21282 ( .A(n18356), .ZN(n18539) );
  NOR2_X1 U21283 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18752), .ZN(
        n18514) );
  NOR2_X1 U21284 ( .A1(n18539), .A2(n18514), .ZN(n18587) );
  NOR2_X1 U21285 ( .A1(n18587), .A2(n18298), .ZN(n18642) );
  AOI21_X1 U21286 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18445), .ZN(n18639) );
  INV_X1 U21287 ( .A(n18357), .ZN(n18299) );
  AOI22_X1 U21288 ( .A1(n18678), .A2(n18642), .B1(n18639), .B2(n18299), .ZN(
        n18333) );
  NAND2_X1 U21289 ( .A1(n18301), .A2(n18300), .ZN(n18331) );
  NOR2_X1 U21290 ( .A1(n18932), .A2(n18331), .ZN(n18643) );
  AOI22_X1 U21291 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18333), .B1(
        n18396), .B2(n18643), .ZN(n18302) );
  OAI211_X1 U21292 ( .C1(n18721), .C2(n18646), .A(n18303), .B(n18302), .ZN(
        P3_U2868) );
  NAND2_X1 U21293 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18678), .ZN(n18650) );
  NOR2_X2 U21294 ( .A1(n18445), .A2(n18304), .ZN(n18683) );
  AND2_X1 U21295 ( .A1(n18678), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18685) );
  AOI22_X1 U21296 ( .A1(n18330), .A2(n18683), .B1(n18664), .B2(n18685), .ZN(
        n18307) );
  NOR2_X1 U21297 ( .A1(n18305), .A2(n18331), .ZN(n18647) );
  AOI22_X1 U21298 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18333), .B1(
        n18396), .B2(n18647), .ZN(n18306) );
  OAI211_X1 U21299 ( .C1(n18721), .C2(n18650), .A(n18307), .B(n18306), .ZN(
        P3_U2869) );
  NAND2_X1 U21300 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18678), .ZN(n18695) );
  NOR2_X2 U21301 ( .A1(n18445), .A2(n18308), .ZN(n18690) );
  AND2_X1 U21302 ( .A1(n18678), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18691) );
  AOI22_X1 U21303 ( .A1(n18330), .A2(n18690), .B1(n18664), .B2(n18691), .ZN(
        n18311) );
  NOR2_X1 U21304 ( .A1(n18309), .A2(n18331), .ZN(n18692) );
  AOI22_X1 U21305 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18333), .B1(
        n18396), .B2(n18692), .ZN(n18310) );
  OAI211_X1 U21306 ( .C1(n18721), .C2(n18695), .A(n18311), .B(n18310), .ZN(
        P3_U2870) );
  NAND2_X1 U21307 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18678), .ZN(n18701) );
  NOR2_X2 U21308 ( .A1(n18445), .A2(n18312), .ZN(n18696) );
  NOR2_X2 U21309 ( .A1(n18313), .A2(n20937), .ZN(n18697) );
  AOI22_X1 U21310 ( .A1(n18330), .A2(n18696), .B1(n18664), .B2(n18697), .ZN(
        n18316) );
  NOR2_X1 U21311 ( .A1(n18314), .A2(n18331), .ZN(n18698) );
  AOI22_X1 U21312 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18333), .B1(
        n18396), .B2(n18698), .ZN(n18315) );
  OAI211_X1 U21313 ( .C1(n18721), .C2(n18701), .A(n18316), .B(n18315), .ZN(
        P3_U2871) );
  NAND2_X1 U21314 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18678), .ZN(n18658) );
  NOR2_X2 U21315 ( .A1(n18445), .A2(n18317), .ZN(n18702) );
  NAND2_X1 U21316 ( .A1(n18678), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18707) );
  INV_X1 U21317 ( .A(n18707), .ZN(n18655) );
  AOI22_X1 U21318 ( .A1(n18330), .A2(n18702), .B1(n18664), .B2(n18655), .ZN(
        n18320) );
  NOR2_X2 U21319 ( .A1(n18318), .A2(n18331), .ZN(n18704) );
  AOI22_X1 U21320 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18333), .B1(
        n18396), .B2(n18704), .ZN(n18319) );
  OAI211_X1 U21321 ( .C1(n18721), .C2(n18658), .A(n18320), .B(n18319), .ZN(
        P3_U2872) );
  INV_X1 U21322 ( .A(n18664), .ZN(n18355) );
  NAND2_X1 U21323 ( .A1(n18678), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18662) );
  INV_X1 U21324 ( .A(n18721), .ZN(n18725) );
  NAND2_X1 U21325 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18678), .ZN(n18713) );
  INV_X1 U21326 ( .A(n18713), .ZN(n18659) );
  NOR2_X2 U21327 ( .A1(n18445), .A2(n18321), .ZN(n18708) );
  AOI22_X1 U21328 ( .A1(n18725), .A2(n18659), .B1(n18330), .B2(n18708), .ZN(
        n18324) );
  NOR2_X2 U21329 ( .A1(n18322), .A2(n18331), .ZN(n18710) );
  AOI22_X1 U21330 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18333), .B1(
        n18396), .B2(n18710), .ZN(n18323) );
  OAI211_X1 U21331 ( .C1(n18355), .C2(n18662), .A(n18324), .B(n18323), .ZN(
        P3_U2873) );
  NAND2_X1 U21332 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18678), .ZN(n18606) );
  NOR2_X2 U21333 ( .A1(n18445), .A2(n18325), .ZN(n18714) );
  NAND2_X1 U21334 ( .A1(n18678), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18720) );
  INV_X1 U21335 ( .A(n18720), .ZN(n18602) );
  AOI22_X1 U21336 ( .A1(n18330), .A2(n18714), .B1(n18664), .B2(n18602), .ZN(
        n18328) );
  NOR2_X2 U21337 ( .A1(n18326), .A2(n18331), .ZN(n18717) );
  AOI22_X1 U21338 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18333), .B1(
        n18396), .B2(n18717), .ZN(n18327) );
  OAI211_X1 U21339 ( .C1(n18721), .C2(n18606), .A(n18328), .B(n18327), .ZN(
        P3_U2874) );
  NAND2_X1 U21340 ( .A1(n18678), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18732) );
  NOR2_X2 U21341 ( .A1(n18329), .A2(n18445), .ZN(n18723) );
  NAND2_X1 U21342 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18678), .ZN(n18613) );
  INV_X1 U21343 ( .A(n18613), .ZN(n18724) );
  AOI22_X1 U21344 ( .A1(n18330), .A2(n18723), .B1(n18664), .B2(n18724), .ZN(
        n18335) );
  NOR2_X2 U21345 ( .A1(n18332), .A2(n18331), .ZN(n18726) );
  AOI22_X1 U21346 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18333), .B1(
        n18396), .B2(n18726), .ZN(n18334) );
  OAI211_X1 U21347 ( .C1(n18721), .C2(n18732), .A(n18335), .B(n18334), .ZN(
        P3_U2875) );
  INV_X1 U21348 ( .A(n18643), .ZN(n18682) );
  INV_X1 U21349 ( .A(n18377), .ZN(n18379) );
  NAND2_X1 U21350 ( .A1(n18514), .A2(n18379), .ZN(n18414) );
  INV_X1 U21351 ( .A(n18646), .ZN(n18674) );
  NAND2_X1 U21352 ( .A1(n18754), .A2(n18637), .ZN(n18515) );
  NOR2_X1 U21353 ( .A1(n18377), .A2(n18515), .ZN(n18351) );
  AOI22_X1 U21354 ( .A1(n18674), .A2(n18664), .B1(n18673), .B2(n18351), .ZN(
        n18338) );
  INV_X1 U21355 ( .A(n18672), .ZN(n18676) );
  NOR2_X1 U21356 ( .A1(n18445), .A2(n18336), .ZN(n18675) );
  INV_X1 U21357 ( .A(n18675), .ZN(n18378) );
  NOR2_X1 U21358 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18378), .ZN(
        n18422) );
  AOI22_X1 U21359 ( .A1(n18678), .A2(n18676), .B1(n18379), .B2(n18422), .ZN(
        n18352) );
  AOI22_X1 U21360 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18352), .B1(
        n18727), .B2(n18679), .ZN(n18337) );
  OAI211_X1 U21361 ( .C1(n18682), .C2(n18414), .A(n18338), .B(n18337), .ZN(
        P3_U2876) );
  AOI22_X1 U21362 ( .A1(n18727), .A2(n18685), .B1(n18683), .B2(n18351), .ZN(
        n18340) );
  INV_X1 U21363 ( .A(n18414), .ZN(n18418) );
  AOI22_X1 U21364 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18352), .B1(
        n18647), .B2(n18418), .ZN(n18339) );
  OAI211_X1 U21365 ( .C1(n18355), .C2(n18650), .A(n18340), .B(n18339), .ZN(
        P3_U2877) );
  INV_X1 U21366 ( .A(n18692), .ZN(n18524) );
  INV_X1 U21367 ( .A(n18695), .ZN(n18521) );
  AOI22_X1 U21368 ( .A1(n18664), .A2(n18521), .B1(n18690), .B2(n18351), .ZN(
        n18342) );
  AOI22_X1 U21369 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18352), .B1(
        n18727), .B2(n18691), .ZN(n18341) );
  OAI211_X1 U21370 ( .C1(n18524), .C2(n18414), .A(n18342), .B(n18341), .ZN(
        P3_U2878) );
  INV_X1 U21371 ( .A(n18698), .ZN(n18624) );
  INV_X1 U21372 ( .A(n18701), .ZN(n18621) );
  AOI22_X1 U21373 ( .A1(n18664), .A2(n18621), .B1(n18696), .B2(n18351), .ZN(
        n18344) );
  AOI22_X1 U21374 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18352), .B1(
        n18727), .B2(n18697), .ZN(n18343) );
  OAI211_X1 U21375 ( .C1(n18624), .C2(n18414), .A(n18344), .B(n18343), .ZN(
        P3_U2879) );
  AOI22_X1 U21376 ( .A1(n18727), .A2(n18655), .B1(n18702), .B2(n18351), .ZN(
        n18346) );
  AOI22_X1 U21377 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18352), .B1(
        n18704), .B2(n18418), .ZN(n18345) );
  OAI211_X1 U21378 ( .C1(n18355), .C2(n18658), .A(n18346), .B(n18345), .ZN(
        P3_U2880) );
  INV_X1 U21379 ( .A(n18727), .ZN(n18689) );
  AOI22_X1 U21380 ( .A1(n18664), .A2(n18659), .B1(n18708), .B2(n18351), .ZN(
        n18348) );
  AOI22_X1 U21381 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18352), .B1(
        n18710), .B2(n18418), .ZN(n18347) );
  OAI211_X1 U21382 ( .C1(n18689), .C2(n18662), .A(n18348), .B(n18347), .ZN(
        P3_U2881) );
  INV_X1 U21383 ( .A(n18606), .ZN(n18716) );
  AOI22_X1 U21384 ( .A1(n18664), .A2(n18716), .B1(n18714), .B2(n18351), .ZN(
        n18350) );
  AOI22_X1 U21385 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18352), .B1(
        n18717), .B2(n18418), .ZN(n18349) );
  OAI211_X1 U21386 ( .C1(n18689), .C2(n18720), .A(n18350), .B(n18349), .ZN(
        P3_U2882) );
  AOI22_X1 U21387 ( .A1(n18727), .A2(n18724), .B1(n18723), .B2(n18351), .ZN(
        n18354) );
  AOI22_X1 U21388 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18352), .B1(
        n18726), .B2(n18418), .ZN(n18353) );
  OAI211_X1 U21389 ( .C1(n18355), .C2(n18732), .A(n18354), .B(n18353), .ZN(
        P3_U2883) );
  NOR2_X1 U21390 ( .A1(n18418), .A2(n18434), .ZN(n18400) );
  NOR2_X1 U21391 ( .A1(n18794), .A2(n18400), .ZN(n18373) );
  AOI22_X1 U21392 ( .A1(n18396), .A2(n18679), .B1(n18673), .B2(n18373), .ZN(
        n18360) );
  INV_X1 U21393 ( .A(n18641), .ZN(n18540) );
  OAI21_X1 U21394 ( .B1(n18357), .B2(n18540), .A(n18400), .ZN(n18358) );
  OAI211_X1 U21395 ( .C1(n18434), .C2(n18887), .A(n18589), .B(n18358), .ZN(
        n18374) );
  AOI22_X1 U21396 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18374), .B1(
        n18643), .B2(n18434), .ZN(n18359) );
  OAI211_X1 U21397 ( .C1(n18646), .C2(n18689), .A(n18360), .B(n18359), .ZN(
        P3_U2884) );
  INV_X1 U21398 ( .A(n18647), .ZN(n18688) );
  INV_X1 U21399 ( .A(n18434), .ZN(n18443) );
  INV_X1 U21400 ( .A(n18650), .ZN(n18684) );
  AOI22_X1 U21401 ( .A1(n18727), .A2(n18684), .B1(n18683), .B2(n18373), .ZN(
        n18362) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18374), .B1(
        n18396), .B2(n18685), .ZN(n18361) );
  OAI211_X1 U21403 ( .C1(n18688), .C2(n18443), .A(n18362), .B(n18361), .ZN(
        P3_U2885) );
  AOI22_X1 U21404 ( .A1(n18396), .A2(n18691), .B1(n18690), .B2(n18373), .ZN(
        n18364) );
  AOI22_X1 U21405 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18374), .B1(
        n18692), .B2(n18434), .ZN(n18363) );
  OAI211_X1 U21406 ( .C1(n18689), .C2(n18695), .A(n18364), .B(n18363), .ZN(
        P3_U2886) );
  AOI22_X1 U21407 ( .A1(n18396), .A2(n18697), .B1(n18696), .B2(n18373), .ZN(
        n18366) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18374), .B1(
        n18698), .B2(n18434), .ZN(n18365) );
  OAI211_X1 U21409 ( .C1(n18689), .C2(n18701), .A(n18366), .B(n18365), .ZN(
        P3_U2887) );
  AOI22_X1 U21410 ( .A1(n18396), .A2(n18655), .B1(n18702), .B2(n18373), .ZN(
        n18368) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18374), .B1(
        n18704), .B2(n18434), .ZN(n18367) );
  OAI211_X1 U21412 ( .C1(n18689), .C2(n18658), .A(n18368), .B(n18367), .ZN(
        P3_U2888) );
  INV_X1 U21413 ( .A(n18396), .ZN(n18392) );
  AOI22_X1 U21414 ( .A1(n18727), .A2(n18659), .B1(n18708), .B2(n18373), .ZN(
        n18370) );
  AOI22_X1 U21415 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18374), .B1(
        n18710), .B2(n18434), .ZN(n18369) );
  OAI211_X1 U21416 ( .C1(n18392), .C2(n18662), .A(n18370), .B(n18369), .ZN(
        P3_U2889) );
  AOI22_X1 U21417 ( .A1(n18396), .A2(n18602), .B1(n18714), .B2(n18373), .ZN(
        n18372) );
  AOI22_X1 U21418 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18374), .B1(
        n18717), .B2(n18434), .ZN(n18371) );
  OAI211_X1 U21419 ( .C1(n18689), .C2(n18606), .A(n18372), .B(n18371), .ZN(
        P3_U2890) );
  AOI22_X1 U21420 ( .A1(n18396), .A2(n18724), .B1(n18723), .B2(n18373), .ZN(
        n18376) );
  AOI22_X1 U21421 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18374), .B1(
        n18726), .B2(n18434), .ZN(n18375) );
  OAI211_X1 U21422 ( .C1(n18689), .C2(n18732), .A(n18376), .B(n18375), .ZN(
        P3_U2891) );
  NOR2_X1 U21423 ( .A1(n18754), .A2(n18377), .ZN(n18423) );
  AND2_X1 U21424 ( .A1(n18637), .A2(n18423), .ZN(n18395) );
  AOI22_X1 U21425 ( .A1(n18673), .A2(n18395), .B1(n18679), .B2(n18418), .ZN(
        n18381) );
  AOI21_X1 U21426 ( .B1(n18754), .B2(n18540), .A(n18378), .ZN(n18469) );
  NAND2_X1 U21427 ( .A1(n18379), .A2(n18469), .ZN(n18397) );
  NAND2_X1 U21428 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18423), .ZN(
        n18467) );
  INV_X1 U21429 ( .A(n18467), .ZN(n18456) );
  AOI22_X1 U21430 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18397), .B1(
        n18643), .B2(n18456), .ZN(n18380) );
  OAI211_X1 U21431 ( .C1(n18646), .C2(n18392), .A(n18381), .B(n18380), .ZN(
        P3_U2892) );
  AOI22_X1 U21432 ( .A1(n18396), .A2(n18684), .B1(n18683), .B2(n18395), .ZN(
        n18383) );
  AOI22_X1 U21433 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18397), .B1(
        n18685), .B2(n18418), .ZN(n18382) );
  OAI211_X1 U21434 ( .C1(n18688), .C2(n18467), .A(n18383), .B(n18382), .ZN(
        P3_U2893) );
  AOI22_X1 U21435 ( .A1(n18396), .A2(n18521), .B1(n18690), .B2(n18395), .ZN(
        n18385) );
  AOI22_X1 U21436 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18397), .B1(
        n18691), .B2(n18418), .ZN(n18384) );
  OAI211_X1 U21437 ( .C1(n18524), .C2(n18467), .A(n18385), .B(n18384), .ZN(
        P3_U2894) );
  AOI22_X1 U21438 ( .A1(n18396), .A2(n18621), .B1(n18696), .B2(n18395), .ZN(
        n18387) );
  AOI22_X1 U21439 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18397), .B1(
        n18697), .B2(n18418), .ZN(n18386) );
  OAI211_X1 U21440 ( .C1(n18624), .C2(n18467), .A(n18387), .B(n18386), .ZN(
        P3_U2895) );
  AOI22_X1 U21441 ( .A1(n18655), .A2(n18418), .B1(n18702), .B2(n18395), .ZN(
        n18389) );
  AOI22_X1 U21442 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18397), .B1(
        n18704), .B2(n18456), .ZN(n18388) );
  OAI211_X1 U21443 ( .C1(n18392), .C2(n18658), .A(n18389), .B(n18388), .ZN(
        P3_U2896) );
  INV_X1 U21444 ( .A(n18662), .ZN(n18709) );
  AOI22_X1 U21445 ( .A1(n18709), .A2(n18418), .B1(n18708), .B2(n18395), .ZN(
        n18391) );
  AOI22_X1 U21446 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18397), .B1(
        n18710), .B2(n18456), .ZN(n18390) );
  OAI211_X1 U21447 ( .C1(n18392), .C2(n18713), .A(n18391), .B(n18390), .ZN(
        P3_U2897) );
  AOI22_X1 U21448 ( .A1(n18396), .A2(n18716), .B1(n18714), .B2(n18395), .ZN(
        n18394) );
  AOI22_X1 U21449 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18397), .B1(
        n18717), .B2(n18456), .ZN(n18393) );
  OAI211_X1 U21450 ( .C1(n18720), .C2(n18414), .A(n18394), .B(n18393), .ZN(
        P3_U2898) );
  INV_X1 U21451 ( .A(n18732), .ZN(n18609) );
  AOI22_X1 U21452 ( .A1(n18396), .A2(n18609), .B1(n18723), .B2(n18395), .ZN(
        n18399) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18397), .B1(
        n18726), .B2(n18456), .ZN(n18398) );
  OAI211_X1 U21454 ( .C1(n18613), .C2(n18414), .A(n18399), .B(n18398), .ZN(
        P3_U2899) );
  INV_X1 U21455 ( .A(n18755), .ZN(n18491) );
  NAND2_X1 U21456 ( .A1(n18491), .A2(n18470), .ZN(n18483) );
  AOI21_X1 U21457 ( .B1(n18467), .B2(n18483), .A(n18794), .ZN(n18417) );
  AOI22_X1 U21458 ( .A1(n18674), .A2(n18418), .B1(n18673), .B2(n18417), .ZN(
        n18403) );
  INV_X1 U21459 ( .A(n18483), .ZN(n18487) );
  AOI221_X1 U21460 ( .B1(n18400), .B2(n18467), .C1(n18540), .C2(n18467), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18401) );
  OAI21_X1 U21461 ( .B1(n18487), .B2(n18401), .A(n18589), .ZN(n18419) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18419), .B1(
        n18679), .B2(n18434), .ZN(n18402) );
  OAI211_X1 U21463 ( .C1(n18682), .C2(n18483), .A(n18403), .B(n18402), .ZN(
        P3_U2900) );
  AOI22_X1 U21464 ( .A1(n18685), .A2(n18434), .B1(n18683), .B2(n18417), .ZN(
        n18405) );
  AOI22_X1 U21465 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18419), .B1(
        n18647), .B2(n18487), .ZN(n18404) );
  OAI211_X1 U21466 ( .C1(n18650), .C2(n18414), .A(n18405), .B(n18404), .ZN(
        P3_U2901) );
  AOI22_X1 U21467 ( .A1(n18521), .A2(n18418), .B1(n18690), .B2(n18417), .ZN(
        n18407) );
  AOI22_X1 U21468 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18419), .B1(
        n18691), .B2(n18434), .ZN(n18406) );
  OAI211_X1 U21469 ( .C1(n18524), .C2(n18483), .A(n18407), .B(n18406), .ZN(
        P3_U2902) );
  AOI22_X1 U21470 ( .A1(n18621), .A2(n18418), .B1(n18696), .B2(n18417), .ZN(
        n18409) );
  AOI22_X1 U21471 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18419), .B1(
        n18697), .B2(n18434), .ZN(n18408) );
  OAI211_X1 U21472 ( .C1(n18624), .C2(n18483), .A(n18409), .B(n18408), .ZN(
        P3_U2903) );
  AOI22_X1 U21473 ( .A1(n18655), .A2(n18434), .B1(n18702), .B2(n18417), .ZN(
        n18411) );
  AOI22_X1 U21474 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18419), .B1(
        n18704), .B2(n18487), .ZN(n18410) );
  OAI211_X1 U21475 ( .C1(n18658), .C2(n18414), .A(n18411), .B(n18410), .ZN(
        P3_U2904) );
  AOI22_X1 U21476 ( .A1(n18709), .A2(n18434), .B1(n18708), .B2(n18417), .ZN(
        n18413) );
  AOI22_X1 U21477 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18419), .B1(
        n18710), .B2(n18487), .ZN(n18412) );
  OAI211_X1 U21478 ( .C1(n18713), .C2(n18414), .A(n18413), .B(n18412), .ZN(
        P3_U2905) );
  AOI22_X1 U21479 ( .A1(n18716), .A2(n18418), .B1(n18714), .B2(n18417), .ZN(
        n18416) );
  AOI22_X1 U21480 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18419), .B1(
        n18717), .B2(n18487), .ZN(n18415) );
  OAI211_X1 U21481 ( .C1(n18720), .C2(n18443), .A(n18416), .B(n18415), .ZN(
        P3_U2906) );
  AOI22_X1 U21482 ( .A1(n18609), .A2(n18418), .B1(n18723), .B2(n18417), .ZN(
        n18421) );
  AOI22_X1 U21483 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18419), .B1(
        n18726), .B2(n18487), .ZN(n18420) );
  OAI211_X1 U21484 ( .C1(n18613), .C2(n18443), .A(n18421), .B(n18420), .ZN(
        P3_U2907) );
  NAND2_X1 U21485 ( .A1(n18470), .A2(n18514), .ZN(n18508) );
  INV_X1 U21486 ( .A(n18470), .ZN(n18468) );
  NOR2_X1 U21487 ( .A1(n18468), .A2(n18515), .ZN(n18439) );
  AOI22_X1 U21488 ( .A1(n18674), .A2(n18434), .B1(n18673), .B2(n18439), .ZN(
        n18425) );
  AOI22_X1 U21489 ( .A1(n18678), .A2(n18423), .B1(n18470), .B2(n18422), .ZN(
        n18440) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18440), .B1(
        n18679), .B2(n18456), .ZN(n18424) );
  OAI211_X1 U21491 ( .C1(n18682), .C2(n18508), .A(n18425), .B(n18424), .ZN(
        P3_U2908) );
  AOI22_X1 U21492 ( .A1(n18685), .A2(n18456), .B1(n18683), .B2(n18439), .ZN(
        n18427) );
  AOI22_X1 U21493 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18440), .B1(
        n18684), .B2(n18434), .ZN(n18426) );
  OAI211_X1 U21494 ( .C1(n18688), .C2(n18508), .A(n18427), .B(n18426), .ZN(
        P3_U2909) );
  AOI22_X1 U21495 ( .A1(n18521), .A2(n18434), .B1(n18690), .B2(n18439), .ZN(
        n18429) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18440), .B1(
        n18691), .B2(n18456), .ZN(n18428) );
  OAI211_X1 U21497 ( .C1(n18524), .C2(n18508), .A(n18429), .B(n18428), .ZN(
        P3_U2910) );
  AOI22_X1 U21498 ( .A1(n18697), .A2(n18456), .B1(n18696), .B2(n18439), .ZN(
        n18431) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18440), .B1(
        n18621), .B2(n18434), .ZN(n18430) );
  OAI211_X1 U21500 ( .C1(n18624), .C2(n18508), .A(n18431), .B(n18430), .ZN(
        P3_U2911) );
  AOI22_X1 U21501 ( .A1(n18655), .A2(n18456), .B1(n18702), .B2(n18439), .ZN(
        n18433) );
  INV_X1 U21502 ( .A(n18508), .ZN(n18510) );
  AOI22_X1 U21503 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18440), .B1(
        n18704), .B2(n18510), .ZN(n18432) );
  OAI211_X1 U21504 ( .C1(n18658), .C2(n18443), .A(n18433), .B(n18432), .ZN(
        P3_U2912) );
  AOI22_X1 U21505 ( .A1(n18659), .A2(n18434), .B1(n18708), .B2(n18439), .ZN(
        n18436) );
  AOI22_X1 U21506 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18440), .B1(
        n18710), .B2(n18510), .ZN(n18435) );
  OAI211_X1 U21507 ( .C1(n18662), .C2(n18467), .A(n18436), .B(n18435), .ZN(
        P3_U2913) );
  AOI22_X1 U21508 ( .A1(n18602), .A2(n18456), .B1(n18714), .B2(n18439), .ZN(
        n18438) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18440), .B1(
        n18717), .B2(n18510), .ZN(n18437) );
  OAI211_X1 U21510 ( .C1(n18606), .C2(n18443), .A(n18438), .B(n18437), .ZN(
        P3_U2914) );
  AOI22_X1 U21511 ( .A1(n18724), .A2(n18456), .B1(n18723), .B2(n18439), .ZN(
        n18442) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18440), .B1(
        n18726), .B2(n18510), .ZN(n18441) );
  OAI211_X1 U21513 ( .C1(n18732), .C2(n18443), .A(n18442), .B(n18441), .ZN(
        P3_U2915) );
  NAND2_X1 U21514 ( .A1(n18470), .A2(n18539), .ZN(n18538) );
  NAND2_X1 U21515 ( .A1(n18467), .A2(n18483), .ZN(n18444) );
  NAND2_X1 U21516 ( .A1(n18508), .A2(n18538), .ZN(n18492) );
  AOI21_X1 U21517 ( .B1(n18641), .B2(n18444), .A(n18492), .ZN(n18446) );
  AOI211_X1 U21518 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(n18538), .A(n18446), 
        .B(n18445), .ZN(n18449) );
  AND2_X1 U21519 ( .A1(n18637), .A2(n18492), .ZN(n18463) );
  AOI22_X1 U21520 ( .A1(n18673), .A2(n18463), .B1(n18679), .B2(n18487), .ZN(
        n18448) );
  INV_X1 U21521 ( .A(n18538), .ZN(n18529) );
  AOI22_X1 U21522 ( .A1(n18674), .A2(n18456), .B1(n18643), .B2(n18529), .ZN(
        n18447) );
  OAI211_X1 U21523 ( .C1(n18449), .C2(n21100), .A(n18448), .B(n18447), .ZN(
        P3_U2916) );
  AOI22_X1 U21524 ( .A1(n18685), .A2(n18487), .B1(n18683), .B2(n18463), .ZN(
        n18451) );
  INV_X1 U21525 ( .A(n18449), .ZN(n18464) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18464), .B1(
        n18647), .B2(n18529), .ZN(n18450) );
  OAI211_X1 U21527 ( .C1(n18650), .C2(n18467), .A(n18451), .B(n18450), .ZN(
        P3_U2917) );
  AOI22_X1 U21528 ( .A1(n18691), .A2(n18487), .B1(n18690), .B2(n18463), .ZN(
        n18453) );
  AOI22_X1 U21529 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18464), .B1(
        n18692), .B2(n18529), .ZN(n18452) );
  OAI211_X1 U21530 ( .C1(n18695), .C2(n18467), .A(n18453), .B(n18452), .ZN(
        P3_U2918) );
  AOI22_X1 U21531 ( .A1(n18621), .A2(n18456), .B1(n18696), .B2(n18463), .ZN(
        n18455) );
  AOI22_X1 U21532 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18464), .B1(
        n18697), .B2(n18487), .ZN(n18454) );
  OAI211_X1 U21533 ( .C1(n18624), .C2(n18538), .A(n18455), .B(n18454), .ZN(
        P3_U2919) );
  INV_X1 U21534 ( .A(n18658), .ZN(n18703) );
  AOI22_X1 U21535 ( .A1(n18703), .A2(n18456), .B1(n18702), .B2(n18463), .ZN(
        n18458) );
  AOI22_X1 U21536 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18464), .B1(
        n18704), .B2(n18529), .ZN(n18457) );
  OAI211_X1 U21537 ( .C1(n18707), .C2(n18483), .A(n18458), .B(n18457), .ZN(
        P3_U2920) );
  AOI22_X1 U21538 ( .A1(n18709), .A2(n18487), .B1(n18708), .B2(n18463), .ZN(
        n18460) );
  AOI22_X1 U21539 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18464), .B1(
        n18710), .B2(n18529), .ZN(n18459) );
  OAI211_X1 U21540 ( .C1(n18713), .C2(n18467), .A(n18460), .B(n18459), .ZN(
        P3_U2921) );
  AOI22_X1 U21541 ( .A1(n18602), .A2(n18487), .B1(n18714), .B2(n18463), .ZN(
        n18462) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18464), .B1(
        n18717), .B2(n18529), .ZN(n18461) );
  OAI211_X1 U21543 ( .C1(n18606), .C2(n18467), .A(n18462), .B(n18461), .ZN(
        P3_U2922) );
  AOI22_X1 U21544 ( .A1(n18724), .A2(n18487), .B1(n18723), .B2(n18463), .ZN(
        n18466) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18464), .B1(
        n18726), .B2(n18529), .ZN(n18465) );
  OAI211_X1 U21546 ( .C1(n18732), .C2(n18467), .A(n18466), .B(n18465), .ZN(
        P3_U2923) );
  NOR2_X1 U21547 ( .A1(n18754), .A2(n18468), .ZN(n18516) );
  AND2_X1 U21548 ( .A1(n18637), .A2(n18516), .ZN(n18486) );
  AOI22_X1 U21549 ( .A1(n18673), .A2(n18486), .B1(n18679), .B2(n18510), .ZN(
        n18472) );
  NAND2_X1 U21550 ( .A1(n18470), .A2(n18469), .ZN(n18488) );
  NAND2_X1 U21551 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18516), .ZN(
        n18562) );
  AOI22_X1 U21552 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18488), .B1(
        n18643), .B2(n18553), .ZN(n18471) );
  OAI211_X1 U21553 ( .C1(n18646), .C2(n18483), .A(n18472), .B(n18471), .ZN(
        P3_U2924) );
  AOI22_X1 U21554 ( .A1(n18684), .A2(n18487), .B1(n18683), .B2(n18486), .ZN(
        n18474) );
  AOI22_X1 U21555 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18488), .B1(
        n18685), .B2(n18510), .ZN(n18473) );
  OAI211_X1 U21556 ( .C1(n18688), .C2(n18562), .A(n18474), .B(n18473), .ZN(
        P3_U2925) );
  AOI22_X1 U21557 ( .A1(n18691), .A2(n18510), .B1(n18690), .B2(n18486), .ZN(
        n18476) );
  AOI22_X1 U21558 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18488), .B1(
        n18692), .B2(n18553), .ZN(n18475) );
  OAI211_X1 U21559 ( .C1(n18695), .C2(n18483), .A(n18476), .B(n18475), .ZN(
        P3_U2926) );
  AOI22_X1 U21560 ( .A1(n18621), .A2(n18487), .B1(n18696), .B2(n18486), .ZN(
        n18478) );
  AOI22_X1 U21561 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18488), .B1(
        n18697), .B2(n18510), .ZN(n18477) );
  OAI211_X1 U21562 ( .C1(n18624), .C2(n18562), .A(n18478), .B(n18477), .ZN(
        P3_U2927) );
  AOI22_X1 U21563 ( .A1(n18655), .A2(n18510), .B1(n18702), .B2(n18486), .ZN(
        n18480) );
  AOI22_X1 U21564 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18488), .B1(
        n18704), .B2(n18553), .ZN(n18479) );
  OAI211_X1 U21565 ( .C1(n18658), .C2(n18483), .A(n18480), .B(n18479), .ZN(
        P3_U2928) );
  AOI22_X1 U21566 ( .A1(n18709), .A2(n18510), .B1(n18708), .B2(n18486), .ZN(
        n18482) );
  AOI22_X1 U21567 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18488), .B1(
        n18710), .B2(n18553), .ZN(n18481) );
  OAI211_X1 U21568 ( .C1(n18713), .C2(n18483), .A(n18482), .B(n18481), .ZN(
        P3_U2929) );
  AOI22_X1 U21569 ( .A1(n18716), .A2(n18487), .B1(n18714), .B2(n18486), .ZN(
        n18485) );
  AOI22_X1 U21570 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18488), .B1(
        n18717), .B2(n18553), .ZN(n18484) );
  OAI211_X1 U21571 ( .C1(n18720), .C2(n18508), .A(n18485), .B(n18484), .ZN(
        P3_U2930) );
  AOI22_X1 U21572 ( .A1(n18609), .A2(n18487), .B1(n18723), .B2(n18486), .ZN(
        n18490) );
  AOI22_X1 U21573 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18488), .B1(
        n18726), .B2(n18553), .ZN(n18489) );
  OAI211_X1 U21574 ( .C1(n18613), .C2(n18508), .A(n18490), .B(n18489), .ZN(
        P3_U2931) );
  NAND2_X1 U21575 ( .A1(n18491), .A2(n18585), .ZN(n18579) );
  INV_X1 U21576 ( .A(n18579), .ZN(n18581) );
  NOR2_X1 U21577 ( .A1(n18553), .A2(n18581), .ZN(n18541) );
  NOR2_X1 U21578 ( .A1(n18794), .A2(n18541), .ZN(n18509) );
  AOI22_X1 U21579 ( .A1(n18673), .A2(n18509), .B1(n18679), .B2(n18529), .ZN(
        n18495) );
  INV_X1 U21580 ( .A(n18541), .ZN(n18493) );
  OAI221_X1 U21581 ( .B1(n18493), .B2(n18641), .C1(n18493), .C2(n18492), .A(
        n18639), .ZN(n18511) );
  AOI22_X1 U21582 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18511), .B1(
        n18674), .B2(n18510), .ZN(n18494) );
  OAI211_X1 U21583 ( .C1(n18682), .C2(n18579), .A(n18495), .B(n18494), .ZN(
        P3_U2932) );
  AOI22_X1 U21584 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18511), .B1(
        n18683), .B2(n18509), .ZN(n18497) );
  AOI22_X1 U21585 ( .A1(n18647), .A2(n18581), .B1(n18685), .B2(n18529), .ZN(
        n18496) );
  OAI211_X1 U21586 ( .C1(n18650), .C2(n18508), .A(n18497), .B(n18496), .ZN(
        P3_U2933) );
  AOI22_X1 U21587 ( .A1(n18691), .A2(n18529), .B1(n18690), .B2(n18509), .ZN(
        n18499) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18511), .B1(
        n18692), .B2(n18581), .ZN(n18498) );
  OAI211_X1 U21589 ( .C1(n18695), .C2(n18508), .A(n18499), .B(n18498), .ZN(
        P3_U2934) );
  AOI22_X1 U21590 ( .A1(n18621), .A2(n18510), .B1(n18696), .B2(n18509), .ZN(
        n18501) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18511), .B1(
        n18697), .B2(n18529), .ZN(n18500) );
  OAI211_X1 U21592 ( .C1(n18624), .C2(n18579), .A(n18501), .B(n18500), .ZN(
        P3_U2935) );
  AOI22_X1 U21593 ( .A1(n18703), .A2(n18510), .B1(n18702), .B2(n18509), .ZN(
        n18503) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18511), .B1(
        n18704), .B2(n18581), .ZN(n18502) );
  OAI211_X1 U21595 ( .C1(n18707), .C2(n18538), .A(n18503), .B(n18502), .ZN(
        P3_U2936) );
  AOI22_X1 U21596 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18511), .B1(
        n18708), .B2(n18509), .ZN(n18505) );
  AOI22_X1 U21597 ( .A1(n18710), .A2(n18581), .B1(n18659), .B2(n18510), .ZN(
        n18504) );
  OAI211_X1 U21598 ( .C1(n18662), .C2(n18538), .A(n18505), .B(n18504), .ZN(
        P3_U2937) );
  AOI22_X1 U21599 ( .A1(n18602), .A2(n18529), .B1(n18714), .B2(n18509), .ZN(
        n18507) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18511), .B1(
        n18717), .B2(n18581), .ZN(n18506) );
  OAI211_X1 U21601 ( .C1(n18606), .C2(n18508), .A(n18507), .B(n18506), .ZN(
        P3_U2938) );
  AOI22_X1 U21602 ( .A1(n18609), .A2(n18510), .B1(n18723), .B2(n18509), .ZN(
        n18513) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18511), .B1(
        n18726), .B2(n18581), .ZN(n18512) );
  OAI211_X1 U21604 ( .C1(n18613), .C2(n18538), .A(n18513), .B(n18512), .ZN(
        P3_U2939) );
  NAND2_X1 U21605 ( .A1(n18585), .A2(n18514), .ZN(n18605) );
  INV_X1 U21606 ( .A(n18585), .ZN(n18563) );
  NOR2_X1 U21607 ( .A1(n18563), .A2(n18515), .ZN(n18534) );
  AOI22_X1 U21608 ( .A1(n18674), .A2(n18529), .B1(n18673), .B2(n18534), .ZN(
        n18518) );
  NOR2_X1 U21609 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18563), .ZN(
        n18564) );
  AOI22_X1 U21610 ( .A1(n18678), .A2(n18516), .B1(n18675), .B2(n18564), .ZN(
        n18535) );
  AOI22_X1 U21611 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18535), .B1(
        n18679), .B2(n18553), .ZN(n18517) );
  OAI211_X1 U21612 ( .C1(n18682), .C2(n18605), .A(n18518), .B(n18517), .ZN(
        P3_U2940) );
  AOI22_X1 U21613 ( .A1(n18684), .A2(n18529), .B1(n18683), .B2(n18534), .ZN(
        n18520) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18535), .B1(
        n18685), .B2(n18553), .ZN(n18519) );
  OAI211_X1 U21615 ( .C1(n18688), .C2(n18605), .A(n18520), .B(n18519), .ZN(
        P3_U2941) );
  AOI22_X1 U21616 ( .A1(n18521), .A2(n18529), .B1(n18690), .B2(n18534), .ZN(
        n18523) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18535), .B1(
        n18691), .B2(n18553), .ZN(n18522) );
  OAI211_X1 U21618 ( .C1(n18524), .C2(n18605), .A(n18523), .B(n18522), .ZN(
        P3_U2942) );
  AOI22_X1 U21619 ( .A1(n18621), .A2(n18529), .B1(n18696), .B2(n18534), .ZN(
        n18526) );
  AOI22_X1 U21620 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18535), .B1(
        n18697), .B2(n18553), .ZN(n18525) );
  OAI211_X1 U21621 ( .C1(n18624), .C2(n18605), .A(n18526), .B(n18525), .ZN(
        P3_U2943) );
  AOI22_X1 U21622 ( .A1(n18703), .A2(n18529), .B1(n18702), .B2(n18534), .ZN(
        n18528) );
  INV_X1 U21623 ( .A(n18605), .ZN(n18608) );
  AOI22_X1 U21624 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18535), .B1(
        n18704), .B2(n18608), .ZN(n18527) );
  OAI211_X1 U21625 ( .C1(n18707), .C2(n18562), .A(n18528), .B(n18527), .ZN(
        P3_U2944) );
  AOI22_X1 U21626 ( .A1(n18659), .A2(n18529), .B1(n18708), .B2(n18534), .ZN(
        n18531) );
  AOI22_X1 U21627 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18535), .B1(
        n18710), .B2(n18608), .ZN(n18530) );
  OAI211_X1 U21628 ( .C1(n18662), .C2(n18562), .A(n18531), .B(n18530), .ZN(
        P3_U2945) );
  AOI22_X1 U21629 ( .A1(n18602), .A2(n18553), .B1(n18714), .B2(n18534), .ZN(
        n18533) );
  AOI22_X1 U21630 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18535), .B1(
        n18717), .B2(n18608), .ZN(n18532) );
  OAI211_X1 U21631 ( .C1(n18606), .C2(n18538), .A(n18533), .B(n18532), .ZN(
        P3_U2946) );
  AOI22_X1 U21632 ( .A1(n18724), .A2(n18553), .B1(n18723), .B2(n18534), .ZN(
        n18537) );
  AOI22_X1 U21633 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18535), .B1(
        n18726), .B2(n18608), .ZN(n18536) );
  OAI211_X1 U21634 ( .C1(n18732), .C2(n18538), .A(n18537), .B(n18536), .ZN(
        P3_U2947) );
  NAND2_X1 U21635 ( .A1(n18585), .A2(n18539), .ZN(n18636) );
  AOI21_X1 U21636 ( .B1(n18605), .B2(n18636), .A(n18794), .ZN(n18558) );
  AOI22_X1 U21637 ( .A1(n18674), .A2(n18553), .B1(n18673), .B2(n18558), .ZN(
        n18544) );
  INV_X1 U21638 ( .A(n18636), .ZN(n18629) );
  OAI211_X1 U21639 ( .C1(n18541), .C2(n18540), .A(n18605), .B(n18636), .ZN(
        n18542) );
  OAI211_X1 U21640 ( .C1(n18629), .C2(n18887), .A(n18589), .B(n18542), .ZN(
        n18559) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18559), .B1(
        n18679), .B2(n18581), .ZN(n18543) );
  OAI211_X1 U21642 ( .C1(n18682), .C2(n18636), .A(n18544), .B(n18543), .ZN(
        P3_U2948) );
  AOI22_X1 U21643 ( .A1(n18685), .A2(n18581), .B1(n18683), .B2(n18558), .ZN(
        n18546) );
  AOI22_X1 U21644 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18559), .B1(
        n18647), .B2(n18629), .ZN(n18545) );
  OAI211_X1 U21645 ( .C1(n18650), .C2(n18562), .A(n18546), .B(n18545), .ZN(
        P3_U2949) );
  AOI22_X1 U21646 ( .A1(n18691), .A2(n18581), .B1(n18690), .B2(n18558), .ZN(
        n18548) );
  AOI22_X1 U21647 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18559), .B1(
        n18692), .B2(n18629), .ZN(n18547) );
  OAI211_X1 U21648 ( .C1(n18695), .C2(n18562), .A(n18548), .B(n18547), .ZN(
        P3_U2950) );
  AOI22_X1 U21649 ( .A1(n18621), .A2(n18553), .B1(n18696), .B2(n18558), .ZN(
        n18550) );
  AOI22_X1 U21650 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18559), .B1(
        n18697), .B2(n18581), .ZN(n18549) );
  OAI211_X1 U21651 ( .C1(n18624), .C2(n18636), .A(n18550), .B(n18549), .ZN(
        P3_U2951) );
  AOI22_X1 U21652 ( .A1(n18655), .A2(n18581), .B1(n18702), .B2(n18558), .ZN(
        n18552) );
  AOI22_X1 U21653 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18559), .B1(
        n18704), .B2(n18629), .ZN(n18551) );
  OAI211_X1 U21654 ( .C1(n18658), .C2(n18562), .A(n18552), .B(n18551), .ZN(
        P3_U2952) );
  AOI22_X1 U21655 ( .A1(n18659), .A2(n18553), .B1(n18708), .B2(n18558), .ZN(
        n18555) );
  AOI22_X1 U21656 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18559), .B1(
        n18710), .B2(n18629), .ZN(n18554) );
  OAI211_X1 U21657 ( .C1(n18662), .C2(n18579), .A(n18555), .B(n18554), .ZN(
        P3_U2953) );
  AOI22_X1 U21658 ( .A1(n18602), .A2(n18581), .B1(n18714), .B2(n18558), .ZN(
        n18557) );
  AOI22_X1 U21659 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18559), .B1(
        n18717), .B2(n18629), .ZN(n18556) );
  OAI211_X1 U21660 ( .C1(n18606), .C2(n18562), .A(n18557), .B(n18556), .ZN(
        P3_U2954) );
  AOI22_X1 U21661 ( .A1(n18724), .A2(n18581), .B1(n18723), .B2(n18558), .ZN(
        n18561) );
  AOI22_X1 U21662 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18559), .B1(
        n18726), .B2(n18629), .ZN(n18560) );
  OAI211_X1 U21663 ( .C1(n18732), .C2(n18562), .A(n18561), .B(n18560), .ZN(
        P3_U2955) );
  NOR2_X1 U21664 ( .A1(n18754), .A2(n18563), .ZN(n18614) );
  AND2_X1 U21665 ( .A1(n18637), .A2(n18614), .ZN(n18580) );
  AOI22_X1 U21666 ( .A1(n18673), .A2(n18580), .B1(n18679), .B2(n18608), .ZN(
        n18566) );
  AOI22_X1 U21667 ( .A1(n18678), .A2(n18564), .B1(n18675), .B2(n18614), .ZN(
        n18582) );
  NAND2_X1 U21668 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18614), .ZN(
        n18671) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18582), .B1(
        n18643), .B2(n18663), .ZN(n18565) );
  OAI211_X1 U21670 ( .C1(n18646), .C2(n18579), .A(n18566), .B(n18565), .ZN(
        P3_U2956) );
  AOI22_X1 U21671 ( .A1(n18685), .A2(n18608), .B1(n18683), .B2(n18580), .ZN(
        n18568) );
  AOI22_X1 U21672 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18582), .B1(
        n18647), .B2(n18663), .ZN(n18567) );
  OAI211_X1 U21673 ( .C1(n18650), .C2(n18579), .A(n18568), .B(n18567), .ZN(
        P3_U2957) );
  AOI22_X1 U21674 ( .A1(n18691), .A2(n18608), .B1(n18690), .B2(n18580), .ZN(
        n18570) );
  AOI22_X1 U21675 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18582), .B1(
        n18692), .B2(n18663), .ZN(n18569) );
  OAI211_X1 U21676 ( .C1(n18695), .C2(n18579), .A(n18570), .B(n18569), .ZN(
        P3_U2958) );
  AOI22_X1 U21677 ( .A1(n18697), .A2(n18608), .B1(n18696), .B2(n18580), .ZN(
        n18572) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18582), .B1(
        n18698), .B2(n18663), .ZN(n18571) );
  OAI211_X1 U21679 ( .C1(n18701), .C2(n18579), .A(n18572), .B(n18571), .ZN(
        P3_U2959) );
  AOI22_X1 U21680 ( .A1(n18703), .A2(n18581), .B1(n18702), .B2(n18580), .ZN(
        n18574) );
  AOI22_X1 U21681 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18582), .B1(
        n18704), .B2(n18663), .ZN(n18573) );
  OAI211_X1 U21682 ( .C1(n18707), .C2(n18605), .A(n18574), .B(n18573), .ZN(
        P3_U2960) );
  AOI22_X1 U21683 ( .A1(n18659), .A2(n18581), .B1(n18708), .B2(n18580), .ZN(
        n18576) );
  AOI22_X1 U21684 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18582), .B1(
        n18710), .B2(n18663), .ZN(n18575) );
  OAI211_X1 U21685 ( .C1(n18662), .C2(n18605), .A(n18576), .B(n18575), .ZN(
        P3_U2961) );
  AOI22_X1 U21686 ( .A1(n18602), .A2(n18608), .B1(n18714), .B2(n18580), .ZN(
        n18578) );
  AOI22_X1 U21687 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18582), .B1(
        n18717), .B2(n18663), .ZN(n18577) );
  OAI211_X1 U21688 ( .C1(n18606), .C2(n18579), .A(n18578), .B(n18577), .ZN(
        P3_U2962) );
  AOI22_X1 U21689 ( .A1(n18609), .A2(n18581), .B1(n18723), .B2(n18580), .ZN(
        n18584) );
  AOI22_X1 U21690 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18582), .B1(
        n18726), .B2(n18663), .ZN(n18583) );
  OAI211_X1 U21691 ( .C1(n18613), .C2(n18605), .A(n18584), .B(n18583), .ZN(
        P3_U2963) );
  NAND2_X1 U21692 ( .A1(n18677), .A2(n18752), .ZN(n18731) );
  INV_X1 U21693 ( .A(n18731), .ZN(n18715) );
  NOR2_X1 U21694 ( .A1(n18663), .A2(n18715), .ZN(n18638) );
  NOR2_X1 U21695 ( .A1(n18794), .A2(n18638), .ZN(n18607) );
  AOI22_X1 U21696 ( .A1(n18673), .A2(n18607), .B1(n18679), .B2(n18629), .ZN(
        n18591) );
  NAND2_X1 U21697 ( .A1(n18641), .A2(n18585), .ZN(n18586) );
  OAI21_X1 U21698 ( .B1(n18587), .B2(n18586), .A(n18638), .ZN(n18588) );
  OAI211_X1 U21699 ( .C1(n18715), .C2(n18887), .A(n18589), .B(n18588), .ZN(
        n18610) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18610), .B1(
        n18674), .B2(n18608), .ZN(n18590) );
  OAI211_X1 U21701 ( .C1(n18682), .C2(n18731), .A(n18591), .B(n18590), .ZN(
        P3_U2964) );
  AOI22_X1 U21702 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18610), .B1(
        n18683), .B2(n18607), .ZN(n18593) );
  AOI22_X1 U21703 ( .A1(n18647), .A2(n18715), .B1(n18685), .B2(n18629), .ZN(
        n18592) );
  OAI211_X1 U21704 ( .C1(n18650), .C2(n18605), .A(n18593), .B(n18592), .ZN(
        P3_U2965) );
  AOI22_X1 U21705 ( .A1(n18691), .A2(n18629), .B1(n18690), .B2(n18607), .ZN(
        n18595) );
  AOI22_X1 U21706 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18610), .B1(
        n18692), .B2(n18715), .ZN(n18594) );
  OAI211_X1 U21707 ( .C1(n18695), .C2(n18605), .A(n18595), .B(n18594), .ZN(
        P3_U2966) );
  AOI22_X1 U21708 ( .A1(n18697), .A2(n18629), .B1(n18696), .B2(n18607), .ZN(
        n18597) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18610), .B1(
        n18698), .B2(n18715), .ZN(n18596) );
  OAI211_X1 U21710 ( .C1(n18701), .C2(n18605), .A(n18597), .B(n18596), .ZN(
        P3_U2967) );
  AOI22_X1 U21711 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18610), .B1(
        n18702), .B2(n18607), .ZN(n18599) );
  AOI22_X1 U21712 ( .A1(n18703), .A2(n18608), .B1(n18704), .B2(n18715), .ZN(
        n18598) );
  OAI211_X1 U21713 ( .C1(n18707), .C2(n18636), .A(n18599), .B(n18598), .ZN(
        P3_U2968) );
  AOI22_X1 U21714 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18610), .B1(
        n18708), .B2(n18607), .ZN(n18601) );
  AOI22_X1 U21715 ( .A1(n18710), .A2(n18715), .B1(n18659), .B2(n18608), .ZN(
        n18600) );
  OAI211_X1 U21716 ( .C1(n18662), .C2(n18636), .A(n18601), .B(n18600), .ZN(
        P3_U2969) );
  AOI22_X1 U21717 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18610), .B1(
        n18714), .B2(n18607), .ZN(n18604) );
  AOI22_X1 U21718 ( .A1(n18717), .A2(n18715), .B1(n18602), .B2(n18629), .ZN(
        n18603) );
  OAI211_X1 U21719 ( .C1(n18606), .C2(n18605), .A(n18604), .B(n18603), .ZN(
        P3_U2970) );
  AOI22_X1 U21720 ( .A1(n18609), .A2(n18608), .B1(n18723), .B2(n18607), .ZN(
        n18612) );
  AOI22_X1 U21721 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18610), .B1(
        n18726), .B2(n18715), .ZN(n18611) );
  OAI211_X1 U21722 ( .C1(n18613), .C2(n18636), .A(n18612), .B(n18611), .ZN(
        P3_U2971) );
  AND2_X1 U21723 ( .A1(n18637), .A2(n18677), .ZN(n18632) );
  AOI22_X1 U21724 ( .A1(n18673), .A2(n18632), .B1(n18679), .B2(n18663), .ZN(
        n18616) );
  AOI22_X1 U21725 ( .A1(n18678), .A2(n18614), .B1(n18677), .B2(n18675), .ZN(
        n18633) );
  AOI22_X1 U21726 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18633), .B1(
        n18725), .B2(n18643), .ZN(n18615) );
  OAI211_X1 U21727 ( .C1(n18646), .C2(n18636), .A(n18616), .B(n18615), .ZN(
        P3_U2972) );
  AOI22_X1 U21728 ( .A1(n18684), .A2(n18629), .B1(n18683), .B2(n18632), .ZN(
        n18618) );
  AOI22_X1 U21729 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18633), .B1(
        n18685), .B2(n18663), .ZN(n18617) );
  OAI211_X1 U21730 ( .C1(n18721), .C2(n18688), .A(n18618), .B(n18617), .ZN(
        P3_U2973) );
  AOI22_X1 U21731 ( .A1(n18691), .A2(n18663), .B1(n18690), .B2(n18632), .ZN(
        n18620) );
  AOI22_X1 U21732 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18633), .B1(
        n18725), .B2(n18692), .ZN(n18619) );
  OAI211_X1 U21733 ( .C1(n18695), .C2(n18636), .A(n18620), .B(n18619), .ZN(
        P3_U2974) );
  AOI22_X1 U21734 ( .A1(n18621), .A2(n18629), .B1(n18696), .B2(n18632), .ZN(
        n18623) );
  AOI22_X1 U21735 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18633), .B1(
        n18697), .B2(n18663), .ZN(n18622) );
  OAI211_X1 U21736 ( .C1(n18721), .C2(n18624), .A(n18623), .B(n18622), .ZN(
        P3_U2975) );
  AOI22_X1 U21737 ( .A1(n18703), .A2(n18629), .B1(n18702), .B2(n18632), .ZN(
        n18626) );
  AOI22_X1 U21738 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18633), .B1(
        n18725), .B2(n18704), .ZN(n18625) );
  OAI211_X1 U21739 ( .C1(n18707), .C2(n18671), .A(n18626), .B(n18625), .ZN(
        P3_U2976) );
  AOI22_X1 U21740 ( .A1(n18709), .A2(n18663), .B1(n18708), .B2(n18632), .ZN(
        n18628) );
  AOI22_X1 U21741 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18633), .B1(
        n18725), .B2(n18710), .ZN(n18627) );
  OAI211_X1 U21742 ( .C1(n18713), .C2(n18636), .A(n18628), .B(n18627), .ZN(
        P3_U2977) );
  AOI22_X1 U21743 ( .A1(n18716), .A2(n18629), .B1(n18714), .B2(n18632), .ZN(
        n18631) );
  AOI22_X1 U21744 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18633), .B1(
        n18725), .B2(n18717), .ZN(n18630) );
  OAI211_X1 U21745 ( .C1(n18720), .C2(n18671), .A(n18631), .B(n18630), .ZN(
        P3_U2978) );
  AOI22_X1 U21746 ( .A1(n18724), .A2(n18663), .B1(n18723), .B2(n18632), .ZN(
        n18635) );
  AOI22_X1 U21747 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18633), .B1(
        n18725), .B2(n18726), .ZN(n18634) );
  OAI211_X1 U21748 ( .C1(n18732), .C2(n18636), .A(n18635), .B(n18634), .ZN(
        P3_U2979) );
  AND2_X1 U21749 ( .A1(n18637), .A2(n18642), .ZN(n18667) );
  AOI22_X1 U21750 ( .A1(n18673), .A2(n18667), .B1(n18679), .B2(n18715), .ZN(
        n18645) );
  INV_X1 U21751 ( .A(n18638), .ZN(n18640) );
  OAI221_X1 U21752 ( .B1(n18642), .B2(n18641), .C1(n18642), .C2(n18640), .A(
        n18639), .ZN(n18668) );
  AOI22_X1 U21753 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18668), .B1(
        n18643), .B2(n18664), .ZN(n18644) );
  OAI211_X1 U21754 ( .C1(n18646), .C2(n18671), .A(n18645), .B(n18644), .ZN(
        P3_U2980) );
  AOI22_X1 U21755 ( .A1(n18685), .A2(n18715), .B1(n18683), .B2(n18667), .ZN(
        n18649) );
  AOI22_X1 U21756 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18668), .B1(
        n18664), .B2(n18647), .ZN(n18648) );
  OAI211_X1 U21757 ( .C1(n18650), .C2(n18671), .A(n18649), .B(n18648), .ZN(
        P3_U2981) );
  AOI22_X1 U21758 ( .A1(n18691), .A2(n18715), .B1(n18690), .B2(n18667), .ZN(
        n18652) );
  AOI22_X1 U21759 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18668), .B1(
        n18664), .B2(n18692), .ZN(n18651) );
  OAI211_X1 U21760 ( .C1(n18695), .C2(n18671), .A(n18652), .B(n18651), .ZN(
        P3_U2982) );
  AOI22_X1 U21761 ( .A1(n18697), .A2(n18715), .B1(n18696), .B2(n18667), .ZN(
        n18654) );
  AOI22_X1 U21762 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18668), .B1(
        n18664), .B2(n18698), .ZN(n18653) );
  OAI211_X1 U21763 ( .C1(n18701), .C2(n18671), .A(n18654), .B(n18653), .ZN(
        P3_U2983) );
  AOI22_X1 U21764 ( .A1(n18655), .A2(n18715), .B1(n18702), .B2(n18667), .ZN(
        n18657) );
  AOI22_X1 U21765 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18668), .B1(
        n18664), .B2(n18704), .ZN(n18656) );
  OAI211_X1 U21766 ( .C1(n18658), .C2(n18671), .A(n18657), .B(n18656), .ZN(
        P3_U2984) );
  AOI22_X1 U21767 ( .A1(n18659), .A2(n18663), .B1(n18708), .B2(n18667), .ZN(
        n18661) );
  AOI22_X1 U21768 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18668), .B1(
        n18664), .B2(n18710), .ZN(n18660) );
  OAI211_X1 U21769 ( .C1(n18662), .C2(n18731), .A(n18661), .B(n18660), .ZN(
        P3_U2985) );
  AOI22_X1 U21770 ( .A1(n18716), .A2(n18663), .B1(n18714), .B2(n18667), .ZN(
        n18666) );
  AOI22_X1 U21771 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18668), .B1(
        n18664), .B2(n18717), .ZN(n18665) );
  OAI211_X1 U21772 ( .C1(n18720), .C2(n18731), .A(n18666), .B(n18665), .ZN(
        P3_U2986) );
  AOI22_X1 U21773 ( .A1(n18724), .A2(n18715), .B1(n18723), .B2(n18667), .ZN(
        n18670) );
  AOI22_X1 U21774 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18668), .B1(
        n18664), .B2(n18726), .ZN(n18669) );
  OAI211_X1 U21775 ( .C1(n18732), .C2(n18671), .A(n18670), .B(n18669), .ZN(
        P3_U2987) );
  NOR2_X1 U21776 ( .A1(n18794), .A2(n18672), .ZN(n18722) );
  AOI22_X1 U21777 ( .A1(n18674), .A2(n18715), .B1(n18673), .B2(n18722), .ZN(
        n18681) );
  AOI22_X1 U21778 ( .A1(n18678), .A2(n18677), .B1(n18676), .B2(n18675), .ZN(
        n18728) );
  AOI22_X1 U21779 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18728), .B1(
        n18725), .B2(n18679), .ZN(n18680) );
  OAI211_X1 U21780 ( .C1(n18689), .C2(n18682), .A(n18681), .B(n18680), .ZN(
        P3_U2988) );
  AOI22_X1 U21781 ( .A1(n18684), .A2(n18715), .B1(n18683), .B2(n18722), .ZN(
        n18687) );
  AOI22_X1 U21782 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18728), .B1(
        n18725), .B2(n18685), .ZN(n18686) );
  OAI211_X1 U21783 ( .C1(n18689), .C2(n18688), .A(n18687), .B(n18686), .ZN(
        P3_U2989) );
  AOI22_X1 U21784 ( .A1(n18725), .A2(n18691), .B1(n18690), .B2(n18722), .ZN(
        n18694) );
  AOI22_X1 U21785 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18728), .B1(
        n18727), .B2(n18692), .ZN(n18693) );
  OAI211_X1 U21786 ( .C1(n18695), .C2(n18731), .A(n18694), .B(n18693), .ZN(
        P3_U2990) );
  AOI22_X1 U21787 ( .A1(n18725), .A2(n18697), .B1(n18696), .B2(n18722), .ZN(
        n18700) );
  AOI22_X1 U21788 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18728), .B1(
        n18727), .B2(n18698), .ZN(n18699) );
  OAI211_X1 U21789 ( .C1(n18701), .C2(n18731), .A(n18700), .B(n18699), .ZN(
        P3_U2991) );
  AOI22_X1 U21790 ( .A1(n18703), .A2(n18715), .B1(n18702), .B2(n18722), .ZN(
        n18706) );
  AOI22_X1 U21791 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18728), .B1(
        n18727), .B2(n18704), .ZN(n18705) );
  OAI211_X1 U21792 ( .C1(n18721), .C2(n18707), .A(n18706), .B(n18705), .ZN(
        P3_U2992) );
  AOI22_X1 U21793 ( .A1(n18725), .A2(n18709), .B1(n18708), .B2(n18722), .ZN(
        n18712) );
  AOI22_X1 U21794 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18728), .B1(
        n18727), .B2(n18710), .ZN(n18711) );
  OAI211_X1 U21795 ( .C1(n18713), .C2(n18731), .A(n18712), .B(n18711), .ZN(
        P3_U2993) );
  AOI22_X1 U21796 ( .A1(n18716), .A2(n18715), .B1(n18714), .B2(n18722), .ZN(
        n18719) );
  AOI22_X1 U21797 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18728), .B1(
        n18727), .B2(n18717), .ZN(n18718) );
  OAI211_X1 U21798 ( .C1(n18721), .C2(n18720), .A(n18719), .B(n18718), .ZN(
        P3_U2994) );
  AOI22_X1 U21799 ( .A1(n18725), .A2(n18724), .B1(n18723), .B2(n18722), .ZN(
        n18730) );
  AOI22_X1 U21800 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18728), .B1(
        n18727), .B2(n18726), .ZN(n18729) );
  OAI211_X1 U21801 ( .C1(n18732), .C2(n18731), .A(n18730), .B(n18729), .ZN(
        P3_U2995) );
  NOR3_X1 U21802 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18734), .A3(
        n18733), .ZN(n18743) );
  AOI211_X1 U21803 ( .C1(n18736), .C2(n18735), .A(n18743), .B(n20949), .ZN(
        n18741) );
  OAI21_X1 U21804 ( .B1(n9746), .B2(n18914), .A(n18749), .ZN(n18742) );
  AOI22_X1 U21805 ( .A1(n18738), .A2(n18742), .B1(n18768), .B2(n18740), .ZN(
        n18739) );
  AOI22_X1 U21806 ( .A1(n18741), .A2(n18740), .B1(n18739), .B2(n20949), .ZN(
        n18890) );
  INV_X1 U21807 ( .A(n18757), .ZN(n18779) );
  AOI22_X1 U21808 ( .A1(n18757), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n18890), .B2(n18779), .ZN(n18765) );
  INV_X1 U21809 ( .A(n18742), .ZN(n18750) );
  NOR3_X1 U21810 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18750), .A3(
        n18908), .ZN(n18747) );
  INV_X1 U21811 ( .A(n18743), .ZN(n18745) );
  AOI211_X1 U21812 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n18745), .A(
        n18744), .B(n18900), .ZN(n18746) );
  AOI211_X1 U21813 ( .C1(n18768), .C2(n18894), .A(n18747), .B(n18746), .ZN(
        n18897) );
  AOI22_X1 U21814 ( .A1(n18757), .A2(n18900), .B1(n18897), .B2(n18779), .ZN(
        n18760) );
  NOR2_X1 U21815 ( .A1(n18748), .A2(n9745), .ZN(n18751) );
  AOI22_X1 U21816 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18749), .B1(
        n18751), .B2(n18914), .ZN(n18910) );
  OAI22_X1 U21817 ( .A1(n18751), .A2(n18901), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18750), .ZN(n18906) );
  OR3_X1 U21818 ( .A1(n18910), .A2(n18754), .A3(n18752), .ZN(n18753) );
  AOI22_X1 U21819 ( .A1(n18910), .A2(n18754), .B1(n18906), .B2(n18753), .ZN(
        n18756) );
  OAI21_X1 U21820 ( .B1(n18757), .B2(n18756), .A(n18755), .ZN(n18759) );
  AND2_X1 U21821 ( .A1(n18760), .A2(n18759), .ZN(n18758) );
  OAI221_X1 U21822 ( .B1(n18760), .B2(n18759), .C1(n21008), .C2(n18758), .A(
        n18762), .ZN(n18764) );
  AOI21_X1 U21823 ( .B1(n18762), .B2(n18761), .A(n18760), .ZN(n18763) );
  AOI222_X1 U21824 ( .A1(n18765), .A2(n18764), .B1(n18765), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18764), .C2(n18763), .ZN(
        n18782) );
  INV_X1 U21825 ( .A(n18766), .ZN(n18774) );
  NOR2_X1 U21826 ( .A1(n18768), .A2(n18767), .ZN(n18770) );
  OAI222_X1 U21827 ( .A1(n18774), .A2(n18773), .B1(n18772), .B2(n18771), .C1(
        n18770), .C2(n18769), .ZN(n18926) );
  AOI221_X1 U21828 ( .B1(P3_MORE_REG_SCAN_IN), .B2(n18776), .C1(
        P3_FLUSH_REG_SCAN_IN), .C2(n18776), .A(n18775), .ZN(n18777) );
  OAI211_X1 U21829 ( .C1(n18780), .C2(n18779), .A(n18778), .B(n18777), .ZN(
        n18781) );
  NOR3_X1 U21830 ( .A1(n18782), .A2(n18926), .A3(n18781), .ZN(n18793) );
  AOI22_X1 U21831 ( .A1(n18909), .A2(n18938), .B1(n18933), .B2(n20824), .ZN(
        n18783) );
  INV_X1 U21832 ( .A(n18783), .ZN(n18788) );
  OAI211_X1 U21833 ( .C1(n18785), .C2(n18784), .A(n18930), .B(n18793), .ZN(
        n18886) );
  OAI21_X1 U21834 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18927), .A(n18886), 
        .ZN(n18795) );
  NOR2_X1 U21835 ( .A1(n18786), .A2(n18795), .ZN(n18787) );
  MUX2_X1 U21836 ( .A(n18788), .B(n18787), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18791) );
  INV_X1 U21837 ( .A(n18789), .ZN(n18790) );
  OAI211_X1 U21838 ( .C1(n18793), .C2(n18792), .A(n18791), .B(n18790), .ZN(
        P3_U2996) );
  NAND2_X1 U21839 ( .A1(n18933), .A2(n20824), .ZN(n18798) );
  NAND4_X1 U21840 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(n18933), .A4(n18945), .ZN(n18801) );
  OR3_X1 U21841 ( .A1(n18796), .A2(n18795), .A3(n18794), .ZN(n18797) );
  NAND4_X1 U21842 ( .A1(n18799), .A2(n18798), .A3(n18801), .A4(n18797), .ZN(
        P3_U2997) );
  OAI21_X1 U21843 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18800), .ZN(n18803) );
  INV_X1 U21844 ( .A(n18801), .ZN(n18802) );
  AOI21_X1 U21845 ( .B1(n18804), .B2(n18803), .A(n18802), .ZN(P3_U2998) );
  AND2_X1 U21846 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18882), .ZN(
        P3_U2999) );
  AND2_X1 U21847 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18882), .ZN(
        P3_U3000) );
  AND2_X1 U21848 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18882), .ZN(
        P3_U3001) );
  AND2_X1 U21849 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18882), .ZN(
        P3_U3002) );
  AND2_X1 U21850 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18882), .ZN(
        P3_U3003) );
  AND2_X1 U21851 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18882), .ZN(
        P3_U3004) );
  AND2_X1 U21852 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18882), .ZN(
        P3_U3005) );
  INV_X1 U21853 ( .A(P3_DATAWIDTH_REG_24__SCAN_IN), .ZN(n20850) );
  NOR2_X1 U21854 ( .A1(n20850), .A2(n18884), .ZN(P3_U3006) );
  NOR2_X1 U21855 ( .A1(n20978), .A2(n18884), .ZN(P3_U3007) );
  AND2_X1 U21856 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18882), .ZN(
        P3_U3008) );
  AND2_X1 U21857 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18882), .ZN(
        P3_U3009) );
  AND2_X1 U21858 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18882), .ZN(
        P3_U3010) );
  AND2_X1 U21859 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18882), .ZN(
        P3_U3011) );
  AND2_X1 U21860 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18882), .ZN(
        P3_U3012) );
  AND2_X1 U21861 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18882), .ZN(
        P3_U3013) );
  AND2_X1 U21862 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18882), .ZN(
        P3_U3014) );
  AND2_X1 U21863 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18882), .ZN(
        P3_U3015) );
  AND2_X1 U21864 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18882), .ZN(
        P3_U3016) );
  AND2_X1 U21865 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18882), .ZN(
        P3_U3017) );
  AND2_X1 U21866 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18882), .ZN(
        P3_U3018) );
  AND2_X1 U21867 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18882), .ZN(
        P3_U3019) );
  AND2_X1 U21868 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18882), .ZN(
        P3_U3020) );
  AND2_X1 U21869 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18882), .ZN(P3_U3021) );
  NOR2_X1 U21870 ( .A1(n20919), .A2(n18884), .ZN(P3_U3022) );
  AND2_X1 U21871 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18882), .ZN(P3_U3023) );
  AND2_X1 U21872 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18882), .ZN(P3_U3024) );
  AND2_X1 U21873 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18882), .ZN(P3_U3025) );
  AND2_X1 U21874 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18882), .ZN(P3_U3026) );
  AND2_X1 U21875 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18882), .ZN(P3_U3027) );
  AND2_X1 U21876 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18882), .ZN(P3_U3028) );
  OAI21_X1 U21877 ( .B1(n18805), .B2(n20719), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18806) );
  AOI22_X1 U21878 ( .A1(n18818), .A2(n18820), .B1(n18943), .B2(n18806), .ZN(
        n18807) );
  NAND3_X1 U21879 ( .A1(NA), .A2(n18818), .A3(n18809), .ZN(n18812) );
  OAI211_X1 U21880 ( .C1(n18927), .C2(n18808), .A(n18807), .B(n18812), .ZN(
        P3_U3029) );
  INV_X1 U21881 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18940) );
  NOR2_X1 U21882 ( .A1(n18820), .A2(n20719), .ZN(n18816) );
  OAI22_X1 U21883 ( .A1(n18940), .A2(n18816), .B1(n20719), .B2(n18808), .ZN(
        n18810) );
  NOR2_X1 U21884 ( .A1(n18927), .A2(n18809), .ZN(n18813) );
  AOI211_X1 U21885 ( .C1(n18810), .C2(P3_STATE_REG_0__SCAN_IN), .A(n18813), 
        .B(n18931), .ZN(n18811) );
  INV_X1 U21886 ( .A(n18811), .ZN(P3_U3030) );
  AOI21_X1 U21887 ( .B1(n18818), .B2(n18812), .A(n18813), .ZN(n18819) );
  INV_X1 U21888 ( .A(n18813), .ZN(n18814) );
  OAI22_X1 U21889 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18814), .ZN(n18815) );
  OAI22_X1 U21890 ( .A1(n18816), .A2(n18815), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18817) );
  OAI22_X1 U21891 ( .A1(n18819), .A2(n18820), .B1(n18818), .B2(n18817), .ZN(
        P3_U3031) );
  INV_X1 U21892 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18822) );
  INV_X1 U21893 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18823) );
  NAND2_X1 U21894 ( .A1(n18942), .A2(n18820), .ZN(n18864) );
  CLKBUF_X1 U21895 ( .A(n18864), .Z(n18873) );
  OAI222_X1 U21896 ( .A1(n18822), .A2(n18876), .B1(n18821), .B2(n18942), .C1(
        n18823), .C2(n18873), .ZN(P3_U3032) );
  OAI222_X1 U21897 ( .A1(n18873), .A2(n18825), .B1(n18824), .B2(n18942), .C1(
        n18823), .C2(n18876), .ZN(P3_U3033) );
  OAI222_X1 U21898 ( .A1(n18864), .A2(n18827), .B1(n18826), .B2(n18942), .C1(
        n18825), .C2(n18876), .ZN(P3_U3034) );
  OAI222_X1 U21899 ( .A1(n18864), .A2(n18829), .B1(n18828), .B2(n18942), .C1(
        n18827), .C2(n18876), .ZN(P3_U3035) );
  OAI222_X1 U21900 ( .A1(n18864), .A2(n20920), .B1(n18830), .B2(n18942), .C1(
        n18829), .C2(n18876), .ZN(P3_U3036) );
  OAI222_X1 U21901 ( .A1(n18864), .A2(n18832), .B1(n18831), .B2(n18942), .C1(
        n20920), .C2(n18876), .ZN(P3_U3037) );
  INV_X1 U21902 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18835) );
  OAI222_X1 U21903 ( .A1(n18864), .A2(n18835), .B1(n18833), .B2(n18942), .C1(
        n18832), .C2(n18876), .ZN(P3_U3038) );
  OAI222_X1 U21904 ( .A1(n18835), .A2(n18876), .B1(n18834), .B2(n18942), .C1(
        n18836), .C2(n18873), .ZN(P3_U3039) );
  OAI222_X1 U21905 ( .A1(n18873), .A2(n18838), .B1(n18837), .B2(n18942), .C1(
        n18836), .C2(n18876), .ZN(P3_U3040) );
  OAI222_X1 U21906 ( .A1(n18873), .A2(n18840), .B1(n18839), .B2(n18942), .C1(
        n18838), .C2(n18876), .ZN(P3_U3041) );
  INV_X1 U21907 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18842) );
  OAI222_X1 U21908 ( .A1(n18873), .A2(n18842), .B1(n18841), .B2(n18942), .C1(
        n18840), .C2(n18876), .ZN(P3_U3042) );
  OAI222_X1 U21909 ( .A1(n18873), .A2(n18844), .B1(n18843), .B2(n18942), .C1(
        n18842), .C2(n18876), .ZN(P3_U3043) );
  OAI222_X1 U21910 ( .A1(n18873), .A2(n18847), .B1(n18845), .B2(n18942), .C1(
        n18844), .C2(n18876), .ZN(P3_U3044) );
  OAI222_X1 U21911 ( .A1(n18847), .A2(n18876), .B1(n18846), .B2(n18942), .C1(
        n18848), .C2(n18873), .ZN(P3_U3045) );
  OAI222_X1 U21912 ( .A1(n18873), .A2(n18850), .B1(n18849), .B2(n18942), .C1(
        n18848), .C2(n18876), .ZN(P3_U3046) );
  OAI222_X1 U21913 ( .A1(n18864), .A2(n18852), .B1(n18851), .B2(n18942), .C1(
        n18850), .C2(n18876), .ZN(P3_U3047) );
  OAI222_X1 U21914 ( .A1(n18864), .A2(n18854), .B1(n18853), .B2(n18942), .C1(
        n18852), .C2(n18876), .ZN(P3_U3048) );
  OAI222_X1 U21915 ( .A1(n18864), .A2(n20997), .B1(n20829), .B2(n18942), .C1(
        n18854), .C2(n18876), .ZN(P3_U3049) );
  OAI222_X1 U21916 ( .A1(n18864), .A2(n18856), .B1(n18855), .B2(n18942), .C1(
        n20997), .C2(n18876), .ZN(P3_U3050) );
  OAI222_X1 U21917 ( .A1(n18864), .A2(n21058), .B1(n18857), .B2(n18942), .C1(
        n18856), .C2(n18876), .ZN(P3_U3051) );
  INV_X1 U21918 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20974) );
  OAI222_X1 U21919 ( .A1(n18864), .A2(n20974), .B1(n18858), .B2(n18942), .C1(
        n21058), .C2(n18876), .ZN(P3_U3052) );
  OAI222_X1 U21920 ( .A1(n18873), .A2(n18860), .B1(n18859), .B2(n18942), .C1(
        n20974), .C2(n18876), .ZN(P3_U3053) );
  OAI222_X1 U21921 ( .A1(n18873), .A2(n18862), .B1(n18861), .B2(n18942), .C1(
        n18860), .C2(n18876), .ZN(P3_U3054) );
  OAI222_X1 U21922 ( .A1(n18864), .A2(n18865), .B1(n18863), .B2(n18942), .C1(
        n18862), .C2(n18876), .ZN(P3_U3055) );
  OAI222_X1 U21923 ( .A1(n18873), .A2(n18867), .B1(n18866), .B2(n18942), .C1(
        n18865), .C2(n18876), .ZN(P3_U3056) );
  INV_X1 U21924 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18869) );
  OAI222_X1 U21925 ( .A1(n18873), .A2(n18869), .B1(n18868), .B2(n18942), .C1(
        n18867), .C2(n18876), .ZN(P3_U3057) );
  INV_X1 U21926 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18870) );
  OAI222_X1 U21927 ( .A1(n18873), .A2(n18870), .B1(n20902), .B2(n18942), .C1(
        n18869), .C2(n18876), .ZN(P3_U3058) );
  INV_X1 U21928 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18871) );
  OAI222_X1 U21929 ( .A1(n18873), .A2(n18871), .B1(n20933), .B2(n18942), .C1(
        n18870), .C2(n18876), .ZN(P3_U3059) );
  OAI222_X1 U21930 ( .A1(n18873), .A2(n18875), .B1(n18872), .B2(n18942), .C1(
        n18871), .C2(n18876), .ZN(P3_U3060) );
  OAI222_X1 U21931 ( .A1(n18876), .A2(n18875), .B1(n21036), .B2(n18942), .C1(
        n18874), .C2(n18873), .ZN(P3_U3061) );
  MUX2_X1 U21932 ( .A(P3_BE_N_REG_3__SCAN_IN), .B(P3_BYTEENABLE_REG_3__SCAN_IN), .S(n18942), .Z(P3_U3274) );
  INV_X1 U21933 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20975) );
  INV_X1 U21934 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18877) );
  AOI22_X1 U21935 ( .A1(n18942), .A2(n20975), .B1(n18877), .B2(n18943), .ZN(
        P3_U3275) );
  INV_X1 U21936 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18878) );
  AOI22_X1 U21937 ( .A1(n18942), .A2(n18879), .B1(n18878), .B2(n18943), .ZN(
        P3_U3276) );
  INV_X1 U21938 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18920) );
  INV_X1 U21939 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18880) );
  AOI22_X1 U21940 ( .A1(n18942), .A2(n18920), .B1(n18880), .B2(n18943), .ZN(
        P3_U3277) );
  INV_X1 U21941 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18916) );
  INV_X1 U21942 ( .A(n18883), .ZN(n18881) );
  AOI21_X1 U21943 ( .B1(n18882), .B2(n18916), .A(n18881), .ZN(P3_U3280) );
  OAI21_X1 U21944 ( .B1(n18884), .B2(n20995), .A(n18883), .ZN(P3_U3281) );
  OAI221_X1 U21945 ( .B1(n18887), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18887), 
        .C2(n18886), .A(n18885), .ZN(P3_U3282) );
  INV_X1 U21946 ( .A(n18888), .ZN(n18889) );
  AOI22_X1 U21947 ( .A1(n18946), .A2(n18890), .B1(n18909), .B2(n18889), .ZN(
        n18891) );
  AOI22_X1 U21948 ( .A1(n18915), .A2(n20949), .B1(n18891), .B2(n18912), .ZN(
        P3_U3285) );
  AOI22_X1 U21949 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n10060), .B2(n18892), .ZN(
        n18902) );
  NOR2_X1 U21950 ( .A1(n18893), .A2(n18911), .ZN(n18903) );
  INV_X1 U21951 ( .A(n18909), .ZN(n18895) );
  OAI22_X1 U21952 ( .A1(n18897), .A2(n18896), .B1(n18895), .B2(n18894), .ZN(
        n18898) );
  AOI21_X1 U21953 ( .B1(n18902), .B2(n18903), .A(n18898), .ZN(n18899) );
  AOI22_X1 U21954 ( .A1(n18915), .A2(n18900), .B1(n18899), .B2(n18912), .ZN(
        P3_U3288) );
  INV_X1 U21955 ( .A(n18901), .ZN(n18905) );
  INV_X1 U21956 ( .A(n18902), .ZN(n18904) );
  AOI222_X1 U21957 ( .A1(n18906), .A2(n18946), .B1(n18909), .B2(n18905), .C1(
        n18904), .C2(n18903), .ZN(n18907) );
  AOI22_X1 U21958 ( .A1(n18915), .A2(n18908), .B1(n18907), .B2(n18912), .ZN(
        P3_U3289) );
  AOI222_X1 U21959 ( .A1(n18911), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18946), 
        .B2(n18910), .C1(n18914), .C2(n18909), .ZN(n18913) );
  AOI22_X1 U21960 ( .A1(n18915), .A2(n18914), .B1(n18913), .B2(n18912), .ZN(
        P3_U3290) );
  OAI211_X1 U21961 ( .C1(n18916), .C2(n18922), .A(n20995), .B(n18923), .ZN(
        n18919) );
  NOR2_X1 U21962 ( .A1(n18921), .A2(n18922), .ZN(n18917) );
  AOI22_X1 U21963 ( .A1(P3_BYTEENABLE_REG_2__SCAN_IN), .A2(n18921), .B1(
        P3_REIP_REG_1__SCAN_IN), .B2(n18917), .ZN(n18918) );
  NAND2_X1 U21964 ( .A1(n18919), .A2(n18918), .ZN(P3_U3292) );
  AOI22_X1 U21965 ( .A1(n18923), .A2(n18922), .B1(n18921), .B2(n18920), .ZN(
        P3_U3293) );
  INV_X1 U21966 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18924) );
  AOI22_X1 U21967 ( .A1(n18942), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18924), 
        .B2(n18943), .ZN(P3_U3294) );
  MUX2_X1 U21968 ( .A(P3_MORE_REG_SCAN_IN), .B(n18926), .S(n18925), .Z(
        P3_U3295) );
  AOI21_X1 U21969 ( .B1(n20824), .B2(n18927), .A(n18948), .ZN(n18928) );
  OAI21_X1 U21970 ( .B1(n18930), .B2(n18929), .A(n18928), .ZN(n18941) );
  OAI21_X1 U21971 ( .B1(n18932), .B2(P3_STATEBS16_REG_SCAN_IN), .A(n18931), 
        .ZN(n18934) );
  AOI211_X1 U21972 ( .C1(n18947), .C2(n18934), .A(n18933), .B(n18945), .ZN(
        n18936) );
  NOR2_X1 U21973 ( .A1(n18936), .A2(n18935), .ZN(n18937) );
  OAI21_X1 U21974 ( .B1(n18938), .B2(n18937), .A(n18941), .ZN(n18939) );
  OAI21_X1 U21975 ( .B1(n18941), .B2(n18940), .A(n18939), .ZN(P3_U3296) );
  OAI22_X1 U21976 ( .A1(n18943), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18942), .ZN(n18944) );
  INV_X1 U21977 ( .A(n18944), .ZN(P3_U3297) );
  AOI21_X1 U21978 ( .B1(n18946), .B2(n18945), .A(n18948), .ZN(n18950) );
  INV_X1 U21979 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18949) );
  AOI22_X1 U21980 ( .A1(n18950), .A2(n18949), .B1(n18948), .B2(n18947), .ZN(
        P3_U3298) );
  INV_X1 U21981 ( .A(n18950), .ZN(n18952) );
  OAI21_X1 U21982 ( .B1(n18952), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n18951), 
        .ZN(n18953) );
  INV_X1 U21983 ( .A(n18953), .ZN(P3_U3299) );
  INV_X1 U21984 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n18954) );
  NAND2_X1 U21985 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19838), .ZN(n19829) );
  NAND2_X1 U21986 ( .A1(n18954), .A2(n18956), .ZN(n19826) );
  OAI21_X1 U21987 ( .B1(n18954), .B2(n19829), .A(n19826), .ZN(n19887) );
  OAI21_X1 U21988 ( .B1(n18954), .B2(n20917), .A(n19884), .ZN(P2_U2815) );
  INV_X1 U21989 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n21010) );
  OAI22_X1 U21990 ( .A1(n19953), .A2(n21010), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n18955), .ZN(P2_U2816) );
  OR2_X1 U21991 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n18956), .ZN(n19958) );
  INV_X2 U21992 ( .A(n19958), .ZN(n19960) );
  AOI22_X1 U21993 ( .A1(n19960), .A2(n21010), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n19958), .ZN(n18957) );
  OAI21_X1 U21994 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n19826), .A(n18957), 
        .ZN(P2_U2817) );
  INV_X1 U21995 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19941) );
  OAI21_X1 U21996 ( .B1(n19820), .B2(BS16), .A(n19887), .ZN(n19885) );
  OAI21_X1 U21997 ( .B1(n19887), .B2(n19941), .A(n19885), .ZN(P2_U2818) );
  NOR4_X1 U21998 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18967) );
  NOR4_X1 U21999 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_6__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18966) );
  AOI211_X1 U22000 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n18958) );
  INV_X1 U22001 ( .A(P2_DATAWIDTH_REG_8__SCAN_IN), .ZN(n21051) );
  INV_X1 U22002 ( .A(P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20899) );
  NAND3_X1 U22003 ( .A1(n18958), .A2(n21051), .A3(n20899), .ZN(n18964) );
  NOR4_X1 U22004 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18962) );
  NOR4_X1 U22005 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18961) );
  NOR4_X1 U22006 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18960) );
  NOR4_X1 U22007 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18959) );
  NAND4_X1 U22008 ( .A1(n18962), .A2(n18961), .A3(n18960), .A4(n18959), .ZN(
        n18963) );
  NOR4_X1 U22009 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(n18964), .A4(n18963), .ZN(n18965)
         );
  NAND3_X1 U22010 ( .A1(n18967), .A2(n18966), .A3(n18965), .ZN(n18973) );
  NOR2_X1 U22011 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18973), .ZN(n18968) );
  INV_X1 U22012 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19882) );
  AOI22_X1 U22013 ( .A1(n18968), .A2(n11406), .B1(n18973), .B2(n19882), .ZN(
        P2_U2820) );
  INV_X1 U22014 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20869) );
  INV_X1 U22015 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19886) );
  NAND3_X1 U22016 ( .A1(n11406), .A2(n20869), .A3(n19886), .ZN(n18972) );
  INV_X1 U22017 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19880) );
  AOI22_X1 U22018 ( .A1(n18968), .A2(n18972), .B1(n18973), .B2(n19880), .ZN(
        P2_U2821) );
  NAND2_X1 U22019 ( .A1(n18968), .A2(n19886), .ZN(n18971) );
  INV_X1 U22020 ( .A(n18973), .ZN(n18974) );
  OAI21_X1 U22021 ( .B1(n19839), .B2(n11406), .A(n18974), .ZN(n18969) );
  OAI21_X1 U22022 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18974), .A(n18969), 
        .ZN(n18970) );
  OAI221_X1 U22023 ( .B1(n18971), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18971), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18970), .ZN(P2_U2822) );
  INV_X1 U22024 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19878) );
  OAI221_X1 U22025 ( .B1(n18974), .B2(n19878), .C1(n18973), .C2(n18972), .A(
        n18971), .ZN(P2_U2823) );
  NOR2_X1 U22026 ( .A1(n19098), .A2(n18975), .ZN(n18976) );
  XOR2_X1 U22027 ( .A(n18977), .B(n18976), .Z(n18988) );
  NAND2_X1 U22028 ( .A1(n18978), .A2(n19125), .ZN(n18983) );
  INV_X1 U22029 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18979) );
  OAI22_X1 U22030 ( .A1(n19129), .A2(n18980), .B1(n18979), .B2(n18992), .ZN(
        n18981) );
  AOI21_X1 U22031 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(n19126), .A(n18981), .ZN(
        n18982) );
  OAI211_X1 U22032 ( .C1(n19085), .C2(n18984), .A(n18983), .B(n18982), .ZN(
        n18985) );
  AOI21_X1 U22033 ( .B1(n18986), .B2(n19123), .A(n18985), .ZN(n18987) );
  OAI21_X1 U22034 ( .B1(n19090), .B2(n18988), .A(n18987), .ZN(P2_U2835) );
  NAND2_X1 U22035 ( .A1(n9740), .A2(n18989), .ZN(n18990) );
  XOR2_X1 U22036 ( .A(n18991), .B(n18990), .Z(n19002) );
  OAI21_X1 U22037 ( .B1(n12047), .B2(n19129), .A(n9725), .ZN(n18996) );
  OAI22_X1 U22038 ( .A1(n18994), .A2(n19107), .B1(n18993), .B2(n18992), .ZN(
        n18995) );
  AOI211_X1 U22039 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19126), .A(n18996), .B(
        n18995), .ZN(n19001) );
  OAI22_X1 U22040 ( .A1(n18998), .A2(n19085), .B1(n18997), .B2(n19121), .ZN(
        n18999) );
  INV_X1 U22041 ( .A(n18999), .ZN(n19000) );
  OAI211_X1 U22042 ( .C1(n19090), .C2(n19002), .A(n19001), .B(n19000), .ZN(
        P2_U2836) );
  NAND2_X1 U22043 ( .A1(n9740), .A2(n19003), .ZN(n19004) );
  XOR2_X1 U22044 ( .A(n19005), .B(n19004), .Z(n19014) );
  AOI22_X1 U22045 ( .A1(n19006), .A2(n19125), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n9717), .ZN(n19007) );
  OAI211_X1 U22046 ( .C1(n19858), .C2(n19129), .A(n19007), .B(n9725), .ZN(
        n19008) );
  AOI21_X1 U22047 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n19126), .A(n19008), .ZN(
        n19013) );
  INV_X1 U22048 ( .A(n19009), .ZN(n19011) );
  AOI22_X1 U22049 ( .A1(n19011), .A2(n19133), .B1(n19010), .B2(n19123), .ZN(
        n19012) );
  OAI211_X1 U22050 ( .C1(n19090), .C2(n19014), .A(n19013), .B(n19012), .ZN(
        P2_U2838) );
  NAND2_X1 U22051 ( .A1(n9740), .A2(n19015), .ZN(n19017) );
  XOR2_X1 U22052 ( .A(n19017), .B(n19016), .Z(n19024) );
  AOI22_X1 U22053 ( .A1(n19018), .A2(n19125), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n9717), .ZN(n19019) );
  OAI211_X1 U22054 ( .C1(n15617), .C2(n19129), .A(n19019), .B(n9725), .ZN(
        n19022) );
  OAI22_X1 U22055 ( .A1(n19020), .A2(n19085), .B1(n19121), .B2(n19182), .ZN(
        n19021) );
  AOI211_X1 U22056 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n19126), .A(n19022), .B(
        n19021), .ZN(n19023) );
  OAI21_X1 U22057 ( .B1(n19024), .B2(n19090), .A(n19023), .ZN(P2_U2840) );
  NOR2_X1 U22058 ( .A1(n19098), .A2(n19035), .ZN(n19026) );
  XOR2_X1 U22059 ( .A(n19026), .B(n19025), .Z(n19033) );
  AOI22_X1 U22060 ( .A1(n19027), .A2(n19125), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n9717), .ZN(n19028) );
  OAI211_X1 U22061 ( .C1(n12030), .C2(n19129), .A(n19028), .B(n9725), .ZN(
        n19029) );
  AOI21_X1 U22062 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(n19126), .A(n19029), .ZN(
        n19032) );
  AOI22_X1 U22063 ( .A1(n19030), .A2(n19133), .B1(n19183), .B2(n19123), .ZN(
        n19031) );
  OAI211_X1 U22064 ( .C1(n19090), .C2(n19033), .A(n19032), .B(n19031), .ZN(
        P2_U2841) );
  INV_X1 U22065 ( .A(n19034), .ZN(n19137) );
  AOI211_X1 U22066 ( .C1(n19044), .C2(n19036), .A(n19035), .B(n19137), .ZN(
        n19043) );
  NAND2_X1 U22067 ( .A1(n19037), .A2(n19125), .ZN(n19041) );
  AOI22_X1 U22068 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n9717), .B1(
        P2_EBX_REG_13__SCAN_IN), .B2(n19126), .ZN(n19038) );
  OAI211_X1 U22069 ( .C1(n19129), .C2(n15847), .A(n19038), .B(n9725), .ZN(
        n19039) );
  INV_X1 U22070 ( .A(n19039), .ZN(n19040) );
  NAND2_X1 U22071 ( .A1(n19041), .A2(n19040), .ZN(n19042) );
  NOR2_X1 U22072 ( .A1(n19043), .A2(n19042), .ZN(n19047) );
  AOI22_X1 U22073 ( .A1(n19045), .A2(n19133), .B1(n19134), .B2(n19044), .ZN(
        n19046) );
  OAI211_X1 U22074 ( .C1(n19188), .C2(n19121), .A(n19047), .B(n19046), .ZN(
        P2_U2842) );
  AOI22_X1 U22075 ( .A1(n19126), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n9717), .ZN(n19048) );
  OAI21_X1 U22076 ( .B1(n19049), .B2(n19107), .A(n19048), .ZN(n19050) );
  AOI211_X1 U22077 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19060), .A(n19276), 
        .B(n19050), .ZN(n19056) );
  XNOR2_X1 U22078 ( .A(n19052), .B(n19051), .ZN(n19054) );
  AOI22_X1 U22079 ( .A1(n19054), .A2(n19117), .B1(n19053), .B2(n19133), .ZN(
        n19055) );
  OAI211_X1 U22080 ( .C1(n19191), .C2(n19121), .A(n19056), .B(n19055), .ZN(
        P2_U2843) );
  AOI22_X1 U22081 ( .A1(n19126), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n9717), .ZN(n19057) );
  OAI21_X1 U22082 ( .B1(n19058), .B2(n19107), .A(n19057), .ZN(n19059) );
  AOI211_X1 U22083 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n19060), .A(n19276), 
        .B(n19059), .ZN(n19067) );
  NOR2_X1 U22084 ( .A1(n19098), .A2(n19061), .ZN(n19063) );
  XNOR2_X1 U22085 ( .A(n19063), .B(n19062), .ZN(n19065) );
  AOI22_X1 U22086 ( .A1(n19065), .A2(n19117), .B1(n19064), .B2(n19133), .ZN(
        n19066) );
  OAI211_X1 U22087 ( .C1(n19196), .C2(n19121), .A(n19067), .B(n19066), .ZN(
        P2_U2845) );
  NAND2_X1 U22088 ( .A1(n9740), .A2(n19068), .ZN(n19070) );
  XOR2_X1 U22089 ( .A(n19070), .B(n19069), .Z(n19078) );
  AOI22_X1 U22090 ( .A1(n19071), .A2(n19125), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n19126), .ZN(n19072) );
  OAI211_X1 U22091 ( .C1(n12010), .C2(n19129), .A(n19072), .B(n9725), .ZN(
        n19076) );
  INV_X1 U22092 ( .A(n19073), .ZN(n19074) );
  OAI22_X1 U22093 ( .A1(n19074), .A2(n19085), .B1(n19199), .B2(n19121), .ZN(
        n19075) );
  AOI211_X1 U22094 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n9717), .A(
        n19076), .B(n19075), .ZN(n19077) );
  OAI21_X1 U22095 ( .B1(n19078), .B2(n19090), .A(n19077), .ZN(P2_U2846) );
  NAND2_X1 U22096 ( .A1(n9740), .A2(n19079), .ZN(n19081) );
  XOR2_X1 U22097 ( .A(n19081), .B(n19080), .Z(n19091) );
  INV_X1 U22098 ( .A(n19082), .ZN(n19083) );
  AOI22_X1 U22099 ( .A1(n19083), .A2(n19125), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19126), .ZN(n19084) );
  OAI211_X1 U22100 ( .C1(n12005), .C2(n19129), .A(n19084), .B(n9725), .ZN(
        n19088) );
  OAI22_X1 U22101 ( .A1(n19086), .A2(n19085), .B1(n19121), .B2(n19204), .ZN(
        n19087) );
  AOI211_X1 U22102 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n9717), .A(
        n19088), .B(n19087), .ZN(n19089) );
  OAI21_X1 U22103 ( .B1(n19091), .B2(n19090), .A(n19089), .ZN(P2_U2848) );
  OAI21_X1 U22104 ( .B1(n19845), .B2(n19129), .A(n9725), .ZN(n19095) );
  INV_X1 U22105 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19093) );
  OAI22_X1 U22106 ( .A1(n19109), .A2(n19093), .B1(n19092), .B2(n19107), .ZN(
        n19094) );
  AOI211_X1 U22107 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n9717), .A(
        n19095), .B(n19094), .ZN(n19105) );
  NOR2_X1 U22108 ( .A1(n19098), .A2(n19097), .ZN(n19100) );
  XNOR2_X1 U22109 ( .A(n19100), .B(n19099), .ZN(n19103) );
  INV_X1 U22110 ( .A(n19101), .ZN(n19102) );
  AOI22_X1 U22111 ( .A1(n19103), .A2(n19117), .B1(n19133), .B2(n19102), .ZN(
        n19104) );
  OAI211_X1 U22112 ( .C1(n19121), .C2(n19206), .A(n19105), .B(n19104), .ZN(
        P2_U2849) );
  OAI21_X1 U22113 ( .B1(n11998), .B2(n19129), .A(n9725), .ZN(n19111) );
  OAI22_X1 U22114 ( .A1(n19109), .A2(n19108), .B1(n19107), .B2(n19106), .ZN(
        n19110) );
  AOI211_X1 U22115 ( .C1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n9717), .A(
        n19111), .B(n19110), .ZN(n19120) );
  NAND2_X1 U22116 ( .A1(n9740), .A2(n19112), .ZN(n19114) );
  XNOR2_X1 U22117 ( .A(n19115), .B(n19114), .ZN(n19118) );
  AOI22_X1 U22118 ( .A1(n19118), .A2(n19117), .B1(n19133), .B2(n19116), .ZN(
        n19119) );
  OAI211_X1 U22119 ( .C1(n19121), .C2(n19214), .A(n19120), .B(n19119), .ZN(
        P2_U2850) );
  AOI22_X1 U22120 ( .A1(n19125), .A2(n19124), .B1(n19123), .B2(n19122), .ZN(
        n19128) );
  NAND2_X1 U22121 ( .A1(n19126), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n19127) );
  OAI211_X1 U22122 ( .C1(n11406), .C2(n19129), .A(n19128), .B(n19127), .ZN(
        n19132) );
  NOR2_X1 U22123 ( .A1(n19925), .A2(n19130), .ZN(n19131) );
  AOI211_X1 U22124 ( .C1(n19133), .C2(n12816), .A(n19132), .B(n19131), .ZN(
        n19136) );
  OAI21_X1 U22125 ( .B1(n9717), .B2(n19134), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19135) );
  OAI211_X1 U22126 ( .C1(n19138), .C2(n19137), .A(n19136), .B(n19135), .ZN(
        P2_U2855) );
  INV_X1 U22127 ( .A(n13758), .ZN(n19139) );
  AOI21_X1 U22128 ( .B1(n19140), .B2(n13621), .A(n19139), .ZN(n19176) );
  AOI22_X1 U22129 ( .A1(n19176), .A2(n19151), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n19161), .ZN(n19141) );
  OAI21_X1 U22130 ( .B1(n19161), .B2(n19142), .A(n19141), .ZN(P2_U2871) );
  XOR2_X1 U22131 ( .A(n13375), .B(n19143), .Z(n19144) );
  AOI22_X1 U22132 ( .A1(n19144), .A2(n19151), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19161), .ZN(n19145) );
  OAI21_X1 U22133 ( .B1(n19146), .B2(n19161), .A(n19145), .ZN(P2_U2873) );
  XNOR2_X1 U22134 ( .A(n13371), .B(n9816), .ZN(n19147) );
  AOI22_X1 U22135 ( .A1(n19147), .A2(n19151), .B1(P2_EBX_REG_12__SCAN_IN), 
        .B2(n19161), .ZN(n19148) );
  OAI21_X1 U22136 ( .B1(n19149), .B2(n19161), .A(n19148), .ZN(P2_U2875) );
  XNOR2_X1 U22137 ( .A(n13219), .B(n19150), .ZN(n19152) );
  AOI22_X1 U22138 ( .A1(n19152), .A2(n19151), .B1(P2_EBX_REG_10__SCAN_IN), 
        .B2(n19161), .ZN(n19153) );
  OAI21_X1 U22139 ( .B1(n19154), .B2(n19161), .A(n19153), .ZN(P2_U2877) );
  INV_X1 U22140 ( .A(n19155), .ZN(n19157) );
  AOI211_X1 U22141 ( .C1(n19158), .C2(n19157), .A(n19165), .B(n19156), .ZN(
        n19159) );
  AOI21_X1 U22142 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n19161), .A(n19159), .ZN(
        n19160) );
  OAI21_X1 U22143 ( .B1(n19162), .B2(n19161), .A(n19160), .ZN(P2_U2879) );
  OAI22_X1 U22144 ( .A1(n19218), .A2(n19165), .B1(n19164), .B2(n19163), .ZN(
        n19166) );
  INV_X1 U22145 ( .A(n19166), .ZN(n19167) );
  OAI21_X1 U22146 ( .B1(n19161), .B2(n19277), .A(n19167), .ZN(P2_U2883) );
  AOI22_X1 U22147 ( .A1(n19173), .A2(BUF1_REG_31__SCAN_IN), .B1(n19232), .B2(
        n19168), .ZN(n19170) );
  AOI22_X1 U22148 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19231), .B1(n19174), 
        .B2(BUF2_REG_31__SCAN_IN), .ZN(n19169) );
  NAND2_X1 U22149 ( .A1(n19170), .A2(n19169), .ZN(P2_U2888) );
  AOI22_X1 U22150 ( .A1(n19172), .A2(n19171), .B1(n19231), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19179) );
  AOI22_X1 U22151 ( .A1(n19174), .A2(BUF2_REG_16__SCAN_IN), .B1(n19173), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19178) );
  AOI22_X1 U22152 ( .A1(n19176), .A2(n19219), .B1(n19232), .B2(n19175), .ZN(
        n19177) );
  NAND3_X1 U22153 ( .A1(n19179), .A2(n19178), .A3(n19177), .ZN(P2_U2903) );
  OAI222_X1 U22154 ( .A1(n19182), .A2(n19215), .B1(n12809), .B2(n19205), .C1(
        n19181), .C2(n19240), .ZN(P2_U2904) );
  INV_X1 U22155 ( .A(n19183), .ZN(n19186) );
  AOI22_X1 U22156 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19231), .B1(n19184), 
        .B2(n19207), .ZN(n19185) );
  OAI21_X1 U22157 ( .B1(n19215), .B2(n19186), .A(n19185), .ZN(P2_U2905) );
  INV_X1 U22158 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n20993) );
  OAI222_X1 U22159 ( .A1(n19188), .A2(n19215), .B1(n20993), .B2(n19205), .C1(
        n19240), .C2(n19187), .ZN(P2_U2906) );
  AOI22_X1 U22160 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19231), .B1(n19189), 
        .B2(n19207), .ZN(n19190) );
  OAI21_X1 U22161 ( .B1(n19215), .B2(n19191), .A(n19190), .ZN(P2_U2907) );
  INV_X1 U22162 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19248) );
  OAI222_X1 U22163 ( .A1(n19193), .A2(n19215), .B1(n19248), .B2(n19205), .C1(
        n19240), .C2(n19192), .ZN(P2_U2908) );
  AOI22_X1 U22164 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19231), .B1(n19194), 
        .B2(n19207), .ZN(n19195) );
  OAI21_X1 U22165 ( .B1(n19215), .B2(n19196), .A(n19195), .ZN(P2_U2909) );
  AOI22_X1 U22166 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(n19231), .B1(n19197), .B2(
        n19207), .ZN(n19198) );
  OAI21_X1 U22167 ( .B1(n19215), .B2(n19199), .A(n19198), .ZN(P2_U2910) );
  INV_X1 U22168 ( .A(n19215), .ZN(n19201) );
  AOI22_X1 U22169 ( .A1(n19202), .A2(n19201), .B1(n19200), .B2(n19207), .ZN(
        n19203) );
  OAI21_X1 U22170 ( .B1(n19205), .B2(n20992), .A(n19203), .ZN(P2_U2911) );
  INV_X1 U22171 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19255) );
  OAI222_X1 U22172 ( .A1(n19204), .A2(n19215), .B1(n19255), .B2(n19205), .C1(
        n19240), .C2(n19344), .ZN(P2_U2912) );
  INV_X1 U22173 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19257) );
  OAI222_X1 U22174 ( .A1(n19206), .A2(n19215), .B1(n19257), .B2(n19205), .C1(
        n19240), .C2(n19331), .ZN(P2_U2913) );
  AOI22_X1 U22175 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19231), .B1(n19208), .B2(
        n19207), .ZN(n19213) );
  AOI21_X1 U22176 ( .B1(n19905), .B2(n19210), .A(n19209), .ZN(n19226) );
  XNOR2_X1 U22177 ( .A(n19567), .B(n19900), .ZN(n19227) );
  NOR2_X1 U22178 ( .A1(n19226), .A2(n19227), .ZN(n19225) );
  AOI21_X1 U22179 ( .B1(n19900), .B2(n19567), .A(n19225), .ZN(n19211) );
  NOR2_X1 U22180 ( .A1(n19211), .A2(n19216), .ZN(n19217) );
  OR3_X1 U22181 ( .A1(n19217), .A2(n19218), .A3(n19236), .ZN(n19212) );
  OAI211_X1 U22182 ( .C1(n19215), .C2(n19214), .A(n19213), .B(n19212), .ZN(
        P2_U2914) );
  AOI22_X1 U22183 ( .A1(n19232), .A2(n19216), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19231), .ZN(n19222) );
  XOR2_X1 U22184 ( .A(n19218), .B(n19217), .Z(n19220) );
  NAND2_X1 U22185 ( .A1(n19220), .A2(n19219), .ZN(n19221) );
  OAI211_X1 U22186 ( .C1(n19223), .C2(n19240), .A(n19222), .B(n19221), .ZN(
        P2_U2915) );
  AOI22_X1 U22187 ( .A1(n19224), .A2(n19232), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19231), .ZN(n19230) );
  AOI21_X1 U22188 ( .B1(n19227), .B2(n19226), .A(n19225), .ZN(n19228) );
  OR2_X1 U22189 ( .A1(n19228), .A2(n19236), .ZN(n19229) );
  OAI211_X1 U22190 ( .C1(n19320), .C2(n19240), .A(n19230), .B(n19229), .ZN(
        P2_U2916) );
  AOI22_X1 U22191 ( .A1(n19232), .A2(n19920), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19231), .ZN(n19239) );
  AOI21_X1 U22192 ( .B1(n19235), .B2(n19234), .A(n19233), .ZN(n19237) );
  OR2_X1 U22193 ( .A1(n19237), .A2(n19236), .ZN(n19238) );
  OAI211_X1 U22194 ( .C1(n19313), .C2(n19240), .A(n19239), .B(n19238), .ZN(
        P2_U2918) );
  NOR2_X1 U22195 ( .A1(n19261), .A2(n19241), .ZN(P2_U2920) );
  INV_X1 U22196 ( .A(n19259), .ZN(n19271) );
  AOI22_X1 U22197 ( .A1(n19269), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19268), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19242) );
  OAI21_X1 U22198 ( .B1(n12809), .B2(n19271), .A(n19242), .ZN(P2_U2936) );
  AOI22_X1 U22199 ( .A1(n19269), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19268), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19243) );
  OAI21_X1 U22200 ( .B1(n19244), .B2(n19271), .A(n19243), .ZN(P2_U2937) );
  AOI22_X1 U22201 ( .A1(n19269), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19268), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19245) );
  OAI21_X1 U22202 ( .B1(n20993), .B2(n19271), .A(n19245), .ZN(P2_U2938) );
  AOI22_X1 U22203 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19259), .B1(n19269), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n19246) );
  OAI21_X1 U22204 ( .B1(n19261), .B2(n20891), .A(n19246), .ZN(P2_U2939) );
  AOI22_X1 U22205 ( .A1(n19269), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19268), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19247) );
  OAI21_X1 U22206 ( .B1(n19248), .B2(n19271), .A(n19247), .ZN(P2_U2940) );
  AOI22_X1 U22207 ( .A1(n19269), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19268), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19249) );
  OAI21_X1 U22208 ( .B1(n19250), .B2(n19271), .A(n19249), .ZN(P2_U2941) );
  AOI22_X1 U22209 ( .A1(n19269), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19268), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19251) );
  OAI21_X1 U22210 ( .B1(n19252), .B2(n19271), .A(n19251), .ZN(P2_U2942) );
  AOI22_X1 U22211 ( .A1(n19269), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19268), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19253) );
  OAI21_X1 U22212 ( .B1(n20992), .B2(n19271), .A(n19253), .ZN(P2_U2943) );
  AOI22_X1 U22213 ( .A1(n19269), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19268), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19254) );
  OAI21_X1 U22214 ( .B1(n19255), .B2(n19271), .A(n19254), .ZN(P2_U2944) );
  AOI22_X1 U22215 ( .A1(n19269), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19268), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19256) );
  OAI21_X1 U22216 ( .B1(n19257), .B2(n19271), .A(n19256), .ZN(P2_U2945) );
  AOI22_X1 U22217 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19259), .B1(n19269), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n19258) );
  OAI21_X1 U22218 ( .B1(n19261), .B2(n20946), .A(n19258), .ZN(P2_U2946) );
  AOI22_X1 U22219 ( .A1(P2_EAX_REG_4__SCAN_IN), .A2(n19259), .B1(n19269), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n19260) );
  OAI21_X1 U22220 ( .B1(n19261), .B2(n20998), .A(n19260), .ZN(P2_U2947) );
  INV_X1 U22221 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19263) );
  AOI22_X1 U22222 ( .A1(n19269), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19268), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19262) );
  OAI21_X1 U22223 ( .B1(n19263), .B2(n19271), .A(n19262), .ZN(P2_U2948) );
  INV_X1 U22224 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19265) );
  AOI22_X1 U22225 ( .A1(n19269), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19268), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19264) );
  OAI21_X1 U22226 ( .B1(n19265), .B2(n19271), .A(n19264), .ZN(P2_U2949) );
  INV_X1 U22227 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19267) );
  AOI22_X1 U22228 ( .A1(n19269), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19268), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19266) );
  OAI21_X1 U22229 ( .B1(n19267), .B2(n19271), .A(n19266), .ZN(P2_U2950) );
  AOI22_X1 U22230 ( .A1(n19269), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19268), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19270) );
  OAI21_X1 U22231 ( .B1(n12966), .B2(n19271), .A(n19270), .ZN(P2_U2951) );
  AOI22_X1 U22232 ( .A1(n19273), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n19272), .ZN(n19275) );
  NAND2_X1 U22233 ( .A1(n19275), .A2(n19274), .ZN(P2_U2979) );
  AOI22_X1 U22234 ( .A1(n19284), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19276), .ZN(n19282) );
  INV_X1 U22235 ( .A(n19277), .ZN(n19279) );
  AOI222_X1 U22236 ( .A1(n19280), .A2(n19288), .B1(n19294), .B2(n19279), .C1(
        n19285), .C2(n19278), .ZN(n19281) );
  OAI211_X1 U22237 ( .C1(n19291), .C2(n19283), .A(n19282), .B(n19281), .ZN(
        P2_U3010) );
  AOI22_X1 U22238 ( .A1(n19286), .A2(n19285), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19284), .ZN(n19297) );
  AOI21_X1 U22239 ( .B1(n19289), .B2(n19288), .A(n19287), .ZN(n19290) );
  OAI21_X1 U22240 ( .B1(n19292), .B2(n19291), .A(n19290), .ZN(n19293) );
  AOI21_X1 U22241 ( .B1(n19295), .B2(n19294), .A(n19293), .ZN(n19296) );
  NAND2_X1 U22242 ( .A1(n19297), .A2(n19296), .ZN(P2_U3012) );
  INV_X1 U22243 ( .A(n19683), .ZN(n19298) );
  INV_X1 U22244 ( .A(n19712), .ZN(n19895) );
  OR2_X1 U22245 ( .A1(n19395), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19356) );
  NOR2_X1 U22246 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19356), .ZN(
        n19342) );
  AOI22_X1 U22247 ( .A1(n19767), .A2(n19792), .B1(n19759), .B2(n19342), .ZN(
        n19309) );
  AOI21_X1 U22248 ( .B1(n19818), .B2(n19378), .A(n19941), .ZN(n19299) );
  NOR2_X1 U22249 ( .A1(n19299), .A2(n19719), .ZN(n19304) );
  INV_X1 U22250 ( .A(n19810), .ZN(n19302) );
  INV_X1 U22251 ( .A(n19300), .ZN(n19305) );
  AOI21_X1 U22252 ( .B1(n19305), .B2(n19757), .A(n19894), .ZN(n19301) );
  AOI21_X1 U22253 ( .B1(n19304), .B2(n19302), .A(n19301), .ZN(n19303) );
  OAI21_X1 U22254 ( .B1(n19303), .B2(n19342), .A(n19765), .ZN(n19346) );
  OAI21_X1 U22255 ( .B1(n19810), .B2(n19342), .A(n19304), .ZN(n19307) );
  OAI21_X1 U22256 ( .B1(n19305), .B2(n19342), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19306) );
  NAND2_X1 U22257 ( .A1(n19307), .A2(n19306), .ZN(n19345) );
  AOI22_X1 U22258 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19346), .B1(
        n19760), .B2(n19345), .ZN(n19308) );
  OAI211_X1 U22259 ( .C1(n19770), .C2(n19378), .A(n19309), .B(n19308), .ZN(
        P2_U3048) );
  AOI22_X1 U22260 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19335), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19334), .ZN(n19731) );
  OAI22_X1 U22261 ( .A1(n19311), .A2(n19338), .B1(n19310), .B2(n19336), .ZN(
        n19728) );
  INV_X1 U22262 ( .A(n19340), .ZN(n19312) );
  AOI22_X1 U22263 ( .A1(n19728), .A2(n19792), .B1(n19771), .B2(n19342), .ZN(
        n19315) );
  NOR2_X2 U22264 ( .A1(n19313), .A2(n19343), .ZN(n19772) );
  AOI22_X1 U22265 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19346), .B1(
        n19772), .B2(n19345), .ZN(n19314) );
  OAI211_X1 U22266 ( .C1(n19731), .C2(n19378), .A(n19315), .B(n19314), .ZN(
        P2_U3049) );
  AOI22_X1 U22267 ( .A1(n19779), .A2(n19792), .B1(n19777), .B2(n19342), .ZN(
        n19317) );
  AOI22_X1 U22268 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19346), .B1(
        n19778), .B2(n19345), .ZN(n19316) );
  OAI211_X1 U22269 ( .C1(n19782), .C2(n19378), .A(n19317), .B(n19316), .ZN(
        P2_U3050) );
  AOI22_X1 U22270 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19335), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19334), .ZN(n19737) );
  OAI22_X2 U22271 ( .A1(n20947), .A2(n19336), .B1(n19318), .B2(n19338), .ZN(
        n19734) );
  NOR2_X2 U22272 ( .A1(n9852), .A2(n19340), .ZN(n19783) );
  AOI22_X1 U22273 ( .A1(n19734), .A2(n19792), .B1(n19783), .B2(n19342), .ZN(
        n19322) );
  NOR2_X2 U22274 ( .A1(n19320), .A2(n19343), .ZN(n19784) );
  AOI22_X1 U22275 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19346), .B1(
        n19784), .B2(n19345), .ZN(n19321) );
  OAI211_X1 U22276 ( .C1(n19737), .C2(n19378), .A(n19322), .B(n19321), .ZN(
        P2_U3051) );
  AOI22_X1 U22277 ( .A1(n19738), .A2(n19792), .B1(n19789), .B2(n19342), .ZN(
        n19324) );
  AOI22_X1 U22278 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19346), .B1(
        n19790), .B2(n19345), .ZN(n19323) );
  OAI211_X1 U22279 ( .C1(n19741), .C2(n19378), .A(n19324), .B(n19323), .ZN(
        P2_U3052) );
  AOI22_X1 U22280 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19335), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19334), .ZN(n19802) );
  AOI22_X1 U22281 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19335), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19334), .ZN(n19653) );
  NOR2_X2 U22282 ( .A1(n19325), .A2(n19340), .ZN(n19797) );
  AOI22_X1 U22283 ( .A1(n19792), .A2(n19799), .B1(n19797), .B2(n19342), .ZN(
        n19328) );
  NOR2_X2 U22284 ( .A1(n19326), .A2(n19343), .ZN(n19798) );
  AOI22_X1 U22285 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19346), .B1(
        n19798), .B2(n19345), .ZN(n19327) );
  OAI211_X1 U22286 ( .C1(n19802), .C2(n19378), .A(n19328), .B(n19327), .ZN(
        P2_U3053) );
  AOI22_X1 U22287 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19335), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19334), .ZN(n19808) );
  OAI22_X1 U22288 ( .A1(n19330), .A2(n19336), .B1(n19329), .B2(n19338), .ZN(
        n19805) );
  NOR2_X2 U22289 ( .A1(n12955), .A2(n19340), .ZN(n19803) );
  AOI22_X1 U22290 ( .A1(n19805), .A2(n19792), .B1(n19803), .B2(n19342), .ZN(
        n19333) );
  NOR2_X2 U22291 ( .A1(n19331), .A2(n19343), .ZN(n19804) );
  AOI22_X1 U22292 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19346), .B1(
        n19804), .B2(n19345), .ZN(n19332) );
  OAI211_X1 U22293 ( .C1(n19808), .C2(n19378), .A(n19333), .B(n19332), .ZN(
        P2_U3054) );
  AOI22_X1 U22294 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19335), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19334), .ZN(n19819) );
  OAI22_X2 U22295 ( .A1(n19339), .A2(n19338), .B1(n19337), .B2(n19336), .ZN(
        n19813) );
  NOR2_X2 U22296 ( .A1(n19341), .A2(n19340), .ZN(n19809) );
  AOI22_X1 U22297 ( .A1(n19813), .A2(n19792), .B1(n19809), .B2(n19342), .ZN(
        n19348) );
  NOR2_X2 U22298 ( .A1(n19344), .A2(n19343), .ZN(n19811) );
  AOI22_X1 U22299 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19346), .B1(
        n19811), .B2(n19345), .ZN(n19347) );
  OAI211_X1 U22300 ( .C1(n19819), .C2(n19378), .A(n19348), .B(n19347), .ZN(
        P2_U3055) );
  INV_X1 U22301 ( .A(n19767), .ZN(n19640) );
  INV_X1 U22302 ( .A(n19349), .ZN(n19350) );
  NOR2_X1 U22303 ( .A1(n19566), .A2(n19395), .ZN(n19373) );
  NOR3_X1 U22304 ( .A1(n19350), .A2(n19373), .A3(n19685), .ZN(n19355) );
  INV_X1 U22305 ( .A(n19356), .ZN(n19351) );
  AOI21_X1 U22306 ( .B1(n19757), .B2(n19351), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19352) );
  NOR2_X1 U22307 ( .A1(n19355), .A2(n19352), .ZN(n19374) );
  AOI22_X1 U22308 ( .A1(n19374), .A2(n19760), .B1(n19759), .B2(n19373), .ZN(
        n19360) );
  INV_X1 U22309 ( .A(n19896), .ZN(n19354) );
  INV_X1 U22310 ( .A(n19568), .ZN(n19353) );
  NAND2_X1 U22311 ( .A1(n19354), .A2(n19353), .ZN(n19357) );
  AOI21_X1 U22312 ( .B1(n19357), .B2(n19356), .A(n19355), .ZN(n19358) );
  OAI211_X1 U22313 ( .C1(n19373), .C2(n19757), .A(n19358), .B(n19765), .ZN(
        n19375) );
  AOI22_X1 U22314 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19375), .B1(
        n19391), .B2(n19637), .ZN(n19359) );
  OAI211_X1 U22315 ( .C1(n19640), .C2(n19378), .A(n19360), .B(n19359), .ZN(
        P2_U3056) );
  INV_X1 U22316 ( .A(n19728), .ZN(n19776) );
  AOI22_X1 U22317 ( .A1(n19374), .A2(n19772), .B1(n19771), .B2(n19373), .ZN(
        n19362) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19375), .B1(
        n19391), .B2(n19773), .ZN(n19361) );
  OAI211_X1 U22319 ( .C1(n19776), .C2(n19378), .A(n19362), .B(n19361), .ZN(
        P2_U3057) );
  INV_X1 U22320 ( .A(n19779), .ZN(n19646) );
  AOI22_X1 U22321 ( .A1(n19374), .A2(n19778), .B1(n19777), .B2(n19373), .ZN(
        n19364) );
  AOI22_X1 U22322 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19375), .B1(
        n19391), .B2(n19643), .ZN(n19363) );
  OAI211_X1 U22323 ( .C1(n19646), .C2(n19378), .A(n19364), .B(n19363), .ZN(
        P2_U3058) );
  INV_X1 U22324 ( .A(n19734), .ZN(n19788) );
  AOI22_X1 U22325 ( .A1(n19374), .A2(n19784), .B1(n19783), .B2(n19373), .ZN(
        n19366) );
  INV_X1 U22326 ( .A(n19737), .ZN(n19785) );
  AOI22_X1 U22327 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19375), .B1(
        n19391), .B2(n19785), .ZN(n19365) );
  OAI211_X1 U22328 ( .C1(n19788), .C2(n19378), .A(n19366), .B(n19365), .ZN(
        P2_U3059) );
  INV_X1 U22329 ( .A(n19738), .ZN(n19796) );
  AOI22_X1 U22330 ( .A1(n19374), .A2(n19790), .B1(n19789), .B2(n19373), .ZN(
        n19368) );
  AOI22_X1 U22331 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19375), .B1(
        n19391), .B2(n19791), .ZN(n19367) );
  OAI211_X1 U22332 ( .C1(n19796), .C2(n19378), .A(n19368), .B(n19367), .ZN(
        P2_U3060) );
  AOI22_X1 U22333 ( .A1(n19374), .A2(n19798), .B1(n19797), .B2(n19373), .ZN(
        n19370) );
  INV_X1 U22334 ( .A(n19802), .ZN(n19670) );
  AOI22_X1 U22335 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19375), .B1(
        n19391), .B2(n19670), .ZN(n19369) );
  OAI211_X1 U22336 ( .C1(n19653), .C2(n19378), .A(n19370), .B(n19369), .ZN(
        P2_U3061) );
  INV_X1 U22337 ( .A(n19805), .ZN(n19656) );
  AOI22_X1 U22338 ( .A1(n19374), .A2(n19804), .B1(n19803), .B2(n19373), .ZN(
        n19372) );
  AOI22_X1 U22339 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19375), .B1(
        n19391), .B2(n19673), .ZN(n19371) );
  OAI211_X1 U22340 ( .C1(n19656), .C2(n19378), .A(n19372), .B(n19371), .ZN(
        P2_U3062) );
  AOI22_X1 U22341 ( .A1(n19374), .A2(n19811), .B1(n19809), .B2(n19373), .ZN(
        n19377) );
  INV_X1 U22342 ( .A(n19819), .ZN(n19748) );
  AOI22_X1 U22343 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19375), .B1(
        n19391), .B2(n19748), .ZN(n19376) );
  OAI211_X1 U22344 ( .C1(n19754), .C2(n19378), .A(n19377), .B(n19376), .ZN(
        P2_U3063) );
  AOI22_X1 U22345 ( .A1(n19390), .A2(n19772), .B1(n19389), .B2(n19771), .ZN(
        n19380) );
  AOI22_X1 U22346 ( .A1(n19391), .A2(n19728), .B1(n19412), .B2(n19773), .ZN(
        n19379) );
  OAI211_X1 U22347 ( .C1(n19394), .C2(n13731), .A(n19380), .B(n19379), .ZN(
        P2_U3065) );
  AOI22_X1 U22348 ( .A1(n19390), .A2(n19778), .B1(n19389), .B2(n19777), .ZN(
        n19382) );
  AOI22_X1 U22349 ( .A1(n19391), .A2(n19779), .B1(n19412), .B2(n19643), .ZN(
        n19381) );
  OAI211_X1 U22350 ( .C1(n19394), .C2(n13985), .A(n19382), .B(n19381), .ZN(
        P2_U3066) );
  AOI22_X1 U22351 ( .A1(n19390), .A2(n19784), .B1(n19389), .B2(n19783), .ZN(
        n19384) );
  AOI22_X1 U22352 ( .A1(n19391), .A2(n19734), .B1(n19412), .B2(n19785), .ZN(
        n19383) );
  OAI211_X1 U22353 ( .C1(n19394), .C2(n14009), .A(n19384), .B(n19383), .ZN(
        P2_U3067) );
  AOI22_X1 U22354 ( .A1(n19390), .A2(n19798), .B1(n19389), .B2(n19797), .ZN(
        n19386) );
  AOI22_X1 U22355 ( .A1(n19391), .A2(n19799), .B1(n19412), .B2(n19670), .ZN(
        n19385) );
  OAI211_X1 U22356 ( .C1(n19394), .C2(n14104), .A(n19386), .B(n19385), .ZN(
        P2_U3069) );
  AOI22_X1 U22357 ( .A1(n19390), .A2(n19804), .B1(n19389), .B2(n19803), .ZN(
        n19388) );
  AOI22_X1 U22358 ( .A1(n19391), .A2(n19805), .B1(n19412), .B2(n19673), .ZN(
        n19387) );
  OAI211_X1 U22359 ( .C1(n19394), .C2(n14113), .A(n19388), .B(n19387), .ZN(
        P2_U3070) );
  AOI22_X1 U22360 ( .A1(n19390), .A2(n19811), .B1(n19389), .B2(n19809), .ZN(
        n19393) );
  AOI22_X1 U22361 ( .A1(n19391), .A2(n19813), .B1(n19412), .B2(n19748), .ZN(
        n19392) );
  OAI211_X1 U22362 ( .C1(n19394), .C2(n14319), .A(n19393), .B(n19392), .ZN(
        P2_U3071) );
  NOR2_X1 U22363 ( .A1(n19629), .A2(n19395), .ZN(n19419) );
  AOI22_X1 U22364 ( .A1(n19767), .A2(n19412), .B1(n19759), .B2(n19419), .ZN(
        n19405) );
  OAI21_X1 U22365 ( .B1(n19896), .B2(n19888), .A(n19894), .ZN(n19403) );
  NOR2_X1 U22366 ( .A1(n19922), .A2(n19395), .ZN(n19398) );
  INV_X1 U22367 ( .A(n19419), .ZN(n19396) );
  OAI211_X1 U22368 ( .C1(n19399), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19719), 
        .B(n19396), .ZN(n19397) );
  OAI211_X1 U22369 ( .C1(n19403), .C2(n19398), .A(n19765), .B(n19397), .ZN(
        n19421) );
  INV_X1 U22370 ( .A(n19398), .ZN(n19402) );
  INV_X1 U22371 ( .A(n19399), .ZN(n19400) );
  OAI21_X1 U22372 ( .B1(n19400), .B2(n19419), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19401) );
  OAI21_X1 U22373 ( .B1(n19403), .B2(n19402), .A(n19401), .ZN(n19420) );
  AOI22_X1 U22374 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19421), .B1(
        n19760), .B2(n19420), .ZN(n19404) );
  OAI211_X1 U22375 ( .C1(n19770), .C2(n19457), .A(n19405), .B(n19404), .ZN(
        P2_U3072) );
  AOI22_X1 U22376 ( .A1(n19447), .A2(n19773), .B1(n19419), .B2(n19771), .ZN(
        n19407) );
  AOI22_X1 U22377 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19421), .B1(
        n19772), .B2(n19420), .ZN(n19406) );
  OAI211_X1 U22378 ( .C1(n19776), .C2(n19424), .A(n19407), .B(n19406), .ZN(
        P2_U3073) );
  AOI22_X1 U22379 ( .A1(n19779), .A2(n19412), .B1(n19777), .B2(n19419), .ZN(
        n19409) );
  AOI22_X1 U22380 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19421), .B1(
        n19778), .B2(n19420), .ZN(n19408) );
  OAI211_X1 U22381 ( .C1(n19782), .C2(n19457), .A(n19409), .B(n19408), .ZN(
        P2_U3074) );
  AOI22_X1 U22382 ( .A1(n19734), .A2(n19412), .B1(n19419), .B2(n19783), .ZN(
        n19411) );
  AOI22_X1 U22383 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19421), .B1(
        n19784), .B2(n19420), .ZN(n19410) );
  OAI211_X1 U22384 ( .C1(n19737), .C2(n19457), .A(n19411), .B(n19410), .ZN(
        P2_U3075) );
  AOI22_X1 U22385 ( .A1(n19738), .A2(n19412), .B1(n19789), .B2(n19419), .ZN(
        n19414) );
  AOI22_X1 U22386 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19421), .B1(
        n19790), .B2(n19420), .ZN(n19413) );
  OAI211_X1 U22387 ( .C1(n19741), .C2(n19457), .A(n19414), .B(n19413), .ZN(
        P2_U3076) );
  AOI22_X1 U22388 ( .A1(n19670), .A2(n19447), .B1(n19419), .B2(n19797), .ZN(
        n19416) );
  AOI22_X1 U22389 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19421), .B1(
        n19798), .B2(n19420), .ZN(n19415) );
  OAI211_X1 U22390 ( .C1(n19653), .C2(n19424), .A(n19416), .B(n19415), .ZN(
        P2_U3077) );
  AOI22_X1 U22391 ( .A1(n19447), .A2(n19673), .B1(n19419), .B2(n19803), .ZN(
        n19418) );
  AOI22_X1 U22392 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19421), .B1(
        n19804), .B2(n19420), .ZN(n19417) );
  OAI211_X1 U22393 ( .C1(n19656), .C2(n19424), .A(n19418), .B(n19417), .ZN(
        P2_U3078) );
  AOI22_X1 U22394 ( .A1(n19748), .A2(n19447), .B1(n19419), .B2(n19809), .ZN(
        n19423) );
  AOI22_X1 U22395 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19421), .B1(
        n19811), .B2(n19420), .ZN(n19422) );
  OAI211_X1 U22396 ( .C1(n19754), .C2(n19424), .A(n19423), .B(n19422), .ZN(
        P2_U3079) );
  NOR2_X1 U22397 ( .A1(n19490), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19459) );
  INV_X1 U22398 ( .A(n19459), .ZN(n19465) );
  NOR2_X1 U22399 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19465), .ZN(
        n19452) );
  INV_X1 U22400 ( .A(n19452), .ZN(n19428) );
  NAND2_X1 U22401 ( .A1(n19426), .A2(n19903), .ZN(n19432) );
  OAI21_X1 U22402 ( .B1(n19482), .B2(n19447), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19429) );
  AOI22_X1 U22403 ( .A1(n19432), .A2(n19429), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19428), .ZN(n19430) );
  NAND2_X1 U22404 ( .A1(n19765), .A2(n19430), .ZN(n19431) );
  INV_X1 U22405 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n19437) );
  OR2_X1 U22406 ( .A1(n19432), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19434) );
  AOI21_X1 U22407 ( .B1(n19685), .B2(n19434), .A(n19433), .ZN(n19453) );
  AOI22_X1 U22408 ( .A1(n19453), .A2(n19760), .B1(n19759), .B2(n19452), .ZN(
        n19436) );
  AOI22_X1 U22409 ( .A1(n19447), .A2(n19767), .B1(n19482), .B2(n19637), .ZN(
        n19435) );
  OAI211_X1 U22410 ( .C1(n19438), .C2(n19437), .A(n19436), .B(n19435), .ZN(
        P2_U3080) );
  AOI22_X1 U22411 ( .A1(n19453), .A2(n19772), .B1(n19771), .B2(n19452), .ZN(
        n19440) );
  AOI22_X1 U22412 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19454), .B1(
        n19482), .B2(n19773), .ZN(n19439) );
  OAI211_X1 U22413 ( .C1(n19776), .C2(n19457), .A(n19440), .B(n19439), .ZN(
        P2_U3081) );
  AOI22_X1 U22414 ( .A1(n19453), .A2(n19778), .B1(n19777), .B2(n19452), .ZN(
        n19442) );
  AOI22_X1 U22415 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19454), .B1(
        n19447), .B2(n19779), .ZN(n19441) );
  OAI211_X1 U22416 ( .C1(n19782), .C2(n19481), .A(n19442), .B(n19441), .ZN(
        P2_U3082) );
  AOI22_X1 U22417 ( .A1(n19453), .A2(n19784), .B1(n19783), .B2(n19452), .ZN(
        n19444) );
  AOI22_X1 U22418 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19454), .B1(
        n19447), .B2(n19734), .ZN(n19443) );
  OAI211_X1 U22419 ( .C1(n19737), .C2(n19481), .A(n19444), .B(n19443), .ZN(
        P2_U3083) );
  AOI22_X1 U22420 ( .A1(n19453), .A2(n19790), .B1(n19789), .B2(n19452), .ZN(
        n19446) );
  AOI22_X1 U22421 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19454), .B1(
        n19447), .B2(n19738), .ZN(n19445) );
  OAI211_X1 U22422 ( .C1(n19741), .C2(n19481), .A(n19446), .B(n19445), .ZN(
        P2_U3084) );
  AOI22_X1 U22423 ( .A1(n19453), .A2(n19798), .B1(n19797), .B2(n19452), .ZN(
        n19449) );
  AOI22_X1 U22424 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19454), .B1(
        n19447), .B2(n19799), .ZN(n19448) );
  OAI211_X1 U22425 ( .C1(n19802), .C2(n19481), .A(n19449), .B(n19448), .ZN(
        P2_U3085) );
  AOI22_X1 U22426 ( .A1(n19453), .A2(n19804), .B1(n19803), .B2(n19452), .ZN(
        n19451) );
  AOI22_X1 U22427 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19454), .B1(
        n19482), .B2(n19673), .ZN(n19450) );
  OAI211_X1 U22428 ( .C1(n19656), .C2(n19457), .A(n19451), .B(n19450), .ZN(
        P2_U3086) );
  AOI22_X1 U22429 ( .A1(n19453), .A2(n19811), .B1(n19809), .B2(n19452), .ZN(
        n19456) );
  AOI22_X1 U22430 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19454), .B1(
        n19482), .B2(n19748), .ZN(n19455) );
  OAI211_X1 U22431 ( .C1(n19754), .C2(n19457), .A(n19456), .B(n19455), .ZN(
        P2_U3087) );
  NOR2_X2 U22432 ( .A1(n19458), .A2(n19687), .ZN(n19511) );
  INV_X1 U22433 ( .A(n19511), .ZN(n19487) );
  NOR2_X1 U22434 ( .A1(n19566), .A2(n19490), .ZN(n19491) );
  AOI22_X1 U22435 ( .A1(n19767), .A2(n19482), .B1(n19759), .B2(n19491), .ZN(
        n19468) );
  OAI21_X1 U22436 ( .B1(n19896), .B2(n19687), .A(n19894), .ZN(n19466) );
  NOR2_X1 U22437 ( .A1(n19466), .A2(n19459), .ZN(n19460) );
  AOI211_X1 U22438 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19462), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19460), .ZN(n19461) );
  OAI21_X1 U22439 ( .B1(n19461), .B2(n19491), .A(n19765), .ZN(n19484) );
  INV_X1 U22440 ( .A(n19462), .ZN(n19463) );
  OAI21_X1 U22441 ( .B1(n19463), .B2(n19491), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19464) );
  OAI21_X1 U22442 ( .B1(n19466), .B2(n19465), .A(n19464), .ZN(n19483) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19484), .B1(
        n19760), .B2(n19483), .ZN(n19467) );
  OAI211_X1 U22444 ( .C1(n19770), .C2(n19487), .A(n19468), .B(n19467), .ZN(
        P2_U3088) );
  AOI22_X1 U22445 ( .A1(n19728), .A2(n19482), .B1(n19771), .B2(n19491), .ZN(
        n19470) );
  AOI22_X1 U22446 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19484), .B1(
        n19772), .B2(n19483), .ZN(n19469) );
  OAI211_X1 U22447 ( .C1(n19731), .C2(n19487), .A(n19470), .B(n19469), .ZN(
        P2_U3089) );
  AOI22_X1 U22448 ( .A1(n19643), .A2(n19511), .B1(n19777), .B2(n19491), .ZN(
        n19472) );
  AOI22_X1 U22449 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19484), .B1(
        n19778), .B2(n19483), .ZN(n19471) );
  OAI211_X1 U22450 ( .C1(n19646), .C2(n19481), .A(n19472), .B(n19471), .ZN(
        P2_U3090) );
  AOI22_X1 U22451 ( .A1(n19785), .A2(n19511), .B1(n19491), .B2(n19783), .ZN(
        n19474) );
  AOI22_X1 U22452 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19484), .B1(
        n19784), .B2(n19483), .ZN(n19473) );
  OAI211_X1 U22453 ( .C1(n19788), .C2(n19481), .A(n19474), .B(n19473), .ZN(
        P2_U3091) );
  AOI22_X1 U22454 ( .A1(n19738), .A2(n19482), .B1(n19789), .B2(n19491), .ZN(
        n19476) );
  AOI22_X1 U22455 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19484), .B1(
        n19790), .B2(n19483), .ZN(n19475) );
  OAI211_X1 U22456 ( .C1(n19741), .C2(n19487), .A(n19476), .B(n19475), .ZN(
        P2_U3092) );
  AOI22_X1 U22457 ( .A1(n19482), .A2(n19799), .B1(n19797), .B2(n19491), .ZN(
        n19478) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19484), .B1(
        n19798), .B2(n19483), .ZN(n19477) );
  OAI211_X1 U22459 ( .C1(n19802), .C2(n19487), .A(n19478), .B(n19477), .ZN(
        P2_U3093) );
  AOI22_X1 U22460 ( .A1(n19511), .A2(n19673), .B1(n19803), .B2(n19491), .ZN(
        n19480) );
  AOI22_X1 U22461 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19484), .B1(
        n19804), .B2(n19483), .ZN(n19479) );
  OAI211_X1 U22462 ( .C1(n19656), .C2(n19481), .A(n19480), .B(n19479), .ZN(
        P2_U3094) );
  AOI22_X1 U22463 ( .A1(n19813), .A2(n19482), .B1(n19809), .B2(n19491), .ZN(
        n19486) );
  AOI22_X1 U22464 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19484), .B1(
        n19811), .B2(n19483), .ZN(n19485) );
  OAI211_X1 U22465 ( .C1(n19819), .C2(n19487), .A(n19486), .B(n19485), .ZN(
        P2_U3095) );
  INV_X1 U22466 ( .A(n11612), .ZN(n19488) );
  NOR2_X1 U22467 ( .A1(n19598), .A2(n19490), .ZN(n19509) );
  OAI21_X1 U22468 ( .B1(n19488), .B2(n19509), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19489) );
  OAI21_X1 U22469 ( .B1(n19490), .B2(n19601), .A(n19489), .ZN(n19510) );
  AOI22_X1 U22470 ( .A1(n19510), .A2(n19760), .B1(n19759), .B2(n19509), .ZN(
        n19496) );
  AOI221_X1 U22471 ( .B1(n19511), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19492), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19491), .ZN(n19493) );
  AOI211_X1 U22472 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n11612), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19493), .ZN(n19494) );
  AOI22_X1 U22473 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19512), .B1(
        n19511), .B2(n19767), .ZN(n19495) );
  OAI211_X1 U22474 ( .C1(n19770), .C2(n19529), .A(n19496), .B(n19495), .ZN(
        P2_U3096) );
  AOI22_X1 U22475 ( .A1(n19510), .A2(n19772), .B1(n19771), .B2(n19509), .ZN(
        n19498) );
  AOI22_X1 U22476 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19512), .B1(
        n19511), .B2(n19728), .ZN(n19497) );
  OAI211_X1 U22477 ( .C1(n19731), .C2(n19529), .A(n19498), .B(n19497), .ZN(
        P2_U3097) );
  AOI22_X1 U22478 ( .A1(n19510), .A2(n19778), .B1(n19777), .B2(n19509), .ZN(
        n19500) );
  AOI22_X1 U22479 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19512), .B1(
        n19511), .B2(n19779), .ZN(n19499) );
  OAI211_X1 U22480 ( .C1(n19782), .C2(n19529), .A(n19500), .B(n19499), .ZN(
        P2_U3098) );
  AOI22_X1 U22481 ( .A1(n19510), .A2(n19784), .B1(n19783), .B2(n19509), .ZN(
        n19502) );
  AOI22_X1 U22482 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19512), .B1(
        n19511), .B2(n19734), .ZN(n19501) );
  OAI211_X1 U22483 ( .C1(n19737), .C2(n19529), .A(n19502), .B(n19501), .ZN(
        P2_U3099) );
  AOI22_X1 U22484 ( .A1(n19510), .A2(n19790), .B1(n19789), .B2(n19509), .ZN(
        n19504) );
  AOI22_X1 U22485 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19512), .B1(
        n19511), .B2(n19738), .ZN(n19503) );
  OAI211_X1 U22486 ( .C1(n19741), .C2(n19529), .A(n19504), .B(n19503), .ZN(
        P2_U3100) );
  AOI22_X1 U22487 ( .A1(n19510), .A2(n19798), .B1(n19797), .B2(n19509), .ZN(
        n19506) );
  AOI22_X1 U22488 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19512), .B1(
        n19511), .B2(n19799), .ZN(n19505) );
  OAI211_X1 U22489 ( .C1(n19802), .C2(n19529), .A(n19506), .B(n19505), .ZN(
        P2_U3101) );
  AOI22_X1 U22490 ( .A1(n19510), .A2(n19804), .B1(n19803), .B2(n19509), .ZN(
        n19508) );
  AOI22_X1 U22491 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19512), .B1(
        n19511), .B2(n19805), .ZN(n19507) );
  OAI211_X1 U22492 ( .C1(n19808), .C2(n19529), .A(n19508), .B(n19507), .ZN(
        P2_U3102) );
  AOI22_X1 U22493 ( .A1(n19510), .A2(n19811), .B1(n19809), .B2(n19509), .ZN(
        n19514) );
  AOI22_X1 U22494 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19512), .B1(
        n19511), .B2(n19813), .ZN(n19513) );
  OAI211_X1 U22495 ( .C1(n19819), .C2(n19529), .A(n19514), .B(n19513), .ZN(
        P2_U3103) );
  AOI22_X1 U22496 ( .A1(n19525), .A2(n19772), .B1(n19533), .B2(n19771), .ZN(
        n19516) );
  AOI22_X1 U22497 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19526), .B1(
        n19560), .B2(n19773), .ZN(n19515) );
  OAI211_X1 U22498 ( .C1(n19776), .C2(n19529), .A(n19516), .B(n19515), .ZN(
        P2_U3105) );
  AOI22_X1 U22499 ( .A1(n19525), .A2(n19784), .B1(n19533), .B2(n19783), .ZN(
        n19518) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19526), .B1(
        n19560), .B2(n19785), .ZN(n19517) );
  OAI211_X1 U22501 ( .C1(n19788), .C2(n19529), .A(n19518), .B(n19517), .ZN(
        P2_U3107) );
  AOI22_X1 U22502 ( .A1(n19525), .A2(n19790), .B1(n19789), .B2(n19533), .ZN(
        n19520) );
  AOI22_X1 U22503 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19526), .B1(
        n19560), .B2(n19791), .ZN(n19519) );
  OAI211_X1 U22504 ( .C1(n19796), .C2(n19529), .A(n19520), .B(n19519), .ZN(
        P2_U3108) );
  AOI22_X1 U22505 ( .A1(n19525), .A2(n19798), .B1(n19533), .B2(n19797), .ZN(
        n19522) );
  AOI22_X1 U22506 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19526), .B1(
        n19560), .B2(n19670), .ZN(n19521) );
  OAI211_X1 U22507 ( .C1(n19653), .C2(n19529), .A(n19522), .B(n19521), .ZN(
        P2_U3109) );
  AOI22_X1 U22508 ( .A1(n19525), .A2(n19804), .B1(n19533), .B2(n19803), .ZN(
        n19524) );
  AOI22_X1 U22509 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19526), .B1(
        n19560), .B2(n19673), .ZN(n19523) );
  OAI211_X1 U22510 ( .C1(n19656), .C2(n19529), .A(n19524), .B(n19523), .ZN(
        P2_U3110) );
  AOI22_X1 U22511 ( .A1(n19525), .A2(n19811), .B1(n19533), .B2(n19809), .ZN(
        n19528) );
  AOI22_X1 U22512 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19526), .B1(
        n19560), .B2(n19748), .ZN(n19527) );
  OAI211_X1 U22513 ( .C1(n19754), .C2(n19529), .A(n19528), .B(n19527), .ZN(
        P2_U3111) );
  NOR2_X2 U22514 ( .A1(n19713), .A2(n19568), .ZN(n19592) );
  INV_X1 U22515 ( .A(n19560), .ZN(n19530) );
  NAND2_X1 U22516 ( .A1(n19894), .A2(n19530), .ZN(n19531) );
  NAND2_X1 U22517 ( .A1(n19894), .A2(n19941), .ZN(n19890) );
  INV_X1 U22518 ( .A(n19541), .ZN(n19536) );
  NAND2_X1 U22519 ( .A1(n19912), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19628) );
  NOR2_X1 U22520 ( .A1(n19628), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19571) );
  INV_X1 U22521 ( .A(n19571), .ZN(n19575) );
  NOR2_X1 U22522 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19575), .ZN(
        n19559) );
  NOR2_X1 U22523 ( .A1(n19559), .A2(n19533), .ZN(n19539) );
  AOI21_X1 U22524 ( .B1(n19537), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19534) );
  OAI21_X1 U22525 ( .B1(n19534), .B2(n19559), .A(n19765), .ZN(n19535) );
  INV_X1 U22526 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n19544) );
  AOI22_X1 U22527 ( .A1(n19637), .A2(n19592), .B1(n19759), .B2(n19559), .ZN(
        n19543) );
  INV_X1 U22528 ( .A(n19537), .ZN(n19538) );
  OAI21_X1 U22529 ( .B1(n19538), .B2(n19559), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19540) );
  AOI22_X1 U22530 ( .A1(n19541), .A2(n19540), .B1(n19539), .B2(n19685), .ZN(
        n19561) );
  AOI22_X1 U22531 ( .A1(n19760), .A2(n19561), .B1(n19560), .B2(n19767), .ZN(
        n19542) );
  OAI211_X1 U22532 ( .C1(n19565), .C2(n19544), .A(n19543), .B(n19542), .ZN(
        P2_U3112) );
  AOI22_X1 U22533 ( .A1(n19592), .A2(n19773), .B1(n19771), .B2(n19559), .ZN(
        n19546) );
  AOI22_X1 U22534 ( .A1(n19772), .A2(n19561), .B1(n19560), .B2(n19728), .ZN(
        n19545) );
  OAI211_X1 U22535 ( .C1(n19565), .C2(n12169), .A(n19546), .B(n19545), .ZN(
        P2_U3113) );
  INV_X1 U22536 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n19549) );
  AOI22_X1 U22537 ( .A1(n19643), .A2(n19592), .B1(n19777), .B2(n19559), .ZN(
        n19548) );
  AOI22_X1 U22538 ( .A1(n19778), .A2(n19561), .B1(n19560), .B2(n19779), .ZN(
        n19547) );
  OAI211_X1 U22539 ( .C1(n19565), .C2(n19549), .A(n19548), .B(n19547), .ZN(
        P2_U3114) );
  AOI22_X1 U22540 ( .A1(n19785), .A2(n19592), .B1(n19783), .B2(n19559), .ZN(
        n19551) );
  AOI22_X1 U22541 ( .A1(n19784), .A2(n19561), .B1(n19560), .B2(n19734), .ZN(
        n19550) );
  OAI211_X1 U22542 ( .C1(n19565), .C2(n12203), .A(n19551), .B(n19550), .ZN(
        P2_U3115) );
  AOI22_X1 U22543 ( .A1(n19791), .A2(n19592), .B1(n19789), .B2(n19559), .ZN(
        n19553) );
  AOI22_X1 U22544 ( .A1(n19790), .A2(n19561), .B1(n19560), .B2(n19738), .ZN(
        n19552) );
  OAI211_X1 U22545 ( .C1(n19565), .C2(n19554), .A(n19553), .B(n19552), .ZN(
        P2_U3116) );
  AOI22_X1 U22546 ( .A1(n19670), .A2(n19592), .B1(n19797), .B2(n19559), .ZN(
        n19556) );
  AOI22_X1 U22547 ( .A1(n19798), .A2(n19561), .B1(n19560), .B2(n19799), .ZN(
        n19555) );
  OAI211_X1 U22548 ( .C1(n19565), .C2(n12242), .A(n19556), .B(n19555), .ZN(
        P2_U3117) );
  AOI22_X1 U22549 ( .A1(n19592), .A2(n19673), .B1(n19803), .B2(n19559), .ZN(
        n19558) );
  AOI22_X1 U22550 ( .A1(n19804), .A2(n19561), .B1(n19560), .B2(n19805), .ZN(
        n19557) );
  OAI211_X1 U22551 ( .C1(n19565), .C2(n12263), .A(n19558), .B(n19557), .ZN(
        P2_U3118) );
  AOI22_X1 U22552 ( .A1(n19592), .A2(n19748), .B1(n19809), .B2(n19559), .ZN(
        n19563) );
  AOI22_X1 U22553 ( .A1(n19811), .A2(n19561), .B1(n19560), .B2(n19813), .ZN(
        n19562) );
  OAI211_X1 U22554 ( .C1(n19565), .C2(n19564), .A(n19563), .B(n19562), .ZN(
        P2_U3119) );
  NOR2_X2 U22555 ( .A1(n19683), .A2(n19568), .ZN(n19623) );
  INV_X1 U22556 ( .A(n19623), .ZN(n19597) );
  NOR2_X1 U22557 ( .A1(n19566), .A2(n19628), .ZN(n19602) );
  AOI22_X1 U22558 ( .A1(n19767), .A2(n19592), .B1(n19759), .B2(n19602), .ZN(
        n19578) );
  INV_X1 U22559 ( .A(n19567), .ZN(n19892) );
  NAND2_X1 U22560 ( .A1(n19892), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19688) );
  OAI21_X1 U22561 ( .B1(n19688), .B2(n19568), .A(n19894), .ZN(n19576) );
  INV_X1 U22562 ( .A(n19602), .ZN(n19569) );
  OAI211_X1 U22563 ( .C1(n19572), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19719), 
        .B(n19569), .ZN(n19570) );
  OAI211_X1 U22564 ( .C1(n19576), .C2(n19571), .A(n19765), .B(n19570), .ZN(
        n19594) );
  INV_X1 U22565 ( .A(n19572), .ZN(n19573) );
  OAI21_X1 U22566 ( .B1(n19573), .B2(n19602), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19574) );
  OAI21_X1 U22567 ( .B1(n19576), .B2(n19575), .A(n19574), .ZN(n19593) );
  AOI22_X1 U22568 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19594), .B1(
        n19760), .B2(n19593), .ZN(n19577) );
  OAI211_X1 U22569 ( .C1(n19770), .C2(n19597), .A(n19578), .B(n19577), .ZN(
        P2_U3120) );
  INV_X1 U22570 ( .A(n19592), .ZN(n19591) );
  AOI22_X1 U22571 ( .A1(n19623), .A2(n19773), .B1(n19771), .B2(n19602), .ZN(
        n19580) );
  AOI22_X1 U22572 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19594), .B1(
        n19772), .B2(n19593), .ZN(n19579) );
  OAI211_X1 U22573 ( .C1(n19776), .C2(n19591), .A(n19580), .B(n19579), .ZN(
        P2_U3121) );
  AOI22_X1 U22574 ( .A1(n19643), .A2(n19623), .B1(n19777), .B2(n19602), .ZN(
        n19582) );
  AOI22_X1 U22575 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19594), .B1(
        n19778), .B2(n19593), .ZN(n19581) );
  OAI211_X1 U22576 ( .C1(n19646), .C2(n19591), .A(n19582), .B(n19581), .ZN(
        P2_U3122) );
  AOI22_X1 U22577 ( .A1(n19734), .A2(n19592), .B1(n19783), .B2(n19602), .ZN(
        n19584) );
  AOI22_X1 U22578 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19594), .B1(
        n19784), .B2(n19593), .ZN(n19583) );
  OAI211_X1 U22579 ( .C1(n19737), .C2(n19597), .A(n19584), .B(n19583), .ZN(
        P2_U3123) );
  AOI22_X1 U22580 ( .A1(n19738), .A2(n19592), .B1(n19789), .B2(n19602), .ZN(
        n19586) );
  AOI22_X1 U22581 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19594), .B1(
        n19790), .B2(n19593), .ZN(n19585) );
  OAI211_X1 U22582 ( .C1(n19741), .C2(n19597), .A(n19586), .B(n19585), .ZN(
        P2_U3124) );
  AOI22_X1 U22583 ( .A1(n19670), .A2(n19623), .B1(n19797), .B2(n19602), .ZN(
        n19588) );
  AOI22_X1 U22584 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19594), .B1(
        n19798), .B2(n19593), .ZN(n19587) );
  OAI211_X1 U22585 ( .C1(n19653), .C2(n19591), .A(n19588), .B(n19587), .ZN(
        P2_U3125) );
  AOI22_X1 U22586 ( .A1(n19623), .A2(n19673), .B1(n19803), .B2(n19602), .ZN(
        n19590) );
  AOI22_X1 U22587 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19594), .B1(
        n19804), .B2(n19593), .ZN(n19589) );
  OAI211_X1 U22588 ( .C1(n19656), .C2(n19591), .A(n19590), .B(n19589), .ZN(
        P2_U3126) );
  AOI22_X1 U22589 ( .A1(n19813), .A2(n19592), .B1(n19809), .B2(n19602), .ZN(
        n19596) );
  AOI22_X1 U22590 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19594), .B1(
        n19811), .B2(n19593), .ZN(n19595) );
  OAI211_X1 U22591 ( .C1(n19819), .C2(n19597), .A(n19596), .B(n19595), .ZN(
        P2_U3127) );
  INV_X1 U22592 ( .A(n19605), .ZN(n19599) );
  NOR2_X1 U22593 ( .A1(n19598), .A2(n19628), .ZN(n19621) );
  OAI21_X1 U22594 ( .B1(n19599), .B2(n19621), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19600) );
  OAI21_X1 U22595 ( .B1(n19628), .B2(n19601), .A(n19600), .ZN(n19622) );
  AOI22_X1 U22596 ( .A1(n19622), .A2(n19760), .B1(n19759), .B2(n19621), .ZN(
        n19608) );
  AOI221_X1 U22597 ( .B1(n19623), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19603), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19602), .ZN(n19604) );
  AOI211_X1 U22598 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19605), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19604), .ZN(n19606) );
  AOI22_X1 U22599 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19624), .B1(
        n19623), .B2(n19767), .ZN(n19607) );
  OAI211_X1 U22600 ( .C1(n19770), .C2(n19662), .A(n19608), .B(n19607), .ZN(
        P2_U3128) );
  AOI22_X1 U22601 ( .A1(n19622), .A2(n19772), .B1(n19771), .B2(n19621), .ZN(
        n19610) );
  AOI22_X1 U22602 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19624), .B1(
        n19623), .B2(n19728), .ZN(n19609) );
  OAI211_X1 U22603 ( .C1(n19731), .C2(n19662), .A(n19610), .B(n19609), .ZN(
        P2_U3129) );
  AOI22_X1 U22604 ( .A1(n19622), .A2(n19778), .B1(n19777), .B2(n19621), .ZN(
        n19612) );
  AOI22_X1 U22605 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19624), .B1(
        n19623), .B2(n19779), .ZN(n19611) );
  OAI211_X1 U22606 ( .C1(n19782), .C2(n19662), .A(n19612), .B(n19611), .ZN(
        P2_U3130) );
  AOI22_X1 U22607 ( .A1(n19622), .A2(n19784), .B1(n19783), .B2(n19621), .ZN(
        n19614) );
  AOI22_X1 U22608 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19624), .B1(
        n19623), .B2(n19734), .ZN(n19613) );
  OAI211_X1 U22609 ( .C1(n19737), .C2(n19662), .A(n19614), .B(n19613), .ZN(
        P2_U3131) );
  AOI22_X1 U22610 ( .A1(n19622), .A2(n19790), .B1(n19789), .B2(n19621), .ZN(
        n19616) );
  AOI22_X1 U22611 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19624), .B1(
        n19623), .B2(n19738), .ZN(n19615) );
  OAI211_X1 U22612 ( .C1(n19741), .C2(n19662), .A(n19616), .B(n19615), .ZN(
        P2_U3132) );
  AOI22_X1 U22613 ( .A1(n19622), .A2(n19798), .B1(n19797), .B2(n19621), .ZN(
        n19618) );
  AOI22_X1 U22614 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19624), .B1(
        n19623), .B2(n19799), .ZN(n19617) );
  OAI211_X1 U22615 ( .C1(n19802), .C2(n19662), .A(n19618), .B(n19617), .ZN(
        P2_U3133) );
  AOI22_X1 U22616 ( .A1(n19622), .A2(n19804), .B1(n19803), .B2(n19621), .ZN(
        n19620) );
  AOI22_X1 U22617 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19624), .B1(
        n19623), .B2(n19805), .ZN(n19619) );
  OAI211_X1 U22618 ( .C1(n19808), .C2(n19662), .A(n19620), .B(n19619), .ZN(
        P2_U3134) );
  AOI22_X1 U22619 ( .A1(n19622), .A2(n19811), .B1(n19809), .B2(n19621), .ZN(
        n19626) );
  AOI22_X1 U22620 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19624), .B1(
        n19623), .B2(n19813), .ZN(n19625) );
  OAI211_X1 U22621 ( .C1(n19819), .C2(n19662), .A(n19626), .B(n19625), .ZN(
        P2_U3135) );
  INV_X1 U22622 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19685) );
  OR2_X1 U22623 ( .A1(n19922), .A2(n19628), .ZN(n19634) );
  OR2_X1 U22624 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19634), .ZN(n19631) );
  INV_X1 U22625 ( .A(n19627), .ZN(n19630) );
  NOR2_X1 U22626 ( .A1(n19629), .A2(n19628), .ZN(n19657) );
  NOR3_X1 U22627 ( .A1(n19630), .A2(n19657), .A3(n19685), .ZN(n19633) );
  AOI21_X1 U22628 ( .B1(n19685), .B2(n19631), .A(n19633), .ZN(n19658) );
  AOI22_X1 U22629 ( .A1(n19658), .A2(n19760), .B1(n19759), .B2(n19657), .ZN(
        n19639) );
  INV_X1 U22630 ( .A(n19688), .ZN(n19761) );
  INV_X1 U22631 ( .A(n19888), .ZN(n19632) );
  NAND2_X1 U22632 ( .A1(n19761), .A2(n19632), .ZN(n19635) );
  AOI21_X1 U22633 ( .B1(n19635), .B2(n19634), .A(n19633), .ZN(n19636) );
  OAI211_X1 U22634 ( .C1(n19657), .C2(n19757), .A(n19636), .B(n19765), .ZN(
        n19659) );
  AOI22_X1 U22635 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19659), .B1(
        n19678), .B2(n19637), .ZN(n19638) );
  OAI211_X1 U22636 ( .C1(n19640), .C2(n19662), .A(n19639), .B(n19638), .ZN(
        P2_U3136) );
  AOI22_X1 U22637 ( .A1(n19658), .A2(n19772), .B1(n19771), .B2(n19657), .ZN(
        n19642) );
  AOI22_X1 U22638 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19659), .B1(
        n19678), .B2(n19773), .ZN(n19641) );
  OAI211_X1 U22639 ( .C1(n19776), .C2(n19662), .A(n19642), .B(n19641), .ZN(
        P2_U3137) );
  AOI22_X1 U22640 ( .A1(n19658), .A2(n19778), .B1(n19777), .B2(n19657), .ZN(
        n19645) );
  AOI22_X1 U22641 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19659), .B1(
        n19678), .B2(n19643), .ZN(n19644) );
  OAI211_X1 U22642 ( .C1(n19646), .C2(n19662), .A(n19645), .B(n19644), .ZN(
        P2_U3138) );
  AOI22_X1 U22643 ( .A1(n19658), .A2(n19784), .B1(n19783), .B2(n19657), .ZN(
        n19648) );
  AOI22_X1 U22644 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19659), .B1(
        n19678), .B2(n19785), .ZN(n19647) );
  OAI211_X1 U22645 ( .C1(n19788), .C2(n19662), .A(n19648), .B(n19647), .ZN(
        P2_U3139) );
  AOI22_X1 U22646 ( .A1(n19658), .A2(n19790), .B1(n19789), .B2(n19657), .ZN(
        n19650) );
  AOI22_X1 U22647 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19659), .B1(
        n19678), .B2(n19791), .ZN(n19649) );
  OAI211_X1 U22648 ( .C1(n19796), .C2(n19662), .A(n19650), .B(n19649), .ZN(
        P2_U3140) );
  AOI22_X1 U22649 ( .A1(n19658), .A2(n19798), .B1(n19797), .B2(n19657), .ZN(
        n19652) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19659), .B1(
        n19678), .B2(n19670), .ZN(n19651) );
  OAI211_X1 U22651 ( .C1(n19653), .C2(n19662), .A(n19652), .B(n19651), .ZN(
        P2_U3141) );
  AOI22_X1 U22652 ( .A1(n19658), .A2(n19804), .B1(n19803), .B2(n19657), .ZN(
        n19655) );
  AOI22_X1 U22653 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19659), .B1(
        n19678), .B2(n19673), .ZN(n19654) );
  OAI211_X1 U22654 ( .C1(n19656), .C2(n19662), .A(n19655), .B(n19654), .ZN(
        P2_U3142) );
  AOI22_X1 U22655 ( .A1(n19658), .A2(n19811), .B1(n19809), .B2(n19657), .ZN(
        n19661) );
  AOI22_X1 U22656 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19659), .B1(
        n19678), .B2(n19748), .ZN(n19660) );
  OAI211_X1 U22657 ( .C1(n19754), .C2(n19662), .A(n19661), .B(n19660), .ZN(
        P2_U3143) );
  AOI22_X1 U22658 ( .A1(n19677), .A2(n19772), .B1(n19676), .B2(n19771), .ZN(
        n19664) );
  AOI22_X1 U22659 ( .A1(n19678), .A2(n19728), .B1(n19708), .B2(n19773), .ZN(
        n19663) );
  OAI211_X1 U22660 ( .C1(n19682), .C2(n11490), .A(n19664), .B(n19663), .ZN(
        P2_U3145) );
  AOI22_X1 U22661 ( .A1(n19677), .A2(n19784), .B1(n19676), .B2(n19783), .ZN(
        n19666) );
  AOI22_X1 U22662 ( .A1(n19678), .A2(n19734), .B1(n19708), .B2(n19785), .ZN(
        n19665) );
  OAI211_X1 U22663 ( .C1(n19682), .C2(n11562), .A(n19666), .B(n19665), .ZN(
        P2_U3147) );
  AOI22_X1 U22664 ( .A1(n19677), .A2(n19790), .B1(n19789), .B2(n19676), .ZN(
        n19668) );
  AOI22_X1 U22665 ( .A1(n19678), .A2(n19738), .B1(n19708), .B2(n19791), .ZN(
        n19667) );
  OAI211_X1 U22666 ( .C1(n19682), .C2(n19669), .A(n19668), .B(n19667), .ZN(
        P2_U3148) );
  AOI22_X1 U22667 ( .A1(n19677), .A2(n19798), .B1(n19676), .B2(n19797), .ZN(
        n19672) );
  AOI22_X1 U22668 ( .A1(n19678), .A2(n19799), .B1(n19708), .B2(n19670), .ZN(
        n19671) );
  OAI211_X1 U22669 ( .C1(n19682), .C2(n11604), .A(n19672), .B(n19671), .ZN(
        P2_U3149) );
  AOI22_X1 U22670 ( .A1(n19677), .A2(n19804), .B1(n19676), .B2(n19803), .ZN(
        n19675) );
  AOI22_X1 U22671 ( .A1(n19678), .A2(n19805), .B1(n19708), .B2(n19673), .ZN(
        n19674) );
  OAI211_X1 U22672 ( .C1(n19682), .C2(n11716), .A(n19675), .B(n19674), .ZN(
        P2_U3150) );
  INV_X1 U22673 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n19681) );
  AOI22_X1 U22674 ( .A1(n19677), .A2(n19811), .B1(n19676), .B2(n19809), .ZN(
        n19680) );
  AOI22_X1 U22675 ( .A1(n19678), .A2(n19813), .B1(n19708), .B2(n19748), .ZN(
        n19679) );
  OAI211_X1 U22676 ( .C1(n19682), .C2(n19681), .A(n19680), .B(n19679), .ZN(
        P2_U3151) );
  NOR2_X1 U22677 ( .A1(n19931), .A2(n19689), .ZN(n19717) );
  INV_X1 U22678 ( .A(n19717), .ZN(n19684) );
  NAND3_X1 U22679 ( .A1(n11616), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19684), 
        .ZN(n19690) );
  OAI21_X1 U22680 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19689), .A(n19685), 
        .ZN(n19686) );
  AND2_X1 U22681 ( .A1(n19690), .A2(n19686), .ZN(n19707) );
  AOI22_X1 U22682 ( .A1(n19707), .A2(n19760), .B1(n19759), .B2(n19717), .ZN(
        n19694) );
  NOR3_X1 U22683 ( .A1(n19688), .A2(P2_STATE2_REG_3__SCAN_IN), .A3(n19687), 
        .ZN(n19692) );
  AOI21_X1 U22684 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19931), .A(n19689), 
        .ZN(n19691) );
  OAI211_X1 U22685 ( .C1(n19692), .C2(n19691), .A(n19765), .B(n19690), .ZN(
        n19709) );
  AOI22_X1 U22686 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19767), .ZN(n19693) );
  OAI211_X1 U22687 ( .C1(n19770), .C2(n19753), .A(n19694), .B(n19693), .ZN(
        P2_U3152) );
  AOI22_X1 U22688 ( .A1(n19707), .A2(n19772), .B1(n19771), .B2(n19717), .ZN(
        n19696) );
  AOI22_X1 U22689 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19728), .ZN(n19695) );
  OAI211_X1 U22690 ( .C1(n19731), .C2(n19753), .A(n19696), .B(n19695), .ZN(
        P2_U3153) );
  AOI22_X1 U22691 ( .A1(n19707), .A2(n19778), .B1(n19777), .B2(n19717), .ZN(
        n19698) );
  AOI22_X1 U22692 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19779), .ZN(n19697) );
  OAI211_X1 U22693 ( .C1(n19782), .C2(n19753), .A(n19698), .B(n19697), .ZN(
        P2_U3154) );
  AOI22_X1 U22694 ( .A1(n19707), .A2(n19784), .B1(n19783), .B2(n19717), .ZN(
        n19700) );
  AOI22_X1 U22695 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19734), .ZN(n19699) );
  OAI211_X1 U22696 ( .C1(n19737), .C2(n19753), .A(n19700), .B(n19699), .ZN(
        P2_U3155) );
  AOI22_X1 U22697 ( .A1(n19707), .A2(n19790), .B1(n19789), .B2(n19717), .ZN(
        n19702) );
  AOI22_X1 U22698 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19738), .ZN(n19701) );
  OAI211_X1 U22699 ( .C1(n19741), .C2(n19753), .A(n19702), .B(n19701), .ZN(
        P2_U3156) );
  AOI22_X1 U22700 ( .A1(n19707), .A2(n19798), .B1(n19797), .B2(n19717), .ZN(
        n19704) );
  AOI22_X1 U22701 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19799), .ZN(n19703) );
  OAI211_X1 U22702 ( .C1(n19802), .C2(n19753), .A(n19704), .B(n19703), .ZN(
        P2_U3157) );
  AOI22_X1 U22703 ( .A1(n19707), .A2(n19804), .B1(n19803), .B2(n19717), .ZN(
        n19706) );
  AOI22_X1 U22704 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19805), .ZN(n19705) );
  OAI211_X1 U22705 ( .C1(n19808), .C2(n19753), .A(n19706), .B(n19705), .ZN(
        P2_U3158) );
  AOI22_X1 U22706 ( .A1(n19707), .A2(n19811), .B1(n19809), .B2(n19717), .ZN(
        n19711) );
  AOI22_X1 U22707 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19813), .ZN(n19710) );
  OAI211_X1 U22708 ( .C1(n19819), .C2(n19753), .A(n19711), .B(n19710), .ZN(
        P2_U3159) );
  NAND2_X1 U22709 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19714), .ZN(
        n19763) );
  NOR2_X1 U22710 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19763), .ZN(
        n19747) );
  AOI22_X1 U22711 ( .A1(n19767), .A2(n19744), .B1(n19759), .B2(n19747), .ZN(
        n19727) );
  NOR3_X1 U22712 ( .A1(n19814), .A2(n19744), .A3(n19719), .ZN(n19716) );
  INV_X1 U22713 ( .A(n19890), .ZN(n19715) );
  NOR2_X1 U22714 ( .A1(n19716), .A2(n19715), .ZN(n19725) );
  NOR2_X1 U22715 ( .A1(n19747), .A2(n19717), .ZN(n19724) );
  INV_X1 U22716 ( .A(n19724), .ZN(n19721) );
  INV_X1 U22717 ( .A(n19747), .ZN(n19718) );
  OAI211_X1 U22718 ( .C1(n11615), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19719), 
        .B(n19718), .ZN(n19720) );
  OAI211_X1 U22719 ( .C1(n19725), .C2(n19721), .A(n19765), .B(n19720), .ZN(
        n19750) );
  INV_X1 U22720 ( .A(n11615), .ZN(n19722) );
  OAI21_X1 U22721 ( .B1(n19722), .B2(n19747), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19723) );
  OAI21_X1 U22722 ( .B1(n19725), .B2(n19724), .A(n19723), .ZN(n19749) );
  AOI22_X1 U22723 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19750), .B1(
        n19760), .B2(n19749), .ZN(n19726) );
  OAI211_X1 U22724 ( .C1(n19770), .C2(n19795), .A(n19727), .B(n19726), .ZN(
        P2_U3160) );
  AOI22_X1 U22725 ( .A1(n19728), .A2(n19744), .B1(n19771), .B2(n19747), .ZN(
        n19730) );
  AOI22_X1 U22726 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19750), .B1(
        n19772), .B2(n19749), .ZN(n19729) );
  OAI211_X1 U22727 ( .C1(n19731), .C2(n19795), .A(n19730), .B(n19729), .ZN(
        P2_U3161) );
  AOI22_X1 U22728 ( .A1(n19779), .A2(n19744), .B1(n19777), .B2(n19747), .ZN(
        n19733) );
  AOI22_X1 U22729 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19750), .B1(
        n19778), .B2(n19749), .ZN(n19732) );
  OAI211_X1 U22730 ( .C1(n19782), .C2(n19795), .A(n19733), .B(n19732), .ZN(
        P2_U3162) );
  AOI22_X1 U22731 ( .A1(n19734), .A2(n19744), .B1(n19783), .B2(n19747), .ZN(
        n19736) );
  AOI22_X1 U22732 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19750), .B1(
        n19784), .B2(n19749), .ZN(n19735) );
  OAI211_X1 U22733 ( .C1(n19737), .C2(n19795), .A(n19736), .B(n19735), .ZN(
        P2_U3163) );
  AOI22_X1 U22734 ( .A1(n19738), .A2(n19744), .B1(n19789), .B2(n19747), .ZN(
        n19740) );
  AOI22_X1 U22735 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19750), .B1(
        n19790), .B2(n19749), .ZN(n19739) );
  OAI211_X1 U22736 ( .C1(n19741), .C2(n19795), .A(n19740), .B(n19739), .ZN(
        P2_U3164) );
  AOI22_X1 U22737 ( .A1(n19744), .A2(n19799), .B1(n19797), .B2(n19747), .ZN(
        n19743) );
  AOI22_X1 U22738 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19750), .B1(
        n19798), .B2(n19749), .ZN(n19742) );
  OAI211_X1 U22739 ( .C1(n19802), .C2(n19795), .A(n19743), .B(n19742), .ZN(
        P2_U3165) );
  AOI22_X1 U22740 ( .A1(n19805), .A2(n19744), .B1(n19803), .B2(n19747), .ZN(
        n19746) );
  AOI22_X1 U22741 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19750), .B1(
        n19804), .B2(n19749), .ZN(n19745) );
  OAI211_X1 U22742 ( .C1(n19808), .C2(n19795), .A(n19746), .B(n19745), .ZN(
        P2_U3166) );
  AOI22_X1 U22743 ( .A1(n19814), .A2(n19748), .B1(n19809), .B2(n19747), .ZN(
        n19752) );
  AOI22_X1 U22744 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19750), .B1(
        n19811), .B2(n19749), .ZN(n19751) );
  OAI211_X1 U22745 ( .C1(n19754), .C2(n19753), .A(n19752), .B(n19751), .ZN(
        P2_U3167) );
  INV_X1 U22746 ( .A(n11608), .ZN(n19755) );
  NOR3_X1 U22747 ( .A1(n19755), .A2(n19810), .A3(n19685), .ZN(n19762) );
  INV_X1 U22748 ( .A(n19763), .ZN(n19756) );
  AOI21_X1 U22749 ( .B1(n19757), .B2(n19756), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19758) );
  NOR2_X1 U22750 ( .A1(n19762), .A2(n19758), .ZN(n19812) );
  AOI22_X1 U22751 ( .A1(n19812), .A2(n19760), .B1(n19810), .B2(n19759), .ZN(
        n19769) );
  NAND2_X1 U22752 ( .A1(n19761), .A2(n19895), .ZN(n19764) );
  AOI21_X1 U22753 ( .B1(n19764), .B2(n19763), .A(n19762), .ZN(n19766) );
  OAI211_X1 U22754 ( .C1(n19810), .C2(n19757), .A(n19766), .B(n19765), .ZN(
        n19815) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n19767), .ZN(n19768) );
  OAI211_X1 U22756 ( .C1(n19770), .C2(n19818), .A(n19769), .B(n19768), .ZN(
        P2_U3168) );
  AOI22_X1 U22757 ( .A1(n19812), .A2(n19772), .B1(n19810), .B2(n19771), .ZN(
        n19775) );
  AOI22_X1 U22758 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19815), .B1(
        n19792), .B2(n19773), .ZN(n19774) );
  OAI211_X1 U22759 ( .C1(n19776), .C2(n19795), .A(n19775), .B(n19774), .ZN(
        P2_U3169) );
  AOI22_X1 U22760 ( .A1(n19812), .A2(n19778), .B1(n19810), .B2(n19777), .ZN(
        n19781) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n19779), .ZN(n19780) );
  OAI211_X1 U22762 ( .C1(n19782), .C2(n19818), .A(n19781), .B(n19780), .ZN(
        P2_U3170) );
  AOI22_X1 U22763 ( .A1(n19812), .A2(n19784), .B1(n19810), .B2(n19783), .ZN(
        n19787) );
  AOI22_X1 U22764 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19815), .B1(
        n19792), .B2(n19785), .ZN(n19786) );
  OAI211_X1 U22765 ( .C1(n19788), .C2(n19795), .A(n19787), .B(n19786), .ZN(
        P2_U3171) );
  AOI22_X1 U22766 ( .A1(n19812), .A2(n19790), .B1(n19810), .B2(n19789), .ZN(
        n19794) );
  AOI22_X1 U22767 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19815), .B1(
        n19792), .B2(n19791), .ZN(n19793) );
  OAI211_X1 U22768 ( .C1(n19796), .C2(n19795), .A(n19794), .B(n19793), .ZN(
        P2_U3172) );
  AOI22_X1 U22769 ( .A1(n19812), .A2(n19798), .B1(n19810), .B2(n19797), .ZN(
        n19801) );
  AOI22_X1 U22770 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n19799), .ZN(n19800) );
  OAI211_X1 U22771 ( .C1(n19802), .C2(n19818), .A(n19801), .B(n19800), .ZN(
        P2_U3173) );
  AOI22_X1 U22772 ( .A1(n19812), .A2(n19804), .B1(n19810), .B2(n19803), .ZN(
        n19807) );
  AOI22_X1 U22773 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n19805), .ZN(n19806) );
  OAI211_X1 U22774 ( .C1(n19808), .C2(n19818), .A(n19807), .B(n19806), .ZN(
        P2_U3174) );
  AOI22_X1 U22775 ( .A1(n19812), .A2(n19811), .B1(n19810), .B2(n19809), .ZN(
        n19817) );
  AOI22_X1 U22776 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n19813), .ZN(n19816) );
  OAI211_X1 U22777 ( .C1(n19819), .C2(n19818), .A(n19817), .B(n19816), .ZN(
        P2_U3175) );
  AND2_X1 U22778 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19884), .ZN(
        P2_U3179) );
  AND2_X1 U22779 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19884), .ZN(
        P2_U3180) );
  AND2_X1 U22780 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19884), .ZN(
        P2_U3181) );
  INV_X1 U22781 ( .A(P2_DATAWIDTH_REG_28__SCAN_IN), .ZN(n20903) );
  NOR2_X1 U22782 ( .A1(n20903), .A2(n19887), .ZN(P2_U3182) );
  AND2_X1 U22783 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19884), .ZN(
        P2_U3183) );
  AND2_X1 U22784 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19884), .ZN(
        P2_U3184) );
  AND2_X1 U22785 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19884), .ZN(
        P2_U3185) );
  AND2_X1 U22786 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19884), .ZN(
        P2_U3186) );
  AND2_X1 U22787 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19884), .ZN(
        P2_U3187) );
  AND2_X1 U22788 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19884), .ZN(
        P2_U3188) );
  AND2_X1 U22789 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19884), .ZN(
        P2_U3189) );
  AND2_X1 U22790 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19884), .ZN(
        P2_U3190) );
  AND2_X1 U22791 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19884), .ZN(
        P2_U3191) );
  AND2_X1 U22792 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19884), .ZN(
        P2_U3192) );
  AND2_X1 U22793 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19884), .ZN(
        P2_U3193) );
  AND2_X1 U22794 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19884), .ZN(
        P2_U3194) );
  AND2_X1 U22795 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19884), .ZN(
        P2_U3195) );
  AND2_X1 U22796 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19884), .ZN(
        P2_U3196) );
  AND2_X1 U22797 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19884), .ZN(
        P2_U3197) );
  AND2_X1 U22798 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19884), .ZN(
        P2_U3198) );
  AND2_X1 U22799 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19884), .ZN(
        P2_U3199) );
  AND2_X1 U22800 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19884), .ZN(
        P2_U3200) );
  NOR2_X1 U22801 ( .A1(n20899), .A2(n19887), .ZN(P2_U3201) );
  NOR2_X1 U22802 ( .A1(n21051), .A2(n19887), .ZN(P2_U3202) );
  AND2_X1 U22803 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19884), .ZN(P2_U3203) );
  AND2_X1 U22804 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19884), .ZN(P2_U3204) );
  INV_X1 U22805 ( .A(P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n21037) );
  NOR2_X1 U22806 ( .A1(n21037), .A2(n19887), .ZN(P2_U3205) );
  AND2_X1 U22807 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19884), .ZN(P2_U3206) );
  AND2_X1 U22808 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19884), .ZN(P2_U3207) );
  AND2_X1 U22809 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19884), .ZN(P2_U3208) );
  NAND2_X1 U22810 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19952), .ZN(n19832) );
  NAND3_X1 U22811 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19832), .ZN(n19822) );
  AOI211_X1 U22812 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20719), .A(
        n19820), .B(n19960), .ZN(n19821) );
  INV_X1 U22813 ( .A(NA), .ZN(n20727) );
  NOR2_X1 U22814 ( .A1(n20727), .A2(n19826), .ZN(n19837) );
  AOI211_X1 U22815 ( .C1(n19838), .C2(n19822), .A(n19821), .B(n19837), .ZN(
        n19823) );
  INV_X1 U22816 ( .A(n19823), .ZN(P2_U3209) );
  INV_X1 U22817 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19824) );
  AOI21_X1 U22818 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20719), .A(n19838), 
        .ZN(n19830) );
  NOR2_X1 U22819 ( .A1(n19824), .A2(n19830), .ZN(n19827) );
  AOI21_X1 U22820 ( .B1(n19827), .B2(n19826), .A(n19825), .ZN(n19828) );
  OAI211_X1 U22821 ( .C1(n20719), .C2(n19829), .A(n19828), .B(n19832), .ZN(
        P2_U3210) );
  AOI21_X1 U22822 ( .B1(n19952), .B2(n19831), .A(n19830), .ZN(n19836) );
  OAI22_X1 U22823 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19833), .B1(NA), 
        .B2(n19832), .ZN(n19834) );
  OAI211_X1 U22824 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19834), .ZN(n19835) );
  OAI21_X1 U22825 ( .B1(n19837), .B2(n19836), .A(n19835), .ZN(P2_U3211) );
  OAI222_X1 U22826 ( .A1(n19876), .A2(n11428), .B1(n19840), .B2(n19960), .C1(
        n19839), .C2(n19875), .ZN(P2_U3212) );
  OAI222_X1 U22827 ( .A1(n19876), .A2(n11446), .B1(n19841), .B2(n19960), .C1(
        n11428), .C2(n19875), .ZN(P2_U3213) );
  OAI222_X1 U22828 ( .A1(n19876), .A2(n11992), .B1(n19842), .B2(n19960), .C1(
        n11446), .C2(n19875), .ZN(P2_U3214) );
  OAI222_X1 U22829 ( .A1(n19876), .A2(n11998), .B1(n19843), .B2(n19960), .C1(
        n11992), .C2(n19875), .ZN(P2_U3215) );
  OAI222_X1 U22830 ( .A1(n19876), .A2(n19845), .B1(n19844), .B2(n19960), .C1(
        n11998), .C2(n19875), .ZN(P2_U3216) );
  OAI222_X1 U22831 ( .A1(n19876), .A2(n12005), .B1(n19846), .B2(n19960), .C1(
        n19845), .C2(n19875), .ZN(P2_U3217) );
  OAI222_X1 U22832 ( .A1(n19876), .A2(n15340), .B1(n19847), .B2(n19960), .C1(
        n12005), .C2(n19875), .ZN(P2_U3218) );
  OAI222_X1 U22833 ( .A1(n19876), .A2(n12010), .B1(n19848), .B2(n19960), .C1(
        n15340), .C2(n19875), .ZN(P2_U3219) );
  OAI222_X1 U22834 ( .A1(n19876), .A2(n12015), .B1(n19849), .B2(n19960), .C1(
        n12010), .C2(n19875), .ZN(P2_U3220) );
  OAI222_X1 U22835 ( .A1(n19876), .A2(n12021), .B1(n19850), .B2(n19960), .C1(
        n12015), .C2(n19875), .ZN(P2_U3221) );
  OAI222_X1 U22836 ( .A1(n19876), .A2(n12024), .B1(n19851), .B2(n19960), .C1(
        n12021), .C2(n19875), .ZN(P2_U3222) );
  OAI222_X1 U22837 ( .A1(n19876), .A2(n15847), .B1(n19852), .B2(n19960), .C1(
        n12024), .C2(n19875), .ZN(P2_U3223) );
  OAI222_X1 U22838 ( .A1(n19876), .A2(n12030), .B1(n19853), .B2(n19960), .C1(
        n15847), .C2(n19875), .ZN(P2_U3224) );
  OAI222_X1 U22839 ( .A1(n19876), .A2(n15617), .B1(n19854), .B2(n19960), .C1(
        n12030), .C2(n19875), .ZN(P2_U3225) );
  OAI222_X1 U22840 ( .A1(n19876), .A2(n19856), .B1(n19855), .B2(n19960), .C1(
        n15617), .C2(n19875), .ZN(P2_U3226) );
  OAI222_X1 U22841 ( .A1(n19876), .A2(n19858), .B1(n19857), .B2(n19960), .C1(
        n19856), .C2(n19875), .ZN(P2_U3227) );
  OAI222_X1 U22842 ( .A1(n19876), .A2(n15287), .B1(n19859), .B2(n19960), .C1(
        n19858), .C2(n19875), .ZN(P2_U3228) );
  OAI222_X1 U22843 ( .A1(n19876), .A2(n12047), .B1(n19860), .B2(n19960), .C1(
        n15287), .C2(n19875), .ZN(P2_U3229) );
  OAI222_X1 U22844 ( .A1(n19876), .A2(n18980), .B1(n19861), .B2(n19960), .C1(
        n12047), .C2(n19875), .ZN(P2_U3230) );
  OAI222_X1 U22845 ( .A1(n19876), .A2(n20953), .B1(n19862), .B2(n19960), .C1(
        n18980), .C2(n19875), .ZN(P2_U3231) );
  OAI222_X1 U22846 ( .A1(n19876), .A2(n12056), .B1(n19863), .B2(n19960), .C1(
        n20953), .C2(n19875), .ZN(P2_U3232) );
  OAI222_X1 U22847 ( .A1(n19876), .A2(n12060), .B1(n19864), .B2(n19960), .C1(
        n12056), .C2(n19875), .ZN(P2_U3233) );
  OAI222_X1 U22848 ( .A1(n19876), .A2(n12064), .B1(n19865), .B2(n19960), .C1(
        n12060), .C2(n19875), .ZN(P2_U3234) );
  OAI222_X1 U22849 ( .A1(n19876), .A2(n19867), .B1(n19866), .B2(n19960), .C1(
        n12064), .C2(n19875), .ZN(P2_U3235) );
  OAI222_X1 U22850 ( .A1(n19876), .A2(n19869), .B1(n19868), .B2(n19960), .C1(
        n19867), .C2(n19875), .ZN(P2_U3236) );
  OAI222_X1 U22851 ( .A1(n19876), .A2(n19871), .B1(n20936), .B2(n19960), .C1(
        n19869), .C2(n19875), .ZN(P2_U3237) );
  OAI222_X1 U22852 ( .A1(n19875), .A2(n19871), .B1(n19870), .B2(n19960), .C1(
        n12332), .C2(n19876), .ZN(P2_U3238) );
  OAI222_X1 U22853 ( .A1(n19876), .A2(n19873), .B1(n19872), .B2(n19960), .C1(
        n12332), .C2(n19875), .ZN(P2_U3239) );
  OAI222_X1 U22854 ( .A1(n19876), .A2(n12346), .B1(n19874), .B2(n19960), .C1(
        n19873), .C2(n19875), .ZN(P2_U3240) );
  OAI222_X1 U22855 ( .A1(n19876), .A2(n21076), .B1(n20965), .B2(n19960), .C1(
        n12346), .C2(n19875), .ZN(P2_U3241) );
  INV_X1 U22856 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19877) );
  AOI22_X1 U22857 ( .A1(n19960), .A2(n19878), .B1(n19877), .B2(n19958), .ZN(
        P2_U3585) );
  MUX2_X1 U22858 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19960), .Z(P2_U3586) );
  INV_X1 U22859 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19879) );
  AOI22_X1 U22860 ( .A1(n19960), .A2(n19880), .B1(n19879), .B2(n19958), .ZN(
        P2_U3587) );
  INV_X1 U22861 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19881) );
  AOI22_X1 U22862 ( .A1(n19960), .A2(n19882), .B1(n19881), .B2(n19958), .ZN(
        P2_U3588) );
  INV_X1 U22863 ( .A(n19885), .ZN(n19883) );
  AOI21_X1 U22864 ( .B1(n19884), .B2(n20869), .A(n19883), .ZN(P2_U3591) );
  OAI21_X1 U22865 ( .B1(n19887), .B2(n19886), .A(n19885), .ZN(P2_U3592) );
  NAND2_X1 U22866 ( .A1(n19894), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19918) );
  OR2_X1 U22867 ( .A1(n19888), .A2(n19918), .ZN(n19910) );
  NAND2_X1 U22868 ( .A1(n19890), .A2(n19889), .ZN(n19891) );
  AOI21_X1 U22869 ( .B1(n19915), .B2(n19894), .A(n19891), .ZN(n19904) );
  NAND2_X1 U22870 ( .A1(n19910), .A2(n19904), .ZN(n19893) );
  NAND2_X1 U22871 ( .A1(n19893), .A2(n19892), .ZN(n19899) );
  NAND2_X1 U22872 ( .A1(n19895), .A2(n19894), .ZN(n19897) );
  OR2_X1 U22873 ( .A1(n19897), .A2(n19896), .ZN(n19898) );
  OAI211_X1 U22874 ( .C1(n19757), .C2(n19900), .A(n19899), .B(n19898), .ZN(
        n19901) );
  INV_X1 U22875 ( .A(n19901), .ZN(n19902) );
  INV_X1 U22876 ( .A(n19932), .ZN(n19929) );
  AOI22_X1 U22877 ( .A1(n19932), .A2(n19903), .B1(n19902), .B2(n19929), .ZN(
        P2_U3602) );
  INV_X1 U22878 ( .A(n19904), .ZN(n19908) );
  NOR2_X1 U22879 ( .A1(n19905), .A2(n19757), .ZN(n19906) );
  AOI21_X1 U22880 ( .B1(n19908), .B2(n19907), .A(n19906), .ZN(n19909) );
  AND2_X1 U22881 ( .A1(n19910), .A2(n19909), .ZN(n19911) );
  AOI22_X1 U22882 ( .A1(n19932), .A2(n19912), .B1(n19911), .B2(n19929), .ZN(
        P2_U3603) );
  INV_X1 U22883 ( .A(n19913), .ZN(n19924) );
  AND2_X1 U22884 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19914) );
  OR3_X1 U22885 ( .A1(n19915), .A2(n19924), .A3(n19914), .ZN(n19916) );
  OAI21_X1 U22886 ( .B1(n19918), .B2(n19917), .A(n19916), .ZN(n19919) );
  AOI21_X1 U22887 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19920), .A(n19919), 
        .ZN(n19921) );
  AOI22_X1 U22888 ( .A1(n19932), .A2(n19922), .B1(n19921), .B2(n19929), .ZN(
        P2_U3604) );
  NAND2_X1 U22889 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19931), .ZN(n19923) );
  OAI21_X1 U22890 ( .B1(n19925), .B2(n19924), .A(n19923), .ZN(n19926) );
  AOI21_X1 U22891 ( .B1(n19928), .B2(n19927), .A(n19926), .ZN(n19930) );
  AOI22_X1 U22892 ( .A1(n19932), .A2(n19931), .B1(n19930), .B2(n19929), .ZN(
        P2_U3605) );
  AOI22_X1 U22893 ( .A1(n19960), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19933), 
        .B2(n19958), .ZN(P2_U3608) );
  INV_X1 U22894 ( .A(n19934), .ZN(n19940) );
  AOI21_X1 U22895 ( .B1(n19937), .B2(n19936), .A(n19935), .ZN(n19939) );
  NAND2_X1 U22896 ( .A1(n19940), .A2(P2_MORE_REG_SCAN_IN), .ZN(n19938) );
  OAI21_X1 U22897 ( .B1(n19940), .B2(n19939), .A(n19938), .ZN(P2_U3609) );
  OAI21_X1 U22898 ( .B1(n19941), .B2(n19942), .A(n11376), .ZN(n19946) );
  NAND3_X1 U22899 ( .A1(n19943), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n19942), 
        .ZN(n19945) );
  MUX2_X1 U22900 ( .A(n19946), .B(n19945), .S(n19944), .Z(n19950) );
  INV_X1 U22901 ( .A(n19947), .ZN(n19948) );
  OAI21_X1 U22902 ( .B1(n19952), .B2(n19685), .A(n19948), .ZN(n19949) );
  NAND2_X1 U22903 ( .A1(n19950), .A2(n19949), .ZN(n19957) );
  NOR2_X1 U22904 ( .A1(n19952), .A2(n19951), .ZN(n19954) );
  AOI211_X1 U22905 ( .C1(n19757), .C2(n19955), .A(n19954), .B(n19953), .ZN(
        n19956) );
  MUX2_X1 U22906 ( .A(n19957), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n19956), 
        .Z(P2_U3610) );
  INV_X1 U22907 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n19959) );
  AOI22_X1 U22908 ( .A1(n19960), .A2(n21023), .B1(n19959), .B2(n19958), .ZN(
        P2_U3611) );
  AND2_X1 U22909 ( .A1(n20723), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n19962) );
  INV_X1 U22910 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19961) );
  NAND2_X1 U22911 ( .A1(n12916), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20807) );
  INV_X2 U22912 ( .A(n20807), .ZN(n20809) );
  AOI21_X1 U22913 ( .B1(n19962), .B2(n19961), .A(n20809), .ZN(P1_U2802) );
  INV_X1 U22914 ( .A(n19963), .ZN(n19965) );
  OAI21_X1 U22915 ( .B1(n19965), .B2(n19964), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19966) );
  OAI21_X1 U22916 ( .B1(n19967), .B2(n20815), .A(n19966), .ZN(P1_U2803) );
  NOR2_X1 U22917 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19969) );
  OAI21_X1 U22918 ( .B1(n19969), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20807), .ZN(
        n19968) );
  OAI21_X1 U22919 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20807), .A(n19968), 
        .ZN(P1_U2804) );
  AOI21_X1 U22920 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20723), .A(n20809), 
        .ZN(n20798) );
  OAI21_X1 U22921 ( .B1(BS16), .B2(n19969), .A(n20798), .ZN(n20796) );
  OAI21_X1 U22922 ( .B1(n20798), .B2(n20812), .A(n20796), .ZN(P1_U2805) );
  OAI21_X1 U22923 ( .B1(n19972), .B2(n19971), .A(n19970), .ZN(P1_U2806) );
  NOR4_X1 U22924 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19976) );
  NOR4_X1 U22925 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_14__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19975) );
  NOR4_X1 U22926 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_27__SCAN_IN), .A3(P1_DATAWIDTH_REG_28__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_29__SCAN_IN), .ZN(n19974) );
  NOR4_X1 U22927 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19973) );
  NAND4_X1 U22928 ( .A1(n19976), .A2(n19975), .A3(n19974), .A4(n19973), .ZN(
        n19982) );
  NOR4_X1 U22929 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_2__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n19980) );
  AOI211_X1 U22930 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_13__SCAN_IN), .B(
        P1_DATAWIDTH_REG_16__SCAN_IN), .ZN(n19979) );
  NOR4_X1 U22931 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_10__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_12__SCAN_IN), .ZN(n19978) );
  NOR4_X1 U22932 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_6__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(n19977) );
  NAND4_X1 U22933 ( .A1(n19980), .A2(n19979), .A3(n19978), .A4(n19977), .ZN(
        n19981) );
  NOR2_X1 U22934 ( .A1(n19982), .A2(n19981), .ZN(n20806) );
  INV_X1 U22935 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20793) );
  NOR3_X1 U22936 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19984) );
  OAI21_X1 U22937 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19984), .A(n20806), .ZN(
        n19983) );
  OAI21_X1 U22938 ( .B1(n20806), .B2(n20793), .A(n19983), .ZN(P1_U2807) );
  INV_X1 U22939 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20790) );
  NOR2_X1 U22940 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20801) );
  OAI21_X1 U22941 ( .B1(n19984), .B2(n20801), .A(n20806), .ZN(n19985) );
  OAI21_X1 U22942 ( .B1(n20806), .B2(n20790), .A(n19985), .ZN(P1_U2808) );
  NAND2_X1 U22943 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20007) );
  NOR4_X1 U22944 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20745), .A3(n20007), .A4(
        n20028), .ZN(n19992) );
  AOI22_X1 U22945 ( .A1(n19986), .A2(n20039), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n20041), .ZN(n19989) );
  AOI21_X1 U22946 ( .B1(n20042), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n19987), .ZN(n19988) );
  OAI211_X1 U22947 ( .C1(n19990), .C2(n20053), .A(n19989), .B(n19988), .ZN(
        n19991) );
  AOI211_X1 U22948 ( .C1(n19993), .C2(n20018), .A(n19992), .B(n19991), .ZN(
        n19994) );
  OAI21_X1 U22949 ( .B1(n19995), .B2(n20746), .A(n19994), .ZN(P1_U2832) );
  OAI21_X1 U22950 ( .B1(n20007), .B2(n19997), .A(n19996), .ZN(n20022) );
  OAI21_X1 U22951 ( .B1(n19999), .B2(n19998), .A(n20043), .ZN(n20004) );
  OAI22_X1 U22952 ( .A1(n20002), .A2(n20030), .B1(n20001), .B2(n20000), .ZN(
        n20003) );
  AOI211_X1 U22953 ( .C1(n20024), .C2(n20005), .A(n20004), .B(n20003), .ZN(
        n20011) );
  INV_X1 U22954 ( .A(n20006), .ZN(n20009) );
  NOR2_X1 U22955 ( .A1(n20007), .A2(n20028), .ZN(n20008) );
  AOI22_X1 U22956 ( .A1(n20009), .A2(n20018), .B1(n20745), .B2(n20008), .ZN(
        n20010) );
  OAI211_X1 U22957 ( .C1(n20745), .C2(n20022), .A(n20011), .B(n20010), .ZN(
        P1_U2833) );
  INV_X1 U22958 ( .A(n20012), .ZN(n20017) );
  NOR3_X1 U22959 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20742), .A3(n20028), .ZN(
        n20016) );
  AOI22_X1 U22960 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20042), .B1(
        P1_EBX_REG_6__SCAN_IN), .B2(n20041), .ZN(n20013) );
  OAI211_X1 U22961 ( .C1(n20053), .C2(n20014), .A(n20013), .B(n20043), .ZN(
        n20015) );
  AOI211_X1 U22962 ( .C1(n20039), .C2(n20017), .A(n20016), .B(n20015), .ZN(
        n20021) );
  NAND2_X1 U22963 ( .A1(n20019), .A2(n20018), .ZN(n20020) );
  OAI211_X1 U22964 ( .C1(n20022), .C2(n13658), .A(n20021), .B(n20020), .ZN(
        P1_U2834) );
  AOI22_X1 U22965 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n20041), .B1(n20024), .B2(
        n20023), .ZN(n20025) );
  NAND2_X1 U22966 ( .A1(n20043), .A2(n20025), .ZN(n20026) );
  AOI21_X1 U22967 ( .B1(n20042), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n20026), .ZN(n20027) );
  OAI21_X1 U22968 ( .B1(n20028), .B2(P1_REIP_REG_5__SCAN_IN), .A(n20027), .ZN(
        n20032) );
  NOR2_X1 U22969 ( .A1(n20030), .A2(n20029), .ZN(n20031) );
  AOI211_X1 U22970 ( .C1(n20033), .C2(n20048), .A(n20032), .B(n20031), .ZN(
        n20034) );
  OAI21_X1 U22971 ( .B1(n20742), .B2(n20045), .A(n20034), .ZN(P1_U2835) );
  INV_X1 U22972 ( .A(n20035), .ZN(n20038) );
  AOI22_X1 U22973 ( .A1(n20039), .A2(n20038), .B1(n20037), .B2(n20036), .ZN(
        n20051) );
  NOR2_X1 U22974 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20040), .ZN(n20046) );
  AOI22_X1 U22975 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n20042), .B1(
        P1_EBX_REG_4__SCAN_IN), .B2(n20041), .ZN(n20044) );
  OAI211_X1 U22976 ( .C1(n20046), .C2(n20045), .A(n20044), .B(n20043), .ZN(
        n20047) );
  AOI21_X1 U22977 ( .B1(n20049), .B2(n20048), .A(n20047), .ZN(n20050) );
  OAI211_X1 U22978 ( .C1(n20053), .C2(n20052), .A(n20051), .B(n20050), .ZN(
        P1_U2836) );
  AOI22_X1 U22979 ( .A1(n20083), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n13252), .ZN(n20056) );
  INV_X1 U22980 ( .A(n20054), .ZN(n20055) );
  NAND2_X1 U22981 ( .A1(n20071), .A2(n20055), .ZN(n20073) );
  NAND2_X1 U22982 ( .A1(n20056), .A2(n20073), .ZN(P1_U2945) );
  AOI22_X1 U22983 ( .A1(n20083), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n13252), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n20059) );
  INV_X1 U22984 ( .A(n20057), .ZN(n20058) );
  NAND2_X1 U22985 ( .A1(n20071), .A2(n20058), .ZN(n20075) );
  NAND2_X1 U22986 ( .A1(n20059), .A2(n20075), .ZN(P1_U2946) );
  AOI22_X1 U22987 ( .A1(n20083), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n13252), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20062) );
  INV_X1 U22988 ( .A(n20060), .ZN(n20061) );
  NAND2_X1 U22989 ( .A1(n20071), .A2(n20061), .ZN(n20077) );
  NAND2_X1 U22990 ( .A1(n20062), .A2(n20077), .ZN(P1_U2947) );
  AOI22_X1 U22991 ( .A1(n20083), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n13252), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20065) );
  INV_X1 U22992 ( .A(n20063), .ZN(n20064) );
  NAND2_X1 U22993 ( .A1(n20071), .A2(n20064), .ZN(n20079) );
  NAND2_X1 U22994 ( .A1(n20065), .A2(n20079), .ZN(P1_U2949) );
  AOI22_X1 U22995 ( .A1(n20083), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n13252), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20068) );
  INV_X1 U22996 ( .A(n20066), .ZN(n20067) );
  NAND2_X1 U22997 ( .A1(n20071), .A2(n20067), .ZN(n20081) );
  NAND2_X1 U22998 ( .A1(n20068), .A2(n20081), .ZN(P1_U2950) );
  AOI22_X1 U22999 ( .A1(n20083), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n13252), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20072) );
  INV_X1 U23000 ( .A(n20069), .ZN(n20070) );
  NAND2_X1 U23001 ( .A1(n20071), .A2(n20070), .ZN(n20084) );
  NAND2_X1 U23002 ( .A1(n20072), .A2(n20084), .ZN(P1_U2951) );
  AOI22_X1 U23003 ( .A1(n20083), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n13252), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n20074) );
  NAND2_X1 U23004 ( .A1(n20074), .A2(n20073), .ZN(P1_U2960) );
  AOI22_X1 U23005 ( .A1(n20083), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n13252), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20076) );
  NAND2_X1 U23006 ( .A1(n20076), .A2(n20075), .ZN(P1_U2961) );
  AOI22_X1 U23007 ( .A1(n20083), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n13252), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20078) );
  NAND2_X1 U23008 ( .A1(n20078), .A2(n20077), .ZN(P1_U2962) );
  AOI22_X1 U23009 ( .A1(n20083), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n13252), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20080) );
  NAND2_X1 U23010 ( .A1(n20080), .A2(n20079), .ZN(P1_U2964) );
  AOI22_X1 U23011 ( .A1(n20083), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n13252), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20082) );
  NAND2_X1 U23012 ( .A1(n20082), .A2(n20081), .ZN(P1_U2965) );
  AOI22_X1 U23013 ( .A1(n20083), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n13252), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20085) );
  NAND2_X1 U23014 ( .A1(n20085), .A2(n20084), .ZN(P1_U2966) );
  NAND2_X1 U23015 ( .A1(n20086), .A2(n20095), .ZN(n20090) );
  AOI21_X1 U23016 ( .B1(n20088), .B2(n20116), .A(n20087), .ZN(n20089) );
  OAI211_X1 U23017 ( .C1(n20092), .C2(n20091), .A(n20090), .B(n20089), .ZN(
        n20093) );
  INV_X1 U23018 ( .A(n20093), .ZN(n20094) );
  OAI21_X1 U23019 ( .B1(n20096), .B2(n20095), .A(n20094), .ZN(P1_U3028) );
  INV_X1 U23020 ( .A(n20097), .ZN(n20098) );
  AOI21_X1 U23021 ( .B1(n11153), .B2(n20099), .A(n20098), .ZN(n20112) );
  NOR2_X1 U23022 ( .A1(n20100), .A2(n11153), .ZN(n20102) );
  AOI21_X1 U23023 ( .B1(n20102), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n20101), .ZN(n20103) );
  NOR2_X1 U23024 ( .A1(n20104), .A2(n20103), .ZN(n20109) );
  OAI21_X1 U23025 ( .B1(n20107), .B2(n20106), .A(n20105), .ZN(n20108) );
  AOI211_X1 U23026 ( .C1(n20110), .C2(n20117), .A(n20109), .B(n20108), .ZN(
        n20111) );
  OAI221_X1 U23027 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20113), .C1(
        n10996), .C2(n20112), .A(n20111), .ZN(P1_U3029) );
  INV_X1 U23028 ( .A(n20114), .ZN(n20115) );
  AOI22_X1 U23029 ( .A1(n20118), .A2(n20117), .B1(n20116), .B2(n20115), .ZN(
        n20124) );
  INV_X1 U23030 ( .A(n20119), .ZN(n20120) );
  OAI22_X1 U23031 ( .A1(n20122), .A2(n20121), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n20120), .ZN(n20123) );
  OAI211_X1 U23032 ( .C1(n20125), .C2(n16200), .A(n20124), .B(n20123), .ZN(
        P1_U3031) );
  NOR2_X1 U23033 ( .A1(n20127), .A2(n20126), .ZN(P1_U3032) );
  NOR2_X2 U23034 ( .A1(n20129), .A2(n20128), .ZN(n20171) );
  AOI22_X1 U23035 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20171), .B1(DATAI_16_), 
        .B2(n20131), .ZN(n20616) );
  INV_X1 U23036 ( .A(n13485), .ZN(n20132) );
  AOI22_X1 U23037 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20171), .B1(DATAI_24_), 
        .B2(n20131), .ZN(n20666) );
  INV_X1 U23038 ( .A(n20666), .ZN(n20613) );
  NAND2_X1 U23039 ( .A1(n20172), .A2(n20135), .ZN(n20460) );
  NAND3_X1 U23040 ( .A1(n21022), .A2(n20459), .A3(n20541), .ZN(n20181) );
  NOR2_X1 U23041 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20181), .ZN(
        n20173) );
  AOI22_X1 U23042 ( .A1(n20708), .A2(n20613), .B1(n20655), .B2(n20173), .ZN(
        n20150) );
  INV_X1 U23043 ( .A(n20466), .ZN(n20136) );
  NOR2_X1 U23044 ( .A1(n20136), .A2(n20407), .ZN(n20146) );
  NOR2_X1 U23045 ( .A1(n20144), .A2(n20811), .ZN(n20286) );
  INV_X1 U23046 ( .A(n20708), .ZN(n20137) );
  NAND3_X1 U23047 ( .A1(n20137), .A2(n20206), .A3(n20661), .ZN(n20138) );
  NAND2_X1 U23048 ( .A1(n20661), .A2(n20812), .ZN(n20543) );
  NAND2_X1 U23049 ( .A1(n20138), .A2(n20543), .ZN(n20143) );
  OR2_X1 U23050 ( .A1(n20406), .A2(n20139), .ZN(n20179) );
  INV_X1 U23051 ( .A(n20464), .ZN(n20603) );
  OR2_X1 U23052 ( .A1(n20179), .A2(n20603), .ZN(n20147) );
  INV_X1 U23053 ( .A(n20173), .ZN(n20140) );
  AOI22_X1 U23054 ( .A1(n20143), .A2(n20147), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20140), .ZN(n20141) );
  OAI211_X1 U23055 ( .C1(n20146), .C2(n20811), .A(n20469), .B(n20141), .ZN(
        n20176) );
  NOR2_X2 U23056 ( .A1(n20142), .A2(n20291), .ZN(n20654) );
  INV_X1 U23057 ( .A(n20143), .ZN(n20148) );
  INV_X1 U23058 ( .A(n20144), .ZN(n20145) );
  NOR2_X1 U23059 ( .A1(n20145), .A2(n20811), .ZN(n20292) );
  INV_X1 U23060 ( .A(n20292), .ZN(n20472) );
  INV_X1 U23061 ( .A(n20146), .ZN(n20287) );
  AOI22_X1 U23062 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20176), .B1(
        n20654), .B2(n20175), .ZN(n20149) );
  OAI211_X1 U23063 ( .C1(n20616), .C2(n20206), .A(n20150), .B(n20149), .ZN(
        P1_U3033) );
  AOI22_X1 U23064 ( .A1(DATAI_25_), .A2(n20131), .B1(BUF1_REG_25__SCAN_IN), 
        .B2(n20171), .ZN(n20672) );
  INV_X1 U23065 ( .A(n20672), .ZN(n20617) );
  AOI22_X1 U23066 ( .A1(n20708), .A2(n20617), .B1(n20668), .B2(n20173), .ZN(
        n20153) );
  NOR2_X2 U23067 ( .A1(n20151), .A2(n20291), .ZN(n20667) );
  AOI22_X1 U23068 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20176), .B1(
        n20667), .B2(n20175), .ZN(n20152) );
  OAI211_X1 U23069 ( .C1(n20620), .C2(n20206), .A(n20153), .B(n20152), .ZN(
        P1_U3034) );
  AOI22_X1 U23070 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20171), .B1(DATAI_18_), 
        .B2(n20131), .ZN(n20624) );
  AOI22_X1 U23071 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20171), .B1(DATAI_26_), 
        .B2(n20131), .ZN(n20678) );
  INV_X1 U23072 ( .A(n20678), .ZN(n20621) );
  NAND2_X1 U23073 ( .A1(n20172), .A2(n10423), .ZN(n20481) );
  AOI22_X1 U23074 ( .A1(n20708), .A2(n20621), .B1(n20674), .B2(n20173), .ZN(
        n20156) );
  NOR2_X2 U23075 ( .A1(n20154), .A2(n20291), .ZN(n20673) );
  AOI22_X1 U23076 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20176), .B1(
        n20673), .B2(n20175), .ZN(n20155) );
  OAI211_X1 U23077 ( .C1(n20624), .C2(n20206), .A(n20156), .B(n20155), .ZN(
        P1_U3035) );
  AOI22_X1 U23078 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20171), .B1(DATAI_19_), 
        .B2(n20131), .ZN(n20628) );
  AOI22_X1 U23079 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20171), .B1(DATAI_27_), 
        .B2(n20131), .ZN(n20684) );
  INV_X1 U23080 ( .A(n20684), .ZN(n20625) );
  NAND2_X1 U23081 ( .A1(n20172), .A2(n20157), .ZN(n20485) );
  AOI22_X1 U23082 ( .A1(n20708), .A2(n20625), .B1(n20680), .B2(n20173), .ZN(
        n20160) );
  NOR2_X2 U23083 ( .A1(n20158), .A2(n20291), .ZN(n20679) );
  AOI22_X1 U23084 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20176), .B1(
        n20679), .B2(n20175), .ZN(n20159) );
  OAI211_X1 U23085 ( .C1(n20628), .C2(n20206), .A(n20160), .B(n20159), .ZN(
        P1_U3036) );
  AOI22_X1 U23086 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20171), .B1(DATAI_20_), 
        .B2(n20131), .ZN(n20632) );
  AOI22_X1 U23087 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20171), .B1(DATAI_28_), 
        .B2(n20131), .ZN(n20690) );
  INV_X1 U23088 ( .A(n20690), .ZN(n20629) );
  NAND2_X1 U23089 ( .A1(n20172), .A2(n20161), .ZN(n20489) );
  AOI22_X1 U23090 ( .A1(n20708), .A2(n20629), .B1(n20686), .B2(n20173), .ZN(
        n20164) );
  NOR2_X2 U23091 ( .A1(n20291), .A2(n20162), .ZN(n20685) );
  AOI22_X1 U23092 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20176), .B1(
        n20685), .B2(n20175), .ZN(n20163) );
  OAI211_X1 U23093 ( .C1(n20632), .C2(n20206), .A(n20164), .B(n20163), .ZN(
        P1_U3037) );
  AOI22_X1 U23094 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20171), .B1(DATAI_21_), 
        .B2(n20131), .ZN(n20636) );
  AOI22_X1 U23095 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20171), .B1(DATAI_29_), 
        .B2(n20131), .ZN(n20696) );
  INV_X1 U23096 ( .A(n20696), .ZN(n20633) );
  NAND2_X1 U23097 ( .A1(n20172), .A2(n10388), .ZN(n20493) );
  AOI22_X1 U23098 ( .A1(n20708), .A2(n20633), .B1(n20692), .B2(n20173), .ZN(
        n20167) );
  NOR2_X2 U23099 ( .A1(n20291), .A2(n20165), .ZN(n20691) );
  AOI22_X1 U23100 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20176), .B1(
        n20691), .B2(n20175), .ZN(n20166) );
  OAI211_X1 U23101 ( .C1(n20636), .C2(n20206), .A(n20167), .B(n20166), .ZN(
        P1_U3038) );
  AOI22_X1 U23102 ( .A1(DATAI_22_), .A2(n20131), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20171), .ZN(n20640) );
  AOI22_X1 U23103 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20171), .B1(DATAI_30_), 
        .B2(n20131), .ZN(n20702) );
  INV_X1 U23104 ( .A(n20702), .ZN(n20637) );
  NAND2_X1 U23105 ( .A1(n20172), .A2(n21125), .ZN(n20497) );
  AOI22_X1 U23106 ( .A1(n20708), .A2(n20637), .B1(n20698), .B2(n20173), .ZN(
        n20170) );
  NOR2_X2 U23107 ( .A1(n20291), .A2(n20168), .ZN(n20697) );
  AOI22_X1 U23108 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20176), .B1(
        n20697), .B2(n20175), .ZN(n20169) );
  OAI211_X1 U23109 ( .C1(n20640), .C2(n20206), .A(n20170), .B(n20169), .ZN(
        P1_U3039) );
  AOI22_X1 U23110 ( .A1(DATAI_23_), .A2(n20131), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n20171), .ZN(n20648) );
  AOI22_X1 U23111 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20171), .B1(DATAI_31_), 
        .B2(n20131), .ZN(n20713) );
  INV_X1 U23112 ( .A(n20713), .ZN(n20643) );
  NAND2_X1 U23113 ( .A1(n20172), .A2(n10389), .ZN(n20501) );
  AOI22_X1 U23114 ( .A1(n20708), .A2(n20643), .B1(n20706), .B2(n20173), .ZN(
        n20178) );
  NOR2_X2 U23115 ( .A1(n20291), .A2(n20174), .ZN(n20704) );
  AOI22_X1 U23116 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20176), .B1(
        n20704), .B2(n20175), .ZN(n20177) );
  OAI211_X1 U23117 ( .C1(n20648), .C2(n20206), .A(n20178), .B(n20177), .ZN(
        P1_U3040) );
  NOR2_X1 U23118 ( .A1(n20573), .A2(n20181), .ZN(n20201) );
  INV_X1 U23119 ( .A(n20180), .ZN(n20575) );
  AOI21_X1 U23120 ( .B1(n20248), .B2(n20575), .A(n20201), .ZN(n20182) );
  OAI22_X1 U23121 ( .A1(n20182), .A2(n20653), .B1(n20181), .B2(n20811), .ZN(
        n20200) );
  AOI22_X1 U23122 ( .A1(n20655), .A2(n20201), .B1(n20200), .B2(n20654), .ZN(
        n20186) );
  INV_X1 U23123 ( .A(n20181), .ZN(n20184) );
  INV_X1 U23124 ( .A(n20543), .ZN(n20578) );
  OAI21_X1 U23125 ( .B1(n20242), .B2(n20578), .A(n20182), .ZN(n20183) );
  OAI211_X1 U23126 ( .C1(n20661), .C2(n20184), .A(n20660), .B(n20183), .ZN(
        n20203) );
  INV_X1 U23127 ( .A(n20236), .ZN(n20202) );
  INV_X1 U23128 ( .A(n20616), .ZN(n20663) );
  AOI22_X1 U23129 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20663), .ZN(n20185) );
  OAI211_X1 U23130 ( .C1(n20666), .C2(n20206), .A(n20186), .B(n20185), .ZN(
        P1_U3041) );
  AOI22_X1 U23131 ( .A1(n20668), .A2(n20201), .B1(n20200), .B2(n20667), .ZN(
        n20188) );
  INV_X1 U23132 ( .A(n20206), .ZN(n20193) );
  AOI22_X1 U23133 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20203), .B1(
        n20193), .B2(n20617), .ZN(n20187) );
  OAI211_X1 U23134 ( .C1(n20620), .C2(n20236), .A(n20188), .B(n20187), .ZN(
        P1_U3042) );
  AOI22_X1 U23135 ( .A1(n20674), .A2(n20201), .B1(n20200), .B2(n20673), .ZN(
        n20190) );
  AOI22_X1 U23136 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20203), .B1(
        n20193), .B2(n20621), .ZN(n20189) );
  OAI211_X1 U23137 ( .C1(n20624), .C2(n20236), .A(n20190), .B(n20189), .ZN(
        P1_U3043) );
  AOI22_X1 U23138 ( .A1(n20680), .A2(n20201), .B1(n20200), .B2(n20679), .ZN(
        n20192) );
  INV_X1 U23139 ( .A(n20628), .ZN(n20681) );
  AOI22_X1 U23140 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20681), .ZN(n20191) );
  OAI211_X1 U23141 ( .C1(n20684), .C2(n20206), .A(n20192), .B(n20191), .ZN(
        P1_U3044) );
  AOI22_X1 U23142 ( .A1(n20686), .A2(n20201), .B1(n20685), .B2(n20200), .ZN(
        n20195) );
  AOI22_X1 U23143 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20203), .B1(
        n20193), .B2(n20629), .ZN(n20194) );
  OAI211_X1 U23144 ( .C1(n20632), .C2(n20236), .A(n20195), .B(n20194), .ZN(
        P1_U3045) );
  AOI22_X1 U23145 ( .A1(n20692), .A2(n20201), .B1(n20691), .B2(n20200), .ZN(
        n20197) );
  INV_X1 U23146 ( .A(n20636), .ZN(n20693) );
  AOI22_X1 U23147 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20693), .ZN(n20196) );
  OAI211_X1 U23148 ( .C1(n20696), .C2(n20206), .A(n20197), .B(n20196), .ZN(
        P1_U3046) );
  AOI22_X1 U23149 ( .A1(n20698), .A2(n20201), .B1(n20697), .B2(n20200), .ZN(
        n20199) );
  INV_X1 U23150 ( .A(n20640), .ZN(n20699) );
  AOI22_X1 U23151 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20699), .ZN(n20198) );
  OAI211_X1 U23152 ( .C1(n20702), .C2(n20206), .A(n20199), .B(n20198), .ZN(
        P1_U3047) );
  AOI22_X1 U23153 ( .A1(n20706), .A2(n20201), .B1(n20704), .B2(n20200), .ZN(
        n20205) );
  INV_X1 U23154 ( .A(n20648), .ZN(n20707) );
  AOI22_X1 U23155 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20707), .ZN(n20204) );
  OAI211_X1 U23156 ( .C1(n20713), .C2(n20206), .A(n20205), .B(n20204), .ZN(
        P1_U3048) );
  NAND3_X1 U23157 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21022), .A3(
        n20459), .ZN(n20254) );
  OR2_X1 U23158 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20254), .ZN(
        n20235) );
  OAI22_X1 U23159 ( .A1(n20284), .A2(n20616), .B1(n20460), .B2(n20235), .ZN(
        n20209) );
  INV_X1 U23160 ( .A(n20209), .ZN(n20216) );
  NAND2_X1 U23161 ( .A1(n20284), .A2(n20236), .ZN(n20210) );
  AOI21_X1 U23162 ( .B1(n20210), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20653), 
        .ZN(n20212) );
  NAND2_X1 U23163 ( .A1(n20248), .A2(n20603), .ZN(n20213) );
  AOI22_X1 U23164 ( .A1(n20212), .A2(n20213), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20235), .ZN(n20211) );
  OR2_X1 U23165 ( .A1(n20466), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20345) );
  NAND2_X1 U23166 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20345), .ZN(n20342) );
  NAND3_X1 U23167 ( .A1(n20469), .A2(n20211), .A3(n20342), .ZN(n20239) );
  INV_X1 U23168 ( .A(n20212), .ZN(n20214) );
  AOI22_X1 U23169 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20239), .B1(
        n20654), .B2(n20238), .ZN(n20215) );
  OAI211_X1 U23170 ( .C1(n20666), .C2(n20236), .A(n20216), .B(n20215), .ZN(
        P1_U3049) );
  OAI22_X1 U23171 ( .A1(n20284), .A2(n20620), .B1(n20477), .B2(n20235), .ZN(
        n20217) );
  INV_X1 U23172 ( .A(n20217), .ZN(n20219) );
  AOI22_X1 U23173 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20239), .B1(
        n20667), .B2(n20238), .ZN(n20218) );
  OAI211_X1 U23174 ( .C1(n20672), .C2(n20236), .A(n20219), .B(n20218), .ZN(
        P1_U3050) );
  OAI22_X1 U23175 ( .A1(n20284), .A2(n20624), .B1(n20481), .B2(n20235), .ZN(
        n20220) );
  INV_X1 U23176 ( .A(n20220), .ZN(n20222) );
  AOI22_X1 U23177 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20239), .B1(
        n20673), .B2(n20238), .ZN(n20221) );
  OAI211_X1 U23178 ( .C1(n20678), .C2(n20236), .A(n20222), .B(n20221), .ZN(
        P1_U3051) );
  OAI22_X1 U23179 ( .A1(n20284), .A2(n20628), .B1(n20485), .B2(n20235), .ZN(
        n20223) );
  INV_X1 U23180 ( .A(n20223), .ZN(n20225) );
  AOI22_X1 U23181 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20239), .B1(
        n20679), .B2(n20238), .ZN(n20224) );
  OAI211_X1 U23182 ( .C1(n20684), .C2(n20236), .A(n20225), .B(n20224), .ZN(
        P1_U3052) );
  OAI22_X1 U23183 ( .A1(n20284), .A2(n20632), .B1(n20489), .B2(n20235), .ZN(
        n20226) );
  INV_X1 U23184 ( .A(n20226), .ZN(n20228) );
  AOI22_X1 U23185 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20239), .B1(
        n20685), .B2(n20238), .ZN(n20227) );
  OAI211_X1 U23186 ( .C1(n20690), .C2(n20236), .A(n20228), .B(n20227), .ZN(
        P1_U3053) );
  OAI22_X1 U23187 ( .A1(n20236), .A2(n20696), .B1(n20493), .B2(n20235), .ZN(
        n20229) );
  INV_X1 U23188 ( .A(n20229), .ZN(n20231) );
  AOI22_X1 U23189 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20239), .B1(
        n20691), .B2(n20238), .ZN(n20230) );
  OAI211_X1 U23190 ( .C1(n20636), .C2(n20284), .A(n20231), .B(n20230), .ZN(
        P1_U3054) );
  OAI22_X1 U23191 ( .A1(n20236), .A2(n20702), .B1(n20497), .B2(n20235), .ZN(
        n20232) );
  INV_X1 U23192 ( .A(n20232), .ZN(n20234) );
  AOI22_X1 U23193 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20239), .B1(
        n20697), .B2(n20238), .ZN(n20233) );
  OAI211_X1 U23194 ( .C1(n20640), .C2(n20284), .A(n20234), .B(n20233), .ZN(
        P1_U3055) );
  OAI22_X1 U23195 ( .A1(n20236), .A2(n20713), .B1(n20501), .B2(n20235), .ZN(
        n20237) );
  INV_X1 U23196 ( .A(n20237), .ZN(n20241) );
  AOI22_X1 U23197 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20239), .B1(
        n20704), .B2(n20238), .ZN(n20240) );
  OAI211_X1 U23198 ( .C1(n20648), .C2(n20284), .A(n20241), .B(n20240), .ZN(
        P1_U3056) );
  NOR2_X2 U23199 ( .A1(n20242), .A2(n20509), .ZN(n20310) );
  INV_X1 U23200 ( .A(n20310), .ZN(n20277) );
  INV_X1 U23201 ( .A(n20511), .ZN(n20243) );
  NAND2_X1 U23202 ( .A1(n20243), .A2(n21022), .ZN(n20278) );
  OAI22_X1 U23203 ( .A1(n20284), .A2(n20666), .B1(n20460), .B2(n20278), .ZN(
        n20244) );
  INV_X1 U23204 ( .A(n20244), .ZN(n20258) );
  NOR2_X1 U23205 ( .A1(n20246), .A2(n20245), .ZN(n20650) );
  INV_X1 U23206 ( .A(n20278), .ZN(n20247) );
  AOI21_X1 U23207 ( .B1(n20248), .B2(n20650), .A(n20247), .ZN(n20256) );
  INV_X1 U23208 ( .A(n20249), .ZN(n20250) );
  AOI21_X1 U23209 ( .B1(n20251), .B2(n20250), .A(n20653), .ZN(n20253) );
  AOI22_X1 U23210 ( .A1(n20256), .A2(n20253), .B1(n20653), .B2(n20254), .ZN(
        n20252) );
  NAND2_X1 U23211 ( .A1(n20660), .A2(n20252), .ZN(n20281) );
  INV_X1 U23212 ( .A(n20253), .ZN(n20255) );
  OAI22_X1 U23213 ( .A1(n20256), .A2(n20255), .B1(n20811), .B2(n20254), .ZN(
        n20280) );
  AOI22_X1 U23214 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20281), .B1(
        n20654), .B2(n20280), .ZN(n20257) );
  OAI211_X1 U23215 ( .C1(n20616), .C2(n20277), .A(n20258), .B(n20257), .ZN(
        P1_U3057) );
  OAI22_X1 U23216 ( .A1(n20284), .A2(n20672), .B1(n20477), .B2(n20278), .ZN(
        n20259) );
  INV_X1 U23217 ( .A(n20259), .ZN(n20261) );
  AOI22_X1 U23218 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20281), .B1(
        n20667), .B2(n20280), .ZN(n20260) );
  OAI211_X1 U23219 ( .C1(n20620), .C2(n20277), .A(n20261), .B(n20260), .ZN(
        P1_U3058) );
  INV_X1 U23220 ( .A(n20624), .ZN(n20675) );
  NOR2_X1 U23221 ( .A1(n20481), .A2(n20278), .ZN(n20262) );
  AOI21_X1 U23222 ( .B1(n20310), .B2(n20675), .A(n20262), .ZN(n20264) );
  AOI22_X1 U23223 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20281), .B1(
        n20673), .B2(n20280), .ZN(n20263) );
  OAI211_X1 U23224 ( .C1(n20678), .C2(n20284), .A(n20264), .B(n20263), .ZN(
        P1_U3059) );
  OAI22_X1 U23225 ( .A1(n20284), .A2(n20684), .B1(n20485), .B2(n20278), .ZN(
        n20265) );
  INV_X1 U23226 ( .A(n20265), .ZN(n20267) );
  AOI22_X1 U23227 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20281), .B1(
        n20679), .B2(n20280), .ZN(n20266) );
  OAI211_X1 U23228 ( .C1(n20628), .C2(n20277), .A(n20267), .B(n20266), .ZN(
        P1_U3060) );
  INV_X1 U23229 ( .A(n20632), .ZN(n20687) );
  NOR2_X1 U23230 ( .A1(n20489), .A2(n20278), .ZN(n20268) );
  AOI21_X1 U23231 ( .B1(n20310), .B2(n20687), .A(n20268), .ZN(n20270) );
  AOI22_X1 U23232 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20281), .B1(
        n20685), .B2(n20280), .ZN(n20269) );
  OAI211_X1 U23233 ( .C1(n20690), .C2(n20284), .A(n20270), .B(n20269), .ZN(
        P1_U3061) );
  NOR2_X1 U23234 ( .A1(n20493), .A2(n20278), .ZN(n20271) );
  AOI21_X1 U23235 ( .B1(n20310), .B2(n20693), .A(n20271), .ZN(n20273) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20281), .B1(
        n20691), .B2(n20280), .ZN(n20272) );
  OAI211_X1 U23237 ( .C1(n20696), .C2(n20284), .A(n20273), .B(n20272), .ZN(
        P1_U3062) );
  OAI22_X1 U23238 ( .A1(n20284), .A2(n20702), .B1(n20497), .B2(n20278), .ZN(
        n20274) );
  INV_X1 U23239 ( .A(n20274), .ZN(n20276) );
  AOI22_X1 U23240 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20281), .B1(
        n20697), .B2(n20280), .ZN(n20275) );
  OAI211_X1 U23241 ( .C1(n20640), .C2(n20277), .A(n20276), .B(n20275), .ZN(
        P1_U3063) );
  NOR2_X1 U23242 ( .A1(n20501), .A2(n20278), .ZN(n20279) );
  AOI21_X1 U23243 ( .B1(n20310), .B2(n20707), .A(n20279), .ZN(n20283) );
  AOI22_X1 U23244 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20281), .B1(
        n20704), .B2(n20280), .ZN(n20282) );
  OAI211_X1 U23245 ( .C1(n20713), .C2(n20284), .A(n20283), .B(n20282), .ZN(
        P1_U3064) );
  NAND3_X1 U23246 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n21022), .A3(
        n20541), .ZN(n20314) );
  NOR2_X1 U23247 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20314), .ZN(
        n20309) );
  OR2_X1 U23248 ( .A1(n13182), .A2(n20285), .ZN(n20341) );
  NAND2_X1 U23249 ( .A1(n20464), .A2(n20661), .ZN(n20288) );
  INV_X1 U23250 ( .A(n20286), .ZN(n20604) );
  OAI22_X1 U23251 ( .A1(n20341), .A2(n20288), .B1(n20604), .B2(n20287), .ZN(
        n20308) );
  AOI22_X1 U23252 ( .A1(n20655), .A2(n20309), .B1(n20654), .B2(n20308), .ZN(
        n20295) );
  INV_X1 U23253 ( .A(n20338), .ZN(n20289) );
  OAI21_X1 U23254 ( .B1(n20310), .B2(n20289), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20290) );
  OAI21_X1 U23255 ( .B1(n20603), .B2(n20341), .A(n20290), .ZN(n20293) );
  OAI221_X1 U23256 ( .B1(n20309), .B2(n20547), .C1(n20309), .C2(n20293), .A(
        n20611), .ZN(n20311) );
  AOI22_X1 U23257 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20311), .B1(
        n20310), .B2(n20613), .ZN(n20294) );
  OAI211_X1 U23258 ( .C1(n20616), .C2(n20338), .A(n20295), .B(n20294), .ZN(
        P1_U3065) );
  AOI22_X1 U23259 ( .A1(n20668), .A2(n20309), .B1(n20667), .B2(n20308), .ZN(
        n20297) );
  AOI22_X1 U23260 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20311), .B1(
        n20310), .B2(n20617), .ZN(n20296) );
  OAI211_X1 U23261 ( .C1(n20620), .C2(n20338), .A(n20297), .B(n20296), .ZN(
        P1_U3066) );
  AOI22_X1 U23262 ( .A1(n20674), .A2(n20309), .B1(n20673), .B2(n20308), .ZN(
        n20299) );
  AOI22_X1 U23263 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20311), .B1(
        n20310), .B2(n20621), .ZN(n20298) );
  OAI211_X1 U23264 ( .C1(n20624), .C2(n20338), .A(n20299), .B(n20298), .ZN(
        P1_U3067) );
  AOI22_X1 U23265 ( .A1(n20680), .A2(n20309), .B1(n20679), .B2(n20308), .ZN(
        n20301) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20311), .B1(
        n20310), .B2(n20625), .ZN(n20300) );
  OAI211_X1 U23267 ( .C1(n20628), .C2(n20338), .A(n20301), .B(n20300), .ZN(
        P1_U3068) );
  AOI22_X1 U23268 ( .A1(n20686), .A2(n20309), .B1(n20685), .B2(n20308), .ZN(
        n20303) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20311), .B1(
        n20310), .B2(n20629), .ZN(n20302) );
  OAI211_X1 U23270 ( .C1(n20632), .C2(n20338), .A(n20303), .B(n20302), .ZN(
        P1_U3069) );
  AOI22_X1 U23271 ( .A1(n20692), .A2(n20309), .B1(n20691), .B2(n20308), .ZN(
        n20305) );
  AOI22_X1 U23272 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20311), .B1(
        n20310), .B2(n20633), .ZN(n20304) );
  OAI211_X1 U23273 ( .C1(n20636), .C2(n20338), .A(n20305), .B(n20304), .ZN(
        P1_U3070) );
  AOI22_X1 U23274 ( .A1(n20698), .A2(n20309), .B1(n20697), .B2(n20308), .ZN(
        n20307) );
  AOI22_X1 U23275 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20311), .B1(
        n20310), .B2(n20637), .ZN(n20306) );
  OAI211_X1 U23276 ( .C1(n20640), .C2(n20338), .A(n20307), .B(n20306), .ZN(
        P1_U3071) );
  AOI22_X1 U23277 ( .A1(n20706), .A2(n20309), .B1(n20704), .B2(n20308), .ZN(
        n20313) );
  AOI22_X1 U23278 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20311), .B1(
        n20310), .B2(n20643), .ZN(n20312) );
  OAI211_X1 U23279 ( .C1(n20648), .C2(n20338), .A(n20313), .B(n20312), .ZN(
        P1_U3072) );
  NOR2_X1 U23280 ( .A1(n20573), .A2(n20314), .ZN(n20333) );
  INV_X1 U23281 ( .A(n20341), .ZN(n20376) );
  AOI21_X1 U23282 ( .B1(n20376), .B2(n20575), .A(n20333), .ZN(n20315) );
  OAI22_X1 U23283 ( .A1(n20315), .A2(n20653), .B1(n20314), .B2(n20811), .ZN(
        n20332) );
  AOI22_X1 U23284 ( .A1(n20655), .A2(n20333), .B1(n20654), .B2(n20332), .ZN(
        n20319) );
  INV_X1 U23285 ( .A(n20314), .ZN(n20317) );
  NOR2_X1 U23286 ( .A1(n20383), .A2(n20653), .ZN(n20379) );
  OAI21_X1 U23287 ( .B1(n20379), .B2(n20578), .A(n20315), .ZN(n20316) );
  OAI211_X1 U23288 ( .C1(n20661), .C2(n20317), .A(n20660), .B(n20316), .ZN(
        n20335) );
  NAND2_X1 U23289 ( .A1(n20383), .A2(n20572), .ZN(n20374) );
  AOI22_X1 U23290 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20335), .B1(
        n20334), .B2(n20663), .ZN(n20318) );
  OAI211_X1 U23291 ( .C1(n20666), .C2(n20338), .A(n20319), .B(n20318), .ZN(
        P1_U3073) );
  AOI22_X1 U23292 ( .A1(n20668), .A2(n20333), .B1(n20667), .B2(n20332), .ZN(
        n20321) );
  INV_X1 U23293 ( .A(n20620), .ZN(n20669) );
  AOI22_X1 U23294 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20335), .B1(
        n20334), .B2(n20669), .ZN(n20320) );
  OAI211_X1 U23295 ( .C1(n20672), .C2(n20338), .A(n20321), .B(n20320), .ZN(
        P1_U3074) );
  AOI22_X1 U23296 ( .A1(n20674), .A2(n20333), .B1(n20673), .B2(n20332), .ZN(
        n20323) );
  AOI22_X1 U23297 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20335), .B1(
        n20334), .B2(n20675), .ZN(n20322) );
  OAI211_X1 U23298 ( .C1(n20678), .C2(n20338), .A(n20323), .B(n20322), .ZN(
        P1_U3075) );
  AOI22_X1 U23299 ( .A1(n20680), .A2(n20333), .B1(n20679), .B2(n20332), .ZN(
        n20325) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20335), .B1(
        n20334), .B2(n20681), .ZN(n20324) );
  OAI211_X1 U23301 ( .C1(n20684), .C2(n20338), .A(n20325), .B(n20324), .ZN(
        P1_U3076) );
  AOI22_X1 U23302 ( .A1(n20686), .A2(n20333), .B1(n20685), .B2(n20332), .ZN(
        n20327) );
  AOI22_X1 U23303 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20335), .B1(
        n20334), .B2(n20687), .ZN(n20326) );
  OAI211_X1 U23304 ( .C1(n20690), .C2(n20338), .A(n20327), .B(n20326), .ZN(
        P1_U3077) );
  AOI22_X1 U23305 ( .A1(n20692), .A2(n20333), .B1(n20691), .B2(n20332), .ZN(
        n20329) );
  AOI22_X1 U23306 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20335), .B1(
        n20334), .B2(n20693), .ZN(n20328) );
  OAI211_X1 U23307 ( .C1(n20696), .C2(n20338), .A(n20329), .B(n20328), .ZN(
        P1_U3078) );
  AOI22_X1 U23308 ( .A1(n20698), .A2(n20333), .B1(n20697), .B2(n20332), .ZN(
        n20331) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20335), .B1(
        n20334), .B2(n20699), .ZN(n20330) );
  OAI211_X1 U23310 ( .C1(n20702), .C2(n20338), .A(n20331), .B(n20330), .ZN(
        P1_U3079) );
  AOI22_X1 U23311 ( .A1(n20706), .A2(n20333), .B1(n20704), .B2(n20332), .ZN(
        n20337) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20335), .B1(
        n20334), .B2(n20707), .ZN(n20336) );
  OAI211_X1 U23313 ( .C1(n20713), .C2(n20338), .A(n20337), .B(n20336), .ZN(
        P1_U3080) );
  INV_X1 U23314 ( .A(n20381), .ZN(n20377) );
  OR2_X1 U23315 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20377), .ZN(
        n20368) );
  OAI22_X1 U23316 ( .A1(n20374), .A2(n20666), .B1(n20368), .B2(n20460), .ZN(
        n20339) );
  INV_X1 U23317 ( .A(n20339), .ZN(n20349) );
  NAND3_X1 U23318 ( .A1(n20405), .A2(n20374), .A3(n20661), .ZN(n20340) );
  NAND2_X1 U23319 ( .A1(n20340), .A2(n20543), .ZN(n20344) );
  OR2_X1 U23320 ( .A1(n20341), .A2(n20464), .ZN(n20346) );
  AOI22_X1 U23321 ( .A1(n20344), .A2(n20346), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20368), .ZN(n20343) );
  NAND3_X1 U23322 ( .A1(n20611), .A2(n20343), .A3(n20342), .ZN(n20371) );
  INV_X1 U23323 ( .A(n20344), .ZN(n20347) );
  OAI22_X1 U23324 ( .A1(n20347), .A2(n20346), .B1(n20345), .B2(n20604), .ZN(
        n20370) );
  AOI22_X1 U23325 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20371), .B1(
        n20654), .B2(n20370), .ZN(n20348) );
  OAI211_X1 U23326 ( .C1(n20616), .C2(n20405), .A(n20349), .B(n20348), .ZN(
        P1_U3081) );
  OAI22_X1 U23327 ( .A1(n20405), .A2(n20620), .B1(n20477), .B2(n20368), .ZN(
        n20350) );
  INV_X1 U23328 ( .A(n20350), .ZN(n20352) );
  AOI22_X1 U23329 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20371), .B1(
        n20667), .B2(n20370), .ZN(n20351) );
  OAI211_X1 U23330 ( .C1(n20672), .C2(n20374), .A(n20352), .B(n20351), .ZN(
        P1_U3082) );
  OAI22_X1 U23331 ( .A1(n20374), .A2(n20678), .B1(n20481), .B2(n20368), .ZN(
        n20353) );
  INV_X1 U23332 ( .A(n20353), .ZN(n20355) );
  AOI22_X1 U23333 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20371), .B1(
        n20673), .B2(n20370), .ZN(n20354) );
  OAI211_X1 U23334 ( .C1(n20624), .C2(n20405), .A(n20355), .B(n20354), .ZN(
        P1_U3083) );
  OAI22_X1 U23335 ( .A1(n20374), .A2(n20684), .B1(n20485), .B2(n20368), .ZN(
        n20356) );
  INV_X1 U23336 ( .A(n20356), .ZN(n20358) );
  AOI22_X1 U23337 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20371), .B1(
        n20679), .B2(n20370), .ZN(n20357) );
  OAI211_X1 U23338 ( .C1(n20628), .C2(n20405), .A(n20358), .B(n20357), .ZN(
        P1_U3084) );
  OAI22_X1 U23339 ( .A1(n20405), .A2(n20632), .B1(n20368), .B2(n20489), .ZN(
        n20359) );
  INV_X1 U23340 ( .A(n20359), .ZN(n20361) );
  AOI22_X1 U23341 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20371), .B1(
        n20685), .B2(n20370), .ZN(n20360) );
  OAI211_X1 U23342 ( .C1(n20690), .C2(n20374), .A(n20361), .B(n20360), .ZN(
        P1_U3085) );
  OAI22_X1 U23343 ( .A1(n20405), .A2(n20636), .B1(n20368), .B2(n20493), .ZN(
        n20362) );
  INV_X1 U23344 ( .A(n20362), .ZN(n20364) );
  AOI22_X1 U23345 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20371), .B1(
        n20691), .B2(n20370), .ZN(n20363) );
  OAI211_X1 U23346 ( .C1(n20696), .C2(n20374), .A(n20364), .B(n20363), .ZN(
        P1_U3086) );
  OAI22_X1 U23347 ( .A1(n20374), .A2(n20702), .B1(n20497), .B2(n20368), .ZN(
        n20365) );
  INV_X1 U23348 ( .A(n20365), .ZN(n20367) );
  AOI22_X1 U23349 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20371), .B1(
        n20697), .B2(n20370), .ZN(n20366) );
  OAI211_X1 U23350 ( .C1(n20640), .C2(n20405), .A(n20367), .B(n20366), .ZN(
        P1_U3087) );
  OAI22_X1 U23351 ( .A1(n20405), .A2(n20648), .B1(n20368), .B2(n20501), .ZN(
        n20369) );
  INV_X1 U23352 ( .A(n20369), .ZN(n20373) );
  AOI22_X1 U23353 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20371), .B1(
        n20704), .B2(n20370), .ZN(n20372) );
  OAI211_X1 U23354 ( .C1(n20713), .C2(n20374), .A(n20373), .B(n20372), .ZN(
        P1_U3088) );
  INV_X1 U23355 ( .A(n20375), .ZN(n20401) );
  AOI21_X1 U23356 ( .B1(n20376), .B2(n20650), .A(n20401), .ZN(n20378) );
  OAI22_X1 U23357 ( .A1(n20378), .A2(n20653), .B1(n20377), .B2(n20811), .ZN(
        n20400) );
  AOI22_X1 U23358 ( .A1(n20655), .A2(n20401), .B1(n20654), .B2(n20400), .ZN(
        n20385) );
  OAI21_X1 U23359 ( .B1(n20658), .B2(n20379), .A(n20378), .ZN(n20380) );
  OAI211_X1 U23360 ( .C1(n20381), .C2(n20661), .A(n20660), .B(n20380), .ZN(
        n20402) );
  NAND2_X1 U23361 ( .A1(n20383), .A2(n20382), .ZN(n20399) );
  AOI22_X1 U23362 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20402), .B1(
        n20428), .B2(n20663), .ZN(n20384) );
  OAI211_X1 U23363 ( .C1(n20666), .C2(n20405), .A(n20385), .B(n20384), .ZN(
        P1_U3089) );
  AOI22_X1 U23364 ( .A1(n20668), .A2(n20401), .B1(n20667), .B2(n20400), .ZN(
        n20387) );
  INV_X1 U23365 ( .A(n20405), .ZN(n20396) );
  AOI22_X1 U23366 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20402), .B1(
        n20396), .B2(n20617), .ZN(n20386) );
  OAI211_X1 U23367 ( .C1(n20620), .C2(n20399), .A(n20387), .B(n20386), .ZN(
        P1_U3090) );
  AOI22_X1 U23368 ( .A1(n20674), .A2(n20401), .B1(n20673), .B2(n20400), .ZN(
        n20389) );
  AOI22_X1 U23369 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20402), .B1(
        n20396), .B2(n20621), .ZN(n20388) );
  OAI211_X1 U23370 ( .C1(n20624), .C2(n20399), .A(n20389), .B(n20388), .ZN(
        P1_U3091) );
  AOI22_X1 U23371 ( .A1(n20680), .A2(n20401), .B1(n20679), .B2(n20400), .ZN(
        n20391) );
  AOI22_X1 U23372 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20402), .B1(
        n20428), .B2(n20681), .ZN(n20390) );
  OAI211_X1 U23373 ( .C1(n20684), .C2(n20405), .A(n20391), .B(n20390), .ZN(
        P1_U3092) );
  AOI22_X1 U23374 ( .A1(n20686), .A2(n20401), .B1(n20685), .B2(n20400), .ZN(
        n20393) );
  AOI22_X1 U23375 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20402), .B1(
        n20428), .B2(n20687), .ZN(n20392) );
  OAI211_X1 U23376 ( .C1(n20690), .C2(n20405), .A(n20393), .B(n20392), .ZN(
        P1_U3093) );
  AOI22_X1 U23377 ( .A1(n20692), .A2(n20401), .B1(n20691), .B2(n20400), .ZN(
        n20395) );
  AOI22_X1 U23378 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20402), .B1(
        n20396), .B2(n20633), .ZN(n20394) );
  OAI211_X1 U23379 ( .C1(n20636), .C2(n20399), .A(n20395), .B(n20394), .ZN(
        P1_U3094) );
  AOI22_X1 U23380 ( .A1(n20698), .A2(n20401), .B1(n20697), .B2(n20400), .ZN(
        n20398) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20402), .B1(
        n20396), .B2(n20637), .ZN(n20397) );
  OAI211_X1 U23382 ( .C1(n20640), .C2(n20399), .A(n20398), .B(n20397), .ZN(
        P1_U3095) );
  AOI22_X1 U23383 ( .A1(n20706), .A2(n20401), .B1(n20704), .B2(n20400), .ZN(
        n20404) );
  AOI22_X1 U23384 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20402), .B1(
        n20428), .B2(n20707), .ZN(n20403) );
  OAI211_X1 U23385 ( .C1(n20713), .C2(n20405), .A(n20404), .B(n20403), .ZN(
        P1_U3096) );
  INV_X1 U23386 ( .A(n20510), .ZN(n20433) );
  NAND3_X1 U23387 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20459), .A3(
        n20541), .ZN(n20432) );
  NOR2_X1 U23388 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20432), .ZN(
        n20427) );
  NAND2_X1 U23389 ( .A1(n20406), .A2(n13182), .ZN(n20465) );
  INV_X1 U23390 ( .A(n20465), .ZN(n20512) );
  AOI21_X1 U23391 ( .B1(n20512), .B2(n20464), .A(n20427), .ZN(n20409) );
  NAND2_X1 U23392 ( .A1(n20407), .A2(n20466), .ZN(n20549) );
  OAI22_X1 U23393 ( .A1(n20409), .A2(n20653), .B1(n20472), .B2(n20549), .ZN(
        n20426) );
  AOI22_X1 U23394 ( .A1(n20655), .A2(n20427), .B1(n20426), .B2(n20654), .ZN(
        n20413) );
  INV_X1 U23395 ( .A(n20457), .ZN(n20408) );
  OAI21_X1 U23396 ( .B1(n20408), .B2(n20428), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20410) );
  NAND2_X1 U23397 ( .A1(n20410), .A2(n20409), .ZN(n20411) );
  AOI22_X1 U23398 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20429), .B1(
        n20428), .B2(n20613), .ZN(n20412) );
  OAI211_X1 U23399 ( .C1(n20616), .C2(n20457), .A(n20413), .B(n20412), .ZN(
        P1_U3097) );
  AOI22_X1 U23400 ( .A1(n20668), .A2(n20427), .B1(n20426), .B2(n20667), .ZN(
        n20415) );
  AOI22_X1 U23401 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20429), .B1(
        n20428), .B2(n20617), .ZN(n20414) );
  OAI211_X1 U23402 ( .C1(n20620), .C2(n20457), .A(n20415), .B(n20414), .ZN(
        P1_U3098) );
  AOI22_X1 U23403 ( .A1(n20674), .A2(n20427), .B1(n20426), .B2(n20673), .ZN(
        n20417) );
  AOI22_X1 U23404 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20429), .B1(
        n20428), .B2(n20621), .ZN(n20416) );
  OAI211_X1 U23405 ( .C1(n20624), .C2(n20457), .A(n20417), .B(n20416), .ZN(
        P1_U3099) );
  AOI22_X1 U23406 ( .A1(n20680), .A2(n20427), .B1(n20426), .B2(n20679), .ZN(
        n20419) );
  AOI22_X1 U23407 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20429), .B1(
        n20428), .B2(n20625), .ZN(n20418) );
  OAI211_X1 U23408 ( .C1(n20628), .C2(n20457), .A(n20419), .B(n20418), .ZN(
        P1_U3100) );
  AOI22_X1 U23409 ( .A1(n20686), .A2(n20427), .B1(n20685), .B2(n20426), .ZN(
        n20421) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20429), .B1(
        n20428), .B2(n20629), .ZN(n20420) );
  OAI211_X1 U23411 ( .C1(n20632), .C2(n20457), .A(n20421), .B(n20420), .ZN(
        P1_U3101) );
  AOI22_X1 U23412 ( .A1(n20692), .A2(n20427), .B1(n20691), .B2(n20426), .ZN(
        n20423) );
  AOI22_X1 U23413 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20429), .B1(
        n20428), .B2(n20633), .ZN(n20422) );
  OAI211_X1 U23414 ( .C1(n20636), .C2(n20457), .A(n20423), .B(n20422), .ZN(
        P1_U3102) );
  AOI22_X1 U23415 ( .A1(n20698), .A2(n20427), .B1(n20697), .B2(n20426), .ZN(
        n20425) );
  AOI22_X1 U23416 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20429), .B1(
        n20428), .B2(n20637), .ZN(n20424) );
  OAI211_X1 U23417 ( .C1(n20640), .C2(n20457), .A(n20425), .B(n20424), .ZN(
        P1_U3103) );
  AOI22_X1 U23418 ( .A1(n20706), .A2(n20427), .B1(n20704), .B2(n20426), .ZN(
        n20431) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20429), .B1(
        n20428), .B2(n20643), .ZN(n20430) );
  OAI211_X1 U23420 ( .C1(n20648), .C2(n20457), .A(n20431), .B(n20430), .ZN(
        P1_U3104) );
  NOR2_X1 U23421 ( .A1(n20573), .A2(n20432), .ZN(n20453) );
  AOI21_X1 U23422 ( .B1(n20512), .B2(n20575), .A(n20453), .ZN(n20434) );
  OAI22_X1 U23423 ( .A1(n20434), .A2(n20653), .B1(n20432), .B2(n20811), .ZN(
        n20452) );
  AOI22_X1 U23424 ( .A1(n20655), .A2(n20453), .B1(n20452), .B2(n20654), .ZN(
        n20439) );
  INV_X1 U23425 ( .A(n20432), .ZN(n20436) );
  NOR2_X1 U23426 ( .A1(n20433), .A2(n20653), .ZN(n20515) );
  OAI21_X1 U23427 ( .B1(n20515), .B2(n20578), .A(n20434), .ZN(n20435) );
  OAI211_X1 U23428 ( .C1(n20661), .C2(n20436), .A(n20660), .B(n20435), .ZN(
        n20454) );
  INV_X1 U23429 ( .A(n20572), .ZN(n20437) );
  AOI22_X1 U23430 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20454), .B1(
        n20462), .B2(n20663), .ZN(n20438) );
  OAI211_X1 U23431 ( .C1(n20666), .C2(n20457), .A(n20439), .B(n20438), .ZN(
        P1_U3105) );
  AOI22_X1 U23432 ( .A1(n20668), .A2(n20453), .B1(n20452), .B2(n20667), .ZN(
        n20441) );
  AOI22_X1 U23433 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20454), .B1(
        n20462), .B2(n20669), .ZN(n20440) );
  OAI211_X1 U23434 ( .C1(n20672), .C2(n20457), .A(n20441), .B(n20440), .ZN(
        P1_U3106) );
  AOI22_X1 U23435 ( .A1(n20674), .A2(n20453), .B1(n20452), .B2(n20673), .ZN(
        n20443) );
  AOI22_X1 U23436 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20454), .B1(
        n20462), .B2(n20675), .ZN(n20442) );
  OAI211_X1 U23437 ( .C1(n20678), .C2(n20457), .A(n20443), .B(n20442), .ZN(
        P1_U3107) );
  AOI22_X1 U23438 ( .A1(n20680), .A2(n20453), .B1(n20452), .B2(n20679), .ZN(
        n20445) );
  AOI22_X1 U23439 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20454), .B1(
        n20462), .B2(n20681), .ZN(n20444) );
  OAI211_X1 U23440 ( .C1(n20684), .C2(n20457), .A(n20445), .B(n20444), .ZN(
        P1_U3108) );
  AOI22_X1 U23441 ( .A1(n20686), .A2(n20453), .B1(n20685), .B2(n20452), .ZN(
        n20447) );
  AOI22_X1 U23442 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20454), .B1(
        n20462), .B2(n20687), .ZN(n20446) );
  OAI211_X1 U23443 ( .C1(n20690), .C2(n20457), .A(n20447), .B(n20446), .ZN(
        P1_U3109) );
  AOI22_X1 U23444 ( .A1(n20692), .A2(n20453), .B1(n20691), .B2(n20452), .ZN(
        n20449) );
  AOI22_X1 U23445 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20454), .B1(
        n20462), .B2(n20693), .ZN(n20448) );
  OAI211_X1 U23446 ( .C1(n20696), .C2(n20457), .A(n20449), .B(n20448), .ZN(
        P1_U3110) );
  AOI22_X1 U23447 ( .A1(n20698), .A2(n20453), .B1(n20697), .B2(n20452), .ZN(
        n20451) );
  AOI22_X1 U23448 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20454), .B1(
        n20462), .B2(n20699), .ZN(n20450) );
  OAI211_X1 U23449 ( .C1(n20702), .C2(n20457), .A(n20451), .B(n20450), .ZN(
        P1_U3111) );
  AOI22_X1 U23450 ( .A1(n20706), .A2(n20453), .B1(n20704), .B2(n20452), .ZN(
        n20456) );
  AOI22_X1 U23451 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20454), .B1(
        n20462), .B2(n20707), .ZN(n20455) );
  OAI211_X1 U23452 ( .C1(n20713), .C2(n20457), .A(n20456), .B(n20455), .ZN(
        P1_U3112) );
  INV_X1 U23453 ( .A(n20601), .ZN(n20458) );
  NAND3_X1 U23454 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20459), .ZN(n20513) );
  NOR2_X1 U23455 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20513), .ZN(
        n20467) );
  INV_X1 U23456 ( .A(n20467), .ZN(n20502) );
  OAI22_X1 U23457 ( .A1(n20508), .A2(n20666), .B1(n20502), .B2(n20460), .ZN(
        n20461) );
  INV_X1 U23458 ( .A(n20461), .ZN(n20476) );
  OAI21_X1 U23459 ( .B1(n20536), .B2(n20462), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20463) );
  NAND2_X1 U23460 ( .A1(n20463), .A2(n20661), .ZN(n20474) );
  NOR2_X1 U23461 ( .A1(n20465), .A2(n20464), .ZN(n20471) );
  OR2_X1 U23462 ( .A1(n20466), .A2(n21022), .ZN(n20605) );
  NAND2_X1 U23463 ( .A1(n20605), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20610) );
  OAI21_X1 U23464 ( .B1(n20547), .B2(n20467), .A(n20610), .ZN(n20468) );
  INV_X1 U23465 ( .A(n20468), .ZN(n20470) );
  OAI211_X1 U23466 ( .C1(n20474), .C2(n20471), .A(n20470), .B(n20469), .ZN(
        n20505) );
  INV_X1 U23467 ( .A(n20471), .ZN(n20473) );
  OAI22_X1 U23468 ( .A1(n20474), .A2(n20473), .B1(n20472), .B2(n20605), .ZN(
        n20504) );
  AOI22_X1 U23469 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20505), .B1(
        n20654), .B2(n20504), .ZN(n20475) );
  OAI211_X1 U23470 ( .C1(n20616), .C2(n20533), .A(n20476), .B(n20475), .ZN(
        P1_U3113) );
  OAI22_X1 U23471 ( .A1(n20508), .A2(n20672), .B1(n20502), .B2(n20477), .ZN(
        n20478) );
  INV_X1 U23472 ( .A(n20478), .ZN(n20480) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20505), .B1(
        n20667), .B2(n20504), .ZN(n20479) );
  OAI211_X1 U23474 ( .C1(n20620), .C2(n20533), .A(n20480), .B(n20479), .ZN(
        P1_U3114) );
  OAI22_X1 U23475 ( .A1(n20533), .A2(n20624), .B1(n20481), .B2(n20502), .ZN(
        n20482) );
  INV_X1 U23476 ( .A(n20482), .ZN(n20484) );
  AOI22_X1 U23477 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20505), .B1(
        n20673), .B2(n20504), .ZN(n20483) );
  OAI211_X1 U23478 ( .C1(n20678), .C2(n20508), .A(n20484), .B(n20483), .ZN(
        P1_U3115) );
  OAI22_X1 U23479 ( .A1(n20533), .A2(n20628), .B1(n20502), .B2(n20485), .ZN(
        n20486) );
  INV_X1 U23480 ( .A(n20486), .ZN(n20488) );
  AOI22_X1 U23481 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20505), .B1(
        n20679), .B2(n20504), .ZN(n20487) );
  OAI211_X1 U23482 ( .C1(n20684), .C2(n20508), .A(n20488), .B(n20487), .ZN(
        P1_U3116) );
  OAI22_X1 U23483 ( .A1(n20533), .A2(n20632), .B1(n20502), .B2(n20489), .ZN(
        n20490) );
  INV_X1 U23484 ( .A(n20490), .ZN(n20492) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20505), .B1(
        n20685), .B2(n20504), .ZN(n20491) );
  OAI211_X1 U23486 ( .C1(n20690), .C2(n20508), .A(n20492), .B(n20491), .ZN(
        P1_U3117) );
  OAI22_X1 U23487 ( .A1(n20533), .A2(n20636), .B1(n20502), .B2(n20493), .ZN(
        n20494) );
  INV_X1 U23488 ( .A(n20494), .ZN(n20496) );
  AOI22_X1 U23489 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20505), .B1(
        n20691), .B2(n20504), .ZN(n20495) );
  OAI211_X1 U23490 ( .C1(n20696), .C2(n20508), .A(n20496), .B(n20495), .ZN(
        P1_U3118) );
  OAI22_X1 U23491 ( .A1(n20533), .A2(n20640), .B1(n20502), .B2(n20497), .ZN(
        n20498) );
  INV_X1 U23492 ( .A(n20498), .ZN(n20500) );
  AOI22_X1 U23493 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20505), .B1(
        n20697), .B2(n20504), .ZN(n20499) );
  OAI211_X1 U23494 ( .C1(n20702), .C2(n20508), .A(n20500), .B(n20499), .ZN(
        P1_U3119) );
  OAI22_X1 U23495 ( .A1(n20533), .A2(n20648), .B1(n20502), .B2(n20501), .ZN(
        n20503) );
  INV_X1 U23496 ( .A(n20503), .ZN(n20507) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20505), .B1(
        n20704), .B2(n20504), .ZN(n20506) );
  OAI211_X1 U23498 ( .C1(n20713), .C2(n20508), .A(n20507), .B(n20506), .ZN(
        P1_U3120) );
  NOR2_X1 U23499 ( .A1(n20511), .A2(n21022), .ZN(n20535) );
  AOI21_X1 U23500 ( .B1(n20512), .B2(n20650), .A(n20535), .ZN(n20514) );
  OAI22_X1 U23501 ( .A1(n20514), .A2(n20653), .B1(n20513), .B2(n20811), .ZN(
        n20534) );
  AOI22_X1 U23502 ( .A1(n20655), .A2(n20535), .B1(n20534), .B2(n20654), .ZN(
        n20519) );
  INV_X1 U23503 ( .A(n20513), .ZN(n20517) );
  OAI21_X1 U23504 ( .B1(n20658), .B2(n20515), .A(n20514), .ZN(n20516) );
  OAI211_X1 U23505 ( .C1(n20661), .C2(n20517), .A(n20660), .B(n20516), .ZN(
        n20537) );
  AOI22_X1 U23506 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20537), .B1(
        n20536), .B2(n20613), .ZN(n20518) );
  OAI211_X1 U23507 ( .C1(n20616), .C2(n20571), .A(n20519), .B(n20518), .ZN(
        P1_U3121) );
  AOI22_X1 U23508 ( .A1(n20668), .A2(n20535), .B1(n20534), .B2(n20667), .ZN(
        n20521) );
  AOI22_X1 U23509 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20537), .B1(
        n20536), .B2(n20617), .ZN(n20520) );
  OAI211_X1 U23510 ( .C1(n20620), .C2(n20571), .A(n20521), .B(n20520), .ZN(
        P1_U3122) );
  AOI22_X1 U23511 ( .A1(n20674), .A2(n20535), .B1(n20534), .B2(n20673), .ZN(
        n20523) );
  INV_X1 U23512 ( .A(n20571), .ZN(n20530) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20537), .B1(
        n20530), .B2(n20675), .ZN(n20522) );
  OAI211_X1 U23514 ( .C1(n20678), .C2(n20533), .A(n20523), .B(n20522), .ZN(
        P1_U3123) );
  AOI22_X1 U23515 ( .A1(n20680), .A2(n20535), .B1(n20534), .B2(n20679), .ZN(
        n20525) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20537), .B1(
        n20536), .B2(n20625), .ZN(n20524) );
  OAI211_X1 U23517 ( .C1(n20628), .C2(n20571), .A(n20525), .B(n20524), .ZN(
        P1_U3124) );
  AOI22_X1 U23518 ( .A1(n20686), .A2(n20535), .B1(n20534), .B2(n20685), .ZN(
        n20527) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20537), .B1(
        n20530), .B2(n20687), .ZN(n20526) );
  OAI211_X1 U23520 ( .C1(n20690), .C2(n20533), .A(n20527), .B(n20526), .ZN(
        P1_U3125) );
  AOI22_X1 U23521 ( .A1(n20692), .A2(n20535), .B1(n20534), .B2(n20691), .ZN(
        n20529) );
  AOI22_X1 U23522 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20537), .B1(
        n20536), .B2(n20633), .ZN(n20528) );
  OAI211_X1 U23523 ( .C1(n20636), .C2(n20571), .A(n20529), .B(n20528), .ZN(
        P1_U3126) );
  AOI22_X1 U23524 ( .A1(n20698), .A2(n20535), .B1(n20534), .B2(n20697), .ZN(
        n20532) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20537), .B1(
        n20530), .B2(n20699), .ZN(n20531) );
  OAI211_X1 U23526 ( .C1(n20702), .C2(n20533), .A(n20532), .B(n20531), .ZN(
        P1_U3127) );
  AOI22_X1 U23527 ( .A1(n20706), .A2(n20535), .B1(n20534), .B2(n20704), .ZN(
        n20539) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20537), .B1(
        n20536), .B2(n20643), .ZN(n20538) );
  OAI211_X1 U23529 ( .C1(n20648), .C2(n20571), .A(n20539), .B(n20538), .ZN(
        P1_U3128) );
  NAND3_X1 U23530 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20541), .ZN(n20576) );
  NOR2_X1 U23531 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20576), .ZN(
        n20566) );
  AOI22_X1 U23532 ( .A1(n20597), .A2(n20663), .B1(n20655), .B2(n20566), .ZN(
        n20553) );
  INV_X1 U23533 ( .A(n20597), .ZN(n20542) );
  NAND3_X1 U23534 ( .A1(n20542), .A2(n20661), .A3(n20571), .ZN(n20544) );
  NAND2_X1 U23535 ( .A1(n20544), .A2(n20543), .ZN(n20548) );
  OR2_X1 U23536 ( .A1(n13182), .A2(n20545), .ZN(n20574) );
  OR2_X1 U23537 ( .A1(n20574), .A2(n20603), .ZN(n20550) );
  AOI22_X1 U23538 ( .A1(n20548), .A2(n20550), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20549), .ZN(n20546) );
  OAI211_X1 U23539 ( .C1(n20566), .C2(n20547), .A(n20611), .B(n20546), .ZN(
        n20568) );
  INV_X1 U23540 ( .A(n20548), .ZN(n20551) );
  OAI22_X1 U23541 ( .A1(n20551), .A2(n20550), .B1(n20549), .B2(n20604), .ZN(
        n20567) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20568), .B1(
        n20654), .B2(n20567), .ZN(n20552) );
  OAI211_X1 U23543 ( .C1(n20666), .C2(n20571), .A(n20553), .B(n20552), .ZN(
        P1_U3129) );
  AOI22_X1 U23544 ( .A1(n20597), .A2(n20669), .B1(n20668), .B2(n20566), .ZN(
        n20555) );
  AOI22_X1 U23545 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20568), .B1(
        n20667), .B2(n20567), .ZN(n20554) );
  OAI211_X1 U23546 ( .C1(n20672), .C2(n20571), .A(n20555), .B(n20554), .ZN(
        P1_U3130) );
  AOI22_X1 U23547 ( .A1(n20597), .A2(n20675), .B1(n20674), .B2(n20566), .ZN(
        n20557) );
  AOI22_X1 U23548 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20568), .B1(
        n20673), .B2(n20567), .ZN(n20556) );
  OAI211_X1 U23549 ( .C1(n20678), .C2(n20571), .A(n20557), .B(n20556), .ZN(
        P1_U3131) );
  AOI22_X1 U23550 ( .A1(n20597), .A2(n20681), .B1(n20680), .B2(n20566), .ZN(
        n20559) );
  AOI22_X1 U23551 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20568), .B1(
        n20679), .B2(n20567), .ZN(n20558) );
  OAI211_X1 U23552 ( .C1(n20684), .C2(n20571), .A(n20559), .B(n20558), .ZN(
        P1_U3132) );
  AOI22_X1 U23553 ( .A1(n20597), .A2(n20687), .B1(n20686), .B2(n20566), .ZN(
        n20561) );
  AOI22_X1 U23554 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20568), .B1(
        n20685), .B2(n20567), .ZN(n20560) );
  OAI211_X1 U23555 ( .C1(n20690), .C2(n20571), .A(n20561), .B(n20560), .ZN(
        P1_U3133) );
  AOI22_X1 U23556 ( .A1(n20597), .A2(n20693), .B1(n20692), .B2(n20566), .ZN(
        n20563) );
  AOI22_X1 U23557 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20568), .B1(
        n20691), .B2(n20567), .ZN(n20562) );
  OAI211_X1 U23558 ( .C1(n20696), .C2(n20571), .A(n20563), .B(n20562), .ZN(
        P1_U3134) );
  AOI22_X1 U23559 ( .A1(n20597), .A2(n20699), .B1(n20698), .B2(n20566), .ZN(
        n20565) );
  AOI22_X1 U23560 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20568), .B1(
        n20697), .B2(n20567), .ZN(n20564) );
  OAI211_X1 U23561 ( .C1(n20702), .C2(n20571), .A(n20565), .B(n20564), .ZN(
        P1_U3135) );
  AOI22_X1 U23562 ( .A1(n20597), .A2(n20707), .B1(n20706), .B2(n20566), .ZN(
        n20570) );
  AOI22_X1 U23563 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20568), .B1(
        n20704), .B2(n20567), .ZN(n20569) );
  OAI211_X1 U23564 ( .C1(n20713), .C2(n20571), .A(n20570), .B(n20569), .ZN(
        P1_U3136) );
  NAND2_X1 U23565 ( .A1(n20602), .A2(n20572), .ZN(n20606) );
  NOR2_X1 U23566 ( .A1(n20573), .A2(n20576), .ZN(n20596) );
  INV_X1 U23567 ( .A(n20574), .ZN(n20651) );
  AOI21_X1 U23568 ( .B1(n20651), .B2(n20575), .A(n20596), .ZN(n20577) );
  OAI22_X1 U23569 ( .A1(n20577), .A2(n20653), .B1(n20576), .B2(n20811), .ZN(
        n20595) );
  AOI22_X1 U23570 ( .A1(n20655), .A2(n20596), .B1(n20654), .B2(n20595), .ZN(
        n20582) );
  INV_X1 U23571 ( .A(n20576), .ZN(n20580) );
  NOR2_X1 U23572 ( .A1(n20602), .A2(n20653), .ZN(n20657) );
  OAI21_X1 U23573 ( .B1(n20657), .B2(n20578), .A(n20577), .ZN(n20579) );
  OAI211_X1 U23574 ( .C1(n20661), .C2(n20580), .A(n20660), .B(n20579), .ZN(
        n20598) );
  AOI22_X1 U23575 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20613), .ZN(n20581) );
  OAI211_X1 U23576 ( .C1(n20616), .C2(n20606), .A(n20582), .B(n20581), .ZN(
        P1_U3137) );
  AOI22_X1 U23577 ( .A1(n20668), .A2(n20596), .B1(n20667), .B2(n20595), .ZN(
        n20584) );
  AOI22_X1 U23578 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20617), .ZN(n20583) );
  OAI211_X1 U23579 ( .C1(n20620), .C2(n20606), .A(n20584), .B(n20583), .ZN(
        P1_U3138) );
  AOI22_X1 U23580 ( .A1(n20674), .A2(n20596), .B1(n20673), .B2(n20595), .ZN(
        n20586) );
  AOI22_X1 U23581 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20621), .ZN(n20585) );
  OAI211_X1 U23582 ( .C1(n20624), .C2(n20606), .A(n20586), .B(n20585), .ZN(
        P1_U3139) );
  AOI22_X1 U23583 ( .A1(n20680), .A2(n20596), .B1(n20679), .B2(n20595), .ZN(
        n20588) );
  AOI22_X1 U23584 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20625), .ZN(n20587) );
  OAI211_X1 U23585 ( .C1(n20628), .C2(n20606), .A(n20588), .B(n20587), .ZN(
        P1_U3140) );
  AOI22_X1 U23586 ( .A1(n20686), .A2(n20596), .B1(n20685), .B2(n20595), .ZN(
        n20590) );
  AOI22_X1 U23587 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20629), .ZN(n20589) );
  OAI211_X1 U23588 ( .C1(n20632), .C2(n20606), .A(n20590), .B(n20589), .ZN(
        P1_U3141) );
  AOI22_X1 U23589 ( .A1(n20692), .A2(n20596), .B1(n20691), .B2(n20595), .ZN(
        n20592) );
  AOI22_X1 U23590 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20633), .ZN(n20591) );
  OAI211_X1 U23591 ( .C1(n20636), .C2(n20606), .A(n20592), .B(n20591), .ZN(
        P1_U3142) );
  AOI22_X1 U23592 ( .A1(n20698), .A2(n20596), .B1(n20697), .B2(n20595), .ZN(
        n20594) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20637), .ZN(n20593) );
  OAI211_X1 U23594 ( .C1(n20640), .C2(n20606), .A(n20594), .B(n20593), .ZN(
        P1_U3143) );
  AOI22_X1 U23595 ( .A1(n20706), .A2(n20596), .B1(n20704), .B2(n20595), .ZN(
        n20600) );
  AOI22_X1 U23596 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20643), .ZN(n20599) );
  OAI211_X1 U23597 ( .C1(n20648), .C2(n20606), .A(n20600), .B(n20599), .ZN(
        P1_U3144) );
  NOR2_X1 U23598 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20652), .ZN(
        n20642) );
  NAND2_X1 U23599 ( .A1(n20651), .A2(n20603), .ZN(n20608) );
  OAI22_X1 U23600 ( .A1(n20608), .A2(n20653), .B1(n20605), .B2(n20604), .ZN(
        n20641) );
  AOI22_X1 U23601 ( .A1(n20655), .A2(n20642), .B1(n20654), .B2(n20641), .ZN(
        n20615) );
  INV_X1 U23602 ( .A(n20712), .ZN(n20607) );
  OAI21_X1 U23603 ( .B1(n20644), .B2(n20607), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20609) );
  AOI21_X1 U23604 ( .B1(n20609), .B2(n20608), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20612) );
  AOI22_X1 U23605 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20613), .ZN(n20614) );
  OAI211_X1 U23606 ( .C1(n20616), .C2(n20712), .A(n20615), .B(n20614), .ZN(
        P1_U3145) );
  AOI22_X1 U23607 ( .A1(n20668), .A2(n20642), .B1(n20667), .B2(n20641), .ZN(
        n20619) );
  AOI22_X1 U23608 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20617), .ZN(n20618) );
  OAI211_X1 U23609 ( .C1(n20620), .C2(n20712), .A(n20619), .B(n20618), .ZN(
        P1_U3146) );
  AOI22_X1 U23610 ( .A1(n20674), .A2(n20642), .B1(n20673), .B2(n20641), .ZN(
        n20623) );
  AOI22_X1 U23611 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20621), .ZN(n20622) );
  OAI211_X1 U23612 ( .C1(n20624), .C2(n20712), .A(n20623), .B(n20622), .ZN(
        P1_U3147) );
  AOI22_X1 U23613 ( .A1(n20680), .A2(n20642), .B1(n20679), .B2(n20641), .ZN(
        n20627) );
  AOI22_X1 U23614 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20625), .ZN(n20626) );
  OAI211_X1 U23615 ( .C1(n20628), .C2(n20712), .A(n20627), .B(n20626), .ZN(
        P1_U3148) );
  AOI22_X1 U23616 ( .A1(n20686), .A2(n20642), .B1(n20685), .B2(n20641), .ZN(
        n20631) );
  AOI22_X1 U23617 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20629), .ZN(n20630) );
  OAI211_X1 U23618 ( .C1(n20632), .C2(n20712), .A(n20631), .B(n20630), .ZN(
        P1_U3149) );
  AOI22_X1 U23619 ( .A1(n20692), .A2(n20642), .B1(n20691), .B2(n20641), .ZN(
        n20635) );
  AOI22_X1 U23620 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20633), .ZN(n20634) );
  OAI211_X1 U23621 ( .C1(n20636), .C2(n20712), .A(n20635), .B(n20634), .ZN(
        P1_U3150) );
  AOI22_X1 U23622 ( .A1(n20698), .A2(n20642), .B1(n20697), .B2(n20641), .ZN(
        n20639) );
  AOI22_X1 U23623 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20637), .ZN(n20638) );
  OAI211_X1 U23624 ( .C1(n20640), .C2(n20712), .A(n20639), .B(n20638), .ZN(
        P1_U3151) );
  AOI22_X1 U23625 ( .A1(n20706), .A2(n20642), .B1(n20704), .B2(n20641), .ZN(
        n20647) );
  AOI22_X1 U23626 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20643), .ZN(n20646) );
  OAI211_X1 U23627 ( .C1(n20648), .C2(n20712), .A(n20647), .B(n20646), .ZN(
        P1_U3152) );
  INV_X1 U23628 ( .A(n20649), .ZN(n20705) );
  AOI21_X1 U23629 ( .B1(n20651), .B2(n20650), .A(n20705), .ZN(n20656) );
  OAI22_X1 U23630 ( .A1(n20656), .A2(n20653), .B1(n20652), .B2(n20811), .ZN(
        n20703) );
  AOI22_X1 U23631 ( .A1(n20655), .A2(n20705), .B1(n20654), .B2(n20703), .ZN(
        n20665) );
  OAI21_X1 U23632 ( .B1(n20658), .B2(n20657), .A(n20656), .ZN(n20659) );
  OAI211_X1 U23633 ( .C1(n20662), .C2(n20661), .A(n20660), .B(n20659), .ZN(
        n20709) );
  AOI22_X1 U23634 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20709), .B1(
        n20708), .B2(n20663), .ZN(n20664) );
  OAI211_X1 U23635 ( .C1(n20666), .C2(n20712), .A(n20665), .B(n20664), .ZN(
        P1_U3153) );
  AOI22_X1 U23636 ( .A1(n20668), .A2(n20705), .B1(n20667), .B2(n20703), .ZN(
        n20671) );
  AOI22_X1 U23637 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20709), .B1(
        n20708), .B2(n20669), .ZN(n20670) );
  OAI211_X1 U23638 ( .C1(n20672), .C2(n20712), .A(n20671), .B(n20670), .ZN(
        P1_U3154) );
  AOI22_X1 U23639 ( .A1(n20674), .A2(n20705), .B1(n20673), .B2(n20703), .ZN(
        n20677) );
  AOI22_X1 U23640 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20709), .B1(
        n20708), .B2(n20675), .ZN(n20676) );
  OAI211_X1 U23641 ( .C1(n20678), .C2(n20712), .A(n20677), .B(n20676), .ZN(
        P1_U3155) );
  AOI22_X1 U23642 ( .A1(n20680), .A2(n20705), .B1(n20679), .B2(n20703), .ZN(
        n20683) );
  AOI22_X1 U23643 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20709), .B1(
        n20708), .B2(n20681), .ZN(n20682) );
  OAI211_X1 U23644 ( .C1(n20684), .C2(n20712), .A(n20683), .B(n20682), .ZN(
        P1_U3156) );
  AOI22_X1 U23645 ( .A1(n20686), .A2(n20705), .B1(n20685), .B2(n20703), .ZN(
        n20689) );
  AOI22_X1 U23646 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20709), .B1(
        n20708), .B2(n20687), .ZN(n20688) );
  OAI211_X1 U23647 ( .C1(n20690), .C2(n20712), .A(n20689), .B(n20688), .ZN(
        P1_U3157) );
  AOI22_X1 U23648 ( .A1(n20692), .A2(n20705), .B1(n20691), .B2(n20703), .ZN(
        n20695) );
  AOI22_X1 U23649 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20709), .B1(
        n20708), .B2(n20693), .ZN(n20694) );
  OAI211_X1 U23650 ( .C1(n20696), .C2(n20712), .A(n20695), .B(n20694), .ZN(
        P1_U3158) );
  AOI22_X1 U23651 ( .A1(n20698), .A2(n20705), .B1(n20697), .B2(n20703), .ZN(
        n20701) );
  AOI22_X1 U23652 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20709), .B1(
        n20708), .B2(n20699), .ZN(n20700) );
  OAI211_X1 U23653 ( .C1(n20702), .C2(n20712), .A(n20701), .B(n20700), .ZN(
        P1_U3159) );
  AOI22_X1 U23654 ( .A1(n20706), .A2(n20705), .B1(n20704), .B2(n20703), .ZN(
        n20711) );
  AOI22_X1 U23655 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20709), .B1(
        n20708), .B2(n20707), .ZN(n20710) );
  OAI211_X1 U23656 ( .C1(n20713), .C2(n20712), .A(n20711), .B(n20710), .ZN(
        P1_U3160) );
  NOR2_X1 U23657 ( .A1(n20815), .A2(n20714), .ZN(n20717) );
  INV_X1 U23658 ( .A(n20715), .ZN(n20716) );
  OAI21_X1 U23659 ( .B1(n20717), .B2(n20811), .A(n20716), .ZN(P1_U3163) );
  INV_X1 U23660 ( .A(P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20928) );
  NOR2_X1 U23661 ( .A1(n20798), .A2(n20928), .ZN(P1_U3164) );
  AND2_X1 U23662 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20718), .ZN(
        P1_U3165) );
  AND2_X1 U23663 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20718), .ZN(
        P1_U3166) );
  AND2_X1 U23664 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20718), .ZN(
        P1_U3167) );
  AND2_X1 U23665 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20718), .ZN(
        P1_U3168) );
  AND2_X1 U23666 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20718), .ZN(
        P1_U3169) );
  AND2_X1 U23667 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20718), .ZN(
        P1_U3170) );
  AND2_X1 U23668 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20718), .ZN(
        P1_U3171) );
  AND2_X1 U23669 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20718), .ZN(
        P1_U3172) );
  AND2_X1 U23670 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20718), .ZN(
        P1_U3173) );
  AND2_X1 U23671 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20718), .ZN(
        P1_U3174) );
  AND2_X1 U23672 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20718), .ZN(
        P1_U3175) );
  AND2_X1 U23673 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20718), .ZN(
        P1_U3176) );
  AND2_X1 U23674 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20718), .ZN(
        P1_U3177) );
  AND2_X1 U23675 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20718), .ZN(
        P1_U3178) );
  INV_X1 U23676 ( .A(P1_DATAWIDTH_REG_16__SCAN_IN), .ZN(n21054) );
  NOR2_X1 U23677 ( .A1(n20798), .A2(n21054), .ZN(P1_U3179) );
  AND2_X1 U23678 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20718), .ZN(
        P1_U3180) );
  AND2_X1 U23679 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20718), .ZN(
        P1_U3181) );
  INV_X1 U23680 ( .A(P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n20916) );
  NOR2_X1 U23681 ( .A1(n20798), .A2(n20916), .ZN(P1_U3182) );
  AND2_X1 U23682 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20718), .ZN(
        P1_U3183) );
  AND2_X1 U23683 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20718), .ZN(
        P1_U3184) );
  AND2_X1 U23684 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20718), .ZN(
        P1_U3185) );
  AND2_X1 U23685 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20718), .ZN(P1_U3186) );
  AND2_X1 U23686 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20718), .ZN(P1_U3187) );
  AND2_X1 U23687 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20718), .ZN(P1_U3188) );
  AND2_X1 U23688 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20718), .ZN(P1_U3189) );
  AND2_X1 U23689 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20718), .ZN(P1_U3190) );
  AND2_X1 U23690 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20718), .ZN(P1_U3191) );
  AND2_X1 U23691 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20718), .ZN(P1_U3192) );
  AND2_X1 U23692 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20718), .ZN(P1_U3193) );
  AOI21_X1 U23693 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20724), .A(n12916), 
        .ZN(n20730) );
  NOR2_X1 U23694 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20720) );
  NOR2_X1 U23695 ( .A1(n20720), .A2(n20719), .ZN(n20721) );
  AOI211_X1 U23696 ( .C1(NA), .C2(n12916), .A(n20721), .B(n20725), .ZN(n20722)
         );
  OAI22_X1 U23697 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20730), .B1(n20809), 
        .B2(n20722), .ZN(P1_U3194) );
  AOI21_X1 U23698 ( .B1(n20724), .B2(n20727), .A(n20723), .ZN(n20732) );
  OAI211_X1 U23699 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20725), .A(
        P1_STATE_REG_0__SCAN_IN), .B(HOLD), .ZN(n20731) );
  AND2_X1 U23700 ( .A1(n20727), .A2(n20726), .ZN(n20728) );
  OAI22_X1 U23701 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20728), .B1(
        P1_STATE_REG_1__SCAN_IN), .B2(n20727), .ZN(n20729) );
  OAI22_X1 U23702 ( .A1(n20732), .A2(n20731), .B1(n20730), .B2(n20729), .ZN(
        P1_U3196) );
  NAND2_X1 U23703 ( .A1(n20809), .A2(n20733), .ZN(n20784) );
  INV_X1 U23704 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20735) );
  AND2_X1 U23705 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20809), .ZN(n20787) );
  OAI222_X1 U23706 ( .A1(n20784), .A2(n20737), .B1(n20735), .B2(n20809), .C1(
        n20734), .C2(n20780), .ZN(P1_U3197) );
  INV_X1 U23707 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20736) );
  OAI222_X1 U23708 ( .A1(n20780), .A2(n20737), .B1(n20736), .B2(n20809), .C1(
        n20739), .C2(n20784), .ZN(P1_U3198) );
  OAI222_X1 U23709 ( .A1(n20780), .A2(n20739), .B1(n20738), .B2(n20809), .C1(
        n13545), .C2(n20784), .ZN(P1_U3199) );
  INV_X1 U23710 ( .A(n20784), .ZN(n20786) );
  AOI222_X1 U23711 ( .A1(n20786), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20807), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20787), .ZN(n20740) );
  INV_X1 U23712 ( .A(n20740), .ZN(P1_U3200) );
  INV_X1 U23713 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20741) );
  OAI222_X1 U23714 ( .A1(n20780), .A2(n20742), .B1(n20741), .B2(n20809), .C1(
        n13658), .C2(n20784), .ZN(P1_U3201) );
  INV_X1 U23715 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20743) );
  OAI222_X1 U23716 ( .A1(n20780), .A2(n13658), .B1(n20743), .B2(n20809), .C1(
        n20745), .C2(n20784), .ZN(P1_U3202) );
  INV_X1 U23717 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20744) );
  OAI222_X1 U23718 ( .A1(n20780), .A2(n20745), .B1(n20744), .B2(n20809), .C1(
        n20746), .C2(n20784), .ZN(P1_U3203) );
  INV_X1 U23719 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20877) );
  OAI222_X1 U23720 ( .A1(n20780), .A2(n20746), .B1(n20877), .B2(n20809), .C1(
        n20748), .C2(n20784), .ZN(P1_U3204) );
  INV_X1 U23721 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20747) );
  OAI222_X1 U23722 ( .A1(n20780), .A2(n20748), .B1(n20747), .B2(n20809), .C1(
        n20750), .C2(n20784), .ZN(P1_U3205) );
  INV_X1 U23723 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20749) );
  OAI222_X1 U23724 ( .A1(n20780), .A2(n20750), .B1(n20749), .B2(n20809), .C1(
        n14877), .C2(n20784), .ZN(P1_U3206) );
  INV_X1 U23725 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20751) );
  OAI222_X1 U23726 ( .A1(n20780), .A2(n14877), .B1(n20751), .B2(n20809), .C1(
        n20753), .C2(n20784), .ZN(P1_U3207) );
  INV_X1 U23727 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20752) );
  OAI222_X1 U23728 ( .A1(n20780), .A2(n20753), .B1(n20752), .B2(n20809), .C1(
        n20755), .C2(n20784), .ZN(P1_U3208) );
  INV_X1 U23729 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20754) );
  OAI222_X1 U23730 ( .A1(n20780), .A2(n20755), .B1(n20754), .B2(n20809), .C1(
        n20756), .C2(n20784), .ZN(P1_U3209) );
  INV_X1 U23731 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20757) );
  OAI222_X1 U23732 ( .A1(n20784), .A2(n20759), .B1(n20757), .B2(n20809), .C1(
        n20756), .C2(n20780), .ZN(P1_U3210) );
  AOI22_X1 U23733 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n20807), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20786), .ZN(n20758) );
  OAI21_X1 U23734 ( .B1(n20759), .B2(n20780), .A(n20758), .ZN(P1_U3211) );
  AOI22_X1 U23735 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20807), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20786), .ZN(n20760) );
  OAI21_X1 U23736 ( .B1(n14829), .B2(n20780), .A(n20760), .ZN(P1_U3212) );
  AOI22_X1 U23737 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20807), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20787), .ZN(n20761) );
  OAI21_X1 U23738 ( .B1(n20763), .B2(n20784), .A(n20761), .ZN(P1_U3213) );
  INV_X1 U23739 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20762) );
  INV_X1 U23740 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20765) );
  OAI222_X1 U23741 ( .A1(n20780), .A2(n20763), .B1(n20762), .B2(n20809), .C1(
        n20765), .C2(n20784), .ZN(P1_U3214) );
  AOI22_X1 U23742 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20807), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20786), .ZN(n20764) );
  OAI21_X1 U23743 ( .B1(n20765), .B2(n20780), .A(n20764), .ZN(P1_U3215) );
  AOI22_X1 U23744 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20807), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20787), .ZN(n20766) );
  OAI21_X1 U23745 ( .B1(n20768), .B2(n20784), .A(n20766), .ZN(P1_U3216) );
  INV_X1 U23746 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20767) );
  OAI222_X1 U23747 ( .A1(n20780), .A2(n20768), .B1(n20767), .B2(n20809), .C1(
        n20770), .C2(n20784), .ZN(P1_U3217) );
  AOI22_X1 U23748 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20807), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20786), .ZN(n20769) );
  OAI21_X1 U23749 ( .B1(n20770), .B2(n20780), .A(n20769), .ZN(P1_U3218) );
  AOI22_X1 U23750 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20807), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20787), .ZN(n20771) );
  OAI21_X1 U23751 ( .B1(n20773), .B2(n20784), .A(n20771), .ZN(P1_U3219) );
  INV_X1 U23752 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20772) );
  OAI222_X1 U23753 ( .A1(n20780), .A2(n20773), .B1(n20772), .B2(n20809), .C1(
        n20775), .C2(n20784), .ZN(P1_U3220) );
  INV_X1 U23754 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20774) );
  OAI222_X1 U23755 ( .A1(n20780), .A2(n20775), .B1(n20774), .B2(n20809), .C1(
        n20776), .C2(n20784), .ZN(P1_U3221) );
  INV_X1 U23756 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20777) );
  OAI222_X1 U23757 ( .A1(n20784), .A2(n20779), .B1(n20777), .B2(n20809), .C1(
        n20776), .C2(n20780), .ZN(P1_U3222) );
  INV_X1 U23758 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20778) );
  OAI222_X1 U23759 ( .A1(n20780), .A2(n20779), .B1(n20778), .B2(n20809), .C1(
        n20781), .C2(n20784), .ZN(P1_U3223) );
  INV_X1 U23760 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20782) );
  OAI222_X1 U23761 ( .A1(n20784), .A2(n20783), .B1(n20782), .B2(n20809), .C1(
        n20781), .C2(n20780), .ZN(P1_U3224) );
  AOI222_X1 U23762 ( .A1(n20787), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20807), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n20786), .ZN(n20785) );
  INV_X1 U23763 ( .A(n20785), .ZN(P1_U3225) );
  AOI222_X1 U23764 ( .A1(n20787), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20807), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20786), .ZN(n20788) );
  INV_X1 U23765 ( .A(n20788), .ZN(P1_U3226) );
  INV_X1 U23766 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20789) );
  AOI22_X1 U23767 ( .A1(n20809), .A2(n20790), .B1(n20789), .B2(n20807), .ZN(
        P1_U3458) );
  INV_X1 U23768 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20802) );
  INV_X1 U23769 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20791) );
  AOI22_X1 U23770 ( .A1(n20809), .A2(n20802), .B1(n20791), .B2(n20807), .ZN(
        P1_U3459) );
  INV_X1 U23771 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20792) );
  AOI22_X1 U23772 ( .A1(n20809), .A2(n20793), .B1(n20792), .B2(n20807), .ZN(
        P1_U3460) );
  INV_X1 U23773 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20828) );
  INV_X1 U23774 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20794) );
  AOI22_X1 U23775 ( .A1(n20809), .A2(n20828), .B1(n20794), .B2(n20807), .ZN(
        P1_U3461) );
  OAI21_X1 U23776 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20798), .A(n20796), 
        .ZN(n20795) );
  INV_X1 U23777 ( .A(n20795), .ZN(P1_U3464) );
  INV_X1 U23778 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20797) );
  OAI21_X1 U23779 ( .B1(n20798), .B2(n20797), .A(n20796), .ZN(P1_U3465) );
  INV_X1 U23780 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20800) );
  NOR3_X1 U23781 ( .A1(n20800), .A2(P1_REIP_REG_0__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .ZN(n20799) );
  AOI221_X1 U23782 ( .B1(n20801), .B2(n20800), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n20799), .ZN(n20803) );
  INV_X1 U23783 ( .A(n20806), .ZN(n20804) );
  AOI22_X1 U23784 ( .A1(n20806), .A2(n20803), .B1(n20802), .B2(n20804), .ZN(
        P1_U3481) );
  NOR2_X1 U23785 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20805) );
  AOI22_X1 U23786 ( .A1(n20806), .A2(n20805), .B1(n20828), .B2(n20804), .ZN(
        P1_U3482) );
  AOI22_X1 U23787 ( .A1(n20809), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20808), 
        .B2(n20807), .ZN(P1_U3483) );
  AOI211_X1 U23788 ( .C1(n20813), .C2(n20812), .A(n20811), .B(n20810), .ZN(
        n20816) );
  OAI21_X1 U23789 ( .B1(n20816), .B2(n20815), .A(n20814), .ZN(n20822) );
  AOI211_X1 U23790 ( .C1(n20820), .C2(n20819), .A(n20818), .B(n20817), .ZN(
        n20821) );
  MUX2_X1 U23791 ( .A(n20822), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20821), 
        .Z(P1_U3485) );
  MUX2_X1 U23792 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20809), .Z(P1_U3486) );
  AOI222_X1 U23793 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n20825), .B1(n20824), 
        .B2(P3_LWORD_REG_5__SCAN_IN), .C1(n20823), .C2(P3_DATAO_REG_5__SCAN_IN), .ZN(n21074) );
  INV_X1 U23794 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n21101) );
  AOI22_X1 U23795 ( .A1(n21101), .A2(keyinput66), .B1(keyinput106), .B2(n13106), .ZN(n20826) );
  OAI221_X1 U23796 ( .B1(n21101), .B2(keyinput66), .C1(n13106), .C2(
        keyinput106), .A(n20826), .ZN(n20838) );
  AOI22_X1 U23797 ( .A1(n20829), .A2(keyinput17), .B1(keyinput5), .B2(n20828), 
        .ZN(n20827) );
  OAI221_X1 U23798 ( .B1(n20829), .B2(keyinput17), .C1(n20828), .C2(keyinput5), 
        .A(n20827), .ZN(n20837) );
  AOI22_X1 U23799 ( .A1(n20831), .A2(keyinput8), .B1(keyinput88), .B2(n13423), 
        .ZN(n20830) );
  OAI221_X1 U23800 ( .B1(n20831), .B2(keyinput8), .C1(n13423), .C2(keyinput88), 
        .A(n20830), .ZN(n20836) );
  INV_X1 U23801 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20834) );
  AOI22_X1 U23802 ( .A1(n20834), .A2(keyinput100), .B1(keyinput3), .B2(n20833), 
        .ZN(n20832) );
  OAI221_X1 U23803 ( .B1(n20834), .B2(keyinput100), .C1(n20833), .C2(keyinput3), .A(n20832), .ZN(n20835) );
  NOR4_X1 U23804 ( .A1(n20838), .A2(n20837), .A3(n20836), .A4(n20835), .ZN(
        n20885) );
  INV_X1 U23805 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n20840) );
  AOI22_X1 U23806 ( .A1(n20840), .A2(keyinput63), .B1(n21076), .B2(keyinput61), 
        .ZN(n20839) );
  OAI221_X1 U23807 ( .B1(n20840), .B2(keyinput63), .C1(n21076), .C2(keyinput61), .A(n20839), .ZN(n20845) );
  XNOR2_X1 U23808 ( .A(n20841), .B(keyinput109), .ZN(n20844) );
  XNOR2_X1 U23809 ( .A(n20842), .B(keyinput54), .ZN(n20843) );
  OR3_X1 U23810 ( .A1(n20845), .A2(n20844), .A3(n20843), .ZN(n20853) );
  AOI22_X1 U23811 ( .A1(n20848), .A2(keyinput95), .B1(n20847), .B2(keyinput78), 
        .ZN(n20846) );
  OAI221_X1 U23812 ( .B1(n20848), .B2(keyinput95), .C1(n20847), .C2(keyinput78), .A(n20846), .ZN(n20852) );
  AOI22_X1 U23813 ( .A1(n20850), .A2(keyinput124), .B1(n13090), .B2(keyinput53), .ZN(n20849) );
  OAI221_X1 U23814 ( .B1(n20850), .B2(keyinput124), .C1(n13090), .C2(
        keyinput53), .A(n20849), .ZN(n20851) );
  NOR3_X1 U23815 ( .A1(n20853), .A2(n20852), .A3(n20851), .ZN(n20884) );
  AOI22_X1 U23816 ( .A1(n20856), .A2(keyinput58), .B1(keyinput111), .B2(n20855), .ZN(n20854) );
  OAI221_X1 U23817 ( .B1(n20856), .B2(keyinput58), .C1(n20855), .C2(
        keyinput111), .A(n20854), .ZN(n20866) );
  AOI22_X1 U23818 ( .A1(n20859), .A2(keyinput75), .B1(n20858), .B2(keyinput11), 
        .ZN(n20857) );
  OAI221_X1 U23819 ( .B1(n20859), .B2(keyinput75), .C1(n20858), .C2(keyinput11), .A(n20857), .ZN(n20865) );
  INV_X1 U23820 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n21102) );
  XNOR2_X1 U23821 ( .A(n21102), .B(keyinput52), .ZN(n20864) );
  XNOR2_X1 U23822 ( .A(n21077), .B(keyinput41), .ZN(n20862) );
  XNOR2_X1 U23823 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(keyinput96), 
        .ZN(n20861) );
  XNOR2_X1 U23824 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B(keyinput62), .ZN(
        n20860) );
  NAND3_X1 U23825 ( .A1(n20862), .A2(n20861), .A3(n20860), .ZN(n20863) );
  NOR4_X1 U23826 ( .A1(n20866), .A2(n20865), .A3(n20864), .A4(n20863), .ZN(
        n20883) );
  AOI22_X1 U23827 ( .A1(n20869), .A2(keyinput122), .B1(n20868), .B2(keyinput86), .ZN(n20867) );
  OAI221_X1 U23828 ( .B1(n20869), .B2(keyinput122), .C1(n20868), .C2(
        keyinput86), .A(n20867), .ZN(n20881) );
  INV_X1 U23829 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n20871) );
  AOI22_X1 U23830 ( .A1(n20872), .A2(keyinput60), .B1(n20871), .B2(keyinput7), 
        .ZN(n20870) );
  OAI221_X1 U23831 ( .B1(n20872), .B2(keyinput60), .C1(n20871), .C2(keyinput7), 
        .A(n20870), .ZN(n20880) );
  AOI22_X1 U23832 ( .A1(n20877), .A2(keyinput73), .B1(n21075), .B2(keyinput30), 
        .ZN(n20876) );
  OAI221_X1 U23833 ( .B1(n20877), .B2(keyinput73), .C1(n21075), .C2(keyinput30), .A(n20876), .ZN(n20878) );
  NOR4_X1 U23834 ( .A1(n20881), .A2(n20880), .A3(n20879), .A4(n20878), .ZN(
        n20882) );
  NAND4_X1 U23835 ( .A1(n20885), .A2(n20884), .A3(n20883), .A4(n20882), .ZN(
        n21072) );
  AOI22_X1 U23836 ( .A1(n20887), .A2(keyinput104), .B1(n11406), .B2(keyinput89), .ZN(n20886) );
  OAI221_X1 U23837 ( .B1(n20887), .B2(keyinput104), .C1(n11406), .C2(
        keyinput89), .A(n20886), .ZN(n20897) );
  AOI22_X1 U23838 ( .A1(n12005), .A2(keyinput37), .B1(keyinput4), .B2(n20889), 
        .ZN(n20888) );
  OAI221_X1 U23839 ( .B1(n12005), .B2(keyinput37), .C1(n20889), .C2(keyinput4), 
        .A(n20888), .ZN(n20896) );
  AOI22_X1 U23840 ( .A1(n20891), .A2(keyinput76), .B1(n13431), .B2(keyinput26), 
        .ZN(n20890) );
  OAI221_X1 U23841 ( .B1(n20891), .B2(keyinput76), .C1(n13431), .C2(keyinput26), .A(n20890), .ZN(n20895) );
  XOR2_X1 U23842 ( .A(n13403), .B(keyinput101), .Z(n20893) );
  XNOR2_X1 U23843 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B(keyinput27), .ZN(
        n20892) );
  NAND2_X1 U23844 ( .A1(n20893), .A2(n20892), .ZN(n20894) );
  NOR4_X1 U23845 ( .A1(n20897), .A2(n20896), .A3(n20895), .A4(n20894), .ZN(
        n20944) );
  AOI22_X1 U23846 ( .A1(n20899), .A2(keyinput114), .B1(n11461), .B2(keyinput28), .ZN(n20898) );
  OAI221_X1 U23847 ( .B1(n20899), .B2(keyinput114), .C1(n11461), .C2(
        keyinput28), .A(n20898), .ZN(n20910) );
  AOI22_X1 U23848 ( .A1(n13441), .A2(keyinput51), .B1(n13077), .B2(keyinput1), 
        .ZN(n20900) );
  OAI221_X1 U23849 ( .B1(n13441), .B2(keyinput51), .C1(n13077), .C2(keyinput1), 
        .A(n20900), .ZN(n20909) );
  AOI22_X1 U23850 ( .A1(n20903), .A2(keyinput39), .B1(n20902), .B2(keyinput83), 
        .ZN(n20901) );
  OAI221_X1 U23851 ( .B1(n20903), .B2(keyinput39), .C1(n20902), .C2(keyinput83), .A(n20901), .ZN(n20908) );
  INV_X1 U23852 ( .A(P3_UWORD_REG_5__SCAN_IN), .ZN(n20905) );
  AOI22_X1 U23853 ( .A1(n20906), .A2(keyinput110), .B1(keyinput15), .B2(n20905), .ZN(n20904) );
  OAI221_X1 U23854 ( .B1(n20906), .B2(keyinput110), .C1(n20905), .C2(
        keyinput15), .A(n20904), .ZN(n20907) );
  NOR4_X1 U23855 ( .A1(n20910), .A2(n20909), .A3(n20908), .A4(n20907), .ZN(
        n20943) );
  INV_X1 U23856 ( .A(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n20912) );
  AOI22_X1 U23857 ( .A1(n9888), .A2(keyinput115), .B1(keyinput33), .B2(n20912), 
        .ZN(n20911) );
  OAI221_X1 U23858 ( .B1(n9888), .B2(keyinput115), .C1(n20912), .C2(keyinput33), .A(n20911), .ZN(n20924) );
  INV_X1 U23859 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n20914) );
  AOI22_X1 U23860 ( .A1(n20914), .A2(keyinput44), .B1(n9892), .B2(keyinput18), 
        .ZN(n20913) );
  OAI221_X1 U23861 ( .B1(n20914), .B2(keyinput44), .C1(n9892), .C2(keyinput18), 
        .A(n20913), .ZN(n20923) );
  AOI22_X1 U23862 ( .A1(n20917), .A2(keyinput125), .B1(n20916), .B2(keyinput79), .ZN(n20915) );
  OAI221_X1 U23863 ( .B1(n20917), .B2(keyinput125), .C1(n20916), .C2(
        keyinput79), .A(n20915), .ZN(n20922) );
  AOI22_X1 U23864 ( .A1(n20920), .A2(keyinput20), .B1(keyinput64), .B2(n20919), 
        .ZN(n20918) );
  OAI221_X1 U23865 ( .B1(n20920), .B2(keyinput20), .C1(n20919), .C2(keyinput64), .A(n20918), .ZN(n20921) );
  NOR4_X1 U23866 ( .A1(n20924), .A2(n20923), .A3(n20922), .A4(n20921), .ZN(
        n20942) );
  INV_X1 U23867 ( .A(P3_LWORD_REG_4__SCAN_IN), .ZN(n20927) );
  INV_X1 U23868 ( .A(P3_LWORD_REG_5__SCAN_IN), .ZN(n20926) );
  AOI22_X1 U23869 ( .A1(n20927), .A2(keyinput118), .B1(n20926), .B2(
        keyinput123), .ZN(n20925) );
  OAI221_X1 U23870 ( .B1(n20927), .B2(keyinput118), .C1(n20926), .C2(
        keyinput123), .A(n20925), .ZN(n20931) );
  XNOR2_X1 U23871 ( .A(n20928), .B(keyinput98), .ZN(n20930) );
  XOR2_X1 U23872 ( .A(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B(keyinput107), .Z(
        n20929) );
  OR3_X1 U23873 ( .A1(n20931), .A2(n20930), .A3(n20929), .ZN(n20940) );
  AOI22_X1 U23874 ( .A1(n20934), .A2(keyinput0), .B1(keyinput99), .B2(n20933), 
        .ZN(n20932) );
  OAI221_X1 U23875 ( .B1(n20934), .B2(keyinput0), .C1(n20933), .C2(keyinput99), 
        .A(n20932), .ZN(n20939) );
  AOI22_X1 U23876 ( .A1(n20937), .A2(keyinput14), .B1(n20936), .B2(keyinput36), 
        .ZN(n20935) );
  OAI221_X1 U23877 ( .B1(n20937), .B2(keyinput14), .C1(n20936), .C2(keyinput36), .A(n20935), .ZN(n20938) );
  NOR3_X1 U23878 ( .A1(n20940), .A2(n20939), .A3(n20938), .ZN(n20941) );
  NAND4_X1 U23879 ( .A1(n20944), .A2(n20943), .A3(n20942), .A4(n20941), .ZN(
        n21071) );
  AOI22_X1 U23880 ( .A1(n20947), .A2(keyinput121), .B1(keyinput56), .B2(n20946), .ZN(n20945) );
  OAI221_X1 U23881 ( .B1(n20947), .B2(keyinput121), .C1(n20946), .C2(
        keyinput56), .A(n20945), .ZN(n20959) );
  AOI22_X1 U23882 ( .A1(n20950), .A2(keyinput6), .B1(keyinput91), .B2(n20949), 
        .ZN(n20948) );
  OAI221_X1 U23883 ( .B1(n20950), .B2(keyinput6), .C1(n20949), .C2(keyinput91), 
        .A(n20948), .ZN(n20958) );
  INV_X1 U23884 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n20952) );
  AOI22_X1 U23885 ( .A1(n20953), .A2(keyinput120), .B1(keyinput38), .B2(n20952), .ZN(n20951) );
  OAI221_X1 U23886 ( .B1(n20953), .B2(keyinput120), .C1(n20952), .C2(
        keyinput38), .A(n20951), .ZN(n20957) );
  XOR2_X1 U23887 ( .A(n13105), .B(keyinput80), .Z(n20955) );
  XNOR2_X1 U23888 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput46), 
        .ZN(n20954) );
  NAND2_X1 U23889 ( .A1(n20955), .A2(n20954), .ZN(n20956) );
  NOR4_X1 U23890 ( .A1(n20959), .A2(n20958), .A3(n20957), .A4(n20956), .ZN(
        n21006) );
  AOI22_X1 U23891 ( .A1(n13418), .A2(keyinput72), .B1(keyinput49), .B2(n20961), 
        .ZN(n20960) );
  OAI221_X1 U23892 ( .B1(n13418), .B2(keyinput72), .C1(n20961), .C2(keyinput49), .A(n20960), .ZN(n20972) );
  INV_X1 U23893 ( .A(P3_LWORD_REG_10__SCAN_IN), .ZN(n20963) );
  AOI22_X1 U23894 ( .A1(n20963), .A2(keyinput71), .B1(n21100), .B2(keyinput67), 
        .ZN(n20962) );
  OAI221_X1 U23895 ( .B1(n20963), .B2(keyinput71), .C1(n21100), .C2(keyinput67), .A(n20962), .ZN(n20971) );
  AOI22_X1 U23896 ( .A1(n20966), .A2(keyinput82), .B1(keyinput57), .B2(n20965), 
        .ZN(n20964) );
  OAI221_X1 U23897 ( .B1(n20966), .B2(keyinput82), .C1(n20965), .C2(keyinput57), .A(n20964), .ZN(n20970) );
  INV_X1 U23898 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n20968) );
  AOI22_X1 U23899 ( .A1(n20968), .A2(keyinput103), .B1(n10603), .B2(keyinput90), .ZN(n20967) );
  OAI221_X1 U23900 ( .B1(n20968), .B2(keyinput103), .C1(n10603), .C2(
        keyinput90), .A(n20967), .ZN(n20969) );
  NOR4_X1 U23901 ( .A1(n20972), .A2(n20971), .A3(n20970), .A4(n20969), .ZN(
        n21005) );
  AOI22_X1 U23902 ( .A1(n20975), .A2(keyinput55), .B1(n20974), .B2(keyinput116), .ZN(n20973) );
  OAI221_X1 U23903 ( .B1(n20975), .B2(keyinput55), .C1(n20974), .C2(
        keyinput116), .A(n20973), .ZN(n20987) );
  AOI22_X1 U23904 ( .A1(n20978), .A2(keyinput25), .B1(n20977), .B2(keyinput22), 
        .ZN(n20976) );
  OAI221_X1 U23905 ( .B1(n20978), .B2(keyinput25), .C1(n20977), .C2(keyinput22), .A(n20976), .ZN(n20986) );
  AOI22_X1 U23906 ( .A1(n20981), .A2(keyinput32), .B1(n20980), .B2(keyinput119), .ZN(n20979) );
  OAI221_X1 U23907 ( .B1(n20981), .B2(keyinput32), .C1(n20980), .C2(
        keyinput119), .A(n20979), .ZN(n20985) );
  XNOR2_X1 U23908 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B(keyinput126), .ZN(
        n20983) );
  XNOR2_X1 U23909 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B(keyinput12), 
        .ZN(n20982) );
  NAND2_X1 U23910 ( .A1(n20983), .A2(n20982), .ZN(n20984) );
  NOR4_X1 U23911 ( .A1(n20987), .A2(n20986), .A3(n20985), .A4(n20984), .ZN(
        n21004) );
  AOI22_X1 U23912 ( .A1(n20990), .A2(keyinput112), .B1(keyinput94), .B2(n20989), .ZN(n20988) );
  OAI221_X1 U23913 ( .B1(n20990), .B2(keyinput112), .C1(n20989), .C2(
        keyinput94), .A(n20988), .ZN(n21002) );
  AOI22_X1 U23914 ( .A1(n20993), .A2(keyinput31), .B1(n20992), .B2(keyinput21), 
        .ZN(n20991) );
  OAI221_X1 U23915 ( .B1(n20993), .B2(keyinput31), .C1(n20992), .C2(keyinput21), .A(n20991), .ZN(n21001) );
  AOI22_X1 U23916 ( .A1(n13427), .A2(keyinput23), .B1(keyinput102), .B2(n20995), .ZN(n20994) );
  OAI221_X1 U23917 ( .B1(n13427), .B2(keyinput23), .C1(n20995), .C2(
        keyinput102), .A(n20994), .ZN(n21000) );
  AOI22_X1 U23918 ( .A1(n20998), .A2(keyinput16), .B1(n20997), .B2(keyinput65), 
        .ZN(n20996) );
  OAI221_X1 U23919 ( .B1(n20998), .B2(keyinput16), .C1(n20997), .C2(keyinput65), .A(n20996), .ZN(n20999) );
  NOR4_X1 U23920 ( .A1(n21002), .A2(n21001), .A3(n21000), .A4(n20999), .ZN(
        n21003) );
  NAND4_X1 U23921 ( .A1(n21006), .A2(n21005), .A3(n21004), .A4(n21003), .ZN(
        n21070) );
  AOI22_X1 U23922 ( .A1(n12966), .A2(keyinput113), .B1(keyinput77), .B2(n21008), .ZN(n21007) );
  OAI221_X1 U23923 ( .B1(n12966), .B2(keyinput113), .C1(n21008), .C2(
        keyinput77), .A(n21007), .ZN(n21020) );
  AOI22_X1 U23924 ( .A1(n21011), .A2(keyinput105), .B1(keyinput34), .B2(n21010), .ZN(n21009) );
  OAI221_X1 U23925 ( .B1(n21011), .B2(keyinput105), .C1(n21010), .C2(
        keyinput34), .A(n21009), .ZN(n21019) );
  AOI22_X1 U23926 ( .A1(n21014), .A2(keyinput42), .B1(n21013), .B2(keyinput85), 
        .ZN(n21012) );
  OAI221_X1 U23927 ( .B1(n21014), .B2(keyinput42), .C1(n21013), .C2(keyinput85), .A(n21012), .ZN(n21018) );
  XOR2_X1 U23928 ( .A(n11552), .B(keyinput50), .Z(n21016) );
  XNOR2_X1 U23929 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B(keyinput40), .ZN(
        n21015) );
  NAND2_X1 U23930 ( .A1(n21016), .A2(n21015), .ZN(n21017) );
  NOR4_X1 U23931 ( .A1(n21020), .A2(n21019), .A3(n21018), .A4(n21017), .ZN(
        n21068) );
  AOI22_X1 U23932 ( .A1(n21022), .A2(keyinput2), .B1(keyinput81), .B2(n13098), 
        .ZN(n21021) );
  OAI221_X1 U23933 ( .B1(n21022), .B2(keyinput2), .C1(n13098), .C2(keyinput81), 
        .A(n21021), .ZN(n21026) );
  XOR2_X1 U23934 ( .A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B(keyinput48), .Z(
        n21025) );
  XNOR2_X1 U23935 ( .A(n21023), .B(keyinput74), .ZN(n21024) );
  OR3_X1 U23936 ( .A1(n21026), .A2(n21025), .A3(n21024), .ZN(n21034) );
  INV_X1 U23937 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n21029) );
  INV_X1 U23938 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n21028) );
  AOI22_X1 U23939 ( .A1(n21029), .A2(keyinput117), .B1(keyinput59), .B2(n21028), .ZN(n21027) );
  OAI221_X1 U23940 ( .B1(n21029), .B2(keyinput117), .C1(n21028), .C2(
        keyinput59), .A(n21027), .ZN(n21033) );
  AOI22_X1 U23941 ( .A1(n12242), .A2(keyinput10), .B1(keyinput69), .B2(n21031), 
        .ZN(n21030) );
  OAI221_X1 U23942 ( .B1(n12242), .B2(keyinput10), .C1(n21031), .C2(keyinput69), .A(n21030), .ZN(n21032) );
  NOR3_X1 U23943 ( .A1(n21034), .A2(n21033), .A3(n21032), .ZN(n21067) );
  AOI22_X1 U23944 ( .A1(n21037), .A2(keyinput47), .B1(n21036), .B2(keyinput9), 
        .ZN(n21035) );
  OAI221_X1 U23945 ( .B1(n21037), .B2(keyinput47), .C1(n21036), .C2(keyinput9), 
        .A(n21035), .ZN(n21049) );
  AOI22_X1 U23946 ( .A1(n21040), .A2(keyinput70), .B1(n21039), .B2(keyinput35), 
        .ZN(n21038) );
  OAI221_X1 U23947 ( .B1(n21040), .B2(keyinput70), .C1(n21039), .C2(keyinput35), .A(n21038), .ZN(n21048) );
  INV_X1 U23948 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n21043) );
  AOI22_X1 U23949 ( .A1(n21043), .A2(keyinput68), .B1(n21042), .B2(keyinput29), 
        .ZN(n21041) );
  OAI221_X1 U23950 ( .B1(n21043), .B2(keyinput68), .C1(n21042), .C2(keyinput29), .A(n21041), .ZN(n21047) );
  AOI22_X1 U23951 ( .A1(n12030), .A2(keyinput92), .B1(keyinput93), .B2(n21045), 
        .ZN(n21044) );
  OAI221_X1 U23952 ( .B1(n12030), .B2(keyinput92), .C1(n21045), .C2(keyinput93), .A(n21044), .ZN(n21046) );
  NOR4_X1 U23953 ( .A1(n21049), .A2(n21048), .A3(n21047), .A4(n21046), .ZN(
        n21066) );
  INV_X1 U23954 ( .A(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n21052) );
  AOI22_X1 U23955 ( .A1(n21052), .A2(keyinput97), .B1(keyinput13), .B2(n21051), 
        .ZN(n21050) );
  OAI221_X1 U23956 ( .B1(n21052), .B2(keyinput97), .C1(n21051), .C2(keyinput13), .A(n21050), .ZN(n21064) );
  INV_X1 U23957 ( .A(P3_MORE_REG_SCAN_IN), .ZN(n21055) );
  AOI22_X1 U23958 ( .A1(n21055), .A2(keyinput127), .B1(keyinput19), .B2(n21054), .ZN(n21053) );
  OAI221_X1 U23959 ( .B1(n21055), .B2(keyinput127), .C1(n21054), .C2(
        keyinput19), .A(n21053), .ZN(n21063) );
  INV_X1 U23960 ( .A(READY21_REG_SCAN_IN), .ZN(n21057) );
  AOI22_X1 U23961 ( .A1(n21058), .A2(keyinput87), .B1(n21057), .B2(keyinput43), 
        .ZN(n21056) );
  OAI221_X1 U23962 ( .B1(n21058), .B2(keyinput87), .C1(n21057), .C2(keyinput43), .A(n21056), .ZN(n21062) );
  AOI22_X1 U23963 ( .A1(n13262), .A2(keyinput84), .B1(keyinput45), .B2(n21060), 
        .ZN(n21059) );
  OAI221_X1 U23964 ( .B1(n13262), .B2(keyinput84), .C1(n21060), .C2(keyinput45), .A(n21059), .ZN(n21061) );
  NOR4_X1 U23965 ( .A1(n21064), .A2(n21063), .A3(n21062), .A4(n21061), .ZN(
        n21065) );
  NAND4_X1 U23966 ( .A1(n21068), .A2(n21067), .A3(n21066), .A4(n21065), .ZN(
        n21069) );
  NOR4_X1 U23967 ( .A1(n21072), .A2(n21071), .A3(n21070), .A4(n21069), .ZN(
        n21073) );
  XNOR2_X1 U23968 ( .A(n21074), .B(n21073), .ZN(n21124) );
  NAND4_X1 U23969 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(
        P2_DATAO_REG_12__SCAN_IN), .A3(P2_DATAO_REG_5__SCAN_IN), .A4(
        P2_ADS_N_REG_SCAN_IN), .ZN(n21087) );
  NAND4_X1 U23970 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(
        P3_ADDRESS_REG_27__SCAN_IN), .A3(n21076), .A4(n21075), .ZN(n21086) );
  NOR4_X1 U23971 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A4(P1_EBX_REG_12__SCAN_IN), .ZN(
        n21084) );
  NOR4_X1 U23972 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_3__6__SCAN_IN), .A3(P1_INSTQUEUE_REG_15__7__SCAN_IN), 
        .A4(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n21083) );
  NAND4_X1 U23973 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(P1_UWORD_REG_13__SCAN_IN), .A3(P1_LWORD_REG_6__SCAN_IN), .A4(P1_DATAO_REG_7__SCAN_IN), .ZN(n21081) );
  NAND4_X1 U23974 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_MORE_REG_SCAN_IN), .A3(P1_LWORD_REG_5__SCAN_IN), .A4(
        P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21080) );
  NAND4_X1 U23975 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(P2_REIP_REG_14__SCAN_IN), .A4(
        P2_EAX_REG_8__SCAN_IN), .ZN(n21079) );
  NAND4_X1 U23976 ( .A1(n21077), .A2(READY21_REG_SCAN_IN), .A3(
        BUF1_REG_9__SCAN_IN), .A4(P2_LWORD_REG_2__SCAN_IN), .ZN(n21078) );
  NOR4_X1 U23977 ( .A1(n21081), .A2(n21080), .A3(n21079), .A4(n21078), .ZN(
        n21082) );
  NAND3_X1 U23978 ( .A1(n21084), .A2(n21083), .A3(n21082), .ZN(n21085) );
  NOR3_X1 U23979 ( .A1(n21087), .A2(n21086), .A3(n21085), .ZN(n21122) );
  NAND4_X1 U23980 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_5__1__SCAN_IN), .A3(P1_INSTQUEUE_REG_8__4__SCAN_IN), 
        .A4(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n21091) );
  NAND4_X1 U23981 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_12__2__SCAN_IN), .A3(P2_INSTQUEUE_REG_8__5__SCAN_IN), 
        .A4(BUF2_REG_19__SCAN_IN), .ZN(n21090) );
  NAND4_X1 U23982 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_10__6__SCAN_IN), .A3(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A4(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n21089) );
  NAND4_X1 U23983 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_14__5__SCAN_IN), .A3(P1_INSTQUEUE_REG_4__2__SCAN_IN), 
        .A4(BUF1_REG_26__SCAN_IN), .ZN(n21088) );
  NOR4_X1 U23984 ( .A1(n21091), .A2(n21090), .A3(n21089), .A4(n21088), .ZN(
        n21121) );
  NAND4_X1 U23985 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_23__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_24__SCAN_IN), .ZN(n21095) );
  NAND4_X1 U23986 ( .A1(P2_EBX_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n21094) );
  NAND4_X1 U23987 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        BUF1_REG_21__SCAN_IN), .A3(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A4(
        P1_DATAO_REG_24__SCAN_IN), .ZN(n21093) );
  NAND4_X1 U23988 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_EAX_REG_16__SCAN_IN), .A3(P3_EAX_REG_8__SCAN_IN), .A4(
        P3_DATAO_REG_19__SCAN_IN), .ZN(n21092) );
  NOR4_X1 U23989 ( .A1(n21095), .A2(n21094), .A3(n21093), .A4(n21092), .ZN(
        n21120) );
  NOR4_X1 U23990 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(
        P1_LWORD_REG_13__SCAN_IN), .A3(P1_DATAO_REG_12__SCAN_IN), .A4(
        P1_DATAO_REG_2__SCAN_IN), .ZN(n21099) );
  NOR4_X1 U23991 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_EBX_REG_2__SCAN_IN), .A3(P1_ADDRESS_REG_7__SCAN_IN), .A4(
        P3_ADDRESS_REG_29__SCAN_IN), .ZN(n21098) );
  NOR4_X1 U23992 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(P2_EAX_REG_0__SCAN_IN), .A4(
        P2_EAX_REG_17__SCAN_IN), .ZN(n21097) );
  NOR4_X1 U23993 ( .A1(P1_EBX_REG_3__SCAN_IN), .A2(P1_LWORD_REG_14__SCAN_IN), 
        .A3(P1_DATAO_REG_15__SCAN_IN), .A4(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(
        n21096) );
  NAND4_X1 U23994 ( .A1(n21099), .A2(n21098), .A3(n21097), .A4(n21096), .ZN(
        n21118) );
  NOR4_X1 U23995 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .A3(P3_INSTQUEUE_REG_8__3__SCAN_IN), 
        .A4(n21100), .ZN(n21106) );
  NOR4_X1 U23996 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_16__SCAN_IN), .A4(
        n21101), .ZN(n21105) );
  NOR4_X1 U23997 ( .A1(P2_ADDRESS_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_31__SCAN_IN), .A3(P3_LWORD_REG_10__SCAN_IN), .A4(
        P3_ADDRESS_REG_26__SCAN_IN), .ZN(n21104) );
  NOR4_X1 U23998 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_LWORD_REG_5__SCAN_IN), .A3(P3_ADDRESS_REG_17__SCAN_IN), .A4(n21102), 
        .ZN(n21103) );
  NAND4_X1 U23999 ( .A1(n21106), .A2(n21105), .A3(n21104), .A4(n21103), .ZN(
        n21117) );
  NOR4_X1 U24000 ( .A1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_5__1__SCAN_IN), .A3(P2_REIP_REG_7__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n21110) );
  NOR4_X1 U24001 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .A3(P3_REIP_REG_21__SCAN_IN), .A4(P3_REIP_REG_19__SCAN_IN), .ZN(n21109) );
  NOR4_X1 U24002 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_EAX_REG_28__SCAN_IN), .A3(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21108) );
  NOR4_X1 U24003 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_6__4__SCAN_IN), .A3(P2_INSTQUEUE_REG_11__3__SCAN_IN), 
        .A4(BUF2_REG_27__SCAN_IN), .ZN(n21107) );
  NAND4_X1 U24004 ( .A1(n21110), .A2(n21109), .A3(n21108), .A4(n21107), .ZN(
        n21116) );
  NOR4_X1 U24005 ( .A1(P3_MORE_REG_SCAN_IN), .A2(P2_DATAWIDTH_REG_28__SCAN_IN), 
        .A3(P2_CODEFETCH_REG_SCAN_IN), .A4(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21114) );
  NOR4_X1 U24006 ( .A1(P2_EBX_REG_3__SCAN_IN), .A2(P2_REIP_REG_21__SCAN_IN), 
        .A3(P2_EAX_REG_13__SCAN_IN), .A4(P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(
        n21113) );
  NOR4_X1 U24007 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_4__SCAN_IN), 
        .A3(P3_DATAO_REG_20__SCAN_IN), .A4(P3_UWORD_REG_5__SCAN_IN), .ZN(
        n21112) );
  NOR4_X1 U24008 ( .A1(P3_BYTEENABLE_REG_2__SCAN_IN), .A2(
        P3_LWORD_REG_4__SCAN_IN), .A3(P3_DATAO_REG_13__SCAN_IN), .A4(
        P3_DATAO_REG_18__SCAN_IN), .ZN(n21111) );
  NAND4_X1 U24009 ( .A1(n21114), .A2(n21113), .A3(n21112), .A4(n21111), .ZN(
        n21115) );
  NOR4_X1 U24010 ( .A1(n21118), .A2(n21117), .A3(n21116), .A4(n21115), .ZN(
        n21119) );
  NAND4_X1 U24011 ( .A1(n21122), .A2(n21121), .A3(n21120), .A4(n21119), .ZN(
        n21123) );
  XNOR2_X1 U24012 ( .A(n21124), .B(n21123), .ZN(P3_U2762) );
  AND2_X1 U13034 ( .A1(n10172), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10180) );
  AND2_X2 U13043 ( .A1(n10178), .A2(n10179), .ZN(n10320) );
  NAND2_X1 U13265 ( .A1(n10415), .A2(n10387), .ZN(n10429) );
  BUF_X1 U11375 ( .A(n10416), .Z(n14049) );
  BUF_X1 U11383 ( .A(n10419), .Z(n11073) );
  CLKBUF_X1 U11189 ( .A(n11381), .Z(n15348) );
  CLKBUF_X1 U11249 ( .A(n11354), .Z(n14265) );
  CLKBUF_X1 U11462 ( .A(n14140), .Z(n14311) );
  CLKBUF_X2 U11475 ( .A(n14030), .Z(n13860) );
  CLKBUF_X1 U11477 ( .A(n11233), .Z(n11224) );
  CLKBUF_X1 U11486 ( .A(n14629), .Z(n9738) );
  CLKBUF_X1 U11500 ( .A(n11380), .Z(n13682) );
  CLKBUF_X1 U11659 ( .A(n11246), .Z(n11233) );
  CLKBUF_X1 U11736 ( .A(n13582), .Z(n20464) );
  INV_X1 U12045 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10094) );
  CLKBUF_X1 U12304 ( .A(n16651), .Z(n16656) );
  NAND2_X2 U12469 ( .A1(n10165), .A2(n10328), .ZN(n21125) );
endmodule

