

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4944, n4946, n4947, n4948, n4949, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852;

  OR2_X1 U5008 ( .A1(n5228), .A2(n10162), .ZN(n5157) );
  AND2_X1 U5009 ( .A1(n8815), .A2(n8816), .ZN(n9388) );
  OR2_X1 U5010 ( .A1(n8093), .A2(n5399), .ZN(n5397) );
  OR2_X1 U5011 ( .A1(n7326), .A2(n8313), .ZN(n7462) );
  CLKBUF_X2 U5012 ( .A(n7006), .Z(n8975) );
  INV_X2 U5013 ( .A(n8647), .ZN(n6601) );
  CLKBUF_X2 U5014 ( .A(n9256), .Z(n4947) );
  BUF_X1 U5015 ( .A(n5750), .Z(n8294) );
  NAND2_X2 U5016 ( .A1(n6249), .A2(n9620), .ZN(n8649) );
  NAND2_X2 U5017 ( .A1(n6242), .A2(n6245), .ZN(n8645) );
  CLKBUF_X1 U5018 ( .A(n9759), .Z(n4944) );
  OAI21_X1 U5019 ( .B1(n7025), .B2(n7577), .A(n10729), .ZN(n9759) );
  INV_X1 U5020 ( .A(n8842), .ZN(n8849) );
  INV_X1 U5021 ( .A(n6815), .ZN(n5954) );
  OR2_X2 U5022 ( .A1(n7462), .A2(n8374), .ZN(n7501) );
  NOR2_X1 U5023 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5511) );
  OR2_X1 U5025 ( .A1(n6542), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6551) );
  OAI21_X1 U5026 ( .B1(n9072), .B2(n9044), .A(n9043), .ZN(n9042) );
  INV_X1 U5027 ( .A(n8645), .ZN(n6621) );
  CLKBUF_X3 U5028 ( .A(n9256), .Z(n4946) );
  INV_X1 U5029 ( .A(n6727), .ZN(n6113) );
  INV_X2 U5031 ( .A(n6305), .ZN(n8643) );
  OAI211_X1 U5032 ( .C1(n6815), .C2(n6953), .A(n5769), .B(n5768), .ZN(n7276)
         );
  AND2_X1 U5033 ( .A1(n8564), .A2(n8501), .ZN(n9996) );
  NAND2_X1 U5034 ( .A1(n5858), .A2(n5857), .ZN(n7807) );
  INV_X1 U5035 ( .A(n8287), .ZN(n8332) );
  AOI211_X1 U5036 ( .C1(n10208), .C2(n10814), .A(n10000), .B(n9999), .ZN(
        n10001) );
  AND2_X1 U5037 ( .A1(n5514), .A2(n5513), .ZN(n6744) );
  NAND2_X1 U5038 ( .A1(n6262), .A2(n6261), .ZN(n9256) );
  MUX2_X2 U5039 ( .A(n6627), .B(n8690), .S(n6626), .Z(n8594) );
  NOR2_X2 U5040 ( .A1(n6610), .A2(n8836), .ZN(n9297) );
  NOR2_X2 U5041 ( .A1(n9307), .A2(n8837), .ZN(n6610) );
  NAND2_X2 U5042 ( .A1(n9723), .A2(n9722), .ZN(n9721) );
  NOR2_X2 U5043 ( .A1(n8621), .A2(n8620), .ZN(n8623) );
  AND2_X2 U5044 ( .A1(n4960), .A2(n4961), .ZN(n8621) );
  XNOR2_X2 U5045 ( .A(n6672), .B(n6671), .ZN(n6703) );
  NAND2_X2 U5046 ( .A1(n6176), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6130) );
  XNOR2_X2 U5047 ( .A(n5596), .B(n10522), .ZN(n5757) );
  AOI21_X2 U5048 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n9191), .A(n9190), .ZN(
        n9212) );
  NAND2_X2 U5049 ( .A1(n6136), .A2(n8576), .ZN(n7574) );
  AOI21_X2 U5050 ( .B1(n10027), .B2(n10026), .A(n5075), .ZN(n10003) );
  OAI21_X2 U5051 ( .B1(n10039), .B2(n8472), .A(n8484), .ZN(n10027) );
  INV_X2 U5052 ( .A(n6137), .ZN(n9946) );
  NAND2_X2 U5053 ( .A1(n6252), .A2(n6251), .ZN(n9151) );
  NOR2_X1 U5054 ( .A1(n6248), .A2(n6247), .ZN(n6252) );
  NAND2_X2 U5055 ( .A1(n6099), .A2(n6098), .ZN(n9990) );
  INV_X1 U5056 ( .A(n6242), .ZN(n6249) );
  XNOR2_X2 U5057 ( .A(n6180), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6198) );
  NAND2_X2 U5058 ( .A1(n6179), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6180) );
  XNOR2_X2 U5060 ( .A(n5284), .B(P2_IR_REG_1__SCAN_IN), .ZN(n10655) );
  AOI21_X1 U5061 ( .B1(n9751), .B2(n9754), .A(n9753), .ZN(n9667) );
  NAND2_X2 U5062 ( .A1(n9356), .A2(n9355), .ZN(n9357) );
  AND2_X1 U5063 ( .A1(n5397), .A2(n5035), .ZN(n8879) );
  NAND2_X1 U5064 ( .A1(n6159), .A2(n6158), .ZN(n10790) );
  INV_X2 U5065 ( .A(n10846), .ZN(n4949) );
  NAND2_X1 U5066 ( .A1(n6998), .A2(n7006), .ZN(n7269) );
  NAND2_X2 U5067 ( .A1(n8341), .A2(n8528), .ZN(n8453) );
  CLKBUF_X2 U5069 ( .A(n7006), .Z(n8963) );
  NAND2_X1 U5070 ( .A1(n6991), .A2(n7028), .ZN(n6998) );
  NAND3_X1 U5071 ( .A1(n6995), .A2(n7028), .A3(n7574), .ZN(n7006) );
  INV_X1 U5072 ( .A(n7689), .ZN(n10756) );
  INV_X2 U5073 ( .A(n8916), .ZN(n8903) );
  INV_X1 U5074 ( .A(n7706), .ZN(n10743) );
  INV_X1 U5075 ( .A(n6292), .ZN(n6305) );
  NAND2_X1 U5076 ( .A1(n6679), .A2(n6704), .ZN(n6682) );
  NAND2_X1 U5077 ( .A1(n6245), .A2(n6249), .ZN(n8647) );
  XNOR2_X1 U5078 ( .A(n5578), .B(n10342), .ZN(n5583) );
  AND2_X1 U5079 ( .A1(n5404), .A2(n4988), .ZN(n9654) );
  NAND2_X1 U5080 ( .A1(n10062), .A2(n10063), .ZN(n10061) );
  NAND2_X1 U5081 ( .A1(n5126), .A2(n6651), .ZN(n9303) );
  AND2_X1 U5082 ( .A1(n8438), .A2(n8334), .ZN(n8499) );
  OR2_X1 U5083 ( .A1(n6734), .A2(n9979), .ZN(n8438) );
  AOI22_X1 U5084 ( .A1(n10344), .A2(n8333), .B1(n8332), .B2(
        P2_DATAO_REG_31__SCAN_IN), .ZN(n10302) );
  CLKBUF_X1 U5085 ( .A(n9692), .Z(n5069) );
  XNOR2_X1 U5086 ( .A(n8331), .B(n8330), .ZN(n10344) );
  NAND2_X1 U5087 ( .A1(n6720), .A2(n6719), .ZN(n6734) );
  OR2_X1 U5088 ( .A1(n9990), .A2(n8983), .ZN(n8564) );
  OR2_X1 U5089 ( .A1(n9483), .A2(n9295), .ZN(n6608) );
  XNOR2_X1 U5090 ( .A(n8282), .B(SI_29_), .ZN(n9619) );
  NOR2_X1 U5091 ( .A1(n9326), .A2(n5505), .ZN(n5504) );
  NAND2_X1 U5092 ( .A1(n6077), .A2(n6076), .ZN(n10214) );
  XNOR2_X1 U5093 ( .A(n5062), .B(n9158), .ZN(n8147) );
  NAND2_X1 U5094 ( .A1(n8103), .A2(n8102), .ZN(n8241) );
  OAI21_X1 U5095 ( .B1(n7780), .B2(n5410), .A(n5408), .ZN(n7961) );
  OR2_X1 U5096 ( .A1(n9519), .A2(n9407), .ZN(n8815) );
  NAND2_X1 U5097 ( .A1(n5076), .A2(n5238), .ZN(n5234) );
  AND2_X1 U5098 ( .A1(n6606), .A2(n6605), .ZN(n9305) );
  NAND2_X1 U5099 ( .A1(n6511), .A2(n6510), .ZN(n9523) );
  NOR2_X1 U5100 ( .A1(n7922), .A2(n5211), .ZN(n7923) );
  AND2_X2 U5101 ( .A1(n7665), .A2(n7664), .ZN(n4965) );
  AOI21_X1 U5102 ( .B1(n5237), .B2(n5238), .A(n5236), .ZN(n5235) );
  NAND2_X1 U5103 ( .A1(n5698), .A2(n5697), .ZN(n8188) );
  NAND2_X1 U5104 ( .A1(n5688), .A2(n5687), .ZN(n8213) );
  NAND2_X1 U5105 ( .A1(n5883), .A2(n5882), .ZN(n10810) );
  NAND2_X1 U5106 ( .A1(n5721), .A2(n5720), .ZN(n7969) );
  NAND2_X1 U5107 ( .A1(n6375), .A2(n6374), .ZN(n10769) );
  AND2_X1 U5108 ( .A1(n5214), .A2(n7350), .ZN(n7522) );
  NAND2_X2 U5109 ( .A1(n7573), .A2(n10729), .ZN(n10732) );
  NAND2_X1 U5110 ( .A1(n5847), .A2(n5846), .ZN(n8374) );
  NAND2_X1 U5111 ( .A1(n6359), .A2(n6358), .ZN(n8004) );
  CLKBUF_X3 U5112 ( .A(n7269), .Z(n8977) );
  NAND2_X2 U5113 ( .A1(n7192), .A2(n10838), .ZN(n10846) );
  NAND2_X1 U5114 ( .A1(n6345), .A2(n6344), .ZN(n8705) );
  NOR2_X1 U5115 ( .A1(n6459), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6460) );
  INV_X2 U5116 ( .A(n7071), .ZN(P1_U3973) );
  INV_X2 U5117 ( .A(n9151), .ZN(n6839) );
  INV_X2 U5118 ( .A(n5766), .ZN(n8333) );
  XNOR2_X1 U5119 ( .A(n6177), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U5120 ( .A1(n8864), .A2(n4946), .ZN(n6272) );
  NAND2_X1 U5121 ( .A1(n5261), .A2(n5262), .ZN(n7151) );
  AND2_X1 U5122 ( .A1(n5582), .A2(n10352), .ZN(n6100) );
  BUF_X2 U5123 ( .A(n5583), .Z(n8991) );
  OAI21_X1 U5124 ( .B1(n6176), .B2(n6175), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6177) );
  NAND2_X1 U5125 ( .A1(n6258), .A2(n6257), .ZN(n8864) );
  XNOR2_X1 U5126 ( .A(n6227), .B(n6226), .ZN(n8712) );
  INV_X1 U5127 ( .A(n9620), .ZN(n6245) );
  AND2_X2 U5128 ( .A1(n6239), .A2(n6240), .ZN(n9620) );
  NAND2_X1 U5129 ( .A1(n6146), .A2(n8304), .ZN(n5731) );
  OR2_X1 U5130 ( .A1(n6254), .A2(n6253), .ZN(n6258) );
  XNOR2_X1 U5131 ( .A(n6307), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7134) );
  MUX2_X1 U5132 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6237), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n6239) );
  XNOR2_X1 U5133 ( .A(n6338), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7231) );
  MUX2_X1 U5134 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6260), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n6262) );
  OR2_X1 U5135 ( .A1(n7110), .A2(n5264), .ZN(n5261) );
  NAND2_X1 U5136 ( .A1(n10349), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5578) );
  NOR2_X1 U5137 ( .A1(n5299), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n5300) );
  INV_X2 U5138 ( .A(n10343), .ZN(n10354) );
  NAND2_X1 U5139 ( .A1(n6240), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6241) );
  AND2_X1 U5140 ( .A1(n6306), .A2(n6297), .ZN(n6919) );
  XNOR2_X1 U5141 ( .A(n5581), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U5142 ( .A1(n6706), .A2(n6670), .ZN(n6709) );
  NAND2_X2 U5143 ( .A1(n6269), .A2(P2_U3151), .ZN(n9625) );
  AND2_X2 U5144 ( .A1(n6233), .A2(n6232), .ZN(n6706) );
  OR3_X1 U5145 ( .A1(n6320), .A2(P2_IR_REG_4__SCAN_IN), .A3(
        P2_IR_REG_3__SCAN_IN), .ZN(n6326) );
  AND2_X1 U5146 ( .A1(n5496), .A2(n6232), .ZN(n5493) );
  AND2_X1 U5147 ( .A1(n6236), .A2(n5031), .ZN(n5496) );
  AND2_X1 U5148 ( .A1(n6212), .A2(n5550), .ZN(n5079) );
  AND4_X1 U5149 ( .A1(n5084), .A2(n5083), .A3(n6924), .A4(n5082), .ZN(n5080)
         );
  AND2_X1 U5150 ( .A1(n5566), .A2(n5670), .ZN(n5416) );
  AND2_X1 U5151 ( .A1(n6210), .A2(n6211), .ZN(n6212) );
  AND2_X1 U5152 ( .A1(n6470), .A2(n6453), .ZN(n5083) );
  AND4_X1 U5153 ( .A1(n5088), .A2(n5086), .A3(n5087), .A4(n5085), .ZN(n6213)
         );
  AND2_X1 U5154 ( .A1(n6322), .A2(n6208), .ZN(n5084) );
  INV_X1 U5155 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6322) );
  INV_X1 U5156 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6208) );
  INV_X2 U5157 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U5158 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5082) );
  INV_X1 U5159 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6218) );
  INV_X1 U5160 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6226) );
  NOR2_X2 U5161 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5754) );
  NOR2_X1 U5162 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5563) );
  NOR2_X1 U5163 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5561) );
  INV_X1 U5164 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6453) );
  INV_X1 U5165 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6470) );
  NOR2_X1 U5166 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n6211) );
  NOR2_X1 U5167 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n6210) );
  INV_X2 U5168 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U5169 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5085) );
  NOR2_X1 U5170 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5086) );
  NOR2_X1 U5171 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5562) );
  NOR2_X1 U5172 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5087) );
  NOR2_X1 U5173 ( .A1(n10193), .A2(n10722), .ZN(n7705) );
  NAND2_X1 U5174 ( .A1(n4952), .A2(n9030), .ZN(n4951) );
  NAND2_X1 U5175 ( .A1(n9089), .A2(n9090), .ZN(n4952) );
  NAND2_X1 U5176 ( .A1(n9029), .A2(n9030), .ZN(n8614) );
  NAND2_X1 U5177 ( .A1(n9089), .A2(n9090), .ZN(n9029) );
  NAND2_X1 U5178 ( .A1(n8610), .A2(n8609), .ZN(n9089) );
  OR2_X2 U5179 ( .A1(n6759), .A2(n9570), .ZN(n6764) );
  NOR2_X2 U5180 ( .A1(n7940), .A2(n10680), .ZN(n7944) );
  NOR2_X1 U5181 ( .A1(n9234), .A2(n9246), .ZN(n10700) );
  NAND2_X1 U5182 ( .A1(n8949), .A2(n4956), .ZN(n4953) );
  AND2_X2 U5183 ( .A1(n4953), .A2(n4954), .ZN(n9763) );
  OR2_X1 U5184 ( .A1(n4955), .A2(n9684), .ZN(n4954) );
  INV_X1 U5185 ( .A(n8960), .ZN(n4955) );
  AND2_X1 U5186 ( .A1(n9713), .A2(n8960), .ZN(n4956) );
  INV_X1 U5187 ( .A(n5037), .ZN(n4957) );
  AND2_X1 U5188 ( .A1(n4958), .A2(n5685), .ZN(n6122) );
  NOR2_X1 U5189 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(n4957), .ZN(n4958) );
  NAND4_X4 U5190 ( .A1(n5776), .A2(n5775), .A3(n5774), .A4(n5773), .ZN(n9805)
         );
  AOI21_X2 U5191 ( .B1(n9998), .B2(n10162), .A(n5057), .ZN(n10210) );
  OAI21_X2 U5192 ( .B1(n5299), .B2(n5667), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5669) );
  NOR2_X2 U5193 ( .A1(n8043), .A2(n9649), .ZN(n8044) );
  AND2_X2 U5194 ( .A1(n8044), .A2(n10341), .ZN(n10171) );
  NOR2_X2 U5195 ( .A1(n10009), .A2(n9990), .ZN(n5302) );
  NAND2_X1 U5196 ( .A1(n5234), .A2(n5232), .ZN(n8119) );
  NAND2_X1 U5197 ( .A1(n7268), .A2(n7267), .ZN(n7400) );
  NAND2_X1 U5198 ( .A1(n9733), .A2(n9734), .ZN(n9732) );
  INV_X1 U5199 ( .A(n7412), .ZN(n7411) );
  AND2_X1 U5200 ( .A1(n5685), .A2(n5566), .ZN(n5671) );
  MUX2_X2 U5201 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10355), .S(n6815), .Z(n10722)
         );
  NAND2_X1 U5202 ( .A1(n6868), .A2(n6869), .ZN(n4959) );
  NAND2_X1 U5203 ( .A1(n8614), .A2(n4963), .ZN(n4960) );
  OR2_X1 U5204 ( .A1(n4962), .A2(n5006), .ZN(n4961) );
  INV_X1 U5205 ( .A(n8619), .ZN(n4962) );
  AND2_X1 U5206 ( .A1(n9031), .A2(n8619), .ZN(n4963) );
  NOR2_X1 U5207 ( .A1(n8622), .A2(n8623), .ZN(n4964) );
  NAND2_X1 U5208 ( .A1(n6868), .A2(n6869), .ZN(n6884) );
  NOR2_X1 U5209 ( .A1(n8622), .A2(n8623), .ZN(n9003) );
  NAND2_X2 U5210 ( .A1(n9946), .A2(n8576), .ZN(n8577) );
  NAND2_X1 U5211 ( .A1(n9667), .A2(n9668), .ZN(n9666) );
  OAI21_X2 U5212 ( .B1(n9641), .B2(n9642), .A(n9639), .ZN(n9777) );
  INV_X1 U5213 ( .A(n4965), .ZN(n7666) );
  NAND2_X1 U5214 ( .A1(n9077), .A2(n7207), .ZN(n7288) );
  MUX2_X1 U5215 ( .A(n8302), .B(n7292), .S(n7194), .Z(n6869) );
  NAND2_X2 U5216 ( .A1(n6865), .A2(n6864), .ZN(n6867) );
  NAND2_X1 U5217 ( .A1(n6867), .A2(n6866), .ZN(n4966) );
  NAND2_X1 U5218 ( .A1(n6867), .A2(n6866), .ZN(n4967) );
  OAI21_X2 U5219 ( .B1(n6682), .B2(P2_D_REG_0__SCAN_IN), .A(n6680), .ZN(n6681)
         );
  INV_X1 U5220 ( .A(n5521), .ZN(n5520) );
  OAI21_X1 U5221 ( .B1(n10065), .B2(n5522), .A(n6033), .ZN(n5521) );
  NAND2_X1 U5222 ( .A1(n9426), .A2(n6639), .ZN(n6641) );
  NAND2_X1 U5223 ( .A1(n5854), .A2(n5553), .ZN(n5626) );
  NAND2_X1 U5224 ( .A1(n6272), .A2(n6269), .ZN(n6319) );
  OR2_X1 U5225 ( .A1(n6712), .A2(n6625), .ZN(n8852) );
  NOR2_X1 U5226 ( .A1(n6655), .A2(n5384), .ZN(n5383) );
  INV_X1 U5227 ( .A(n6653), .ZN(n5384) );
  INV_X1 U5228 ( .A(n5385), .ZN(n5381) );
  NAND2_X1 U5229 ( .A1(n9483), .A2(n9295), .ZN(n6611) );
  NOR2_X1 U5230 ( .A1(n9308), .A2(n9317), .ZN(n8836) );
  OR2_X1 U5231 ( .A1(n9314), .A2(n6652), .ZN(n5126) );
  OR2_X1 U5232 ( .A1(n9366), .A2(n4982), .ZN(n9348) );
  OR2_X1 U5233 ( .A1(n9375), .A2(n9391), .ZN(n8702) );
  OR2_X1 U5234 ( .A1(n9388), .A2(n9386), .ZN(n9367) );
  OR2_X1 U5235 ( .A1(n9538), .A2(n9458), .ZN(n8795) );
  OR2_X1 U5236 ( .A1(n9545), .A2(n10576), .ZN(n8786) );
  NAND2_X1 U5237 ( .A1(n10769), .A2(n8013), .ZN(n8708) );
  INV_X1 U5238 ( .A(n4983), .ZN(n5111) );
  OR4_X1 U5239 ( .A1(n8477), .A2(n8476), .A3(n8475), .A4(n8474), .ZN(n8479) );
  NAND2_X1 U5240 ( .A1(n9963), .A2(n8439), .ZN(n8567) );
  NOR2_X1 U5241 ( .A1(n6064), .A2(n5175), .ZN(n5174) );
  INV_X1 U5242 ( .A(n5518), .ZN(n5175) );
  OR2_X1 U5243 ( .A1(n10214), .A2(n9634), .ZN(n8483) );
  OR2_X1 U5244 ( .A1(n10227), .A2(n9660), .ZN(n8484) );
  OR2_X1 U5245 ( .A1(n10220), .A2(n10224), .ZN(n8488) );
  NAND2_X1 U5246 ( .A1(n10787), .A2(n8386), .ZN(n6162) );
  XNOR2_X1 U5247 ( .A(n8280), .B(n8279), .ZN(n8282) );
  OAI21_X1 U5248 ( .B1(n5912), .B2(n5911), .A(n5658), .ZN(n5927) );
  INV_X1 U5249 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U5250 ( .A1(n5328), .A2(n5630), .ZN(n5327) );
  INV_X1 U5251 ( .A(n5878), .ZN(n5328) );
  XNOR2_X1 U5252 ( .A(n5628), .B(SI_10_), .ZN(n5713) );
  NOR2_X1 U5253 ( .A1(n5842), .A2(n5308), .ZN(n5307) );
  INV_X1 U5254 ( .A(n5614), .ZN(n5308) );
  NAND2_X1 U5255 ( .A1(n5355), .A2(n5354), .ZN(n6292) );
  NAND2_X1 U5256 ( .A1(n6258), .A2(n4994), .ZN(n5355) );
  AOI21_X1 U5257 ( .B1(n5432), .B2(n5431), .A(n8634), .ZN(n5430) );
  INV_X1 U5258 ( .A(n9121), .ZN(n5431) );
  INV_X1 U5259 ( .A(n8856), .ZN(n5193) );
  OAI21_X1 U5260 ( .B1(n5481), .B2(n5480), .A(n5485), .ZN(n5479) );
  NOR2_X1 U5261 ( .A1(n5486), .A2(n5484), .ZN(n5480) );
  NAND2_X1 U5262 ( .A1(n8692), .A2(n5000), .ZN(n5481) );
  NAND2_X1 U5263 ( .A1(n7110), .A2(n7111), .ZN(n7109) );
  XNOR2_X1 U5264 ( .A(n7225), .B(n7137), .ZN(n7136) );
  AOI22_X1 U5265 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(n4948), .B1(n7349), .B2(
        n6330), .ZN(n7228) );
  XNOR2_X1 U5266 ( .A(n7522), .B(n7537), .ZN(n7351) );
  INV_X1 U5267 ( .A(n7753), .ZN(n5276) );
  AND2_X1 U5268 ( .A1(n7938), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U5269 ( .A1(n5061), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5068) );
  INV_X1 U5270 ( .A(n10685), .ZN(n5061) );
  NAND2_X1 U5271 ( .A1(n5218), .A2(n5217), .ZN(n5216) );
  INV_X1 U5272 ( .A(n7924), .ZN(n5217) );
  OAI21_X1 U5273 ( .B1(n9314), .B2(n5016), .A(n5118), .ZN(n5117) );
  NAND2_X1 U5274 ( .A1(n5120), .A2(n5119), .ZN(n5118) );
  INV_X1 U5275 ( .A(n5123), .ZN(n5122) );
  NAND2_X1 U5276 ( .A1(n5502), .A2(n5501), .ZN(n5500) );
  AND2_X1 U5277 ( .A1(n5499), .A2(n8661), .ZN(n5498) );
  AOI21_X1 U5278 ( .B1(n9337), .B2(n6647), .A(n6646), .ZN(n9327) );
  AND2_X1 U5279 ( .A1(n8702), .A2(n9364), .ZN(n9349) );
  XNOR2_X1 U5280 ( .A(n9101), .B(n9373), .ZN(n9352) );
  NAND2_X1 U5281 ( .A1(n6638), .A2(n6637), .ZN(n9426) );
  AOI21_X1 U5282 ( .B1(n5350), .B2(n5352), .A(n5349), .ZN(n5348) );
  AND2_X1 U5283 ( .A1(n8791), .A2(n6450), .ZN(n9549) );
  NAND2_X1 U5284 ( .A1(n5473), .A2(n5471), .ZN(n8054) );
  AOI21_X1 U5285 ( .B1(n5021), .B2(n5474), .A(n5472), .ZN(n5471) );
  INV_X1 U5286 ( .A(n8762), .ZN(n5472) );
  INV_X1 U5287 ( .A(n6272), .ZN(n6484) );
  NOR2_X1 U5288 ( .A1(n8669), .A2(n5368), .ZN(n5367) );
  NOR2_X1 U5289 ( .A1(n7795), .A2(n4970), .ZN(n5368) );
  NAND2_X1 U5290 ( .A1(n6633), .A2(n6632), .ZN(n7796) );
  OR2_X1 U5291 ( .A1(n9146), .A2(n7293), .ZN(n6632) );
  OAI21_X1 U5292 ( .B1(n7383), .B2(n5106), .A(n5104), .ZN(n6633) );
  AOI21_X1 U5293 ( .B1(n5108), .B2(n5105), .A(n5012), .ZN(n5104) );
  NAND2_X1 U5294 ( .A1(n6597), .A2(n6596), .ZN(n8632) );
  NAND2_X1 U5296 ( .A1(n8991), .A2(n5584), .ZN(n5771) );
  OR2_X1 U5297 ( .A1(n5771), .A2(n6950), .ZN(n5724) );
  NAND2_X1 U5298 ( .A1(n10214), .A2(n9634), .ZN(n9995) );
  AOI21_X1 U5299 ( .B1(n5555), .B2(n5544), .A(n5011), .ZN(n5543) );
  AOI21_X1 U5300 ( .B1(n5170), .B2(n10115), .A(n5013), .ZN(n5169) );
  NAND2_X1 U5301 ( .A1(n5530), .A2(n5528), .ZN(n10116) );
  AOI21_X1 U5302 ( .B1(n5533), .B2(n5002), .A(n5529), .ZN(n5528) );
  NOR2_X1 U5303 ( .A1(n10331), .A2(n10279), .ZN(n5529) );
  AND2_X1 U5304 ( .A1(n5180), .A2(n5517), .ZN(n5179) );
  NAND2_X1 U5305 ( .A1(n10825), .A2(n10795), .ZN(n5517) );
  INV_X1 U5306 ( .A(n8290), .ZN(n8289) );
  XNOR2_X1 U5307 ( .A(n6089), .B(n6088), .ZN(n8228) );
  OAI21_X1 U5308 ( .B1(n6071), .B2(n6070), .A(n6069), .ZN(n6089) );
  INV_X1 U5309 ( .A(n6020), .ZN(n6019) );
  AND2_X1 U5310 ( .A1(n8605), .A2(n9427), .ZN(n8606) );
  AND2_X1 U5311 ( .A1(n5213), .A2(n5212), .ZN(n7922) );
  INV_X1 U5312 ( .A(n7737), .ZN(n5212) );
  NAND2_X1 U5313 ( .A1(n6668), .A2(n5375), .ZN(n8587) );
  INV_X1 U5314 ( .A(n8475), .ZN(n6721) );
  OAI22_X1 U5315 ( .A1(n6718), .A2(n6717), .B1(n5301), .B2(n10205), .ZN(n6722)
         );
  NAND2_X1 U5316 ( .A1(n5132), .A2(n5042), .ZN(n5249) );
  NAND2_X1 U5317 ( .A1(n5258), .A2(n8445), .ZN(n5257) );
  NAND2_X1 U5318 ( .A1(n5260), .A2(n8442), .ZN(n5259) );
  NAND2_X1 U5319 ( .A1(n8406), .A2(n8408), .ZN(n5258) );
  AND2_X1 U5320 ( .A1(n9403), .A2(n8809), .ZN(n5199) );
  NAND2_X1 U5321 ( .A1(n9421), .A2(n8806), .ZN(n5200) );
  AOI21_X1 U5322 ( .B1(n8799), .B2(n8798), .A(n8797), .ZN(n8804) );
  NAND2_X1 U5323 ( .A1(n5127), .A2(n10040), .ZN(n8431) );
  NAND2_X1 U5324 ( .A1(n5128), .A2(n5256), .ZN(n5127) );
  INV_X1 U5325 ( .A(n8423), .ZN(n5256) );
  AND2_X1 U5326 ( .A1(n9308), .A2(n9317), .ZN(n8837) );
  NOR2_X1 U5327 ( .A1(n7951), .A2(n5412), .ZN(n5411) );
  INV_X1 U5328 ( .A(n5414), .ZN(n5412) );
  INV_X1 U5329 ( .A(n5415), .ZN(n5409) );
  NAND2_X1 U5330 ( .A1(n5142), .A2(n5140), .ZN(n5139) );
  NOR2_X1 U5331 ( .A1(n5141), .A2(n8476), .ZN(n5140) );
  NAND2_X1 U5332 ( .A1(n5144), .A2(n5143), .ZN(n5142) );
  INV_X1 U5333 ( .A(n8434), .ZN(n5141) );
  INV_X1 U5334 ( .A(n6009), .ZN(n5522) );
  NOR2_X1 U5335 ( .A1(n10091), .A2(n10110), .ZN(n5288) );
  NOR2_X1 U5336 ( .A1(n5631), .A2(n5326), .ZN(n5325) );
  INV_X1 U5337 ( .A(n5713), .ZN(n5631) );
  INV_X1 U5338 ( .A(n5625), .ZN(n5326) );
  INV_X1 U5339 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5344) );
  INV_X1 U5340 ( .A(n7882), .ZN(n5421) );
  AND2_X1 U5341 ( .A1(n7513), .A2(n7510), .ZN(n5437) );
  INV_X1 U5342 ( .A(n8691), .ZN(n5485) );
  AND2_X1 U5343 ( .A1(n7938), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5275) );
  NOR2_X1 U5344 ( .A1(n9285), .A2(n8839), .ZN(n5489) );
  INV_X1 U5345 ( .A(n5383), .ZN(n5382) );
  INV_X1 U5346 ( .A(n5007), .ZN(n5377) );
  NOR2_X1 U5347 ( .A1(n6598), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6588) );
  NOR2_X1 U5348 ( .A1(n6654), .A2(n4976), .ZN(n5385) );
  OR2_X1 U5349 ( .A1(n9523), .A2(n9113), .ZN(n8810) );
  OR2_X1 U5350 ( .A1(n9530), .A2(n9406), .ZN(n8807) );
  NAND2_X1 U5351 ( .A1(n5458), .A2(n5461), .ZN(n5456) );
  AND2_X1 U5352 ( .A1(n9567), .A2(n8239), .ZN(n8774) );
  AOI21_X1 U5353 ( .B1(n5101), .B2(n5099), .A(n8060), .ZN(n5097) );
  AOI21_X1 U5354 ( .B1(n8009), .B2(n5099), .A(n9141), .ZN(n5098) );
  OR2_X1 U5355 ( .A1(n6360), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6380) );
  INV_X1 U5356 ( .A(n8746), .ZN(n5469) );
  AOI21_X1 U5357 ( .B1(n8665), .B2(n5470), .A(n5469), .ZN(n5468) );
  INV_X1 U5358 ( .A(n8745), .ZN(n5470) );
  NAND2_X1 U5359 ( .A1(n7284), .A2(n7096), .ZN(n8725) );
  NAND2_X1 U5360 ( .A1(n6839), .A2(n7359), .ZN(n8716) );
  OR2_X1 U5361 ( .A1(n6782), .A2(n8328), .ZN(n5094) );
  OAI22_X1 U5362 ( .A1(n5094), .A2(n4947), .B1(n5093), .B2(n5092), .ZN(n5091)
         );
  NAND2_X1 U5363 ( .A1(n4946), .A2(n6922), .ZN(n5092) );
  NAND2_X1 U5364 ( .A1(n5074), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6219) );
  NOR2_X1 U5365 ( .A1(n5078), .A2(n5077), .ZN(n9692) );
  NOR2_X1 U5366 ( .A1(n9777), .A2(n9774), .ZN(n5078) );
  AOI21_X1 U5367 ( .B1(n9777), .B2(n9774), .A(n9775), .ZN(n5077) );
  NAND2_X1 U5368 ( .A1(n6996), .A2(n6997), .ZN(n7002) );
  INV_X1 U5369 ( .A(n5583), .ZN(n5582) );
  OR2_X1 U5370 ( .A1(n10077), .A2(n9677), .ZN(n8421) );
  NAND2_X1 U5371 ( .A1(n10282), .A2(n10266), .ZN(n5539) );
  NOR2_X1 U5372 ( .A1(n10282), .A2(n10176), .ZN(n5298) );
  OR2_X1 U5373 ( .A1(n10176), .A2(n10278), .ZN(n8553) );
  OR2_X1 U5374 ( .A1(n9786), .A2(n9695), .ZN(n8518) );
  NOR2_X1 U5375 ( .A1(n4968), .A2(n9797), .ZN(n5176) );
  OR2_X1 U5376 ( .A1(n5294), .A2(n7969), .ZN(n5293) );
  NAND2_X1 U5377 ( .A1(n10785), .A2(n5295), .ZN(n5294) );
  OR2_X1 U5378 ( .A1(n7969), .A2(n10797), .ZN(n8540) );
  INV_X1 U5379 ( .A(n10193), .ZN(n5164) );
  NOR2_X1 U5380 ( .A1(n7704), .A2(n7276), .ZN(n7044) );
  NAND2_X1 U5381 ( .A1(n5329), .A2(n5333), .ZN(n6110) );
  AOI21_X1 U5382 ( .B1(n5337), .B2(n5335), .A(n5334), .ZN(n5333) );
  INV_X1 U5383 ( .A(n6094), .ZN(n5334) );
  BUF_X1 U5384 ( .A(n5664), .Z(n5299) );
  NAND2_X1 U5385 ( .A1(n6054), .A2(n6053), .ZN(n6071) );
  NAND2_X1 U5386 ( .A1(n6035), .A2(n6034), .ZN(n6052) );
  AND2_X1 U5387 ( .A1(n5928), .A2(n5661), .ZN(n5926) );
  AOI21_X1 U5388 ( .B1(n5314), .B2(n5885), .A(n5044), .ZN(n5313) );
  INV_X1 U5389 ( .A(n5322), .ZN(n5321) );
  OAI21_X1 U5390 ( .B1(n5641), .B2(n5323), .A(n5640), .ZN(n5322) );
  NAND2_X1 U5391 ( .A1(n5638), .A2(n5637), .ZN(n5878) );
  NAND2_X1 U5392 ( .A1(n5629), .A2(SI_10_), .ZN(n5630) );
  XNOR2_X1 U5393 ( .A(n5613), .B(SI_7_), .ZN(n5826) );
  INV_X1 U5394 ( .A(n5808), .ZN(n5608) );
  INV_X1 U5395 ( .A(n5591), .ZN(n6771) );
  NOR2_X1 U5396 ( .A1(n7973), .A2(n5421), .ZN(n5420) );
  INV_X1 U5397 ( .A(n5430), .ZN(n5427) );
  NAND2_X1 U5398 ( .A1(n9120), .A2(n9121), .ZN(n5433) );
  NAND2_X1 U5399 ( .A1(n5438), .A2(n9014), .ZN(n9077) );
  AND2_X1 U5400 ( .A1(n9078), .A2(n7205), .ZN(n5438) );
  NOR2_X1 U5401 ( .A1(n6512), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6522) );
  NAND2_X1 U5402 ( .A1(n4951), .A2(n9031), .ZN(n9034) );
  AOI21_X1 U5403 ( .B1(n8853), .B2(n8851), .A(n8689), .ZN(n5194) );
  NAND2_X1 U5404 ( .A1(n5485), .A2(n5483), .ZN(n5482) );
  NOR2_X1 U5405 ( .A1(n5488), .A2(n5484), .ZN(n5483) );
  NOR2_X1 U5406 ( .A1(n8655), .A2(n8654), .ZN(n8856) );
  NOR2_X1 U5407 ( .A1(n6238), .A2(n6256), .ZN(n6257) );
  NOR2_X1 U5408 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6256) );
  INV_X1 U5409 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6253) );
  AND3_X1 U5410 ( .A1(n6494), .A2(n6493), .A3(n6492), .ZN(n9060) );
  NAND2_X1 U5411 ( .A1(n5025), .A2(n7109), .ZN(n5265) );
  INV_X1 U5412 ( .A(n5263), .ZN(n5262) );
  OAI21_X1 U5413 ( .B1(n7156), .B2(n7158), .A(n7157), .ZN(n7160) );
  OR2_X1 U5414 ( .A1(n7226), .A2(n7228), .ZN(n5273) );
  NAND2_X1 U5415 ( .A1(n7136), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7227) );
  NOR2_X1 U5416 ( .A1(n5073), .A2(n8002), .ZN(n5072) );
  NAND2_X1 U5417 ( .A1(n5216), .A2(n5215), .ZN(n5062) );
  NAND2_X1 U5418 ( .A1(n8154), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5215) );
  XNOR2_X1 U5419 ( .A(n9212), .B(n9213), .ZN(n9192) );
  NOR2_X1 U5420 ( .A1(n9224), .A2(n5551), .ZN(n9245) );
  NOR2_X1 U5421 ( .A1(n9246), .A2(n9245), .ZN(n9248) );
  AOI21_X1 U5422 ( .B1(n5489), .B2(n8840), .A(n5487), .ZN(n5486) );
  INV_X1 U5423 ( .A(n6611), .ZN(n5487) );
  INV_X1 U5424 ( .A(n5489), .ZN(n5488) );
  AND2_X1 U5425 ( .A1(n8852), .A2(n8688), .ZN(n8686) );
  AND4_X1 U5426 ( .A1(n6594), .A2(n6593), .A3(n6592), .A4(n6591), .ZN(n9295)
         );
  INV_X1 U5427 ( .A(n9137), .ZN(n9317) );
  NAND2_X1 U5428 ( .A1(n6650), .A2(n6649), .ZN(n9314) );
  AOI21_X1 U5429 ( .B1(n5504), .B2(n8828), .A(n5024), .ZN(n5502) );
  OR2_X1 U5430 ( .A1(n8832), .A2(n8831), .ZN(n9321) );
  INV_X1 U5431 ( .A(n9341), .ZN(n5508) );
  OR2_X1 U5432 ( .A1(n9355), .A2(n9349), .ZN(n6645) );
  NAND2_X1 U5433 ( .A1(n6641), .A2(n5374), .ZN(n5373) );
  AND2_X1 U5434 ( .A1(n4992), .A2(n6640), .ZN(n5374) );
  INV_X1 U5435 ( .A(n9352), .ZN(n9355) );
  OR2_X1 U5436 ( .A1(n4982), .A2(n6644), .ZN(n9364) );
  AND2_X1 U5437 ( .A1(n9368), .A2(n9367), .ZN(n9389) );
  AOI21_X1 U5438 ( .B1(n9421), .B2(n5449), .A(n5448), .ZN(n5447) );
  INV_X1 U5439 ( .A(n6495), .ZN(n5449) );
  INV_X1 U5440 ( .A(n8807), .ZN(n5448) );
  INV_X1 U5441 ( .A(n9421), .ZN(n5450) );
  NAND2_X1 U5442 ( .A1(n6641), .A2(n6640), .ZN(n9347) );
  AOI21_X1 U5443 ( .B1(n6481), .B2(n9455), .A(n5453), .ZN(n5452) );
  INV_X1 U5444 ( .A(n8795), .ZN(n5453) );
  NAND2_X1 U5445 ( .A1(n9435), .A2(n9434), .ZN(n9433) );
  NAND2_X1 U5446 ( .A1(n5454), .A2(n5352), .ZN(n9445) );
  INV_X1 U5447 ( .A(n9454), .ZN(n5454) );
  AOI21_X1 U5448 ( .B1(n9455), .B2(n5351), .A(n5043), .ZN(n5350) );
  INV_X1 U5449 ( .A(n8791), .ZN(n5351) );
  OAI21_X1 U5450 ( .B1(n6636), .B2(n8239), .A(n6635), .ZN(n9550) );
  OAI21_X1 U5451 ( .B1(n9467), .B2(n9554), .A(n9567), .ZN(n6635) );
  NAND2_X1 U5452 ( .A1(n6416), .A2(n10545), .ZN(n6434) );
  INV_X1 U5453 ( .A(n6417), .ZN(n6416) );
  OR2_X1 U5454 ( .A1(n5459), .A2(n8774), .ZN(n9466) );
  NAND2_X1 U5455 ( .A1(n6415), .A2(n6414), .ZN(n8768) );
  NAND2_X1 U5456 ( .A1(n6409), .A2(n8763), .ZN(n8132) );
  AND2_X1 U5457 ( .A1(n8765), .A2(n8763), .ZN(n8675) );
  INV_X1 U5458 ( .A(n5477), .ZN(n5476) );
  AOI21_X1 U5459 ( .B1(n5477), .B2(n5475), .A(n8703), .ZN(n5474) );
  INV_X1 U5460 ( .A(n8756), .ZN(n5475) );
  AOI21_X1 U5461 ( .B1(n4974), .B2(n5365), .A(n5017), .ZN(n5361) );
  AOI21_X1 U5462 ( .B1(n5367), .B2(n4970), .A(n5019), .ZN(n5366) );
  AND2_X1 U5463 ( .A1(n7988), .A2(n8707), .ZN(n5477) );
  AND2_X1 U5464 ( .A1(n8756), .A2(n8707), .ZN(n8669) );
  AND2_X1 U5465 ( .A1(n7770), .A2(n8751), .ZN(n7794) );
  OR2_X1 U5466 ( .A1(n6331), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6349) );
  INV_X1 U5467 ( .A(n9145), .ZN(n8704) );
  NOR2_X1 U5468 ( .A1(n5111), .A2(n5369), .ZN(n5109) );
  NAND2_X1 U5469 ( .A1(n5110), .A2(n5113), .ZN(n5108) );
  NAND2_X1 U5470 ( .A1(n7550), .A2(n7775), .ZN(n5370) );
  INV_X1 U5471 ( .A(n9147), .ZN(n7775) );
  NAND2_X1 U5472 ( .A1(n7097), .A2(n6629), .ZN(n7282) );
  INV_X1 U5473 ( .A(n9553), .ZN(n9471) );
  NAND2_X1 U5474 ( .A1(n8658), .A2(n8657), .ZN(n9278) );
  NAND2_X1 U5475 ( .A1(n6620), .A2(n6619), .ZN(n6712) );
  NAND2_X1 U5476 ( .A1(n6541), .A2(n6540), .ZN(n9101) );
  NAND2_X1 U5477 ( .A1(n9763), .A2(n5059), .ZN(n9629) );
  AND2_X1 U5478 ( .A1(n9630), .A2(n9631), .ZN(n5059) );
  INV_X1 U5479 ( .A(n10004), .ZN(n8983) );
  OR2_X1 U5480 ( .A1(n8919), .A2(n8918), .ZN(n8920) );
  NAND2_X1 U5481 ( .A1(n5069), .A2(n9693), .ZN(n9691) );
  XNOR2_X1 U5482 ( .A(n7272), .B(n8975), .ZN(n7395) );
  NAND2_X1 U5483 ( .A1(n7271), .A2(n7270), .ZN(n7272) );
  NAND2_X1 U5484 ( .A1(n7779), .A2(n7778), .ZN(n5414) );
  OR2_X1 U5485 ( .A1(n7779), .A2(n7778), .ZN(n5415) );
  NAND2_X1 U5486 ( .A1(n7254), .A2(n10194), .ZN(n7001) );
  INV_X1 U5487 ( .A(n9794), .ZN(n9782) );
  OAI21_X1 U5488 ( .B1(n8446), .B2(n8573), .A(n5149), .ZN(n8447) );
  AOI21_X1 U5489 ( .B1(n8573), .B2(n8442), .A(n8519), .ZN(n5149) );
  MUX2_X1 U5490 ( .A(n8508), .B(n8482), .S(n8442), .Z(n8443) );
  NAND2_X1 U5491 ( .A1(n5341), .A2(n5049), .ZN(n8571) );
  NOR2_X1 U5492 ( .A1(n10302), .A2(n9790), .ZN(n8573) );
  INV_X1 U5493 ( .A(n5771), .ZN(n8292) );
  NAND2_X1 U5494 ( .A1(n6100), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U5495 ( .A1(n8990), .A2(n8333), .ZN(n5341) );
  NOR2_X1 U5496 ( .A1(n6735), .A2(n6734), .ZN(n8290) );
  AND2_X1 U5497 ( .A1(n5174), .A2(n5544), .ZN(n5173) );
  NAND2_X1 U5498 ( .A1(n5542), .A2(n5540), .ZN(n9987) );
  AND2_X1 U5499 ( .A1(n5543), .A2(n5541), .ZN(n5540) );
  INV_X1 U5500 ( .A(n9996), .ZN(n5541) );
  INV_X1 U5501 ( .A(n10007), .ZN(n5544) );
  OR2_X1 U5502 ( .A1(n6066), .A2(n5555), .ZN(n5545) );
  AND2_X1 U5503 ( .A1(n5519), .A2(n5174), .ZN(n6066) );
  AND2_X1 U5504 ( .A1(n8483), .A2(n9995), .ZN(n10007) );
  INV_X1 U5505 ( .A(n8488), .ZN(n5075) );
  NOR2_X1 U5506 ( .A1(n10220), .A2(n10033), .ZN(n10022) );
  NAND2_X1 U5507 ( .A1(n10053), .A2(n8487), .ZN(n10039) );
  OR2_X1 U5508 ( .A1(n10227), .A2(n10046), .ZN(n10033) );
  AND2_X1 U5509 ( .A1(n8424), .A2(n8487), .ZN(n10054) );
  NAND2_X1 U5510 ( .A1(n10066), .A2(n10065), .ZN(n10064) );
  NAND2_X1 U5511 ( .A1(n5168), .A2(n5166), .ZN(n10080) );
  AOI21_X1 U5512 ( .B1(n5169), .B2(n5171), .A(n5167), .ZN(n5166) );
  OR2_X1 U5513 ( .A1(n10282), .A2(n10137), .ZN(n10128) );
  NAND2_X1 U5514 ( .A1(n4971), .A2(n5539), .ZN(n5535) );
  NAND2_X1 U5515 ( .A1(n5534), .A2(n5539), .ZN(n5533) );
  INV_X1 U5516 ( .A(n5536), .ZN(n5534) );
  NOR2_X1 U5517 ( .A1(n10147), .A2(n5537), .ZN(n5536) );
  NOR2_X1 U5518 ( .A1(n5538), .A2(n6165), .ZN(n5537) );
  AND2_X1 U5519 ( .A1(n10128), .A2(n8407), .ZN(n10147) );
  NAND2_X1 U5520 ( .A1(n8113), .A2(n5552), .ZN(n10170) );
  NAND2_X1 U5521 ( .A1(n8114), .A2(n8467), .ZN(n8113) );
  OR2_X1 U5522 ( .A1(n7899), .A2(n8213), .ZN(n8043) );
  AND2_X1 U5523 ( .A1(n8545), .A2(n8393), .ZN(n8464) );
  NAND2_X1 U5524 ( .A1(n7556), .A2(n4969), .ZN(n5884) );
  NAND2_X1 U5525 ( .A1(n10790), .A2(n6161), .ZN(n10787) );
  NAND2_X1 U5526 ( .A1(n6162), .A2(n8463), .ZN(n7893) );
  NAND2_X1 U5527 ( .A1(n8374), .A2(n8373), .ZN(n8369) );
  NAND2_X1 U5528 ( .A1(n6153), .A2(n8369), .ZN(n8359) );
  NAND2_X1 U5529 ( .A1(n7323), .A2(n8358), .ZN(n7322) );
  AND2_X1 U5530 ( .A1(n7044), .A2(n5290), .ZN(n7687) );
  NAND2_X1 U5531 ( .A1(n5290), .A2(n7415), .ZN(n5790) );
  OAI21_X1 U5532 ( .B1(n7051), .B2(n5163), .A(n5161), .ZN(n7683) );
  INV_X1 U5533 ( .A(n5162), .ZN(n5161) );
  OAI21_X1 U5534 ( .B1(n8454), .B2(n5163), .A(n8455), .ZN(n5162) );
  INV_X1 U5535 ( .A(n5790), .ZN(n5163) );
  NAND2_X1 U5536 ( .A1(n7051), .A2(n8454), .ZN(n7050) );
  NAND2_X1 U5537 ( .A1(n8438), .A2(n8503), .ZN(n8475) );
  INV_X1 U5538 ( .A(n10796), .ZN(n10267) );
  OAI21_X1 U5539 ( .B1(n8282), .B2(n10487), .A(n8281), .ZN(n8327) );
  NAND2_X1 U5540 ( .A1(n5671), .A2(n5575), .ZN(n5664) );
  NAND2_X1 U5541 ( .A1(n5156), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5581) );
  AND2_X1 U5542 ( .A1(n5038), .A2(n5575), .ZN(n5155) );
  AND2_X1 U5543 ( .A1(n5575), .A2(n5580), .ZN(n5241) );
  XNOR2_X1 U5544 ( .A(n6071), .B(n6067), .ZN(n8051) );
  XNOR2_X1 U5545 ( .A(n6052), .B(n6051), .ZN(n8033) );
  NAND2_X1 U5546 ( .A1(n6012), .A2(n6011), .ZN(n5310) );
  NAND2_X1 U5547 ( .A1(n5982), .A2(n5981), .ZN(n5995) );
  NAND2_X1 U5548 ( .A1(n5312), .A2(n5650), .ZN(n5900) );
  OR2_X1 U5549 ( .A1(n5886), .A2(n5885), .ZN(n5312) );
  NAND2_X1 U5550 ( .A1(n5626), .A2(n5625), .ZN(n5714) );
  NAND2_X1 U5552 ( .A1(n6444), .A2(n6443), .ZN(n8780) );
  NAND2_X1 U5553 ( .A1(n6550), .A2(n6549), .ZN(n9503) );
  NAND2_X1 U5554 ( .A1(n6586), .A2(n6585), .ZN(n9483) );
  INV_X1 U5555 ( .A(n9338), .ZN(n9373) );
  INV_X1 U5556 ( .A(n5441), .ZN(n5440) );
  OAI22_X1 U5557 ( .A1(n5442), .A2(n5444), .B1(n9428), .B2(n9051), .ZN(n5441)
         );
  OR2_X1 U5558 ( .A1(n8599), .A2(n5443), .ZN(n5442) );
  AND2_X1 U5559 ( .A1(n6558), .A2(n6557), .ZN(n9330) );
  AND2_X1 U5560 ( .A1(n7883), .A2(n7882), .ZN(n7974) );
  INV_X1 U5561 ( .A(n9330), .ZN(n9353) );
  AND2_X1 U5562 ( .A1(n6342), .A2(n6355), .ZN(n7537) );
  OR2_X1 U5563 ( .A1(n7734), .A2(n7735), .ZN(n5213) );
  INV_X1 U5564 ( .A(n5277), .ZN(n7754) );
  NAND2_X1 U5565 ( .A1(n5068), .A2(n4984), .ZN(n5218) );
  INV_X1 U5566 ( .A(n5216), .ZN(n8146) );
  NOR2_X1 U5567 ( .A1(n8147), .A2(n6431), .ZN(n9153) );
  XNOR2_X1 U5568 ( .A(n9199), .B(n9213), .ZN(n9181) );
  XNOR2_X1 U5569 ( .A(n9245), .B(n9246), .ZN(n9225) );
  NOR2_X1 U5570 ( .A1(n9225), .A2(n9226), .ZN(n9247) );
  NAND2_X1 U5571 ( .A1(n5490), .A2(n8660), .ZN(n9286) );
  OR2_X1 U5572 ( .A1(n9297), .A2(n8840), .ZN(n5490) );
  AND2_X1 U5573 ( .A1(n5067), .A2(n5066), .ZN(n9486) );
  AOI22_X1 U5574 ( .A1(n9283), .A2(n9553), .B1(n9282), .B2(n9552), .ZN(n5066)
         );
  NAND2_X1 U5575 ( .A1(n9284), .A2(n9547), .ZN(n5067) );
  AOI22_X1 U5576 ( .A1(n10344), .A2(n8656), .B1(n8643), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n9573) );
  INV_X1 U5577 ( .A(n6712), .ZN(n8589) );
  NOR2_X1 U5578 ( .A1(n8587), .A2(n6669), .ZN(n6759) );
  CLKBUF_X1 U5579 ( .A(n7780), .Z(n7727) );
  OR2_X1 U5580 ( .A1(n8911), .A2(n8910), .ZN(n8912) );
  NAND2_X1 U5581 ( .A1(n8228), .A2(n8333), .ZN(n6077) );
  NAND2_X1 U5582 ( .A1(n5889), .A2(n5888), .ZN(n9649) );
  AND2_X1 U5583 ( .A1(n10732), .A2(n7575), .ZN(n10189) );
  NAND2_X1 U5584 ( .A1(n7024), .A2(n7023), .ZN(n10729) );
  NOR2_X1 U5585 ( .A1(n5230), .A2(n6732), .ZN(n5158) );
  INV_X1 U5586 ( .A(n9969), .ZN(n5230) );
  NOR2_X1 U5587 ( .A1(n6747), .A2(n10340), .ZN(n6737) );
  NAND2_X1 U5588 ( .A1(n8993), .A2(n8333), .ZN(n6112) );
  INV_X1 U5589 ( .A(n8359), .ZN(n8363) );
  OAI21_X1 U5590 ( .B1(n5255), .B2(n5253), .A(n5022), .ZN(n5252) );
  AND2_X1 U5591 ( .A1(n8386), .A2(n8445), .ZN(n5254) );
  OAI21_X1 U5592 ( .B1(n8357), .B2(n8445), .A(n5153), .ZN(n5152) );
  NOR2_X1 U5593 ( .A1(n8358), .A2(n5154), .ZN(n5153) );
  NOR2_X1 U5594 ( .A1(n8457), .A2(n8442), .ZN(n5154) );
  NAND2_X1 U5595 ( .A1(n8760), .A2(n5196), .ZN(n8711) );
  AOI21_X1 U5596 ( .B1(n5198), .B2(n8842), .A(n5197), .ZN(n5196) );
  NAND2_X1 U5597 ( .A1(n8708), .A2(n8707), .ZN(n5198) );
  NOR2_X1 U5598 ( .A1(n8756), .A2(n8842), .ZN(n5197) );
  NAND2_X1 U5599 ( .A1(n5251), .A2(n5150), .ZN(n8384) );
  NAND2_X1 U5600 ( .A1(n5152), .A2(n5151), .ZN(n5150) );
  AOI21_X1 U5601 ( .B1(n5254), .B2(n8371), .A(n5252), .ZN(n5251) );
  NOR2_X1 U5602 ( .A1(n8364), .A2(n5253), .ZN(n5151) );
  AND2_X1 U5603 ( .A1(n8391), .A2(n8545), .ZN(n5250) );
  AND2_X1 U5604 ( .A1(n8765), .A2(n8842), .ZN(n5190) );
  NAND2_X1 U5605 ( .A1(n5189), .A2(n5187), .ZN(n8773) );
  AND2_X1 U5606 ( .A1(n5188), .A2(n8767), .ZN(n5187) );
  NAND2_X1 U5607 ( .A1(n5191), .A2(n5190), .ZN(n5189) );
  OR2_X1 U5608 ( .A1(n8766), .A2(n8842), .ZN(n5188) );
  NAND2_X1 U5609 ( .A1(n5249), .A2(n4991), .ZN(n8403) );
  NAND2_X1 U5610 ( .A1(n8420), .A2(n8445), .ZN(n5129) );
  AOI21_X1 U5611 ( .B1(n8416), .B2(n8559), .A(n8412), .ZN(n8414) );
  NAND2_X1 U5612 ( .A1(n8419), .A2(n8442), .ZN(n5131) );
  NOR2_X1 U5613 ( .A1(n10051), .A2(n4990), .ZN(n5130) );
  OAI21_X1 U5614 ( .B1(n8804), .B2(n5200), .A(n5199), .ZN(n8813) );
  NOR2_X1 U5615 ( .A1(n8436), .A2(n5145), .ZN(n5144) );
  AND2_X1 U5616 ( .A1(n8429), .A2(n8445), .ZN(n5145) );
  NAND2_X1 U5617 ( .A1(n8428), .A2(n8442), .ZN(n5143) );
  OAI21_X1 U5618 ( .B1(n8431), .B2(n8425), .A(n5010), .ZN(n8426) );
  OAI21_X1 U5619 ( .B1(n8830), .B2(n8829), .A(n9333), .ZN(n5186) );
  INV_X1 U5620 ( .A(n8838), .ZN(n5184) );
  NAND2_X1 U5621 ( .A1(n6859), .A2(n9151), .ZN(n8717) );
  NAND2_X1 U5622 ( .A1(n6706), .A2(n6236), .ZN(n6259) );
  NOR2_X1 U5623 ( .A1(n6326), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n6371) );
  AND2_X1 U5624 ( .A1(n5972), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5985) );
  NOR2_X1 U5625 ( .A1(n5834), .A2(n5833), .ZN(n5832) );
  AND3_X1 U5626 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5798) );
  NOR2_X1 U5627 ( .A1(n5336), .A2(n5331), .ZN(n5330) );
  INV_X1 U5628 ( .A(n6053), .ZN(n5331) );
  INV_X1 U5629 ( .A(n5337), .ZN(n5336) );
  INV_X1 U5630 ( .A(n5339), .ZN(n5335) );
  NAND2_X1 U5631 ( .A1(n6052), .A2(n6051), .ZN(n6054) );
  NOR2_X1 U5632 ( .A1(n5653), .A2(n5315), .ZN(n5314) );
  INV_X1 U5633 ( .A(n5650), .ZN(n5315) );
  NAND2_X1 U5634 ( .A1(n5327), .A2(n5638), .ZN(n5323) );
  NOR2_X1 U5635 ( .A1(n5324), .A2(n5318), .ZN(n5317) );
  INV_X1 U5636 ( .A(n5325), .ZN(n5318) );
  NAND2_X1 U5637 ( .A1(n5689), .A2(n5638), .ZN(n5324) );
  NAND2_X1 U5638 ( .A1(n5616), .A2(n10374), .ZN(n5619) );
  OAI21_X1 U5639 ( .B1(n5185), .B2(n5183), .A(n5182), .ZN(n8845) );
  NAND2_X1 U5640 ( .A1(n9296), .A2(n5184), .ZN(n5183) );
  INV_X1 U5641 ( .A(n8841), .ZN(n5182) );
  AOI211_X1 U5642 ( .C1(n5186), .C2(n8835), .A(n8833), .B(n8834), .ZN(n5185)
         );
  INV_X1 U5643 ( .A(n8852), .ZN(n5484) );
  INV_X1 U5644 ( .A(n6282), .ZN(n6293) );
  NAND2_X1 U5645 ( .A1(n7122), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5205) );
  INV_X1 U5646 ( .A(n6928), .ZN(n5264) );
  OAI21_X1 U5647 ( .B1(n5264), .B2(n7111), .A(n7126), .ZN(n5263) );
  NAND2_X1 U5648 ( .A1(n5204), .A2(n7126), .ZN(n5201) );
  NOR2_X1 U5649 ( .A1(n8153), .A2(n5071), .ZN(n9166) );
  NOR2_X1 U5650 ( .A1(n7941), .A2(n8134), .ZN(n5071) );
  XNOR2_X1 U5651 ( .A(n9166), .B(n9167), .ZN(n8155) );
  INV_X1 U5652 ( .A(n5268), .ZN(n5272) );
  INV_X1 U5653 ( .A(n10700), .ZN(n5270) );
  AOI21_X1 U5654 ( .B1(n5124), .B2(n6652), .A(n4976), .ZN(n5123) );
  NAND2_X1 U5655 ( .A1(n9293), .A2(n5123), .ZN(n5119) );
  NAND2_X1 U5656 ( .A1(n9296), .A2(n5121), .ZN(n5120) );
  NAND2_X1 U5657 ( .A1(n5123), .A2(n5125), .ZN(n5121) );
  OR2_X1 U5658 ( .A1(n6578), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6598) );
  INV_X1 U5659 ( .A(n8832), .ZN(n5501) );
  OR2_X1 U5660 ( .A1(n8836), .A2(n8837), .ZN(n8833) );
  OR2_X1 U5661 ( .A1(n9385), .A2(n9388), .ZN(n9366) );
  NOR2_X1 U5662 ( .A1(n8774), .A2(n5463), .ZN(n5462) );
  NAND2_X1 U5663 ( .A1(n5366), .A2(n5364), .ZN(n5363) );
  INV_X1 U5664 ( .A(n5367), .ZN(n5364) );
  INV_X1 U5665 ( .A(n5366), .ZN(n5365) );
  NAND2_X1 U5666 ( .A1(n6348), .A2(n6347), .ZN(n6360) );
  INV_X1 U5667 ( .A(n5109), .ZN(n5105) );
  INV_X1 U5668 ( .A(n5108), .ZN(n5106) );
  INV_X1 U5669 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10456) );
  INV_X1 U5670 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6209) );
  INV_X1 U5671 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6410) );
  OR2_X1 U5672 ( .A1(n6371), .A2(n9613), .ZN(n6338) );
  NAND2_X1 U5673 ( .A1(n6209), .A2(n6208), .ZN(n6282) );
  AOI21_X1 U5674 ( .B1(n5411), .B2(n5409), .A(n4995), .ZN(n5408) );
  INV_X1 U5675 ( .A(n5411), .ZN(n5410) );
  NOR2_X1 U5676 ( .A1(n5871), .A2(n5870), .ZN(n5700) );
  AND2_X1 U5677 ( .A1(n5890), .A2(n5556), .ZN(n5557) );
  AOI21_X1 U5678 ( .B1(n5138), .B2(n8441), .A(n5137), .ZN(n8444) );
  OR2_X1 U5679 ( .A1(n8508), .A2(n8482), .ZN(n5137) );
  NAND2_X1 U5680 ( .A1(n5139), .A2(n5003), .ZN(n5138) );
  OR2_X1 U5681 ( .A1(n9983), .A2(n10205), .ZN(n8334) );
  AOI21_X1 U5682 ( .B1(n5520), .B2(n5522), .A(n5015), .ZN(n5518) );
  AND2_X1 U5683 ( .A1(n5533), .A2(n4985), .ZN(n5531) );
  NAND2_X1 U5684 ( .A1(n5557), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5935) );
  OR2_X1 U5685 ( .A1(n5702), .A2(n5676), .ZN(n5892) );
  OR2_X1 U5686 ( .A1(n5860), .A2(n5859), .ZN(n5862) );
  INV_X1 U5687 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U5688 ( .A1(n5798), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U5689 ( .A1(n8523), .A2(n8452), .ZN(n8339) );
  NAND2_X1 U5690 ( .A1(n5302), .A2(n5301), .ZN(n6735) );
  NAND2_X1 U5691 ( .A1(n10120), .A2(n5288), .ZN(n10089) );
  NAND2_X1 U5692 ( .A1(n10120), .A2(n10323), .ZN(n10107) );
  NAND2_X1 U5693 ( .A1(n10171), .A2(n5296), .ZN(n10140) );
  NOR2_X1 U5694 ( .A1(n10143), .A2(n5297), .ZN(n5296) );
  INV_X1 U5695 ( .A(n5298), .ZN(n5297) );
  NOR2_X1 U5696 ( .A1(n7501), .A2(n7807), .ZN(n7560) );
  NAND2_X1 U5697 ( .A1(n6617), .A2(n6616), .ZN(n8280) );
  NAND2_X1 U5698 ( .A1(n6613), .A2(n6612), .ZN(n6617) );
  NAND2_X1 U5699 ( .A1(n6110), .A2(n6109), .ZN(n6613) );
  AOI21_X1 U5700 ( .B1(n5339), .B2(n6070), .A(n5338), .ZN(n5337) );
  INV_X1 U5701 ( .A(n6087), .ZN(n5338) );
  NOR2_X1 U5702 ( .A1(n6088), .A2(n5340), .ZN(n5339) );
  INV_X1 U5703 ( .A(n6069), .ZN(n5340) );
  INV_X1 U5704 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6195) );
  OR2_X1 U5705 ( .A1(n5855), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U5706 ( .A1(n5622), .A2(n5621), .ZN(n5625) );
  NAND2_X1 U5707 ( .A1(n5827), .A2(n5612), .ZN(n5309) );
  XNOR2_X1 U5708 ( .A(n5609), .B(SI_6_), .ZN(n5808) );
  INV_X1 U5709 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5560) );
  INV_X1 U5710 ( .A(SI_3_), .ZN(n10411) );
  INV_X1 U5711 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5346) );
  AND2_X1 U5712 ( .A1(n5436), .A2(n7606), .ZN(n5435) );
  OR2_X1 U5713 ( .A1(n5437), .A2(n5052), .ZN(n5436) );
  NOR2_X1 U5714 ( .A1(n6475), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6490) );
  INV_X1 U5715 ( .A(n8597), .ZN(n5443) );
  NAND2_X1 U5716 ( .A1(n9003), .A2(n9330), .ZN(n9070) );
  AND2_X1 U5717 ( .A1(n9030), .A2(n8613), .ZN(n9090) );
  OR2_X1 U5718 ( .A1(n6502), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6512) );
  AND2_X1 U5719 ( .A1(n8271), .A2(n8269), .ZN(n5444) );
  OR2_X1 U5720 ( .A1(n6436), .A2(n6275), .ZN(n6279) );
  OAI21_X1 U5721 ( .B1(n6244), .B2(n8647), .A(n6243), .ZN(n6248) );
  NOR2_X1 U5722 ( .A1(n6920), .A2(n6287), .ZN(n7156) );
  INV_X1 U5723 ( .A(n5201), .ZN(n7158) );
  NOR2_X1 U5724 ( .A1(n7220), .A2(n5548), .ZN(n7222) );
  OR2_X1 U5725 ( .A1(n7750), .A2(n7751), .ZN(n5277) );
  OAI21_X1 U5726 ( .B1(n8155), .B2(n5279), .A(n5278), .ZN(n9190) );
  NAND2_X1 U5727 ( .A1(n5280), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5279) );
  NAND2_X1 U5728 ( .A1(n9169), .A2(n5280), .ZN(n5278) );
  INV_X1 U5729 ( .A(n9172), .ZN(n5280) );
  NOR2_X1 U5730 ( .A1(n8155), .A2(n6430), .ZN(n9168) );
  NAND2_X1 U5731 ( .A1(n5283), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U5732 ( .A1(n9215), .A2(n5283), .ZN(n5281) );
  INV_X1 U5733 ( .A(n9217), .ZN(n5283) );
  NOR2_X1 U5734 ( .A1(n9192), .A2(n9461), .ZN(n9214) );
  OR2_X1 U5735 ( .A1(n10700), .A2(n5272), .ZN(n9235) );
  NOR2_X1 U5736 ( .A1(n5272), .A2(n5269), .ZN(n10699) );
  NAND2_X1 U5737 ( .A1(n5270), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5269) );
  OAI21_X1 U5738 ( .B1(n9303), .B2(n5023), .A(n5379), .ZN(n6656) );
  AOI21_X1 U5739 ( .B1(n5383), .B2(n5381), .A(n5380), .ZN(n5379) );
  NOR2_X1 U5740 ( .A1(n9287), .A2(n9295), .ZN(n5380) );
  NAND2_X1 U5741 ( .A1(n5378), .A2(n6653), .ZN(n9281) );
  NAND2_X1 U5742 ( .A1(n5126), .A2(n5124), .ZN(n5386) );
  INV_X1 U5743 ( .A(n8833), .ZN(n9306) );
  NAND2_X1 U5744 ( .A1(n6569), .A2(n6568), .ZN(n6578) );
  NOR2_X1 U5745 ( .A1(n6561), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6569) );
  OR2_X1 U5746 ( .A1(n6551), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6561) );
  NAND2_X1 U5747 ( .A1(n5371), .A2(n5373), .ZN(n9337) );
  NOR2_X1 U5748 ( .A1(n5372), .A2(n5001), .ZN(n5371) );
  INV_X1 U5749 ( .A(n6645), .ZN(n5372) );
  NAND2_X1 U5750 ( .A1(n6532), .A2(n10544), .ZN(n6542) );
  AND2_X1 U5751 ( .A1(n6522), .A2(n9093), .ZN(n6532) );
  AOI21_X1 U5752 ( .B1(n5447), .B2(n5450), .A(n8607), .ZN(n5445) );
  AND2_X1 U5753 ( .A1(n9557), .A2(n5456), .ZN(n5455) );
  INV_X1 U5754 ( .A(n5462), .ZN(n5461) );
  AOI21_X1 U5755 ( .B1(n5462), .B2(n5460), .A(n5459), .ZN(n5458) );
  INV_X1 U5756 ( .A(n9549), .ZN(n9557) );
  NAND2_X1 U5757 ( .A1(n6433), .A2(n6432), .ZN(n6459) );
  NAND2_X1 U5758 ( .A1(n8127), .A2(n6634), .ZN(n9467) );
  NAND2_X1 U5759 ( .A1(n5096), .A2(n5095), .ZN(n8126) );
  AOI22_X1 U5760 ( .A1(n5097), .A2(n5102), .B1(n5098), .B2(n5100), .ZN(n5095)
         );
  INV_X1 U5761 ( .A(n8009), .ZN(n5100) );
  OR2_X1 U5762 ( .A1(n8126), .A2(n8767), .ZN(n8127) );
  OR2_X1 U5763 ( .A1(n6402), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6417) );
  NAND2_X1 U5764 ( .A1(n6379), .A2(n6378), .ZN(n6392) );
  INV_X1 U5765 ( .A(n6380), .ZN(n6379) );
  OR2_X1 U5766 ( .A1(n6392), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U5767 ( .A1(n6311), .A2(n10459), .ZN(n6331) );
  INV_X1 U5768 ( .A(n6312), .ZN(n6311) );
  INV_X1 U5769 ( .A(n5465), .ZN(n5466) );
  OAI21_X1 U5770 ( .B1(n8665), .B2(n5469), .A(n8668), .ZN(n5465) );
  NAND2_X1 U5771 ( .A1(n7387), .A2(n8745), .ZN(n7481) );
  NAND2_X1 U5772 ( .A1(n7481), .A2(n8665), .ZN(n7771) );
  NAND2_X1 U5773 ( .A1(n10466), .A2(n10456), .ZN(n6312) );
  NAND2_X1 U5774 ( .A1(n5112), .A2(n8729), .ZN(n5114) );
  INV_X1 U5775 ( .A(n7383), .ZN(n5112) );
  INV_X1 U5776 ( .A(n9148), .ZN(n7484) );
  AND2_X1 U5777 ( .A1(n8748), .A2(n8732), .ZN(n8663) );
  OAI21_X1 U5778 ( .B1(n7100), .B2(n7099), .A(n7098), .ZN(n7097) );
  AND4_X1 U5779 ( .A1(n6291), .A2(n6290), .A3(n6289), .A4(n6288), .ZN(n7384)
         );
  INV_X1 U5780 ( .A(n7098), .ZN(n8722) );
  NAND2_X1 U5781 ( .A1(n6292), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6284) );
  NOR2_X1 U5782 ( .A1(n5091), .A2(n5090), .ZN(n5089) );
  NOR2_X1 U5783 ( .A1(n5094), .A2(n8864), .ZN(n5090) );
  NAND2_X1 U5784 ( .A1(n6292), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5358) );
  NOR2_X1 U5785 ( .A1(n6783), .A2(n8328), .ZN(n5356) );
  AND2_X1 U5786 ( .A1(n6628), .A2(n5353), .ZN(n7100) );
  INV_X1 U5787 ( .A(n7076), .ZN(n5353) );
  CLKBUF_X1 U5788 ( .A(n6865), .Z(n7182) );
  OR2_X1 U5789 ( .A1(n6386), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n6398) );
  OR2_X1 U5790 ( .A1(n5935), .A2(n5934), .ZN(n5958) );
  NOR2_X1 U5791 ( .A1(n9673), .A2(n5406), .ZN(n5405) );
  INV_X1 U5792 ( .A(n8920), .ZN(n5406) );
  INV_X1 U5793 ( .A(n5396), .ZN(n5395) );
  OAI21_X1 U5794 ( .B1(n9693), .B2(n8890), .A(n9702), .ZN(n5396) );
  NAND2_X1 U5795 ( .A1(n4973), .A2(n5402), .ZN(n5398) );
  NAND2_X1 U5796 ( .A1(n4973), .A2(n5400), .ZN(n5399) );
  INV_X1 U5797 ( .A(n8094), .ZN(n5400) );
  CLKBUF_X1 U5798 ( .A(n6998), .Z(n8902) );
  AND2_X1 U5799 ( .A1(n6057), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6078) );
  AND2_X1 U5800 ( .A1(n9765), .A2(n9762), .ZN(n8960) );
  INV_X1 U5801 ( .A(n8564), .ZN(n5239) );
  AND2_X1 U5802 ( .A1(n9996), .A2(n9995), .ZN(n5240) );
  INV_X2 U5803 ( .A(n8292), .ZN(n6141) );
  NAND2_X1 U5804 ( .A1(n9987), .A2(n6108), .ZN(n6718) );
  NAND2_X1 U5805 ( .A1(n8264), .A2(n8333), .ZN(n6099) );
  NAND2_X1 U5806 ( .A1(n5519), .A2(n5518), .ZN(n10017) );
  NAND2_X1 U5807 ( .A1(n10061), .A2(n5004), .ZN(n10053) );
  NAND2_X1 U5808 ( .A1(n10120), .A2(n5285), .ZN(n10046) );
  NOR2_X1 U5809 ( .A1(n5287), .A2(n10232), .ZN(n5285) );
  NAND2_X1 U5810 ( .A1(n10171), .A2(n5298), .ZN(n10138) );
  NAND2_X1 U5811 ( .A1(n10163), .A2(n8553), .ZN(n10146) );
  NAND2_X1 U5812 ( .A1(n10171), .A2(n10336), .ZN(n10172) );
  NAND2_X1 U5813 ( .A1(n8204), .A2(n5040), .ZN(n8114) );
  INV_X1 U5814 ( .A(n5516), .ZN(n8040) );
  OAI21_X1 U5815 ( .B1(n5179), .B2(n4968), .A(n5177), .ZN(n5516) );
  AOI21_X1 U5816 ( .B1(n10780), .B2(n5176), .A(n5020), .ZN(n5177) );
  NAND2_X1 U5817 ( .A1(n5234), .A2(n5235), .ZN(n8036) );
  AND2_X1 U5818 ( .A1(n5235), .A2(n5233), .ZN(n5232) );
  NOR2_X1 U5819 ( .A1(n8188), .A2(n5293), .ZN(n5292) );
  NOR2_X1 U5820 ( .A1(n7501), .A2(n5293), .ZN(n10781) );
  NOR3_X1 U5821 ( .A1(n7501), .A2(n7969), .A3(n7807), .ZN(n10784) );
  OR2_X1 U5822 ( .A1(n7807), .A2(n9799), .ZN(n5868) );
  NAND2_X1 U5823 ( .A1(n7557), .A2(n8460), .ZN(n7556) );
  NAND2_X1 U5824 ( .A1(n5524), .A2(n5525), .ZN(n7497) );
  AOI21_X1 U5825 ( .B1(n8359), .B2(n5526), .A(n5018), .ZN(n5525) );
  INV_X1 U5826 ( .A(n5841), .ZN(n5526) );
  NAND2_X1 U5827 ( .A1(n7683), .A2(n5807), .ZN(n7170) );
  AND2_X1 U5828 ( .A1(n8340), .A2(n8522), .ZN(n8452) );
  NAND2_X1 U5829 ( .A1(n8520), .A2(n10721), .ZN(n5746) );
  INV_X1 U5830 ( .A(n8452), .ZN(n8342) );
  INV_X1 U5831 ( .A(n5063), .ZN(n10186) );
  NAND2_X1 U5832 ( .A1(n5136), .A2(n5739), .ZN(n10194) );
  AND3_X1 U5833 ( .A1(n5737), .A2(n5740), .A3(n5738), .ZN(n5136) );
  INV_X1 U5834 ( .A(n8451), .ZN(n7064) );
  NAND2_X1 U5835 ( .A1(n7060), .A2(n7064), .ZN(n7059) );
  NOR2_X1 U5836 ( .A1(n8449), .A2(n10194), .ZN(n8450) );
  NAND2_X1 U5837 ( .A1(n6056), .A2(n6055), .ZN(n10220) );
  NAND2_X1 U5838 ( .A1(n8051), .A2(n8333), .ZN(n6056) );
  NAND2_X1 U5839 ( .A1(n5984), .A2(n5983), .ZN(n10091) );
  INV_X1 U5840 ( .A(n9649), .ZN(n8877) );
  OR2_X1 U5841 ( .A1(n7044), .A2(n5290), .ZN(n7052) );
  INV_X1 U5842 ( .A(n10794), .ZN(n10268) );
  XNOR2_X1 U5843 ( .A(n8327), .B(n8326), .ZN(n8990) );
  OR2_X1 U5844 ( .A1(n5666), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n5667) );
  XNOR2_X1 U5845 ( .A(n6613), .B(n6612), .ZN(n8993) );
  NAND2_X1 U5846 ( .A1(n6110), .A2(n6096), .ZN(n8264) );
  OR2_X1 U5847 ( .A1(n6095), .A2(n6094), .ZN(n6096) );
  NAND2_X1 U5848 ( .A1(n5332), .A2(n5337), .ZN(n6095) );
  NAND2_X1 U5849 ( .A1(n6071), .A2(n5339), .ZN(n5332) );
  NAND2_X1 U5850 ( .A1(n5299), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6173) );
  AND2_X1 U5851 ( .A1(n5981), .A2(n5967), .ZN(n5968) );
  OAI21_X1 U5852 ( .B1(n5320), .B2(n5327), .A(n5638), .ZN(n5690) );
  INV_X1 U5853 ( .A(n5319), .ZN(n5320) );
  NAND2_X1 U5854 ( .A1(n5319), .A2(n5630), .ZN(n5879) );
  OR2_X1 U5855 ( .A1(n5843), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5855) );
  XNOR2_X1 U5856 ( .A(n5242), .B(n5842), .ZN(n6796) );
  NAND2_X1 U5857 ( .A1(n5309), .A2(n5614), .ZN(n5242) );
  XNOR2_X1 U5858 ( .A(n5601), .B(n5600), .ZN(n5786) );
  INV_X1 U5859 ( .A(n5757), .ZN(n5305) );
  CLKBUF_X1 U5860 ( .A(n5691), .Z(n5692) );
  INV_X1 U5861 ( .A(n5420), .ZN(n5419) );
  AOI21_X1 U5862 ( .B1(n5420), .B2(n7667), .A(n4975), .ZN(n5418) );
  NOR2_X1 U5863 ( .A1(n8636), .A2(n5427), .ZN(n5423) );
  OAI21_X1 U5864 ( .B1(n8636), .B2(n5426), .A(n5425), .ZN(n5424) );
  NAND2_X1 U5865 ( .A1(n8636), .A2(n5430), .ZN(n5425) );
  NOR2_X1 U5866 ( .A1(n5427), .A2(n5432), .ZN(n5426) );
  NAND2_X1 U5867 ( .A1(n8636), .A2(n5432), .ZN(n5428) );
  NAND2_X1 U5868 ( .A1(n5434), .A2(n5005), .ZN(n8103) );
  NAND2_X1 U5869 ( .A1(n5434), .A2(n8023), .ZN(n8024) );
  NAND2_X1 U5870 ( .A1(n8598), .A2(n8597), .ZN(n9053) );
  AND2_X1 U5871 ( .A1(n9014), .A2(n7205), .ZN(n5439) );
  OR2_X1 U5872 ( .A1(n6862), .A2(n6861), .ZN(n9094) );
  NAND2_X1 U5873 ( .A1(n6429), .A2(n6428), .ZN(n9567) );
  NAND2_X1 U5874 ( .A1(n9034), .A2(n5006), .ZN(n9104) );
  NAND2_X1 U5875 ( .A1(n9034), .A2(n8616), .ZN(n9103) );
  AND2_X1 U5876 ( .A1(n6519), .A2(n6518), .ZN(n9113) );
  NAND2_X1 U5877 ( .A1(n6577), .A2(n6576), .ZN(n9308) );
  NAND2_X1 U5878 ( .A1(n8228), .A2(n8656), .ZN(n6577) );
  NAND2_X1 U5879 ( .A1(n8270), .A2(n5444), .ZN(n8598) );
  AOI21_X1 U5880 ( .B1(n5195), .B2(n4977), .A(n5192), .ZN(n8858) );
  OAI21_X1 U5881 ( .B1(n5194), .B2(n8855), .A(n5193), .ZN(n5192) );
  OAI21_X1 U5882 ( .B1(n5492), .B2(n5482), .A(n5479), .ZN(n8694) );
  NAND4_X1 U5883 ( .A1(n6337), .A2(n6336), .A3(n6335), .A4(n6334), .ZN(n9146)
         );
  NAND2_X1 U5884 ( .A1(n7151), .A2(n5265), .ZN(n6930) );
  AND2_X1 U5885 ( .A1(n7227), .A2(n7226), .ZN(n7229) );
  NOR2_X1 U5886 ( .A1(n7524), .A2(n7523), .ZN(n7526) );
  INV_X1 U5887 ( .A(n5068), .ZN(n10684) );
  NOR2_X1 U5888 ( .A1(n9153), .A2(n9154), .ZN(n9156) );
  INV_X1 U5889 ( .A(n5062), .ZN(n9152) );
  NOR2_X1 U5890 ( .A1(n9181), .A2(n6461), .ZN(n9201) );
  NAND2_X1 U5891 ( .A1(n5221), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5220) );
  NOR2_X1 U5892 ( .A1(n9247), .A2(n9248), .ZN(n10712) );
  OAI21_X1 U5893 ( .B1(n9225), .B2(n5208), .A(n5207), .ZN(n10715) );
  NAND2_X1 U5894 ( .A1(n5209), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5208) );
  INV_X1 U5895 ( .A(n10711), .ZN(n5209) );
  XNOR2_X1 U5896 ( .A(n5070), .B(n9262), .ZN(n9268) );
  INV_X1 U5897 ( .A(n8686), .ZN(n6626) );
  OAI21_X1 U5898 ( .B1(n5492), .B2(n5488), .A(n5486), .ZN(n8690) );
  AND2_X1 U5899 ( .A1(n8588), .A2(n6589), .ZN(n9288) );
  NAND2_X1 U5900 ( .A1(n5116), .A2(n5115), .ZN(n9294) );
  NAND2_X1 U5901 ( .A1(n9314), .A2(n4978), .ZN(n5115) );
  INV_X1 U5902 ( .A(n5117), .ZN(n5116) );
  NAND2_X1 U5903 ( .A1(n6567), .A2(n6566), .ZN(n9318) );
  NAND2_X1 U5904 ( .A1(n5497), .A2(n5502), .ZN(n9322) );
  NAND2_X1 U5905 ( .A1(n9341), .A2(n5504), .ZN(n5497) );
  NAND2_X1 U5906 ( .A1(n5506), .A2(n8662), .ZN(n9334) );
  NAND2_X1 U5907 ( .A1(n5508), .A2(n5507), .ZN(n5506) );
  AND2_X1 U5908 ( .A1(n5373), .A2(n6645), .ZN(n9350) );
  AND2_X1 U5909 ( .A1(n9371), .A2(n9370), .ZN(n9372) );
  NAND2_X1 U5910 ( .A1(n9376), .A2(n4982), .ZN(n9515) );
  NAND2_X1 U5911 ( .A1(n6531), .A2(n6530), .ZN(n9375) );
  NAND2_X1 U5912 ( .A1(n9422), .A2(n9421), .ZN(n9420) );
  NAND2_X1 U5913 ( .A1(n9433), .A2(n6495), .ZN(n9422) );
  NAND2_X1 U5914 ( .A1(n6501), .A2(n6500), .ZN(n9530) );
  NAND2_X1 U5915 ( .A1(n6486), .A2(n6485), .ZN(n9534) );
  NAND2_X1 U5916 ( .A1(n9445), .A2(n6481), .ZN(n9448) );
  NAND2_X1 U5917 ( .A1(n6474), .A2(n6473), .ZN(n9538) );
  OAI21_X1 U5918 ( .B1(n9548), .B2(n5352), .A(n5350), .ZN(n9439) );
  NAND2_X1 U5919 ( .A1(n6457), .A2(n6456), .ZN(n9545) );
  NAND2_X1 U5920 ( .A1(n9548), .A2(n8791), .ZN(n9456) );
  NAND2_X1 U5921 ( .A1(n8131), .A2(n8769), .ZN(n9465) );
  NAND2_X1 U5922 ( .A1(n8011), .A2(n8008), .ZN(n5103) );
  OAI21_X1 U5923 ( .B1(n6366), .B2(n5476), .A(n5474), .ZN(n8010) );
  NAND2_X1 U5924 ( .A1(n6391), .A2(n6390), .ZN(n8144) );
  NAND2_X1 U5925 ( .A1(n5362), .A2(n5366), .ZN(n7990) );
  NAND2_X1 U5926 ( .A1(n7796), .A2(n5367), .ZN(n5362) );
  AND2_X1 U5927 ( .A1(n5478), .A2(n8707), .ZN(n7989) );
  NAND2_X1 U5928 ( .A1(n6366), .A2(n8756), .ZN(n5478) );
  AOI21_X1 U5929 ( .B1(n7796), .B2(n7795), .A(n4970), .ZN(n7983) );
  INV_X1 U5930 ( .A(n7293), .ZN(n7873) );
  NAND2_X1 U5931 ( .A1(n5107), .A2(n5108), .ZN(n7773) );
  NAND2_X1 U5932 ( .A1(n7383), .A2(n5109), .ZN(n5107) );
  INV_X1 U5933 ( .A(n9278), .ZN(n9576) );
  NAND2_X1 U5934 ( .A1(n9485), .A2(n9486), .ZN(n9577) );
  INV_X1 U5935 ( .A(n9318), .ZN(n9589) );
  OR2_X1 U5936 ( .A1(n9611), .A2(n6800), .ZN(n8278) );
  AND2_X1 U5937 ( .A1(n5496), .A2(n5495), .ZN(n5494) );
  NOR2_X1 U5938 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n5495) );
  INV_X1 U5939 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9613) );
  AND2_X1 U5940 ( .A1(P2_U3151), .A2(n8328), .ZN(n9623) );
  INV_X1 U5941 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6809) );
  INV_X1 U5942 ( .A(n4948), .ZN(n7349) );
  INV_X1 U5943 ( .A(n6922), .ZN(n7122) );
  INV_X1 U5944 ( .A(n9990), .ZN(n10206) );
  NAND2_X1 U5945 ( .A1(n9732), .A2(n8920), .ZN(n9674) );
  NAND2_X1 U5946 ( .A1(n5392), .A2(n7411), .ZN(n7439) );
  INV_X1 U5947 ( .A(n5394), .ZN(n5392) );
  NAND2_X1 U5948 ( .A1(n9691), .A2(n8891), .ZN(n9701) );
  NAND2_X1 U5949 ( .A1(n5674), .A2(n5673), .ZN(n10282) );
  CLKBUF_X1 U5950 ( .A(n9711), .Z(n9715) );
  NAND2_X1 U5951 ( .A1(n6041), .A2(n6040), .ZN(n10227) );
  NAND2_X1 U5952 ( .A1(n8033), .A2(n8333), .ZN(n6041) );
  NAND2_X1 U5953 ( .A1(n7727), .A2(n5415), .ZN(n5413) );
  NAND2_X1 U5954 ( .A1(n7411), .A2(n7437), .ZN(n5388) );
  INV_X1 U5955 ( .A(n9779), .ZN(n9768) );
  NAND2_X1 U5956 ( .A1(n5906), .A2(n5905), .ZN(n9786) );
  AOI21_X1 U5957 ( .B1(n8447), .B2(n5148), .A(n5147), .ZN(n5146) );
  AOI21_X1 U5958 ( .B1(n8575), .B2(n8574), .A(n8573), .ZN(n8580) );
  INV_X1 U5959 ( .A(n10186), .ZN(n9806) );
  OR2_X1 U5960 ( .A1(n6140), .A2(n10190), .ZN(n5725) );
  AND2_X1 U5961 ( .A1(n7081), .A2(n7080), .ZN(n7083) );
  NOR2_X1 U5962 ( .A1(n9956), .A2(n10174), .ZN(n10202) );
  NAND2_X1 U5963 ( .A1(n5341), .A2(n8288), .ZN(n9963) );
  XNOR2_X1 U5964 ( .A(n6718), .B(n8476), .ZN(n9975) );
  AND2_X1 U5965 ( .A1(n10028), .A2(n10267), .ZN(n5057) );
  INV_X1 U5966 ( .A(n9792), .ZN(n10205) );
  NAND2_X1 U5967 ( .A1(n5542), .A2(n5543), .ZN(n9989) );
  INV_X1 U5968 ( .A(n5545), .ZN(n10008) );
  NAND2_X1 U5969 ( .A1(n5545), .A2(n5544), .ZN(n10213) );
  INV_X1 U5970 ( .A(n10220), .ZN(n10025) );
  NAND2_X1 U5971 ( .A1(n10064), .A2(n6009), .ZN(n10045) );
  NAND2_X1 U5972 ( .A1(n5165), .A2(n5169), .ZN(n10081) );
  OR2_X1 U5973 ( .A1(n10116), .A2(n5171), .ZN(n5165) );
  AND2_X1 U5974 ( .A1(n5172), .A2(n4989), .ZN(n10102) );
  NAND2_X1 U5975 ( .A1(n10116), .A2(n10113), .ZN(n5172) );
  NAND2_X1 U5976 ( .A1(n5956), .A2(n5955), .ZN(n10125) );
  NAND2_X1 U5977 ( .A1(n5527), .A2(n5533), .ZN(n10132) );
  OR2_X1 U5978 ( .A1(n10170), .A2(n5535), .ZN(n5527) );
  OR2_X1 U5979 ( .A1(n10170), .A2(n5538), .ZN(n5532) );
  NAND2_X1 U5980 ( .A1(n8040), .A2(n8466), .ZN(n8204) );
  NAND2_X1 U5981 ( .A1(n7893), .A2(n5238), .ZN(n7896) );
  NAND2_X1 U5982 ( .A1(n5178), .A2(n4972), .ZN(n7898) );
  NAND2_X1 U5983 ( .A1(n5179), .A2(n5181), .ZN(n5178) );
  AND2_X1 U5984 ( .A1(n5181), .A2(n5180), .ZN(n7831) );
  INV_X1 U5985 ( .A(n10184), .ZN(n10814) );
  NAND2_X1 U5986 ( .A1(n7458), .A2(n8359), .ZN(n7457) );
  NAND2_X1 U5987 ( .A1(n7322), .A2(n5841), .ZN(n7458) );
  NAND2_X1 U5988 ( .A1(n5831), .A2(n5830), .ZN(n8313) );
  NAND2_X1 U5989 ( .A1(n7050), .A2(n5790), .ZN(n7684) );
  INV_X1 U5990 ( .A(n9805), .ZN(n7657) );
  CLKBUF_X1 U5991 ( .A(n10194), .Z(n5056) );
  INV_X1 U5992 ( .A(n9963), .ZN(n10306) );
  INV_X1 U5993 ( .A(n10125), .ZN(n10327) );
  INV_X1 U5994 ( .A(n9786), .ZN(n10341) );
  INV_X1 U5995 ( .A(n7851), .ZN(n5824) );
  INV_X1 U5996 ( .A(n10193), .ZN(n8520) );
  OAI21_X1 U5997 ( .B1(n8327), .B2(n8326), .A(n8325), .ZN(n8331) );
  NAND2_X1 U5998 ( .A1(n5160), .A2(n4993), .ZN(n10349) );
  INV_X1 U5999 ( .A(n5664), .ZN(n5160) );
  INV_X1 U6000 ( .A(n5584), .ZN(n10352) );
  CLKBUF_X1 U6001 ( .A(n6146), .Z(n8995) );
  XNOR2_X1 U6002 ( .A(n5663), .B(n5665), .ZN(n8304) );
  NAND2_X1 U6003 ( .A1(n5310), .A2(n6014), .ZN(n6021) );
  AND2_X1 U6004 ( .A1(P1_U3086), .A2(n8328), .ZN(n10343) );
  OR2_X1 U6005 ( .A1(n5671), .A2(n6124), .ZN(n5887) );
  AND2_X1 U6006 ( .A1(n5814), .A2(n5828), .ZN(n9887) );
  AND2_X1 U6007 ( .A1(n9002), .A2(n5041), .ZN(n5064) );
  INV_X1 U6008 ( .A(n5213), .ZN(n7738) );
  INV_X1 U6009 ( .A(n5218), .ZN(n7925) );
  OAI21_X1 U6010 ( .B1(n8589), .B2(n9529), .A(n6761), .ZN(n6762) );
  OAI21_X1 U6011 ( .B1(n6759), .B2(n10850), .A(n6716), .ZN(P2_U3456) );
  NOR2_X1 U6012 ( .A1(n8589), .A2(n9606), .ZN(n6714) );
  AND2_X1 U6013 ( .A1(n5229), .A2(n5231), .ZN(n9974) );
  AOI21_X1 U6014 ( .B1(n5226), .B2(n5228), .A(n6748), .ZN(n5225) );
  AND2_X1 U6015 ( .A1(n5157), .A2(n10831), .ZN(n5226) );
  OR2_X1 U6016 ( .A1(n10831), .A2(n6745), .ZN(n5512) );
  AND2_X1 U6017 ( .A1(n5229), .A2(n5227), .ZN(n6749) );
  AOI21_X1 U6018 ( .B1(n9983), .B2(n6205), .A(n6204), .ZN(n6206) );
  INV_X4 U6019 ( .A(n6998), .ZN(n7254) );
  NAND2_X1 U6020 ( .A1(n4972), .A2(n5008), .ZN(n4968) );
  OR2_X1 U6021 ( .A1(n9278), .A2(n8659), .ZN(n8853) );
  AND2_X1 U6022 ( .A1(n5515), .A2(n9797), .ZN(n4969) );
  AND2_X1 U6024 ( .A1(n8745), .A2(n8734), .ZN(n7388) );
  AND2_X1 U6025 ( .A1(n7844), .A2(n8704), .ZN(n4970) );
  NAND2_X1 U6026 ( .A1(n10176), .A2(n9793), .ZN(n4971) );
  INV_X1 U6027 ( .A(n9983), .ZN(n5301) );
  OR2_X1 U6028 ( .A1(n10825), .A2(n10795), .ZN(n4972) );
  INV_X1 U6029 ( .A(n8386), .ZN(n5253) );
  NOR2_X1 U6030 ( .A1(n8218), .A2(n8219), .ZN(n4973) );
  INV_X1 U6031 ( .A(n5171), .ZN(n5170) );
  NAND2_X1 U6032 ( .A1(n10101), .A2(n4989), .ZN(n5171) );
  AND2_X1 U6033 ( .A1(n5363), .A2(n8671), .ZN(n4974) );
  INV_X1 U6034 ( .A(n8008), .ZN(n5099) );
  AND2_X1 U6035 ( .A1(n7973), .A2(n5421), .ZN(n4975) );
  AND2_X1 U6036 ( .A1(n9308), .A2(n9137), .ZN(n4976) );
  AND3_X1 U6037 ( .A1(n8853), .A2(n8852), .A3(n8857), .ZN(n4977) );
  INV_X1 U6038 ( .A(n8828), .ZN(n5507) );
  AND2_X1 U6039 ( .A1(n5124), .A2(n9293), .ZN(n4978) );
  INV_X1 U6040 ( .A(n8775), .ZN(n5459) );
  INV_X1 U6041 ( .A(n5228), .ZN(n5227) );
  NAND2_X1 U6042 ( .A1(n5159), .A2(n5158), .ZN(n5228) );
  INV_X1 U6043 ( .A(n10232), .ZN(n10050) );
  NAND2_X1 U6044 ( .A1(n6024), .A2(n6023), .ZN(n10232) );
  INV_X1 U6045 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6232) );
  INV_X1 U6046 ( .A(n9455), .ZN(n5352) );
  INV_X1 U6047 ( .A(n9246), .ZN(n5210) );
  NAND2_X1 U6048 ( .A1(n7511), .A2(n5437), .ZN(n7605) );
  NAND2_X1 U6049 ( .A1(n7258), .A2(n7257), .ZN(n7259) );
  AND2_X1 U6050 ( .A1(n10701), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4979) );
  OR2_X1 U6051 ( .A1(n8004), .A2(n7673), .ZN(n8756) );
  INV_X1 U6052 ( .A(n9728), .ZN(n5290) );
  AND2_X1 U6053 ( .A1(n5724), .A2(n5726), .ZN(n4980) );
  INV_X1 U6054 ( .A(n8466), .ZN(n5233) );
  OR2_X1 U6055 ( .A1(n5731), .A2(n6949), .ZN(n4981) );
  NAND2_X1 U6056 ( .A1(n8702), .A2(n8701), .ZN(n4982) );
  INV_X2 U6057 ( .A(n6771), .ZN(n8328) );
  AND2_X1 U6058 ( .A1(n8997), .A2(n5433), .ZN(n5432) );
  NAND2_X1 U6059 ( .A1(n9148), .A2(n9082), .ZN(n4983) );
  NAND2_X1 U6060 ( .A1(n5007), .A2(n6651), .ZN(n5125) );
  AND2_X1 U6061 ( .A1(n8887), .A2(n8886), .ZN(n8890) );
  OR2_X1 U6062 ( .A1(n10675), .A2(n7923), .ZN(n4984) );
  OR2_X1 U6063 ( .A1(n10143), .A2(n10257), .ZN(n4985) );
  AND2_X1 U6064 ( .A1(n10025), .A2(n10224), .ZN(n4986) );
  OR2_X1 U6065 ( .A1(n8144), .A2(n8057), .ZN(n4987) );
  NAND2_X1 U6066 ( .A1(n8925), .A2(n8924), .ZN(n4988) );
  OR2_X1 U6067 ( .A1(n10327), .A2(n9756), .ZN(n4989) );
  NAND2_X1 U6068 ( .A1(n5916), .A2(n5915), .ZN(n10176) );
  INV_X1 U6069 ( .A(n8662), .ZN(n5505) );
  AND2_X1 U6070 ( .A1(n8562), .A2(n8442), .ZN(n4990) );
  AND3_X1 U6071 ( .A1(n8518), .A2(n8553), .A3(n8445), .ZN(n4991) );
  NAND2_X1 U6072 ( .A1(n8786), .A2(n8784), .ZN(n9455) );
  NOR2_X1 U6073 ( .A1(n9348), .A2(n9355), .ZN(n4992) );
  NAND2_X1 U6074 ( .A1(n6001), .A2(n6000), .ZN(n10077) );
  NOR2_X1 U6075 ( .A1(n5666), .A2(n5577), .ZN(n4993) );
  INV_X1 U6076 ( .A(n10143), .ZN(n10331) );
  NAND2_X1 U6077 ( .A1(n5933), .A2(n5932), .ZN(n10143) );
  NAND2_X1 U6078 ( .A1(n5754), .A2(n5511), .ZN(n5783) );
  AND2_X1 U6079 ( .A1(n6257), .A2(n8328), .ZN(n4994) );
  AND2_X1 U6080 ( .A1(n7954), .A2(n7953), .ZN(n4995) );
  NOR2_X1 U6081 ( .A1(n7228), .A2(n7490), .ZN(n4996) );
  OR2_X1 U6082 ( .A1(n8632), .A2(n9305), .ZN(n8660) );
  NOR2_X1 U6083 ( .A1(n9168), .A2(n9169), .ZN(n4997) );
  NOR2_X1 U6084 ( .A1(n9201), .A2(n9200), .ZN(n4998) );
  NOR2_X1 U6085 ( .A1(n9214), .A2(n9215), .ZN(n4999) );
  NOR2_X1 U6086 ( .A1(n8689), .A2(n8851), .ZN(n5000) );
  NOR2_X1 U6087 ( .A1(n9101), .A2(n9338), .ZN(n5001) );
  INV_X1 U6088 ( .A(n5504), .ZN(n5503) );
  NAND2_X1 U6089 ( .A1(n6148), .A2(n8413), .ZN(n10084) );
  INV_X1 U6090 ( .A(n10084), .ZN(n5167) );
  AND2_X1 U6091 ( .A1(n4985), .A2(n5535), .ZN(n5002) );
  AND2_X1 U6092 ( .A1(n8437), .A2(n8503), .ZN(n5003) );
  AND2_X1 U6093 ( .A1(n8632), .A2(n9305), .ZN(n8840) );
  INV_X1 U6094 ( .A(n8840), .ZN(n5491) );
  INV_X1 U6095 ( .A(n10110), .ZN(n10323) );
  NAND2_X1 U6096 ( .A1(n5971), .A2(n5970), .ZN(n10110) );
  AND2_X1 U6097 ( .A1(n10054), .A2(n8421), .ZN(n5004) );
  AND2_X1 U6098 ( .A1(n8026), .A2(n8023), .ZN(n5005) );
  AND2_X1 U6099 ( .A1(n8617), .A2(n8616), .ZN(n5006) );
  OR2_X1 U6100 ( .A1(n9308), .A2(n9137), .ZN(n5007) );
  INV_X1 U6101 ( .A(n5102), .ZN(n5101) );
  NAND2_X1 U6102 ( .A1(n8009), .A2(n9141), .ZN(n5102) );
  NAND2_X1 U6103 ( .A1(n6560), .A2(n6559), .ZN(n8698) );
  INV_X1 U6104 ( .A(n8698), .ZN(n5510) );
  NAND2_X1 U6105 ( .A1(n8213), .A2(n9795), .ZN(n5008) );
  AND2_X1 U6106 ( .A1(n5532), .A2(n5536), .ZN(n5009) );
  AND2_X1 U6107 ( .A1(n8495), .A2(n8494), .ZN(n5010) );
  AND2_X1 U6108 ( .A1(n10214), .A2(n10028), .ZN(n5011) );
  AND2_X1 U6109 ( .A1(n8334), .A2(n8502), .ZN(n8435) );
  INV_X1 U6110 ( .A(n8435), .ZN(n8476) );
  AND2_X1 U6111 ( .A1(n8464), .A2(n8391), .ZN(n5238) );
  INV_X1 U6112 ( .A(n5402), .ZN(n5401) );
  INV_X2 U6113 ( .A(n8903), .ZN(n8965) );
  NOR2_X1 U6114 ( .A1(n7483), .A2(n7873), .ZN(n5012) );
  AND2_X1 U6115 ( .A1(n10323), .A2(n9676), .ZN(n5013) );
  NAND2_X1 U6116 ( .A1(n8875), .A2(n8874), .ZN(n5014) );
  INV_X1 U6117 ( .A(n8769), .ZN(n5463) );
  INV_X1 U6118 ( .A(n5287), .ZN(n5286) );
  NAND2_X1 U6119 ( .A1(n5288), .A2(n10315), .ZN(n5287) );
  AND2_X1 U6120 ( .A1(n10050), .A2(n10071), .ZN(n5015) );
  OR2_X1 U6121 ( .A1(n5122), .A2(n9293), .ZN(n5016) );
  NOR2_X1 U6122 ( .A1(n10769), .A2(n9143), .ZN(n5017) );
  NOR2_X1 U6123 ( .A1(n8374), .A2(n9800), .ZN(n5018) );
  NOR2_X1 U6124 ( .A1(n8004), .A2(n9144), .ZN(n5019) );
  OAI22_X1 U6125 ( .A1(n6747), .A2(n10298), .B1(n10831), .B2(n6746), .ZN(n6748) );
  INV_X1 U6126 ( .A(n5369), .ZN(n5113) );
  AND2_X1 U6127 ( .A1(n7492), .A2(n9147), .ZN(n5369) );
  AND2_X1 U6128 ( .A1(n8227), .A2(n9646), .ZN(n5020) );
  INV_X1 U6129 ( .A(n5689), .ZN(n5641) );
  XNOR2_X1 U6130 ( .A(n5639), .B(n10393), .ZN(n5689) );
  AND2_X1 U6131 ( .A1(n5476), .A2(n4987), .ZN(n5021) );
  OR3_X1 U6132 ( .A1(n8374), .A2(n8445), .A3(n8373), .ZN(n5022) );
  AND2_X1 U6133 ( .A1(n5491), .A2(n8660), .ZN(n9296) );
  INV_X1 U6134 ( .A(n9296), .ZN(n9293) );
  OR2_X1 U6135 ( .A1(n5382), .A2(n5377), .ZN(n5023) );
  AND2_X1 U6136 ( .A1(n5510), .A2(n5509), .ZN(n5024) );
  AND2_X1 U6137 ( .A1(n9278), .A2(n8659), .ZN(n8689) );
  AND2_X1 U6138 ( .A1(n6919), .A2(n6928), .ZN(n5025) );
  OAI21_X1 U6139 ( .B1(n8729), .B2(n5111), .A(n5370), .ZN(n5110) );
  INV_X1 U6140 ( .A(n5125), .ZN(n5124) );
  OR2_X1 U6141 ( .A1(n10769), .A2(n8013), .ZN(n8760) );
  NOR2_X1 U6142 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5026) );
  INV_X1 U6143 ( .A(n4971), .ZN(n5538) );
  AND2_X1 U6144 ( .A1(n5474), .A2(n4987), .ZN(n5027) );
  OR2_X1 U6145 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n5666) );
  OR2_X1 U6146 ( .A1(n10025), .A2(n10224), .ZN(n5028) );
  OR2_X1 U6147 ( .A1(n7028), .A2(n10739), .ZN(n5029) );
  AND2_X1 U6148 ( .A1(n8934), .A2(n4988), .ZN(n5030) );
  NOR2_X1 U6149 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n5031) );
  AND2_X1 U6150 ( .A1(n10719), .A2(n10717), .ZN(n5032) );
  OR2_X1 U6151 ( .A1(n9523), .A2(n9415), .ZN(n5033) );
  OR2_X1 U6152 ( .A1(n5097), .A2(n5098), .ZN(n5034) );
  INV_X1 U6153 ( .A(n6919), .ZN(n7126) );
  OR2_X1 U6154 ( .A1(n10091), .A2(n10106), .ZN(n6148) );
  AND2_X1 U6155 ( .A1(n5398), .A2(n5014), .ZN(n5035) );
  AND2_X1 U6156 ( .A1(n7973), .A2(n7668), .ZN(n5036) );
  NAND2_X1 U6157 ( .A1(n5619), .A2(n5618), .ZN(n5842) );
  AND2_X1 U6158 ( .A1(n5026), .A2(n5416), .ZN(n5037) );
  AND2_X1 U6159 ( .A1(n5580), .A2(n5579), .ZN(n5038) );
  INV_X2 U6160 ( .A(n6458), .ZN(n6436) );
  AND2_X1 U6161 ( .A1(n10732), .A2(n7578), .ZN(n10809) );
  NAND2_X1 U6162 ( .A1(n10780), .A2(n8195), .ZN(n5181) );
  INV_X1 U6163 ( .A(n9446), .ZN(n5349) );
  AND2_X1 U6164 ( .A1(n5403), .A2(n5401), .ZN(n5039) );
  INV_X1 U6165 ( .A(n10655), .ZN(n5359) );
  OR2_X1 U6166 ( .A1(n8877), .A2(n9782), .ZN(n5040) );
  NAND2_X1 U6167 ( .A1(n8717), .A2(n8716), .ZN(n6628) );
  OR2_X1 U6168 ( .A1(n9581), .A2(n9114), .ZN(n5041) );
  NAND2_X1 U6169 ( .A1(n8132), .A2(n8767), .ZN(n8131) );
  NAND2_X1 U6170 ( .A1(n5685), .A2(n5416), .ZN(n5901) );
  AND2_X1 U6171 ( .A1(n8400), .A2(n8396), .ZN(n5042) );
  INV_X1 U6172 ( .A(n9141), .ZN(n8021) );
  NAND2_X1 U6173 ( .A1(n10120), .A2(n5286), .ZN(n5289) );
  AND2_X1 U6174 ( .A1(n9545), .A2(n9551), .ZN(n5043) );
  NAND2_X1 U6175 ( .A1(n6112), .A2(n6111), .ZN(n9983) );
  OR2_X1 U6176 ( .A1(n8093), .A2(n8094), .ZN(n5403) );
  AND2_X1 U6177 ( .A1(n5652), .A2(SI_15_), .ZN(n5044) );
  AND2_X1 U6178 ( .A1(n5397), .A2(n5398), .ZN(n5045) );
  AND2_X1 U6179 ( .A1(n5996), .A2(n5981), .ZN(n5046) );
  AND2_X1 U6180 ( .A1(n5549), .A2(n5512), .ZN(n5047) );
  AND2_X1 U6181 ( .A1(n8270), .A2(n8269), .ZN(n5048) );
  INV_X1 U6182 ( .A(n7630), .ZN(n5073) );
  NAND2_X1 U6183 ( .A1(n9721), .A2(n7407), .ZN(n5394) );
  NAND2_X1 U6184 ( .A1(n6135), .A2(n6137), .ZN(n8442) );
  XNOR2_X1 U6185 ( .A(n8768), .B(n9140), .ZN(n8767) );
  INV_X1 U6186 ( .A(n8767), .ZN(n5460) );
  NAND2_X1 U6187 ( .A1(n5931), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5952) );
  NAND2_X1 U6188 ( .A1(n5413), .A2(n5414), .ZN(n7952) );
  NAND2_X1 U6189 ( .A1(n5478), .A2(n5477), .ZN(n7987) );
  AND2_X1 U6190 ( .A1(n7511), .A2(n7510), .ZN(n7512) );
  NAND2_X1 U6191 ( .A1(n5394), .A2(n7412), .ZN(n7438) );
  INV_X1 U6192 ( .A(n8668), .ZN(n5467) );
  AND2_X1 U6193 ( .A1(n9791), .A2(n8288), .ZN(n5049) );
  AND2_X1 U6194 ( .A1(n8391), .A2(n8392), .ZN(n8463) );
  INV_X1 U6195 ( .A(n8463), .ZN(n5237) );
  AND2_X1 U6196 ( .A1(n5114), .A2(n4983), .ZN(n5050) );
  OR2_X1 U6197 ( .A1(n6135), .A2(n6137), .ZN(n6995) );
  AND2_X1 U6198 ( .A1(n6019), .A2(n6014), .ZN(n5051) );
  INV_X1 U6199 ( .A(n5114), .ZN(n7382) );
  INV_X1 U6200 ( .A(n7359), .ZN(n6859) );
  INV_X1 U6201 ( .A(n8864), .ZN(n5093) );
  INV_X1 U6202 ( .A(n7807), .ZN(n5295) );
  AND2_X1 U6203 ( .A1(n7603), .A2(n8704), .ZN(n5052) );
  INV_X1 U6204 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10422) );
  INV_X1 U6205 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5345) );
  NAND2_X1 U6206 ( .A1(n10786), .A2(n10778), .ZN(n5053) );
  OR2_X1 U6207 ( .A1(n8442), .A2(n8515), .ZN(n10778) );
  NAND2_X1 U6208 ( .A1(n9975), .A2(n5053), .ZN(n5514) );
  NAND2_X1 U6209 ( .A1(n9966), .A2(n10828), .ZN(n5159) );
  NAND2_X2 U6210 ( .A1(n5054), .A2(n7296), .ZN(n7511) );
  INV_X1 U6211 ( .A(n7294), .ZN(n5054) );
  NAND2_X1 U6212 ( .A1(n7291), .A2(n7290), .ZN(n7294) );
  NAND2_X1 U6213 ( .A1(n8247), .A2(n8246), .ZN(n8270) );
  OAI211_X1 U6214 ( .C1(n4965), .C2(n5419), .A(n5417), .B(n5418), .ZN(n7972)
         );
  NAND2_X2 U6215 ( .A1(n5342), .A2(n5343), .ZN(n5591) );
  NAND2_X1 U6216 ( .A1(n5969), .A2(n5968), .ZN(n5982) );
  OAI21_X1 U6217 ( .B1(n5946), .B2(n5945), .A(n5944), .ZN(n5964) );
  NAND2_X1 U6218 ( .A1(n5055), .A2(n5602), .ZN(n5793) );
  NAND2_X1 U6219 ( .A1(n5645), .A2(n5644), .ZN(n5886) );
  INV_X1 U6220 ( .A(n8517), .ZN(n5148) );
  INV_X1 U6221 ( .A(n8513), .ZN(n8480) );
  NAND3_X1 U6222 ( .A1(n5243), .A2(n5244), .A3(n5786), .ZN(n5055) );
  NAND2_X1 U6223 ( .A1(n5620), .A2(n5619), .ZN(n5854) );
  INV_X1 U6224 ( .A(n5146), .ZN(n8582) );
  NAND2_X1 U6225 ( .A1(n5929), .A2(n5928), .ZN(n5946) );
  NOR2_X1 U6226 ( .A1(n8479), .A2(n8478), .ZN(n8513) );
  NAND2_X1 U6227 ( .A1(n8516), .A2(n8515), .ZN(n5147) );
  NAND2_X1 U6228 ( .A1(n8085), .A2(n8084), .ZN(n8093) );
  OAI21_X1 U6229 ( .B1(n8308), .B2(n8306), .A(n8305), .ZN(n7720) );
  NAND4_X1 U6230 ( .A1(n10217), .A2(n10218), .A3(n10215), .A4(n10216), .ZN(
        n10308) );
  INV_X1 U6231 ( .A(n6162), .ZN(n5076) );
  NAND2_X1 U6232 ( .A1(n5222), .A2(n8351), .ZN(n7171) );
  INV_X1 U6233 ( .A(n7011), .ZN(n7008) );
  NAND2_X1 U6234 ( .A1(n8317), .A2(n7003), .ZN(n7011) );
  NAND2_X1 U6235 ( .A1(n6733), .A2(n10162), .ZN(n5229) );
  NAND2_X1 U6236 ( .A1(n5058), .A2(n6148), .ZN(n8497) );
  NAND2_X1 U6237 ( .A1(n10003), .A2(n10007), .ZN(n10002) );
  NAND2_X1 U6238 ( .A1(n5060), .A2(n5029), .ZN(n8319) );
  XNOR2_X1 U6239 ( .A(n5669), .B(n5668), .ZN(n6146) );
  INV_X1 U6240 ( .A(n7002), .ZN(n5060) );
  NAND2_X1 U6241 ( .A1(n9629), .A2(n8974), .ZN(n8981) );
  NAND2_X1 U6242 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5284) );
  NOR2_X1 U6243 ( .A1(n7124), .A2(n6314), .ZN(n7220) );
  NAND2_X1 U6244 ( .A1(n5202), .A2(n5201), .ZN(n6920) );
  INV_X1 U6245 ( .A(n5204), .ZN(n5203) );
  NOR2_X1 U6246 ( .A1(n9180), .A2(n9179), .ZN(n9199) );
  NOR2_X1 U6247 ( .A1(n7222), .A2(n7221), .ZN(n7348) );
  XNOR2_X1 U6248 ( .A(n7733), .B(n7749), .ZN(n7643) );
  NAND2_X1 U6249 ( .A1(n7202), .A2(n7201), .ZN(n9014) );
  OAI211_X2 U6250 ( .C1(n6775), .C2(n6319), .A(n6299), .B(n6298), .ZN(n9017)
         );
  NAND2_X1 U6251 ( .A1(n10114), .A2(n10115), .ZN(n6167) );
  NAND2_X1 U6252 ( .A1(n6166), .A2(n8408), .ZN(n10114) );
  NAND2_X1 U6253 ( .A1(n6151), .A2(n8528), .ZN(n7049) );
  INV_X1 U6254 ( .A(n10083), .ZN(n5058) );
  AND2_X2 U6255 ( .A1(n8497), .A2(n8492), .ZN(n10062) );
  INV_X1 U6256 ( .A(n6172), .ZN(n5513) );
  OAI21_X1 U6257 ( .B1(n6744), .B2(n10830), .A(n5047), .ZN(P1_U3550) );
  NAND2_X1 U6258 ( .A1(n7008), .A2(n7009), .ZN(n7256) );
  NAND2_X1 U6259 ( .A1(n5203), .A2(n6919), .ZN(n5202) );
  NAND2_X1 U6260 ( .A1(n9200), .A2(n5221), .ZN(n5219) );
  NAND2_X1 U6261 ( .A1(n9248), .A2(n5209), .ZN(n5207) );
  NOR2_X1 U6262 ( .A1(n7642), .A2(n7641), .ZN(n7733) );
  NAND2_X1 U6263 ( .A1(n7252), .A2(n7251), .ZN(n7253) );
  AOI21_X1 U6264 ( .B1(n7400), .B2(n7399), .A(n7398), .ZN(n9723) );
  NOR2_X2 U6265 ( .A1(n8879), .A2(n8878), .ZN(n9641) );
  NAND4_X1 U6266 ( .A1(n5751), .A2(n5748), .A3(n5747), .A4(n5752), .ZN(n5063)
         );
  NAND2_X1 U6267 ( .A1(n8339), .A2(n8522), .ZN(n7045) );
  NAND2_X1 U6268 ( .A1(n6167), .A2(n8415), .ZN(n10100) );
  NAND2_X1 U6269 ( .A1(n5223), .A2(n6152), .ZN(n7678) );
  NAND2_X1 U6270 ( .A1(n5065), .A2(n5064), .ZN(P2_U3154) );
  OAI211_X1 U6271 ( .C1(n8998), .C2(n8997), .A(n8996), .B(n9091), .ZN(n5065)
         );
  NAND2_X1 U6272 ( .A1(n7972), .A2(n8057), .ZN(n7976) );
  INV_X1 U6273 ( .A(n6681), .ZN(n6865) );
  XNOR2_X2 U6274 ( .A(n6724), .B(n8475), .ZN(n6733) );
  OAI21_X1 U6275 ( .B1(n8594), .B2(n8140), .A(n6667), .ZN(n5376) );
  INV_X1 U6276 ( .A(n5376), .ZN(n5375) );
  OAI21_X1 U6277 ( .B1(n5306), .B2(n5758), .A(n5764), .ZN(n5248) );
  NAND2_X1 U6278 ( .A1(n5611), .A2(n5610), .ZN(n5827) );
  NAND2_X1 U6279 ( .A1(n5386), .A2(n5385), .ZN(n5378) );
  NAND2_X1 U6280 ( .A1(n5316), .A2(n5321), .ZN(n5684) );
  NAND3_X1 U6281 ( .A1(n10716), .A2(n10718), .A3(n5032), .ZN(P2_U3200) );
  NOR2_X1 U6282 ( .A1(n7643), .A2(n6377), .ZN(n7734) );
  INV_X1 U6283 ( .A(n7348), .ZN(n5214) );
  INV_X1 U6284 ( .A(n7112), .ZN(n5206) );
  NAND2_X1 U6285 ( .A1(n5206), .A2(n5205), .ZN(n5204) );
  NOR2_X1 U6286 ( .A1(n7526), .A2(n7525), .ZN(n7642) );
  NOR2_X1 U6287 ( .A1(n7351), .A2(n6346), .ZN(n7523) );
  NOR2_X1 U6288 ( .A1(n9156), .A2(n9155), .ZN(n9180) );
  NOR2_X2 U6289 ( .A1(n8905), .A2(n8904), .ZN(n9753) );
  OAI21_X2 U6290 ( .B1(n7713), .B2(n7712), .A(n7711), .ZN(n8308) );
  INV_X1 U6291 ( .A(n5300), .ZN(n6179) );
  NOR2_X1 U6292 ( .A1(n7343), .A2(n7813), .ZN(n7538) );
  XNOR2_X1 U6293 ( .A(n7536), .B(n7537), .ZN(n7343) );
  NOR2_X1 U6294 ( .A1(n7631), .A2(n6376), .ZN(n7750) );
  AOI21_X2 U6295 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n9233), .A(n9232), .ZN(
        n9234) );
  NAND3_X1 U6296 ( .A1(n5267), .A2(n5266), .A3(n5271), .ZN(n5070) );
  NOR2_X2 U6297 ( .A1(n7629), .A2(n5072), .ZN(n7748) );
  NAND2_X2 U6298 ( .A1(n9042), .A2(n8629), .ZN(n9124) );
  NAND2_X1 U6299 ( .A1(n8020), .A2(n8019), .ZN(n5434) );
  NAND3_X1 U6300 ( .A1(n5080), .A2(n6212), .A3(n6213), .ZN(n5074) );
  NAND2_X1 U6301 ( .A1(n7975), .A2(n7976), .ZN(n8020) );
  NAND2_X1 U6302 ( .A1(n5429), .A2(n5432), .ZN(n8996) );
  NAND2_X1 U6303 ( .A1(n7678), .A2(n8533), .ZN(n5222) );
  NAND2_X1 U6304 ( .A1(n8451), .A2(n8450), .ZN(n5135) );
  NAND2_X1 U6305 ( .A1(n6168), .A2(n8435), .ZN(n6723) );
  INV_X1 U6306 ( .A(n7049), .ZN(n5223) );
  NAND3_X2 U6307 ( .A1(n5733), .A2(n5732), .A3(n4981), .ZN(n10193) );
  NAND3_X2 U6308 ( .A1(n6198), .A2(n6197), .A3(n6199), .ZN(n7028) );
  NAND2_X1 U6309 ( .A1(n5389), .A2(n5388), .ZN(n7713) );
  INV_X1 U6310 ( .A(n6100), .ZN(n5735) );
  AND3_X2 U6311 ( .A1(n5080), .A2(n6213), .A3(n5079), .ZN(n6233) );
  AND3_X1 U6312 ( .A1(n5083), .A2(n5084), .A3(n5081), .ZN(n6214) );
  AND2_X1 U6313 ( .A1(n6209), .A2(n6410), .ZN(n5081) );
  NOR2_X1 U6314 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5088) );
  NAND2_X1 U6315 ( .A1(n5089), .A2(n6284), .ZN(n7096) );
  NAND2_X1 U6316 ( .A1(n8011), .A2(n5034), .ZN(n5096) );
  NAND2_X1 U6317 ( .A1(n5103), .A2(n8009), .ZN(n8055) );
  NAND3_X1 U6318 ( .A1(n5131), .A2(n5130), .A3(n5129), .ZN(n5128) );
  NAND2_X1 U6319 ( .A1(n5133), .A2(n5233), .ZN(n5132) );
  NAND2_X1 U6320 ( .A1(n5134), .A2(n8393), .ZN(n5133) );
  NAND2_X1 U6321 ( .A1(n8395), .A2(n5250), .ZN(n5134) );
  NAND2_X2 U6322 ( .A1(n5135), .A2(n6149), .ZN(n8523) );
  XNOR2_X2 U6323 ( .A(n5745), .B(n5164), .ZN(n8451) );
  NAND2_X1 U6324 ( .A1(n5671), .A2(n5155), .ZN(n5156) );
  NOR2_X2 U6325 ( .A1(n5691), .A2(n5565), .ZN(n5685) );
  NAND3_X4 U6326 ( .A1(n4980), .A2(n5723), .A3(n5725), .ZN(n9807) );
  NAND2_X1 U6327 ( .A1(n10116), .A2(n5169), .ZN(n5168) );
  NAND2_X1 U6328 ( .A1(n5519), .A2(n5173), .ZN(n5542) );
  NAND2_X1 U6329 ( .A1(n5884), .A2(n10785), .ZN(n5180) );
  MUX2_X1 U6330 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n6269), .Z(n5598) );
  MUX2_X1 U6331 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n6269), .Z(n5601) );
  MUX2_X1 U6332 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6269), .Z(n5791) );
  MUX2_X1 U6333 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n6269), .Z(n5609) );
  MUX2_X1 U6334 ( .A(n5615), .B(n6799), .S(n6269), .Z(n5616) );
  MUX2_X1 U6335 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6269), .Z(n5613) );
  MUX2_X1 U6336 ( .A(n6810), .B(n6809), .S(n6269), .Z(n5622) );
  MUX2_X1 U6337 ( .A(n5632), .B(n5633), .S(n6269), .Z(n5635) );
  MUX2_X1 U6338 ( .A(n5627), .B(n6813), .S(n6771), .Z(n5628) );
  NAND3_X1 U6339 ( .A1(n8764), .A2(n8762), .A3(n8763), .ZN(n5191) );
  XNOR2_X1 U6340 ( .A(n8850), .B(n8849), .ZN(n5195) );
  OAI21_X1 U6341 ( .B1(n9181), .B2(n5220), .A(n5219), .ZN(n9224) );
  INV_X1 U6342 ( .A(n9203), .ZN(n5221) );
  OR2_X2 U6343 ( .A1(n7171), .A2(n8532), .ZN(n7324) );
  NAND2_X1 U6344 ( .A1(n6733), .A2(n5226), .ZN(n5224) );
  NAND2_X1 U6345 ( .A1(n5225), .A2(n5224), .ZN(P1_U3551) );
  INV_X1 U6346 ( .A(n6732), .ZN(n5231) );
  INV_X1 U6347 ( .A(n8393), .ZN(n5236) );
  AOI21_X2 U6348 ( .B1(n10002), .B2(n5240), .A(n5239), .ZN(n6168) );
  NAND2_X1 U6349 ( .A1(n5241), .A2(n5671), .ZN(n5662) );
  INV_X1 U6350 ( .A(n5248), .ZN(n5247) );
  NAND2_X1 U6351 ( .A1(n5248), .A2(n5599), .ZN(n5243) );
  NAND2_X1 U6352 ( .A1(n5246), .A2(n5599), .ZN(n5244) );
  NAND2_X1 U6353 ( .A1(n5245), .A2(n5599), .ZN(n5787) );
  NAND2_X1 U6354 ( .A1(n5247), .A2(n5304), .ZN(n5245) );
  INV_X1 U6355 ( .A(n5304), .ZN(n5246) );
  AND2_X1 U6356 ( .A1(n8372), .A2(n8540), .ZN(n5255) );
  MUX2_X1 U6357 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n6771), .Z(n5596) );
  NAND3_X1 U6358 ( .A1(n5259), .A2(n5257), .A3(n8415), .ZN(n8416) );
  NAND3_X1 U6359 ( .A1(n8410), .A2(n8411), .A3(n8558), .ZN(n5260) );
  NAND3_X1 U6360 ( .A1(n7151), .A2(P2_REG2_REG_3__SCAN_IN), .A3(n5265), .ZN(
        n7153) );
  NAND2_X1 U6361 ( .A1(n9234), .A2(n9246), .ZN(n5268) );
  OAI21_X1 U6362 ( .B1(n10700), .B2(P2_REG2_REG_18__SCAN_IN), .A(n10705), .ZN(
        n5266) );
  NAND3_X1 U6363 ( .A1(n5268), .A2(n5270), .A3(n4979), .ZN(n5267) );
  NAND2_X1 U6364 ( .A1(n10700), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6365 ( .A1(n7136), .A2(n4996), .ZN(n5274) );
  NAND2_X1 U6366 ( .A1(n5274), .A2(n5273), .ZN(n7342) );
  NOR2_X2 U6367 ( .A1(n7937), .A2(n5275), .ZN(n7939) );
  AND2_X2 U6368 ( .A1(n5277), .A2(n5276), .ZN(n7937) );
  OAI21_X1 U6369 ( .B1(n9192), .B2(n5282), .A(n5281), .ZN(n9232) );
  INV_X1 U6370 ( .A(n5289), .ZN(n10074) );
  INV_X1 U6371 ( .A(n7501), .ZN(n5291) );
  NAND2_X1 U6372 ( .A1(n5291), .A2(n5292), .ZN(n7899) );
  INV_X1 U6373 ( .A(n10138), .ZN(n10149) );
  NAND2_X1 U6374 ( .A1(n5303), .A2(n5597), .ZN(n5765) );
  NAND2_X1 U6375 ( .A1(n5758), .A2(n5757), .ZN(n5303) );
  NAND2_X1 U6376 ( .A1(n5305), .A2(n5597), .ZN(n5304) );
  INV_X1 U6377 ( .A(n5597), .ZN(n5306) );
  NAND2_X1 U6378 ( .A1(n5595), .A2(n5594), .ZN(n5758) );
  NAND2_X1 U6379 ( .A1(n5309), .A2(n5307), .ZN(n5620) );
  NAND2_X1 U6380 ( .A1(n5310), .A2(n5051), .ZN(n6035) );
  NAND2_X1 U6381 ( .A1(n5886), .A2(n5314), .ZN(n5311) );
  NAND2_X1 U6382 ( .A1(n5311), .A2(n5313), .ZN(n5912) );
  NAND2_X1 U6383 ( .A1(n5982), .A2(n5046), .ZN(n5999) );
  NAND2_X1 U6384 ( .A1(n5626), .A2(n5317), .ZN(n5316) );
  NAND2_X1 U6385 ( .A1(n5626), .A2(n5325), .ZN(n5319) );
  NAND2_X1 U6386 ( .A1(n6054), .A2(n5330), .ZN(n5329) );
  NAND3_X1 U6387 ( .A1(n10422), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n5342) );
  NAND3_X1 U6388 ( .A1(n5346), .A2(n5345), .A3(n5344), .ZN(n5343) );
  NAND2_X1 U6389 ( .A1(n9548), .A2(n5350), .ZN(n5347) );
  NAND2_X1 U6390 ( .A1(n5347), .A2(n5348), .ZN(n6638) );
  NAND3_X1 U6391 ( .A1(n6262), .A2(n6261), .A3(n8328), .ZN(n5354) );
  NAND2_X1 U6392 ( .A1(n6272), .A2(n5356), .ZN(n5357) );
  OAI211_X2 U6393 ( .C1(n6272), .C2(n5359), .A(n5358), .B(n5357), .ZN(n7359)
         );
  NAND2_X1 U6394 ( .A1(n7796), .A2(n4974), .ZN(n5360) );
  NAND2_X1 U6395 ( .A1(n5360), .A2(n5361), .ZN(n8011) );
  NAND3_X1 U6396 ( .A1(n7258), .A2(n5387), .A3(n7257), .ZN(n7268) );
  INV_X1 U6397 ( .A(n7261), .ZN(n5387) );
  XNOR2_X1 U6398 ( .A(n7266), .B(n7265), .ZN(n7261) );
  NAND2_X1 U6399 ( .A1(n9721), .A2(n5390), .ZN(n5389) );
  NOR2_X1 U6400 ( .A1(n5393), .A2(n5391), .ZN(n5390) );
  INV_X1 U6401 ( .A(n7407), .ZN(n5391) );
  NOR2_X1 U6402 ( .A1(n7411), .A2(n7437), .ZN(n5393) );
  OAI21_X2 U6403 ( .B1(n9692), .B2(n8890), .A(n5395), .ZN(n9700) );
  INV_X1 U6404 ( .A(n5403), .ZN(n8191) );
  OR2_X1 U6405 ( .A1(n8189), .A2(n8190), .ZN(n5402) );
  NAND2_X1 U6406 ( .A1(n5407), .A2(n5030), .ZN(n8939) );
  NAND2_X1 U6407 ( .A1(n9732), .A2(n5405), .ZN(n5407) );
  CLKBUF_X1 U6408 ( .A(n5407), .Z(n5404) );
  NAND2_X1 U6409 ( .A1(n5685), .A2(n5037), .ZN(n5930) );
  NAND2_X1 U6410 ( .A1(n4965), .A2(n7668), .ZN(n7883) );
  NAND2_X1 U6411 ( .A1(n4965), .A2(n5036), .ZN(n5417) );
  NAND2_X1 U6412 ( .A1(n9124), .A2(n5423), .ZN(n5422) );
  OAI211_X1 U6413 ( .C1(n9124), .C2(n5428), .A(n5424), .B(n5422), .ZN(n8642)
         );
  NAND2_X1 U6414 ( .A1(n9124), .A2(n9121), .ZN(n5429) );
  OAI21_X1 U6415 ( .B1(n9124), .B2(n9120), .A(n9121), .ZN(n8998) );
  OAI21_X2 U6416 ( .B1(n7511), .B2(n5052), .A(n5435), .ZN(n7665) );
  OAI21_X1 U6417 ( .B1(n9078), .B2(n5439), .A(n9077), .ZN(n9079) );
  OAI21_X2 U6418 ( .B1(n8270), .B2(n5442), .A(n5440), .ZN(n9059) );
  NAND3_X1 U6419 ( .A1(n6214), .A2(n6213), .A3(n6212), .ZN(n6496) );
  OAI21_X1 U6420 ( .B1(n9433), .B2(n5450), .A(n5447), .ZN(n9397) );
  NAND2_X1 U6421 ( .A1(n5446), .A2(n5445), .ZN(n9399) );
  NAND2_X1 U6422 ( .A1(n9433), .A2(n5447), .ZN(n5446) );
  NAND2_X1 U6423 ( .A1(n5451), .A2(n5452), .ZN(n9435) );
  NAND2_X1 U6424 ( .A1(n9454), .A2(n6481), .ZN(n5451) );
  OAI21_X1 U6425 ( .B1(n8132), .B2(n5461), .A(n5458), .ZN(n9558) );
  NAND2_X1 U6426 ( .A1(n5457), .A2(n5455), .ZN(n6452) );
  NAND2_X1 U6427 ( .A1(n8132), .A2(n5458), .ZN(n5457) );
  NAND2_X1 U6428 ( .A1(n7387), .A2(n5468), .ZN(n5464) );
  NAND2_X1 U6429 ( .A1(n5464), .A2(n5466), .ZN(n7770) );
  NAND2_X1 U6430 ( .A1(n6366), .A2(n5027), .ZN(n5473) );
  INV_X1 U6431 ( .A(n9297), .ZN(n5492) );
  AND2_X1 U6432 ( .A1(n6233), .A2(n5493), .ZN(n6238) );
  NAND2_X1 U6433 ( .A1(n6215), .A2(n5494), .ZN(n6240) );
  OAI21_X2 U6434 ( .B1(n9341), .B2(n5500), .A(n5498), .ZN(n9307) );
  NAND3_X1 U6435 ( .A1(n5502), .A2(n5503), .A3(n5501), .ZN(n5499) );
  INV_X1 U6436 ( .A(n9316), .ZN(n5509) );
  NAND3_X1 U6437 ( .A1(n5754), .A2(n5511), .A3(n5560), .ZN(n5691) );
  NAND2_X1 U6438 ( .A1(n7556), .A2(n5515), .ZN(n10780) );
  OR2_X1 U6439 ( .A1(n7969), .A2(n9798), .ZN(n5515) );
  NAND2_X1 U6440 ( .A1(n10066), .A2(n5520), .ZN(n5519) );
  NAND2_X1 U6441 ( .A1(n7323), .A2(n5523), .ZN(n5524) );
  AND2_X1 U6442 ( .A1(n8358), .A2(n8359), .ZN(n5523) );
  NAND2_X1 U6443 ( .A1(n10170), .A2(n5531), .ZN(n5530) );
  AOI21_X1 U6444 ( .B1(n10170), .B2(n6165), .A(n5538), .ZN(n10148) );
  AND2_X1 U6445 ( .A1(n8621), .A2(n8620), .ZN(n8622) );
  XNOR2_X1 U6446 ( .A(n7096), .B(n4967), .ZN(n7198) );
  INV_X1 U6447 ( .A(n8600), .ZN(n7292) );
  NAND2_X1 U6448 ( .A1(n5952), .A2(n5951), .ZN(n5953) );
  XNOR2_X1 U6449 ( .A(n6130), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6136) );
  AOI21_X1 U6450 ( .B1(n6130), .B2(n6125), .A(n6124), .ZN(n6128) );
  NOR2_X2 U6451 ( .A1(n10140), .A2(n10125), .ZN(n10120) );
  OR2_X1 U6452 ( .A1(n8649), .A2(n6917), .ZN(n6277) );
  OR2_X1 U6453 ( .A1(n6436), .A2(n7193), .ZN(n6267) );
  INV_X1 U6454 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5730) );
  AOI21_X1 U6455 ( .B1(n9989), .B2(n9996), .A(n9988), .ZN(n10211) );
  OR2_X1 U6456 ( .A1(n9150), .A2(n7096), .ZN(n6629) );
  AOI21_X2 U6457 ( .B1(n9070), .B2(n9069), .A(n9068), .ZN(n9072) );
  INV_X1 U6458 ( .A(n10340), .ZN(n6205) );
  OR2_X1 U6459 ( .A1(n7276), .A2(n9805), .ZN(n5546) );
  OR2_X1 U6460 ( .A1(n7706), .A2(n9806), .ZN(n5547) );
  AND2_X1 U6461 ( .A1(n7219), .A2(n7224), .ZN(n5548) );
  OR2_X1 U6462 ( .A1(n5301), .A2(n10298), .ZN(n5549) );
  AND3_X1 U6463 ( .A1(n6218), .A2(n6222), .A3(n6226), .ZN(n5550) );
  AND2_X1 U6464 ( .A1(n9233), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5551) );
  OR2_X1 U6465 ( .A1(n10341), .A2(n9695), .ZN(n5552) );
  AND2_X1 U6466 ( .A1(n5625), .A2(n5624), .ZN(n5553) );
  NAND2_X1 U6467 ( .A1(n9387), .A2(n9386), .ZN(n5554) );
  NAND2_X1 U6468 ( .A1(n6575), .A2(n6574), .ZN(n9138) );
  NOR2_X1 U6469 ( .A1(n4986), .A2(n6065), .ZN(n5555) );
  INV_X1 U6470 ( .A(n5666), .ZN(n5580) );
  INV_X1 U6471 ( .A(n7960), .ZN(n7958) );
  INV_X1 U6472 ( .A(n9022), .ZN(n8608) );
  NAND2_X1 U6473 ( .A1(n6922), .A2(n6917), .ZN(n6918) );
  INV_X1 U6474 ( .A(n6434), .ZN(n6433) );
  INV_X1 U6475 ( .A(n6349), .ZN(n6348) );
  INV_X1 U6476 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6294) );
  OR2_X1 U6477 ( .A1(n8507), .A2(n8573), .ZN(n8478) );
  NOR2_X1 U6478 ( .A1(n5958), .A2(n5957), .ZN(n5972) );
  OR2_X1 U6479 ( .A1(n6025), .A2(n9659), .ZN(n6042) );
  NOR2_X1 U6480 ( .A1(n5892), .A2(n5891), .ZN(n5890) );
  INV_X1 U6481 ( .A(n9807), .ZN(n5745) );
  INV_X1 U6482 ( .A(n5683), .ZN(n5642) );
  INV_X1 U6483 ( .A(n5826), .ZN(n5612) );
  XNOR2_X1 U6484 ( .A(n4966), .B(n7359), .ZN(n6880) );
  NAND2_X1 U6485 ( .A1(n8608), .A2(n9113), .ZN(n8609) );
  NAND2_X1 U6486 ( .A1(n6490), .A2(n10457), .ZN(n6502) );
  INV_X1 U6487 ( .A(n8250), .ZN(n8246) );
  NOR2_X1 U6488 ( .A1(n7539), .A2(n7538), .ZN(n7542) );
  NOR2_X1 U6489 ( .A1(n9318), .A2(n9329), .ZN(n8832) );
  INV_X1 U6490 ( .A(n8607), .ZN(n9403) );
  INV_X1 U6491 ( .A(n9146), .ZN(n7483) );
  AND2_X1 U6492 ( .A1(n8736), .A2(n8751), .ZN(n8668) );
  INV_X1 U6493 ( .A(n8713), .ZN(n6273) );
  NAND2_X1 U6494 ( .A1(n5985), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6002) );
  NOR2_X1 U6495 ( .A1(n6042), .A2(n9716), .ZN(n6057) );
  OR2_X1 U6496 ( .A1(n6002), .A2(n9746), .ZN(n6025) );
  OR2_X1 U6497 ( .A1(n5862), .A2(n5707), .ZN(n5871) );
  INV_X1 U6498 ( .A(n6102), .ZN(n6114) );
  OR2_X1 U6499 ( .A1(n8313), .A2(n9801), .ZN(n5841) );
  OR2_X1 U6500 ( .A1(n7689), .A2(n9803), .ZN(n5807) );
  AND2_X1 U6501 ( .A1(n8481), .A2(n6136), .ZN(n7016) );
  OR2_X1 U6502 ( .A1(n8280), .A2(n8279), .ZN(n8281) );
  NAND2_X1 U6503 ( .A1(n5647), .A2(n10504), .ZN(n5650) );
  NAND2_X1 U6504 ( .A1(n5635), .A2(n5634), .ZN(n5638) );
  INV_X1 U6505 ( .A(n9144), .ZN(n7673) );
  NAND2_X1 U6506 ( .A1(n8628), .A2(n9329), .ZN(n8629) );
  NAND2_X1 U6507 ( .A1(n6460), .A2(n8272), .ZN(n6475) );
  NOR2_X1 U6508 ( .A1(n8645), .A2(n6246), .ZN(n6247) );
  INV_X1 U6509 ( .A(n9138), .ZN(n9329) );
  AND2_X1 U6510 ( .A1(n6529), .A2(n6528), .ZN(n9407) );
  OR2_X1 U6511 ( .A1(n8144), .A2(n9142), .ZN(n8009) );
  OR2_X1 U6512 ( .A1(n9561), .A2(n6760), .ZN(n6761) );
  AND2_X1 U6513 ( .A1(n8807), .A2(n8808), .ZN(n9421) );
  INV_X1 U6514 ( .A(n9143), .ZN(n8013) );
  AND2_X1 U6515 ( .A1(n8746), .A2(n8733), .ZN(n8665) );
  INV_X1 U6516 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6222) );
  NAND2_X1 U6517 ( .A1(n6282), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6283) );
  NOR2_X1 U6518 ( .A1(n9654), .A2(n9653), .ZN(n9743) );
  CLKBUF_X3 U6519 ( .A(n5735), .Z(n6727) );
  OR2_X1 U6520 ( .A1(n6947), .A2(n6948), .ZN(n7081) );
  INV_X1 U6521 ( .A(n9799), .ZN(n7966) );
  INV_X1 U6522 ( .A(n6734), .ZN(n6747) );
  XNOR2_X1 U6523 ( .A(n9649), .B(n9782), .ZN(n8466) );
  INV_X1 U6524 ( .A(n9800), .ZN(n8373) );
  NAND2_X1 U6525 ( .A1(n7059), .A2(n5746), .ZN(n7703) );
  AND2_X1 U6526 ( .A1(n6202), .A2(n6827), .ZN(n7571) );
  OAI21_X1 U6527 ( .B1(n5964), .B2(n5963), .A(n5962), .ZN(n5969) );
  XNOR2_X1 U6528 ( .A(n5643), .B(SI_13_), .ZN(n5683) );
  AND2_X1 U6529 ( .A1(n6860), .A2(n6861), .ZN(n9081) );
  OR2_X1 U6530 ( .A1(n6436), .A2(n8588), .ZN(n8653) );
  AOI21_X1 U6531 ( .B1(n9332), .B2(n6458), .A(n6565), .ZN(n9316) );
  AND4_X1 U6532 ( .A1(n6440), .A2(n6439), .A3(n6438), .A4(n6437), .ZN(n8239)
         );
  AND4_X1 U6533 ( .A1(n6397), .A2(n6396), .A3(n6395), .A4(n6394), .ZN(n8057)
         );
  OR2_X1 U6534 ( .A1(n6436), .A2(n7872), .ZN(n6335) );
  NAND2_X1 U6535 ( .A1(n6857), .A2(n8859), .ZN(n10838) );
  INV_X1 U6536 ( .A(n9360), .ZN(n10768) );
  AND2_X1 U6537 ( .A1(n10846), .A2(n10844), .ZN(n9377) );
  AND2_X1 U6538 ( .A1(n8092), .A2(n8091), .ZN(n8190) );
  OR2_X1 U6539 ( .A1(n6975), .A2(n6944), .ZN(n9906) );
  AND2_X1 U6540 ( .A1(n8488), .A2(n8495), .ZN(n10026) );
  NAND2_X1 U6541 ( .A1(n8418), .A2(n10082), .ZN(n10101) );
  NAND2_X1 U6542 ( .A1(n8411), .A2(n8415), .ZN(n10113) );
  NAND2_X1 U6543 ( .A1(n8518), .A2(n8400), .ZN(n8467) );
  AND2_X1 U6544 ( .A1(n10723), .A2(n8577), .ZN(n10283) );
  AND2_X1 U6545 ( .A1(n6183), .A2(n6182), .ZN(n7014) );
  AND2_X1 U6546 ( .A1(n5719), .A2(n5880), .ZN(n7309) );
  XNOR2_X1 U6547 ( .A(n5598), .B(n10411), .ZN(n5764) );
  INV_X1 U6548 ( .A(n9131), .ZN(n9114) );
  NAND2_X1 U6549 ( .A1(n6584), .A2(n6583), .ZN(n9137) );
  INV_X1 U6550 ( .A(n8057), .ZN(n9142) );
  INV_X1 U6551 ( .A(n7384), .ZN(n9149) );
  OAI21_X1 U6552 ( .B1(n10715), .B2(n10714), .A(n10661), .ZN(n10716) );
  INV_X1 U6553 ( .A(n9377), .ZN(n9479) );
  INV_X1 U6554 ( .A(n9561), .ZN(n9570) );
  INV_X1 U6555 ( .A(n8632), .ZN(n9581) );
  INV_X1 U6556 ( .A(n10852), .ZN(n10850) );
  AND2_X1 U6557 ( .A1(n6685), .A2(n6684), .ZN(n9612) );
  INV_X1 U6558 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6813) );
  INV_X1 U6559 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6799) );
  INV_X1 U6560 ( .A(n8188), .ZN(n10825) );
  AND4_X1 U6561 ( .A1(n6145), .A2(n6144), .A3(n6143), .A4(n6142), .ZN(n9979)
         );
  AND2_X1 U6562 ( .A1(n7083), .A2(n7082), .ZN(n7308) );
  INV_X1 U6563 ( .A(n10831), .ZN(n10830) );
  INV_X1 U6564 ( .A(n10834), .ZN(n6207) );
  INV_X1 U6565 ( .A(n10091), .ZN(n10319) );
  INV_X1 U6566 ( .A(n7019), .ZN(n7023) );
  NAND2_X1 U6567 ( .A1(n5832), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5860) );
  INV_X1 U6568 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5859) );
  INV_X1 U6569 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5707) );
  INV_X1 U6570 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U6571 ( .A1(n5700), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5702) );
  INV_X1 U6572 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5676) );
  INV_X1 U6573 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5891) );
  AND2_X1 U6574 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n5556) );
  INV_X1 U6575 ( .A(n5557), .ZN(n5920) );
  INV_X1 U6576 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U6577 ( .A1(n5920), .A2(n5558), .ZN(n5559) );
  NAND2_X1 U6578 ( .A1(n5935), .A2(n5559), .ZN(n10150) );
  NOR2_X1 U6579 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5564) );
  NAND4_X1 U6580 ( .A1(n5564), .A2(n5563), .A3(n5562), .A4(n5561), .ZN(n5565)
         );
  NOR2_X1 U6581 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n6174) );
  NOR2_X1 U6582 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5569) );
  NOR2_X1 U6583 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5568) );
  INV_X1 U6584 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5567) );
  NAND4_X1 U6585 ( .A1(n6174), .A2(n5569), .A3(n5568), .A4(n5567), .ZN(n5574)
         );
  INV_X1 U6586 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5572) );
  INV_X1 U6587 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5571) );
  INV_X1 U6588 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5570) );
  NAND4_X1 U6589 ( .A1(n6195), .A2(n5572), .A3(n5571), .A4(n5570), .ZN(n5573)
         );
  NOR2_X1 U6590 ( .A1(n5574), .A2(n5573), .ZN(n5575) );
  NOR2_X1 U6591 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5579) );
  INV_X1 U6592 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U6593 ( .A1(n5579), .A2(n5576), .ZN(n5577) );
  INV_X1 U6594 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10342) );
  NAND2_X4 U6595 ( .A1(n5582), .A2(n5584), .ZN(n6140) );
  OR2_X1 U6596 ( .A1(n10150), .A2(n6140), .ZN(n5588) );
  NAND2_X1 U6597 ( .A1(n6113), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U6598 ( .A1(n8292), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U6599 ( .A1(n8991), .A2(n10352), .ZN(n5750) );
  INV_X2 U6600 ( .A(n8294), .ZN(n6139) );
  NAND2_X1 U6601 ( .A1(n6139), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5585) );
  NAND4_X1 U6602 ( .A1(n5588), .A2(n5587), .A3(n5586), .A4(n5585), .ZN(n10266)
         );
  INV_X2 U6603 ( .A(n5591), .ZN(n6269) );
  INV_X1 U6604 ( .A(SI_2_), .ZN(n10522) );
  AND2_X1 U6605 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U6606 ( .A1(n5591), .A2(n5589), .ZN(n5743) );
  NAND3_X1 U6607 ( .A1(n6269), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n5590) );
  NAND2_X1 U6608 ( .A1(n5743), .A2(n5590), .ZN(n5728) );
  MUX2_X1 U6609 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5591), .Z(n5593) );
  INV_X1 U6610 ( .A(SI_1_), .ZN(n5592) );
  XNOR2_X1 U6611 ( .A(n5593), .B(n5592), .ZN(n5727) );
  NAND2_X1 U6612 ( .A1(n5728), .A2(n5727), .ZN(n5595) );
  NAND2_X1 U6613 ( .A1(n5593), .A2(SI_1_), .ZN(n5594) );
  NAND2_X1 U6614 ( .A1(n5596), .A2(SI_2_), .ZN(n5597) );
  NAND2_X1 U6615 ( .A1(n5598), .A2(SI_3_), .ZN(n5599) );
  INV_X1 U6616 ( .A(SI_4_), .ZN(n5600) );
  NAND2_X1 U6617 ( .A1(n5601), .A2(SI_4_), .ZN(n5602) );
  INV_X1 U6618 ( .A(n5791), .ZN(n5604) );
  INV_X1 U6619 ( .A(SI_5_), .ZN(n5603) );
  NAND2_X1 U6620 ( .A1(n5604), .A2(n5603), .ZN(n5605) );
  NAND2_X1 U6621 ( .A1(n5793), .A2(n5605), .ZN(n5607) );
  NAND2_X1 U6622 ( .A1(n5791), .A2(SI_5_), .ZN(n5606) );
  NAND2_X1 U6623 ( .A1(n5607), .A2(n5606), .ZN(n5809) );
  NAND2_X1 U6624 ( .A1(n5809), .A2(n5608), .ZN(n5611) );
  NAND2_X1 U6625 ( .A1(n5609), .A2(SI_6_), .ZN(n5610) );
  NAND2_X1 U6626 ( .A1(n5613), .A2(SI_7_), .ZN(n5614) );
  INV_X1 U6627 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5615) );
  INV_X1 U6628 ( .A(SI_8_), .ZN(n10374) );
  INV_X1 U6629 ( .A(n5616), .ZN(n5617) );
  NAND2_X1 U6630 ( .A1(n5617), .A2(SI_8_), .ZN(n5618) );
  INV_X1 U6631 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6810) );
  INV_X1 U6632 ( .A(SI_9_), .ZN(n5621) );
  INV_X1 U6633 ( .A(n5622), .ZN(n5623) );
  NAND2_X1 U6634 ( .A1(n5623), .A2(SI_9_), .ZN(n5624) );
  INV_X1 U6635 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5627) );
  INV_X1 U6636 ( .A(n5628), .ZN(n5629) );
  INV_X1 U6637 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5633) );
  INV_X1 U6638 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5632) );
  INV_X1 U6639 ( .A(SI_11_), .ZN(n5634) );
  INV_X1 U6640 ( .A(n5635), .ZN(n5636) );
  NAND2_X1 U6641 ( .A1(n5636), .A2(SI_11_), .ZN(n5637) );
  MUX2_X1 U6642 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n8328), .Z(n5639) );
  INV_X1 U6643 ( .A(SI_12_), .ZN(n10393) );
  NAND2_X1 U6644 ( .A1(n5639), .A2(SI_12_), .ZN(n5640) );
  MUX2_X1 U6645 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n8328), .Z(n5643) );
  NAND2_X1 U6646 ( .A1(n5684), .A2(n5642), .ZN(n5645) );
  NAND2_X1 U6647 ( .A1(n5643), .A2(SI_13_), .ZN(n5644) );
  INV_X1 U6648 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6989) );
  INV_X1 U6649 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5646) );
  MUX2_X1 U6650 ( .A(n6989), .B(n5646), .S(n8328), .Z(n5647) );
  INV_X1 U6651 ( .A(SI_14_), .ZN(n10504) );
  INV_X1 U6652 ( .A(n5647), .ZN(n5648) );
  NAND2_X1 U6653 ( .A1(n5648), .A2(SI_14_), .ZN(n5649) );
  NAND2_X1 U6654 ( .A1(n5650), .A2(n5649), .ZN(n5885) );
  MUX2_X1 U6655 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n8328), .Z(n5652) );
  INV_X1 U6656 ( .A(SI_15_), .ZN(n5651) );
  XNOR2_X1 U6657 ( .A(n5652), .B(n5651), .ZN(n5899) );
  INV_X1 U6658 ( .A(n5899), .ZN(n5653) );
  INV_X1 U6659 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7321) );
  INV_X1 U6660 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7319) );
  MUX2_X1 U6661 ( .A(n7321), .B(n7319), .S(n8328), .Z(n5655) );
  INV_X1 U6662 ( .A(SI_16_), .ZN(n5654) );
  NAND2_X1 U6663 ( .A1(n5655), .A2(n5654), .ZN(n5658) );
  INV_X1 U6664 ( .A(n5655), .ZN(n5656) );
  NAND2_X1 U6665 ( .A1(n5656), .A2(SI_16_), .ZN(n5657) );
  NAND2_X1 U6666 ( .A1(n5658), .A2(n5657), .ZN(n5911) );
  INV_X1 U6667 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7366) );
  INV_X1 U6668 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7368) );
  MUX2_X1 U6669 ( .A(n7366), .B(n7368), .S(n8328), .Z(n5659) );
  INV_X1 U6670 ( .A(SI_17_), .ZN(n10500) );
  NAND2_X1 U6671 ( .A1(n5659), .A2(n10500), .ZN(n5928) );
  INV_X1 U6672 ( .A(n5659), .ZN(n5660) );
  NAND2_X1 U6673 ( .A1(n5660), .A2(SI_17_), .ZN(n5661) );
  XNOR2_X1 U6674 ( .A(n5927), .B(n5926), .ZN(n7365) );
  NAND2_X1 U6675 ( .A1(n5662), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5663) );
  INV_X1 U6676 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5665) );
  INV_X1 U6677 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U6678 ( .A1(n5731), .A2(n8328), .ZN(n5766) );
  NAND2_X1 U6679 ( .A1(n7365), .A2(n8333), .ZN(n5674) );
  NAND2_X1 U6680 ( .A1(n5731), .A2(n6771), .ZN(n5767) );
  INV_X1 U6681 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U6682 ( .A1(n5930), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5672) );
  XNOR2_X1 U6683 ( .A(n5672), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9922) );
  AOI22_X1 U6684 ( .A1(n8332), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5954), .B2(
        n9922), .ZN(n5673) );
  NAND2_X1 U6685 ( .A1(n6113), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5682) );
  INV_X1 U6686 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n5675) );
  OR2_X1 U6687 ( .A1(n6141), .A2(n5675), .ZN(n5681) );
  NAND2_X1 U6688 ( .A1(n5702), .A2(n5676), .ZN(n5677) );
  NAND2_X1 U6689 ( .A1(n5892), .A2(n5677), .ZN(n8222) );
  OR2_X1 U6690 ( .A1(n6140), .A2(n8222), .ZN(n5680) );
  INV_X1 U6691 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5678) );
  OR2_X1 U6692 ( .A1(n8294), .A2(n5678), .ZN(n5679) );
  NAND4_X1 U6693 ( .A1(n5682), .A2(n5681), .A3(n5680), .A4(n5679), .ZN(n9795)
         );
  INV_X1 U6694 ( .A(n9795), .ZN(n9646) );
  XNOR2_X1 U6695 ( .A(n5684), .B(n5683), .ZN(n6898) );
  NAND2_X1 U6696 ( .A1(n6898), .A2(n8333), .ZN(n5688) );
  OR2_X1 U6697 ( .A1(n5685), .A2(n6124), .ZN(n5686) );
  XNOR2_X1 U6698 ( .A(n5686), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7823) );
  AOI22_X1 U6699 ( .A1(n8332), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5954), .B2(
        n7823), .ZN(n5687) );
  INV_X1 U6700 ( .A(n8213), .ZN(n8227) );
  XNOR2_X1 U6701 ( .A(n5690), .B(n5689), .ZN(n6893) );
  NAND2_X1 U6702 ( .A1(n6893), .A2(n8333), .ZN(n5698) );
  NOR2_X1 U6703 ( .A1(n5692), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5810) );
  NOR2_X1 U6704 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5693) );
  NAND2_X1 U6705 ( .A1(n5810), .A2(n5693), .ZN(n5843) );
  INV_X1 U6706 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5717) );
  INV_X1 U6707 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U6708 ( .A1(n5717), .A2(n5694), .ZN(n5695) );
  OAI21_X1 U6709 ( .B1(n5715), .B2(n5695), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5696) );
  XNOR2_X1 U6710 ( .A(n5696), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7621) );
  AOI22_X1 U6711 ( .A1(n8332), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5954), .B2(
        n7621), .ZN(n5697) );
  NAND2_X1 U6712 ( .A1(n6139), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5706) );
  INV_X1 U6713 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7835) );
  OR2_X1 U6714 ( .A1(n6727), .A2(n7835), .ZN(n5705) );
  INV_X1 U6715 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5699) );
  OR2_X1 U6716 ( .A1(n6141), .A2(n5699), .ZN(n5704) );
  INV_X1 U6717 ( .A(n5700), .ZN(n5873) );
  INV_X1 U6718 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7426) );
  NAND2_X1 U6719 ( .A1(n5873), .A2(n7426), .ZN(n5701) );
  NAND2_X1 U6720 ( .A1(n5702), .A2(n5701), .ZN(n8194) );
  OR2_X1 U6721 ( .A1(n6140), .A2(n8194), .ZN(n5703) );
  NAND4_X1 U6722 ( .A1(n5706), .A2(n5705), .A3(n5704), .A4(n5703), .ZN(n9796)
         );
  INV_X1 U6723 ( .A(n9796), .ZN(n10795) );
  NAND2_X1 U6724 ( .A1(n6139), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5712) );
  INV_X1 U6725 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7590) );
  OR2_X1 U6726 ( .A1(n6727), .A2(n7590), .ZN(n5711) );
  NAND2_X1 U6727 ( .A1(n5862), .A2(n5707), .ZN(n5708) );
  NAND2_X1 U6728 ( .A1(n5871), .A2(n5708), .ZN(n7965) );
  OR2_X1 U6729 ( .A1(n6140), .A2(n7965), .ZN(n5710) );
  INV_X1 U6730 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7084) );
  OR2_X1 U6731 ( .A1(n6141), .A2(n7084), .ZN(n5709) );
  NAND4_X1 U6732 ( .A1(n5712), .A2(n5711), .A3(n5710), .A4(n5709), .ZN(n9798)
         );
  XNOR2_X1 U6733 ( .A(n5714), .B(n5713), .ZN(n6806) );
  NAND2_X1 U6734 ( .A1(n6806), .A2(n8333), .ZN(n5721) );
  NAND2_X1 U6735 ( .A1(n5715), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5718) );
  INV_X1 U6736 ( .A(n5718), .ZN(n5716) );
  NAND2_X1 U6737 ( .A1(n5716), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U6738 ( .A1(n5718), .A2(n5717), .ZN(n5880) );
  AOI22_X1 U6739 ( .A1(n8332), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5954), .B2(
        n7309), .ZN(n5720) );
  INV_X1 U6740 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10190) );
  INV_X1 U6741 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6950) );
  INV_X1 U6742 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5722) );
  OR2_X1 U6743 ( .A1(n5750), .A2(n5722), .ZN(n5723) );
  XNOR2_X1 U6744 ( .A(n5727), .B(n5728), .ZN(n6783) );
  OR2_X1 U6745 ( .A1(n5766), .A2(n6783), .ZN(n5733) );
  INV_X1 U6746 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6784) );
  OR2_X1 U6747 ( .A1(n5767), .A2(n6784), .ZN(n5732) );
  NAND2_X1 U6748 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5729) );
  XNOR2_X1 U6749 ( .A(n5730), .B(n5729), .ZN(n6949) );
  NAND2_X1 U6750 ( .A1(n8292), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5740) );
  INV_X1 U6751 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10728) );
  OR2_X1 U6752 ( .A1(n6140), .A2(n10728), .ZN(n5739) );
  INV_X1 U6753 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5734) );
  OR2_X1 U6754 ( .A1(n5735), .A2(n5734), .ZN(n5738) );
  INV_X1 U6755 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5736) );
  OR2_X1 U6756 ( .A1(n5750), .A2(n5736), .ZN(n5737) );
  NAND2_X1 U6757 ( .A1(n8328), .A2(SI_0_), .ZN(n5742) );
  INV_X1 U6758 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5741) );
  NAND2_X1 U6759 ( .A1(n5742), .A2(n5741), .ZN(n5744) );
  AND2_X1 U6760 ( .A1(n5744), .A2(n5743), .ZN(n10355) );
  NAND2_X1 U6761 ( .A1(n5056), .A2(n10722), .ZN(n7060) );
  INV_X1 U6762 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6952) );
  OR2_X1 U6763 ( .A1(n5771), .A2(n6952), .ZN(n5748) );
  NAND2_X1 U6764 ( .A1(n6100), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5747) );
  INV_X1 U6765 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9825) );
  OR2_X1 U6766 ( .A1(n6140), .A2(n9825), .ZN(n5752) );
  INV_X1 U6767 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5749) );
  OR2_X1 U6768 ( .A1(n5750), .A2(n5749), .ZN(n5751) );
  OR2_X1 U6769 ( .A1(n5754), .A2(n6124), .ZN(n5756) );
  INV_X1 U6770 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5755) );
  NAND2_X1 U6771 ( .A1(n5756), .A2(n5755), .ZN(n5761) );
  OAI21_X1 U6772 ( .B1(n5756), .B2(n5755), .A(n5761), .ZN(n6951) );
  XNOR2_X1 U6773 ( .A(n5758), .B(n5757), .ZN(n6782) );
  OR2_X1 U6774 ( .A1(n5766), .A2(n6782), .ZN(n5760) );
  INV_X1 U6775 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6781) );
  OR2_X1 U6776 ( .A1(n5767), .A2(n6781), .ZN(n5759) );
  OAI211_X2 U6777 ( .C1(n6815), .C2(n6951), .A(n5760), .B(n5759), .ZN(n7706)
         );
  NAND2_X1 U6778 ( .A1(n10186), .A2(n7706), .ZN(n8522) );
  NAND2_X1 U6779 ( .A1(n10743), .A2(n9806), .ZN(n8340) );
  NAND2_X1 U6780 ( .A1(n7703), .A2(n8342), .ZN(n7702) );
  NAND2_X1 U6781 ( .A1(n7702), .A2(n5547), .ZN(n7043) );
  NAND2_X1 U6782 ( .A1(n5761), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5763) );
  INV_X1 U6783 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5762) );
  XNOR2_X1 U6784 ( .A(n5763), .B(n5762), .ZN(n6953) );
  XNOR2_X1 U6785 ( .A(n5765), .B(n5764), .ZN(n6775) );
  OR2_X1 U6786 ( .A1(n5766), .A2(n6775), .ZN(n5769) );
  INV_X1 U6787 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6770) );
  OR2_X1 U6788 ( .A1(n5767), .A2(n6770), .ZN(n5768) );
  INV_X1 U6789 ( .A(n7276), .ZN(n7765) );
  INV_X1 U6790 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5770) );
  OR2_X2 U6791 ( .A1(n6727), .A2(n5770), .ZN(n5776) );
  OR2_X1 U6792 ( .A1(n6140), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5775) );
  INV_X1 U6793 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6954) );
  OR2_X1 U6794 ( .A1(n5771), .A2(n6954), .ZN(n5774) );
  INV_X1 U6795 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5772) );
  OR2_X1 U6796 ( .A1(n8294), .A2(n5772), .ZN(n5773) );
  NAND2_X1 U6797 ( .A1(n7765), .A2(n9805), .ZN(n8341) );
  NAND2_X1 U6798 ( .A1(n7657), .A2(n7276), .ZN(n8528) );
  NAND2_X1 U6799 ( .A1(n7043), .A2(n8453), .ZN(n7042) );
  NAND2_X1 U6800 ( .A1(n7042), .A2(n5546), .ZN(n7051) );
  NAND2_X1 U6801 ( .A1(n6139), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5782) );
  INV_X1 U6802 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5777) );
  OR2_X1 U6803 ( .A1(n6727), .A2(n5777), .ZN(n5781) );
  XNOR2_X1 U6804 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n9724) );
  OR2_X1 U6805 ( .A1(n6140), .A2(n9724), .ZN(n5780) );
  INV_X1 U6806 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5778) );
  OR2_X1 U6807 ( .A1(n6141), .A2(n5778), .ZN(n5779) );
  NAND4_X1 U6808 ( .A1(n5782), .A2(n5781), .A3(n5780), .A4(n5779), .ZN(n9804)
         );
  INV_X1 U6809 ( .A(n9804), .ZN(n7415) );
  NAND2_X1 U6810 ( .A1(n5783), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5784) );
  MUX2_X1 U6811 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5784), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5785) );
  NAND2_X1 U6812 ( .A1(n5785), .A2(n5692), .ZN(n9852) );
  XNOR2_X1 U6813 ( .A(n5787), .B(n5786), .ZN(n6780) );
  OR2_X1 U6814 ( .A1(n5766), .A2(n6780), .ZN(n5789) );
  INV_X1 U6815 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6779) );
  OR2_X1 U6816 ( .A1(n8287), .A2(n6779), .ZN(n5788) );
  OAI211_X1 U6817 ( .C1(n6815), .C2(n9852), .A(n5789), .B(n5788), .ZN(n9728)
         );
  NAND2_X1 U6818 ( .A1(n7415), .A2(n9728), .ZN(n6152) );
  NAND2_X1 U6819 ( .A1(n5290), .A2(n9804), .ZN(n8344) );
  NAND2_X1 U6820 ( .A1(n6152), .A2(n8344), .ZN(n8454) );
  INV_X1 U6821 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6785) );
  XNOR2_X1 U6822 ( .A(n5791), .B(SI_5_), .ZN(n5792) );
  XNOR2_X1 U6823 ( .A(n5793), .B(n5792), .ZN(n6777) );
  NAND2_X1 U6824 ( .A1(n6777), .A2(n8333), .ZN(n5796) );
  NAND2_X1 U6825 ( .A1(n5692), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5794) );
  XNOR2_X1 U6826 ( .A(n5794), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9872) );
  NAND2_X1 U6827 ( .A1(n5954), .A2(n9872), .ZN(n5795) );
  OAI211_X1 U6828 ( .C1(n8287), .C2(n6785), .A(n5796), .B(n5795), .ZN(n7689)
         );
  NAND2_X1 U6829 ( .A1(n6113), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5806) );
  INV_X1 U6830 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5797) );
  OR2_X1 U6831 ( .A1(n6141), .A2(n5797), .ZN(n5805) );
  INV_X1 U6832 ( .A(n5798), .ZN(n5817) );
  INV_X1 U6833 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U6834 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5799) );
  NAND2_X1 U6835 ( .A1(n5800), .A2(n5799), .ZN(n5801) );
  NAND2_X1 U6836 ( .A1(n5817), .A2(n5801), .ZN(n7414) );
  OR2_X1 U6837 ( .A1(n6140), .A2(n7414), .ZN(n5804) );
  INV_X1 U6838 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5802) );
  OR2_X1 U6839 ( .A1(n8294), .A2(n5802), .ZN(n5803) );
  NAND4_X1 U6840 ( .A1(n5806), .A2(n5805), .A3(n5804), .A4(n5803), .ZN(n9803)
         );
  NAND2_X1 U6841 ( .A1(n10756), .A2(n9803), .ZN(n8365) );
  INV_X1 U6842 ( .A(n9803), .ZN(n9726) );
  NAND2_X1 U6843 ( .A1(n9726), .A2(n7689), .ZN(n8351) );
  NAND2_X1 U6844 ( .A1(n8365), .A2(n8351), .ZN(n8455) );
  XNOR2_X1 U6845 ( .A(n5809), .B(n5808), .ZN(n6788) );
  NAND2_X1 U6846 ( .A1(n6788), .A2(n8333), .ZN(n5816) );
  INV_X1 U6847 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6124) );
  NOR2_X1 U6848 ( .A1(n5810), .A2(n6124), .ZN(n5811) );
  NAND2_X1 U6849 ( .A1(n5811), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5814) );
  INV_X1 U6850 ( .A(n5811), .ZN(n5813) );
  INV_X1 U6851 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U6852 ( .A1(n5813), .A2(n5812), .ZN(n5828) );
  AOI22_X1 U6853 ( .A1(n8332), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5954), .B2(
        n9887), .ZN(n5815) );
  NAND2_X1 U6854 ( .A1(n5816), .A2(n5815), .ZN(n7851) );
  NAND2_X1 U6855 ( .A1(n6139), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5822) );
  INV_X1 U6856 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7856) );
  OR2_X1 U6857 ( .A1(n6727), .A2(n7856), .ZN(n5821) );
  INV_X1 U6858 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7452) );
  NAND2_X1 U6859 ( .A1(n5817), .A2(n7452), .ZN(n5818) );
  NAND2_X1 U6860 ( .A1(n5834), .A2(n5818), .ZN(n7848) );
  OR2_X1 U6861 ( .A1(n6140), .A2(n7848), .ZN(n5820) );
  INV_X1 U6862 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6957) );
  OR2_X1 U6863 ( .A1(n6141), .A2(n6957), .ZN(n5819) );
  NAND4_X1 U6864 ( .A1(n5822), .A2(n5821), .A3(n5820), .A4(n5819), .ZN(n9802)
         );
  INV_X1 U6865 ( .A(n9802), .ZN(n5823) );
  OR2_X1 U6866 ( .A1(n7851), .A2(n5823), .ZN(n8354) );
  NAND2_X1 U6867 ( .A1(n7851), .A2(n5823), .ZN(n8457) );
  NAND2_X1 U6868 ( .A1(n8354), .A2(n8457), .ZN(n8353) );
  NAND2_X1 U6869 ( .A1(n7170), .A2(n8353), .ZN(n7169) );
  NAND2_X1 U6870 ( .A1(n5824), .A2(n5823), .ZN(n5825) );
  NAND2_X1 U6871 ( .A1(n7169), .A2(n5825), .ZN(n7323) );
  XNOR2_X1 U6872 ( .A(n5827), .B(n5826), .ZN(n6792) );
  NAND2_X1 U6873 ( .A1(n6792), .A2(n8333), .ZN(n5831) );
  NAND2_X1 U6874 ( .A1(n5828), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5829) );
  XNOR2_X1 U6875 ( .A(n5829), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6978) );
  AOI22_X1 U6876 ( .A1(n8332), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5954), .B2(
        n6978), .ZN(n5830) );
  NAND2_X1 U6877 ( .A1(n6139), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5840) );
  INV_X1 U6878 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7579) );
  OR2_X1 U6879 ( .A1(n6727), .A2(n7579), .ZN(n5839) );
  INV_X1 U6880 ( .A(n5832), .ZN(n5848) );
  NAND2_X1 U6881 ( .A1(n5834), .A2(n5833), .ZN(n5835) );
  NAND2_X1 U6882 ( .A1(n5848), .A2(n5835), .ZN(n8310) );
  OR2_X1 U6883 ( .A1(n6140), .A2(n8310), .ZN(n5838) );
  INV_X1 U6884 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5836) );
  OR2_X1 U6885 ( .A1(n6141), .A2(n5836), .ZN(n5837) );
  NAND4_X1 U6886 ( .A1(n5840), .A2(n5839), .A3(n5838), .A4(n5837), .ZN(n9801)
         );
  INV_X1 U6887 ( .A(n9801), .ZN(n7864) );
  OR2_X1 U6888 ( .A1(n8313), .A2(n7864), .ZN(n8361) );
  NAND2_X1 U6889 ( .A1(n8313), .A2(n7864), .ZN(n8360) );
  NAND2_X1 U6890 ( .A1(n8361), .A2(n8360), .ZN(n8358) );
  NAND2_X1 U6891 ( .A1(n6796), .A2(n8333), .ZN(n5847) );
  NAND2_X1 U6892 ( .A1(n5843), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5844) );
  MUX2_X1 U6893 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5844), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5845) );
  AND2_X1 U6894 ( .A1(n5845), .A2(n5855), .ZN(n9903) );
  AOI22_X1 U6895 ( .A1(n8332), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5954), .B2(
        n9903), .ZN(n5846) );
  NAND2_X1 U6896 ( .A1(n6139), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5853) );
  INV_X1 U6897 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7861) );
  OR2_X1 U6898 ( .A1(n6727), .A2(n7861), .ZN(n5852) );
  INV_X1 U6899 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7728) );
  NAND2_X1 U6900 ( .A1(n5848), .A2(n7728), .ZN(n5849) );
  NAND2_X1 U6901 ( .A1(n5860), .A2(n5849), .ZN(n7860) );
  OR2_X1 U6902 ( .A1(n6140), .A2(n7860), .ZN(n5851) );
  INV_X1 U6903 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6958) );
  OR2_X1 U6904 ( .A1(n6141), .A2(n6958), .ZN(n5850) );
  NAND4_X1 U6905 ( .A1(n5853), .A2(n5852), .A3(n5851), .A4(n5850), .ZN(n9800)
         );
  OR2_X1 U6906 ( .A1(n8374), .A2(n8373), .ZN(n6153) );
  XNOR2_X1 U6907 ( .A(n5854), .B(n5553), .ZN(n6808) );
  NAND2_X1 U6908 ( .A1(n6808), .A2(n8333), .ZN(n5858) );
  NAND2_X1 U6909 ( .A1(n5855), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5856) );
  XNOR2_X1 U6910 ( .A(n5856), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7086) );
  AOI22_X1 U6911 ( .A1(n8332), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5954), .B2(
        n7086), .ZN(n5857) );
  NAND2_X1 U6912 ( .A1(n6113), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5867) );
  INV_X1 U6913 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6959) );
  OR2_X1 U6914 ( .A1(n6141), .A2(n6959), .ZN(n5866) );
  NAND2_X1 U6915 ( .A1(n5860), .A2(n5859), .ZN(n5861) );
  NAND2_X1 U6916 ( .A1(n5862), .A2(n5861), .ZN(n7801) );
  OR2_X1 U6917 ( .A1(n6140), .A2(n7801), .ZN(n5865) );
  INV_X1 U6918 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5863) );
  OR2_X1 U6919 ( .A1(n8294), .A2(n5863), .ZN(n5864) );
  NAND4_X1 U6920 ( .A1(n5867), .A2(n5866), .A3(n5865), .A4(n5864), .ZN(n9799)
         );
  OR2_X1 U6921 ( .A1(n7807), .A2(n7966), .ZN(n8375) );
  NAND2_X1 U6922 ( .A1(n7807), .A2(n7966), .ZN(n8378) );
  NAND2_X1 U6923 ( .A1(n8375), .A2(n8378), .ZN(n7499) );
  NAND2_X1 U6924 ( .A1(n7497), .A2(n7499), .ZN(n7496) );
  NAND2_X1 U6925 ( .A1(n7496), .A2(n5868), .ZN(n7557) );
  INV_X1 U6926 ( .A(n9798), .ZN(n10797) );
  NAND2_X1 U6927 ( .A1(n7969), .A2(n10797), .ZN(n10789) );
  NAND2_X1 U6928 ( .A1(n8540), .A2(n10789), .ZN(n8460) );
  NAND2_X1 U6929 ( .A1(n6139), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5877) );
  INV_X1 U6930 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5869) );
  OR2_X1 U6931 ( .A1(n6727), .A2(n5869), .ZN(n5876) );
  NAND2_X1 U6932 ( .A1(n5871), .A2(n5870), .ZN(n5872) );
  NAND2_X1 U6933 ( .A1(n5873), .A2(n5872), .ZN(n10806) );
  OR2_X1 U6934 ( .A1(n6140), .A2(n10806), .ZN(n5875) );
  INV_X1 U6935 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7305) );
  OR2_X1 U6936 ( .A1(n6141), .A2(n7305), .ZN(n5874) );
  NAND4_X1 U6937 ( .A1(n5877), .A2(n5876), .A3(n5875), .A4(n5874), .ZN(n9797)
         );
  XNOR2_X1 U6938 ( .A(n5879), .B(n5878), .ZN(n6831) );
  NAND2_X1 U6939 ( .A1(n6831), .A2(n8333), .ZN(n5883) );
  NAND2_X1 U6940 ( .A1(n5880), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5881) );
  XNOR2_X1 U6941 ( .A(n5881), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7430) );
  AOI22_X1 U6942 ( .A1(n8332), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5954), .B2(
        n7430), .ZN(n5882) );
  INV_X1 U6943 ( .A(n9797), .ZN(n8195) );
  XNOR2_X1 U6944 ( .A(n5886), .B(n5885), .ZN(n6986) );
  NAND2_X1 U6945 ( .A1(n6986), .A2(n8333), .ZN(n5889) );
  XNOR2_X1 U6946 ( .A(n5887), .B(P1_IR_REG_14__SCAN_IN), .ZN(n8074) );
  AOI22_X1 U6947 ( .A1(n8332), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5954), .B2(
        n8074), .ZN(n5888) );
  NAND2_X1 U6948 ( .A1(n6139), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5898) );
  INV_X1 U6949 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8042) );
  OR2_X1 U6950 ( .A1(n6727), .A2(n8042), .ZN(n5897) );
  INV_X1 U6951 ( .A(n5890), .ZN(n5919) );
  NAND2_X1 U6952 ( .A1(n5892), .A2(n5891), .ZN(n5893) );
  NAND2_X1 U6953 ( .A1(n5919), .A2(n5893), .ZN(n9645) );
  OR2_X1 U6954 ( .A1(n6140), .A2(n9645), .ZN(n5896) );
  INV_X1 U6955 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5894) );
  OR2_X1 U6956 ( .A1(n6141), .A2(n5894), .ZN(n5895) );
  NAND4_X1 U6957 ( .A1(n5898), .A2(n5897), .A3(n5896), .A4(n5895), .ZN(n9794)
         );
  XNOR2_X1 U6958 ( .A(n5900), .B(n5899), .ZN(n7072) );
  NAND2_X1 U6959 ( .A1(n7072), .A2(n8333), .ZN(n5906) );
  NAND2_X1 U6960 ( .A1(n5901), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5903) );
  INV_X1 U6961 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U6962 ( .A1(n5903), .A2(n5902), .ZN(n5913) );
  OR2_X1 U6963 ( .A1(n5903), .A2(n5902), .ZN(n5904) );
  NAND2_X1 U6964 ( .A1(n5913), .A2(n5904), .ZN(n8173) );
  INV_X1 U6965 ( .A(n8173), .ZN(n8076) );
  AOI22_X1 U6966 ( .A1(n8332), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5954), .B2(
        n8076), .ZN(n5905) );
  NAND2_X1 U6967 ( .A1(n6139), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5910) );
  INV_X1 U6968 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8116) );
  OR2_X1 U6969 ( .A1(n6727), .A2(n8116), .ZN(n5909) );
  INV_X1 U6970 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5918) );
  XNOR2_X1 U6971 ( .A(n5919), .B(n5918), .ZN(n9780) );
  OR2_X1 U6972 ( .A1(n6140), .A2(n9780), .ZN(n5908) );
  INV_X1 U6973 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10296) );
  OR2_X1 U6974 ( .A1(n6141), .A2(n10296), .ZN(n5907) );
  NAND4_X1 U6975 ( .A1(n5910), .A2(n5909), .A3(n5908), .A4(n5907), .ZN(n10165)
         );
  INV_X1 U6976 ( .A(n10165), .ZN(n9695) );
  NAND2_X1 U6977 ( .A1(n9786), .A2(n9695), .ZN(n8400) );
  XNOR2_X1 U6978 ( .A(n5912), .B(n5911), .ZN(n7318) );
  NAND2_X1 U6979 ( .A1(n7318), .A2(n8333), .ZN(n5916) );
  NAND2_X1 U6980 ( .A1(n5913), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5914) );
  XNOR2_X1 U6981 ( .A(n5914), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8232) );
  AOI22_X1 U6982 ( .A1(n8332), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5954), .B2(
        n8232), .ZN(n5915) );
  INV_X1 U6983 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5917) );
  OAI21_X1 U6984 ( .B1(n5919), .B2(n5918), .A(n5917), .ZN(n5921) );
  NAND2_X1 U6985 ( .A1(n5921), .A2(n5920), .ZN(n10161) );
  OR2_X1 U6986 ( .A1(n10161), .A2(n6140), .ZN(n5925) );
  INV_X1 U6987 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10177) );
  OR2_X1 U6988 ( .A1(n6727), .A2(n10177), .ZN(n5924) );
  INV_X1 U6989 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10334) );
  OR2_X1 U6990 ( .A1(n8294), .A2(n10334), .ZN(n5923) );
  INV_X1 U6991 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10290) );
  OR2_X1 U6992 ( .A1(n6141), .A2(n10290), .ZN(n5922) );
  NAND4_X1 U6993 ( .A1(n5925), .A2(n5924), .A3(n5923), .A4(n5922), .ZN(n9793)
         );
  INV_X1 U6994 ( .A(n9793), .ZN(n10278) );
  NAND2_X1 U6995 ( .A1(n10176), .A2(n10278), .ZN(n8549) );
  NAND2_X1 U6996 ( .A1(n8553), .A2(n8549), .ZN(n6165) );
  INV_X1 U6997 ( .A(n10266), .ZN(n10137) );
  NAND2_X1 U6998 ( .A1(n10282), .A2(n10137), .ZN(n8407) );
  NAND2_X1 U6999 ( .A1(n5927), .A2(n5926), .ZN(n5929) );
  INV_X1 U7000 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7472) );
  INV_X1 U7001 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7470) );
  MUX2_X1 U7002 ( .A(n7472), .B(n7470), .S(n8328), .Z(n5942) );
  XNOR2_X1 U7003 ( .A(n5942), .B(SI_18_), .ZN(n5941) );
  XNOR2_X1 U7004 ( .A(n5946), .B(n5941), .ZN(n7469) );
  NAND2_X1 U7005 ( .A1(n7469), .A2(n8333), .ZN(n5933) );
  INV_X1 U7006 ( .A(n6122), .ZN(n5931) );
  XNOR2_X1 U7007 ( .A(n5952), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9929) );
  AOI22_X1 U7008 ( .A1(n8332), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5954), .B2(
        n9929), .ZN(n5932) );
  INV_X1 U7009 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U7010 ( .A1(n5935), .A2(n5934), .ZN(n5936) );
  NAND2_X1 U7011 ( .A1(n5958), .A2(n5936), .ZN(n10133) );
  INV_X1 U7012 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10134) );
  OR2_X1 U7013 ( .A1(n6727), .A2(n10134), .ZN(n5938) );
  INV_X1 U7014 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10275) );
  OR2_X1 U7015 ( .A1(n6141), .A2(n10275), .ZN(n5937) );
  AND2_X1 U7016 ( .A1(n5938), .A2(n5937), .ZN(n5940) );
  NAND2_X1 U7017 ( .A1(n6139), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5939) );
  OAI211_X1 U7018 ( .C1(n10133), .C2(n6140), .A(n5940), .B(n5939), .ZN(n10257)
         );
  INV_X1 U7019 ( .A(n10257), .ZN(n10279) );
  INV_X1 U7020 ( .A(n5941), .ZN(n5945) );
  INV_X1 U7021 ( .A(n5942), .ZN(n5943) );
  NAND2_X1 U7022 ( .A1(n5943), .A2(SI_18_), .ZN(n5944) );
  INV_X1 U7023 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7600) );
  INV_X1 U7024 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7601) );
  MUX2_X1 U7025 ( .A(n7600), .B(n7601), .S(n8328), .Z(n5947) );
  INV_X1 U7026 ( .A(SI_19_), .ZN(n10506) );
  NAND2_X1 U7027 ( .A1(n5947), .A2(n10506), .ZN(n5962) );
  INV_X1 U7028 ( .A(n5947), .ZN(n5948) );
  NAND2_X1 U7029 ( .A1(n5948), .A2(SI_19_), .ZN(n5949) );
  NAND2_X1 U7030 ( .A1(n5962), .A2(n5949), .ZN(n5963) );
  XNOR2_X1 U7031 ( .A(n5964), .B(n5963), .ZN(n7599) );
  NAND2_X1 U7032 ( .A1(n7599), .A2(n8333), .ZN(n5956) );
  INV_X1 U7033 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5950) );
  OR2_X1 U7034 ( .A1(n6124), .A2(n5950), .ZN(n5951) );
  XNOR2_X2 U7035 ( .A(n5953), .B(n5571), .ZN(n6137) );
  AOI22_X1 U7036 ( .A1(n8332), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6137), .B2(
        n5954), .ZN(n5955) );
  INV_X1 U7037 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10264) );
  INV_X1 U7038 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5957) );
  INV_X1 U7039 ( .A(n5972), .ZN(n5974) );
  NAND2_X1 U7040 ( .A1(n5958), .A2(n5957), .ZN(n5959) );
  NAND2_X1 U7041 ( .A1(n5974), .A2(n5959), .ZN(n10117) );
  OR2_X1 U7042 ( .A1(n10117), .A2(n6140), .ZN(n5961) );
  AOI22_X1 U7043 ( .A1(n6113), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n6139), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5960) );
  OAI211_X1 U7044 ( .C1(n6141), .C2(n10264), .A(n5961), .B(n5960), .ZN(n10269)
         );
  INV_X1 U7045 ( .A(n10269), .ZN(n9756) );
  OR2_X1 U7046 ( .A1(n10125), .A2(n9756), .ZN(n8411) );
  NAND2_X1 U7047 ( .A1(n10125), .A2(n9756), .ZN(n8415) );
  INV_X1 U7048 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7698) );
  INV_X1 U7049 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7652) );
  MUX2_X1 U7050 ( .A(n7698), .B(n7652), .S(n8328), .Z(n5965) );
  INV_X1 U7051 ( .A(SI_20_), .ZN(n10501) );
  NAND2_X1 U7052 ( .A1(n5965), .A2(n10501), .ZN(n5981) );
  INV_X1 U7053 ( .A(n5965), .ZN(n5966) );
  NAND2_X1 U7054 ( .A1(n5966), .A2(SI_20_), .ZN(n5967) );
  OAI21_X1 U7055 ( .B1(n5969), .B2(n5968), .A(n5982), .ZN(n7695) );
  NAND2_X1 U7056 ( .A1(n7695), .A2(n8333), .ZN(n5971) );
  OR2_X1 U7057 ( .A1(n8287), .A2(n7652), .ZN(n5970) );
  INV_X1 U7058 ( .A(n5985), .ZN(n5987) );
  INV_X1 U7059 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U7060 ( .A1(n5974), .A2(n5973), .ZN(n5975) );
  AND2_X1 U7061 ( .A1(n5987), .A2(n5975), .ZN(n10103) );
  INV_X1 U7062 ( .A(n6140), .ZN(n6080) );
  NAND2_X1 U7063 ( .A1(n10103), .A2(n6080), .ZN(n5980) );
  INV_X1 U7064 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10255) );
  NAND2_X1 U7065 ( .A1(n6113), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U7066 ( .A1(n6139), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5976) );
  OAI211_X1 U7067 ( .C1(n10255), .C2(n6141), .A(n5977), .B(n5976), .ZN(n5978)
         );
  INV_X1 U7068 ( .A(n5978), .ZN(n5979) );
  NAND2_X1 U7069 ( .A1(n5980), .A2(n5979), .ZN(n10258) );
  INV_X1 U7070 ( .A(n10258), .ZN(n9676) );
  OR2_X1 U7071 ( .A1(n10110), .A2(n9676), .ZN(n8418) );
  NAND2_X1 U7072 ( .A1(n10110), .A2(n9676), .ZN(n10082) );
  MUX2_X1 U7073 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n8328), .Z(n5997) );
  INV_X1 U7074 ( .A(SI_21_), .ZN(n10397) );
  XNOR2_X1 U7075 ( .A(n5997), .B(n10397), .ZN(n5996) );
  XNOR2_X1 U7076 ( .A(n5995), .B(n5996), .ZN(n7790) );
  NAND2_X1 U7077 ( .A1(n7790), .A2(n8333), .ZN(n5984) );
  INV_X1 U7078 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7841) );
  OR2_X1 U7079 ( .A1(n8287), .A2(n7841), .ZN(n5983) );
  INV_X1 U7080 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7081 ( .A1(n5987), .A2(n5986), .ZN(n5988) );
  NAND2_X1 U7082 ( .A1(n6002), .A2(n5988), .ZN(n10092) );
  OR2_X1 U7083 ( .A1(n10092), .A2(n6140), .ZN(n5993) );
  INV_X1 U7084 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10247) );
  NAND2_X1 U7085 ( .A1(n6139), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7086 ( .A1(n6113), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5989) );
  OAI211_X1 U7087 ( .C1(n10247), .C2(n6141), .A(n5990), .B(n5989), .ZN(n5991)
         );
  INV_X1 U7088 ( .A(n5991), .ZN(n5992) );
  NAND2_X1 U7089 ( .A1(n5993), .A2(n5992), .ZN(n10249) );
  INV_X1 U7090 ( .A(n10249), .ZN(n10106) );
  NAND2_X1 U7091 ( .A1(n10091), .A2(n10106), .ZN(n8413) );
  NAND2_X1 U7092 ( .A1(n10319), .A2(n10106), .ZN(n5994) );
  NAND2_X1 U7093 ( .A1(n10080), .A2(n5994), .ZN(n10066) );
  NAND2_X1 U7094 ( .A1(n5997), .A2(SI_21_), .ZN(n5998) );
  NAND2_X1 U7095 ( .A1(n5999), .A2(n5998), .ZN(n6012) );
  MUX2_X1 U7096 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n8328), .Z(n6013) );
  XNOR2_X1 U7097 ( .A(n6013), .B(SI_22_), .ZN(n6010) );
  XNOR2_X1 U7098 ( .A(n6012), .B(n6010), .ZN(n7879) );
  NAND2_X1 U7099 ( .A1(n7879), .A2(n8333), .ZN(n6001) );
  INV_X1 U7100 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8988) );
  OR2_X1 U7101 ( .A1(n8287), .A2(n8988), .ZN(n6000) );
  INV_X1 U7102 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9746) );
  NAND2_X1 U7103 ( .A1(n6002), .A2(n9746), .ZN(n6003) );
  NAND2_X1 U7104 ( .A1(n6025), .A2(n6003), .ZN(n10067) );
  OR2_X1 U7105 ( .A1(n10067), .A2(n6140), .ZN(n6008) );
  INV_X1 U7106 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10242) );
  NAND2_X1 U7107 ( .A1(n6139), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U7108 ( .A1(n6113), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6004) );
  OAI211_X1 U7109 ( .C1(n10242), .C2(n6141), .A(n6005), .B(n6004), .ZN(n6006)
         );
  INV_X1 U7110 ( .A(n6006), .ZN(n6007) );
  NAND2_X1 U7111 ( .A1(n6008), .A2(n6007), .ZN(n10086) );
  INV_X1 U7112 ( .A(n10086), .ZN(n9677) );
  NAND2_X1 U7113 ( .A1(n10077), .A2(n9677), .ZN(n8422) );
  NAND2_X1 U7114 ( .A1(n8421), .A2(n8422), .ZN(n10065) );
  INV_X1 U7115 ( .A(n10077), .ZN(n10315) );
  NAND2_X1 U7116 ( .A1(n10315), .A2(n9677), .ZN(n6009) );
  INV_X1 U7117 ( .A(n6010), .ZN(n6011) );
  NAND2_X1 U7118 ( .A1(n6013), .A2(SI_22_), .ZN(n6014) );
  INV_X1 U7119 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n6015) );
  INV_X1 U7120 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7912) );
  MUX2_X1 U7121 ( .A(n6015), .B(n7912), .S(n8328), .Z(n6016) );
  INV_X1 U7122 ( .A(SI_23_), .ZN(n10498) );
  NAND2_X1 U7123 ( .A1(n6016), .A2(n10498), .ZN(n6034) );
  INV_X1 U7124 ( .A(n6016), .ZN(n6017) );
  NAND2_X1 U7125 ( .A1(n6017), .A2(SI_23_), .ZN(n6018) );
  NAND2_X1 U7126 ( .A1(n6034), .A2(n6018), .ZN(n6020) );
  NAND2_X1 U7127 ( .A1(n6021), .A2(n6020), .ZN(n6022) );
  NAND2_X1 U7128 ( .A1(n6035), .A2(n6022), .ZN(n7909) );
  NAND2_X1 U7129 ( .A1(n7909), .A2(n8333), .ZN(n6024) );
  OR2_X1 U7130 ( .A1(n8287), .A2(n7912), .ZN(n6023) );
  INV_X1 U7131 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9659) );
  NAND2_X1 U7132 ( .A1(n6025), .A2(n9659), .ZN(n6026) );
  AND2_X1 U7133 ( .A1(n6042), .A2(n6026), .ZN(n10048) );
  NAND2_X1 U7134 ( .A1(n10048), .A2(n6080), .ZN(n6032) );
  INV_X1 U7135 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7136 ( .A1(n6113), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U7137 ( .A1(n6139), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6027) );
  OAI211_X1 U7138 ( .C1(n6029), .C2(n6141), .A(n6028), .B(n6027), .ZN(n6030)
         );
  INV_X1 U7139 ( .A(n6030), .ZN(n6031) );
  NAND2_X1 U7140 ( .A1(n6032), .A2(n6031), .ZN(n10236) );
  NAND2_X1 U7141 ( .A1(n10232), .A2(n10236), .ZN(n6033) );
  INV_X1 U7142 ( .A(n10236), .ZN(n10071) );
  INV_X1 U7143 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n6036) );
  INV_X1 U7144 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8068) );
  MUX2_X1 U7145 ( .A(n6036), .B(n8068), .S(n8328), .Z(n6037) );
  INV_X1 U7146 ( .A(SI_24_), .ZN(n10379) );
  NAND2_X1 U7147 ( .A1(n6037), .A2(n10379), .ZN(n6053) );
  INV_X1 U7148 ( .A(n6037), .ZN(n6038) );
  NAND2_X1 U7149 ( .A1(n6038), .A2(SI_24_), .ZN(n6039) );
  AND2_X1 U7150 ( .A1(n6053), .A2(n6039), .ZN(n6051) );
  OR2_X1 U7151 ( .A1(n8287), .A2(n8068), .ZN(n6040) );
  INV_X1 U7152 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9716) );
  INV_X1 U7153 ( .A(n6057), .ZN(n6044) );
  NAND2_X1 U7154 ( .A1(n6042), .A2(n9716), .ZN(n6043) );
  NAND2_X1 U7155 ( .A1(n6044), .A2(n6043), .ZN(n10035) );
  OR2_X1 U7156 ( .A1(n10035), .A2(n6140), .ZN(n6050) );
  INV_X1 U7157 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6047) );
  NAND2_X1 U7158 ( .A1(n6113), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U7159 ( .A1(n6139), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6045) );
  OAI211_X1 U7160 ( .C1(n6047), .C2(n6141), .A(n6046), .B(n6045), .ZN(n6048)
         );
  INV_X1 U7161 ( .A(n6048), .ZN(n6049) );
  NAND2_X1 U7162 ( .A1(n6050), .A2(n6049), .ZN(n10056) );
  NOR2_X1 U7163 ( .A1(n10227), .A2(n10056), .ZN(n10018) );
  MUX2_X1 U7164 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n8328), .Z(n6068) );
  INV_X1 U7165 ( .A(SI_25_), .ZN(n10480) );
  XNOR2_X1 U7166 ( .A(n6068), .B(n10480), .ZN(n6067) );
  INV_X1 U7167 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8110) );
  OR2_X1 U7168 ( .A1(n8287), .A2(n8110), .ZN(n6055) );
  NOR2_X1 U7169 ( .A1(n6057), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6058) );
  OR2_X1 U7170 ( .A1(n6078), .A2(n6058), .ZN(n9685) );
  INV_X1 U7171 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7172 ( .A1(n6113), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7173 ( .A1(n6139), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6059) );
  OAI211_X1 U7174 ( .C1(n6061), .C2(n6141), .A(n6060), .B(n6059), .ZN(n6062)
         );
  INV_X1 U7175 ( .A(n6062), .ZN(n6063) );
  OAI21_X1 U7176 ( .B1(n9685), .B2(n6140), .A(n6063), .ZN(n10005) );
  INV_X1 U7177 ( .A(n10005), .ZN(n10224) );
  OR2_X1 U7178 ( .A1(n10018), .A2(n4986), .ZN(n6064) );
  NAND2_X1 U7179 ( .A1(n10227), .A2(n10056), .ZN(n10019) );
  AND2_X1 U7180 ( .A1(n5028), .A2(n10019), .ZN(n6065) );
  INV_X1 U7181 ( .A(n6067), .ZN(n6070) );
  NAND2_X1 U7182 ( .A1(n6068), .A2(SI_25_), .ZN(n6069) );
  INV_X1 U7183 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n6072) );
  INV_X1 U7184 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8261) );
  MUX2_X1 U7185 ( .A(n6072), .B(n8261), .S(n8328), .Z(n6073) );
  INV_X1 U7186 ( .A(SI_26_), .ZN(n10495) );
  NAND2_X1 U7187 ( .A1(n6073), .A2(n10495), .ZN(n6087) );
  INV_X1 U7188 ( .A(n6073), .ZN(n6074) );
  NAND2_X1 U7189 ( .A1(n6074), .A2(SI_26_), .ZN(n6075) );
  NAND2_X1 U7190 ( .A1(n6087), .A2(n6075), .ZN(n6088) );
  OR2_X1 U7191 ( .A1(n8287), .A2(n8261), .ZN(n6076) );
  OR2_X1 U7192 ( .A1(n6078), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7193 ( .A1(n6078), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6102) );
  AND2_X1 U7194 ( .A1(n6079), .A2(n6102), .ZN(n10010) );
  NAND2_X1 U7195 ( .A1(n10010), .A2(n6080), .ZN(n6086) );
  INV_X1 U7196 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U7197 ( .A1(n6113), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6082) );
  NAND2_X1 U7198 ( .A1(n6139), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6081) );
  OAI211_X1 U7199 ( .C1(n6083), .C2(n6141), .A(n6082), .B(n6081), .ZN(n6084)
         );
  INV_X1 U7200 ( .A(n6084), .ZN(n6085) );
  NAND2_X1 U7201 ( .A1(n6086), .A2(n6085), .ZN(n10028) );
  INV_X1 U7202 ( .A(n10028), .ZN(n9634) );
  INV_X1 U7203 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6090) );
  INV_X1 U7204 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n6097) );
  MUX2_X1 U7205 ( .A(n6090), .B(n6097), .S(n8328), .Z(n6091) );
  INV_X1 U7206 ( .A(SI_27_), .ZN(n10486) );
  NAND2_X1 U7207 ( .A1(n6091), .A2(n10486), .ZN(n6109) );
  INV_X1 U7208 ( .A(n6091), .ZN(n6092) );
  NAND2_X1 U7209 ( .A1(n6092), .A2(SI_27_), .ZN(n6093) );
  AND2_X1 U7210 ( .A1(n6109), .A2(n6093), .ZN(n6094) );
  OR2_X1 U7211 ( .A1(n8287), .A2(n6097), .ZN(n6098) );
  NAND2_X1 U7212 ( .A1(n6113), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6107) );
  INV_X1 U7213 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6101) );
  OR2_X1 U7214 ( .A1(n6141), .A2(n6101), .ZN(n6106) );
  XNOR2_X1 U7215 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n6114), .ZN(n9991) );
  OR2_X1 U7216 ( .A1(n6140), .A2(n9991), .ZN(n6105) );
  INV_X1 U7217 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n6103) );
  OR2_X1 U7218 ( .A1(n8294), .A2(n6103), .ZN(n6104) );
  NAND4_X1 U7219 ( .A1(n6107), .A2(n6106), .A3(n6105), .A4(n6104), .ZN(n10004)
         );
  NAND2_X1 U7220 ( .A1(n9990), .A2(n8983), .ZN(n8501) );
  NAND2_X1 U7221 ( .A1(n10206), .A2(n8983), .ZN(n6108) );
  MUX2_X1 U7222 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n8328), .Z(n6614) );
  INV_X1 U7223 ( .A(SI_28_), .ZN(n10491) );
  XNOR2_X1 U7224 ( .A(n6614), .B(n10491), .ZN(n6612) );
  INV_X1 U7225 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8994) );
  OR2_X1 U7226 ( .A1(n8287), .A2(n8994), .ZN(n6111) );
  NAND2_X1 U7227 ( .A1(n6113), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6120) );
  INV_X1 U7228 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6203) );
  OR2_X1 U7229 ( .A1(n8294), .A2(n6203), .ZN(n6119) );
  NAND3_X1 U7230 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .A3(n6114), .ZN(n9967) );
  INV_X1 U7231 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8982) );
  NAND2_X1 U7232 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n6114), .ZN(n6115) );
  NAND2_X1 U7233 ( .A1(n8982), .A2(n6115), .ZN(n6116) );
  NAND2_X1 U7234 ( .A1(n9967), .A2(n6116), .ZN(n9976) );
  OR2_X1 U7235 ( .A1(n6140), .A2(n9976), .ZN(n6118) );
  INV_X1 U7236 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6745) );
  OR2_X1 U7237 ( .A1(n6141), .A2(n6745), .ZN(n6117) );
  NAND4_X1 U7238 ( .A1(n6120), .A2(n6119), .A3(n6118), .A4(n6117), .ZN(n9792)
         );
  NAND2_X1 U7239 ( .A1(n9983), .A2(n10205), .ZN(n8502) );
  NOR2_X1 U7240 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n6121) );
  NAND2_X1 U7241 ( .A1(n6122), .A2(n6121), .ZN(n6131) );
  INV_X1 U7242 ( .A(n6131), .ZN(n6123) );
  NAND2_X1 U7243 ( .A1(n6123), .A2(n6132), .ZN(n6176) );
  INV_X1 U7244 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6125) );
  INV_X1 U7245 ( .A(n6128), .ZN(n6127) );
  INV_X1 U7246 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6126) );
  NAND2_X1 U7247 ( .A1(n6127), .A2(n6126), .ZN(n6194) );
  NAND2_X1 U7248 ( .A1(n6128), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7249 ( .A1(n6194), .A2(n6129), .ZN(n6135) );
  INV_X1 U7250 ( .A(n6995), .ZN(n6134) );
  NAND2_X1 U7251 ( .A1(n6131), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6133) );
  INV_X1 U7252 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6132) );
  XNOR2_X1 U7253 ( .A(n6133), .B(n6132), .ZN(n8576) );
  INV_X1 U7254 ( .A(n7574), .ZN(n6992) );
  NAND2_X1 U7255 ( .A1(n6134), .A2(n6992), .ZN(n7020) );
  INV_X1 U7256 ( .A(n6136), .ZN(n8519) );
  AND2_X1 U7257 ( .A1(n6135), .A2(n8519), .ZN(n10723) );
  INV_X1 U7258 ( .A(n10723), .ZN(n7022) );
  NAND2_X1 U7259 ( .A1(n7020), .A2(n7022), .ZN(n10720) );
  AND2_X1 U7260 ( .A1(n6995), .A2(n8577), .ZN(n6138) );
  OR2_X1 U7261 ( .A1(n10720), .A2(n6138), .ZN(n10786) );
  INV_X1 U7262 ( .A(n8576), .ZN(n8515) );
  NAND2_X1 U7263 ( .A1(n10786), .A2(n10778), .ZN(n10828) );
  NAND2_X1 U7264 ( .A1(n6139), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6145) );
  INV_X1 U7265 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9968) );
  OR2_X1 U7266 ( .A1(n6727), .A2(n9968), .ZN(n6144) );
  OR2_X1 U7267 ( .A1(n6140), .A2(n9967), .ZN(n6143) );
  INV_X1 U7268 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6746) );
  OR2_X1 U7269 ( .A1(n6141), .A2(n6746), .ZN(n6142) );
  INV_X1 U7270 ( .A(n6135), .ZN(n8481) );
  NAND2_X1 U7271 ( .A1(n7016), .A2(n8995), .ZN(n10794) );
  OR2_X1 U7272 ( .A1(n10232), .A2(n10071), .ZN(n8424) );
  NAND2_X1 U7273 ( .A1(n10232), .A2(n10071), .ZN(n8487) );
  INV_X1 U7274 ( .A(n10065), .ZN(n10063) );
  INV_X1 U7275 ( .A(n10082), .ZN(n8412) );
  NAND2_X1 U7276 ( .A1(n6148), .A2(n8412), .ZN(n6147) );
  AND2_X1 U7277 ( .A1(n6147), .A2(n8413), .ZN(n8492) );
  INV_X1 U7278 ( .A(n6148), .ZN(n8562) );
  INV_X1 U7279 ( .A(n10113), .ZN(n10115) );
  INV_X1 U7280 ( .A(n10722), .ZN(n8449) );
  INV_X1 U7281 ( .A(n9807), .ZN(n10721) );
  NAND2_X1 U7282 ( .A1(n10721), .A2(n10193), .ZN(n6149) );
  INV_X1 U7283 ( .A(n8453), .ZN(n6150) );
  NAND2_X1 U7284 ( .A1(n7045), .A2(n6150), .ZN(n6151) );
  INV_X1 U7285 ( .A(n6152), .ZN(n8350) );
  AND2_X1 U7286 ( .A1(n8365), .A2(n8344), .ZN(n8533) );
  INV_X1 U7287 ( .A(n8457), .ZN(n8532) );
  NAND2_X1 U7288 ( .A1(n8375), .A2(n6153), .ZN(n6155) );
  NAND2_X1 U7289 ( .A1(n8361), .A2(n8354), .ZN(n6154) );
  NOR2_X1 U7290 ( .A1(n6155), .A2(n6154), .ZN(n8535) );
  NAND2_X1 U7291 ( .A1(n7324), .A2(n8535), .ZN(n7558) );
  NAND2_X1 U7292 ( .A1(n6155), .A2(n8378), .ZN(n6157) );
  AND2_X1 U7293 ( .A1(n8369), .A2(n8360), .ZN(n6156) );
  NAND2_X1 U7294 ( .A1(n8378), .A2(n6156), .ZN(n8448) );
  NAND2_X1 U7295 ( .A1(n6157), .A2(n8448), .ZN(n8536) );
  NAND2_X1 U7296 ( .A1(n7558), .A2(n8536), .ZN(n6159) );
  INV_X1 U7297 ( .A(n8460), .ZN(n6158) );
  OR2_X1 U7298 ( .A1(n10810), .A2(n8195), .ZN(n8386) );
  NAND2_X1 U7299 ( .A1(n10810), .A2(n8195), .ZN(n8385) );
  NAND2_X1 U7300 ( .A1(n8386), .A2(n8385), .ZN(n10779) );
  INV_X1 U7301 ( .A(n10789), .ZN(n6160) );
  NOR2_X1 U7302 ( .A1(n10779), .A2(n6160), .ZN(n6161) );
  OR2_X1 U7303 ( .A1(n8188), .A2(n10795), .ZN(n8391) );
  NAND2_X1 U7304 ( .A1(n8188), .A2(n10795), .ZN(n8392) );
  OR2_X1 U7305 ( .A1(n8213), .A2(n9646), .ZN(n8545) );
  NAND2_X1 U7306 ( .A1(n8213), .A2(n9646), .ZN(n8393) );
  OR2_X1 U7307 ( .A1(n9649), .A2(n9782), .ZN(n8397) );
  NAND2_X1 U7308 ( .A1(n8119), .A2(n8397), .ZN(n6164) );
  INV_X1 U7309 ( .A(n8467), .ZN(n6163) );
  NAND2_X1 U7310 ( .A1(n6164), .A2(n6163), .ZN(n8121) );
  NAND2_X1 U7311 ( .A1(n8121), .A2(n8518), .ZN(n10164) );
  INV_X1 U7312 ( .A(n6165), .ZN(n10169) );
  NAND2_X1 U7313 ( .A1(n10164), .A2(n10169), .ZN(n10163) );
  NAND2_X1 U7314 ( .A1(n10146), .A2(n8407), .ZN(n10129) );
  OR2_X1 U7315 ( .A1(n10143), .A2(n10279), .ZN(n8558) );
  AND2_X1 U7316 ( .A1(n8558), .A2(n10128), .ZN(n8405) );
  NAND2_X1 U7317 ( .A1(n10129), .A2(n8405), .ZN(n6166) );
  NAND2_X1 U7318 ( .A1(n10143), .A2(n10279), .ZN(n8408) );
  NAND2_X1 U7319 ( .A1(n10100), .A2(n8418), .ZN(n10083) );
  INV_X1 U7320 ( .A(n10056), .ZN(n9660) );
  NAND2_X1 U7321 ( .A1(n10227), .A2(n9660), .ZN(n8494) );
  NAND2_X1 U7322 ( .A1(n8484), .A2(n8494), .ZN(n8472) );
  NAND2_X1 U7323 ( .A1(n10220), .A2(n10224), .ZN(n8495) );
  OAI21_X1 U7324 ( .B1(n8435), .B2(n6168), .A(n6723), .ZN(n6171) );
  OR2_X1 U7325 ( .A1(n6135), .A2(n9946), .ZN(n6170) );
  NAND2_X1 U7326 ( .A1(n6136), .A2(n8515), .ZN(n6169) );
  NAND2_X1 U7327 ( .A1(n6170), .A2(n6169), .ZN(n10162) );
  INV_X1 U7328 ( .A(n8995), .ZN(n9819) );
  NAND2_X1 U7329 ( .A1(n7016), .A2(n9819), .ZN(n10796) );
  AOI22_X1 U7330 ( .A1(n6171), .A2(n10162), .B1(n10267), .B2(n10004), .ZN(
        n9986) );
  INV_X1 U7331 ( .A(n10214), .ZN(n10012) );
  NAND2_X1 U7332 ( .A1(n7705), .A2(n10743), .ZN(n7704) );
  AND2_X1 U7333 ( .A1(n7687), .A2(n10756), .ZN(n7685) );
  NAND2_X1 U7334 ( .A1(n7685), .A2(n5824), .ZN(n7326) );
  INV_X1 U7335 ( .A(n7969), .ZN(n7567) );
  INV_X1 U7336 ( .A(n10810), .ZN(n10785) );
  INV_X1 U7337 ( .A(n10176), .ZN(n10336) );
  NAND2_X1 U7338 ( .A1(n10012), .A2(n10022), .ZN(n10009) );
  AND2_X1 U7339 ( .A1(n10723), .A2(n8576), .ZN(n10782) );
  OAI211_X1 U7340 ( .C1(n5301), .C2(n5302), .A(n10782), .B(n6735), .ZN(n9980)
         );
  OAI211_X1 U7341 ( .C1(n9979), .C2(n10794), .A(n9986), .B(n9980), .ZN(n6172)
         );
  XNOR2_X1 U7342 ( .A(n6173), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6197) );
  INV_X1 U7343 ( .A(n6197), .ZN(n8112) );
  NAND2_X1 U7344 ( .A1(n8112), .A2(P1_B_REG_SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7345 ( .A1(n6174), .A2(n6195), .ZN(n6175) );
  MUX2_X1 U7346 ( .A(n6178), .B(P1_B_REG_SCAN_IN), .S(n6199), .Z(n6181) );
  NAND2_X1 U7347 ( .A1(n6181), .A2(n6198), .ZN(n6826) );
  OR2_X1 U7348 ( .A1(n6826), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6183) );
  INV_X1 U7349 ( .A(n6199), .ZN(n8070) );
  INV_X1 U7350 ( .A(n6198), .ZN(n8263) );
  NAND2_X1 U7351 ( .A1(n8070), .A2(n8263), .ZN(n6182) );
  INV_X1 U7352 ( .A(n7014), .ZN(n6201) );
  NOR4_X1 U7353 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6192) );
  NOR4_X1 U7354 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6191) );
  OR4_X1 U7355 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6189) );
  NOR4_X1 U7356 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6187) );
  NOR4_X1 U7357 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6186) );
  NOR4_X1 U7358 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6185) );
  NOR4_X1 U7359 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6184) );
  NAND4_X1 U7360 ( .A1(n6187), .A2(n6186), .A3(n6185), .A4(n6184), .ZN(n6188)
         );
  NOR4_X1 U7361 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n6189), .A4(n6188), .ZN(n6190) );
  AND3_X1 U7362 ( .A1(n6192), .A2(n6191), .A3(n6190), .ZN(n6193) );
  OR2_X1 U7363 ( .A1(n6826), .A2(n6193), .ZN(n7013) );
  NAND2_X1 U7364 ( .A1(n6194), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6196) );
  XNOR2_X1 U7365 ( .A(n6196), .B(n6195), .ZN(n7910) );
  AND2_X1 U7366 ( .A1(n7028), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7367 ( .A1(n7910), .A2(n6200), .ZN(n7019) );
  NAND2_X1 U7368 ( .A1(n7016), .A2(n8577), .ZN(n7029) );
  AND3_X1 U7369 ( .A1(n7013), .A2(n7023), .A3(n7029), .ZN(n6741) );
  AND2_X1 U7370 ( .A1(n6201), .A2(n6741), .ZN(n7572) );
  OR2_X1 U7371 ( .A1(n6826), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6202) );
  NAND2_X1 U7372 ( .A1(n8263), .A2(n8112), .ZN(n6827) );
  NOR2_X1 U7373 ( .A1(n10778), .A2(n6136), .ZN(n7024) );
  NOR2_X1 U7374 ( .A1(n7571), .A2(n7024), .ZN(n6742) );
  AND2_X2 U7375 ( .A1(n7572), .A2(n6742), .ZN(n10834) );
  NAND2_X1 U7376 ( .A1(n10834), .A2(n10283), .ZN(n10340) );
  NOR2_X1 U7377 ( .A1(n10834), .A2(n6203), .ZN(n6204) );
  OAI21_X1 U7378 ( .B1(n6744), .B2(n6207), .A(n6206), .ZN(P1_U3518) );
  BUF_X1 U7379 ( .A(n6233), .Z(n6215) );
  INV_X1 U7380 ( .A(n6215), .ZN(n6216) );
  NAND2_X1 U7381 ( .A1(n6216), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6217) );
  XNOR2_X1 U7382 ( .A(n6217), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8867) );
  XNOR2_X1 U7383 ( .A(n6219), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9266) );
  INV_X1 U7384 ( .A(n9266), .ZN(n8696) );
  AND2_X1 U7385 ( .A1(n8867), .A2(n8696), .ZN(n6753) );
  NAND2_X1 U7386 ( .A1(n6219), .A2(n6218), .ZN(n6220) );
  NAND2_X1 U7387 ( .A1(n6220), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6223) );
  INV_X1 U7388 ( .A(n6223), .ZN(n6221) );
  NAND2_X1 U7389 ( .A1(n6221), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U7390 ( .A1(n6223), .A2(n6222), .ZN(n6225) );
  NAND2_X1 U7391 ( .A1(n6224), .A2(n6225), .ZN(n7696) );
  AND2_X1 U7392 ( .A1(n7696), .A2(n8696), .ZN(n8860) );
  OR2_X1 U7393 ( .A1(n6753), .A2(n8860), .ZN(n6229) );
  NAND2_X1 U7394 ( .A1(n6225), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6227) );
  INV_X1 U7395 ( .A(n8867), .ZN(n6228) );
  NAND2_X1 U7396 ( .A1(n8712), .A2(n6228), .ZN(n9559) );
  AND2_X1 U7397 ( .A1(n6229), .A2(n9559), .ZN(n6231) );
  INV_X1 U7398 ( .A(n8712), .ZN(n8693) );
  NAND2_X2 U7399 ( .A1(n8693), .A2(n8867), .ZN(n8842) );
  INV_X1 U7400 ( .A(n8860), .ZN(n6230) );
  OR2_X1 U7401 ( .A1(n8842), .A2(n6230), .ZN(n7188) );
  NAND2_X1 U7402 ( .A1(n6231), .A2(n7188), .ZN(n8140) );
  INV_X1 U7403 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6244) );
  NOR2_X1 U7404 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n6235) );
  NOR2_X1 U7405 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n6234) );
  AND2_X1 U7406 ( .A1(n6235), .A2(n6234), .ZN(n6236) );
  INV_X1 U7407 ( .A(n6238), .ZN(n6255) );
  NAND2_X1 U7408 ( .A1(n6255), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6237) );
  XNOR2_X2 U7409 ( .A(n6241), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6242) );
  AND2_X4 U7410 ( .A1(n9620), .A2(n6242), .ZN(n6458) );
  NAND2_X1 U7411 ( .A1(n6458), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6243) );
  INV_X1 U7412 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6246) );
  INV_X1 U7413 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6250) );
  OR2_X1 U7414 ( .A1(n8649), .A2(n6250), .ZN(n6251) );
  OR2_X2 U7415 ( .A1(n6259), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n6261) );
  NAND2_X1 U7416 ( .A1(n6261), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U7417 ( .A1(n6259), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6260) );
  INV_X1 U7418 ( .A(n6628), .ZN(n6274) );
  NAND2_X1 U7419 ( .A1(n6601), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6268) );
  INV_X1 U7420 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7193) );
  INV_X1 U7421 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6263) );
  OR2_X1 U7422 ( .A1(n8645), .A2(n6263), .ZN(n6266) );
  INV_X1 U7423 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6264) );
  OR2_X1 U7424 ( .A1(n8649), .A2(n6264), .ZN(n6265) );
  AND4_X2 U7425 ( .A1(n6268), .A2(n6267), .A3(n6266), .A4(n6265), .ZN(n8302)
         );
  INV_X1 U7426 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6924) );
  NAND2_X1 U7427 ( .A1(n6269), .A2(SI_0_), .ZN(n6271) );
  INV_X1 U7428 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6270) );
  XNOR2_X1 U7429 ( .A(n6271), .B(n6270), .ZN(n9627) );
  MUX2_X1 U7430 ( .A(n6924), .B(n9627), .S(n6272), .Z(n7194) );
  INV_X1 U7431 ( .A(n7194), .ZN(n6838) );
  NAND2_X1 U7432 ( .A1(n8302), .A2(n6838), .ZN(n8713) );
  NAND2_X1 U7433 ( .A1(n6274), .A2(n6273), .ZN(n7075) );
  NAND2_X1 U7434 ( .A1(n7075), .A2(n8716), .ZN(n7095) );
  INV_X1 U7435 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6275) );
  INV_X1 U7436 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6276) );
  OR2_X1 U7437 ( .A1(n8647), .A2(n6276), .ZN(n6278) );
  INV_X1 U7438 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6917) );
  AND3_X1 U7439 ( .A1(n6279), .A2(n6278), .A3(n6277), .ZN(n6281) );
  NAND2_X1 U7440 ( .A1(n6621), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6280) );
  NAND2_X2 U7441 ( .A1(n6281), .A2(n6280), .ZN(n9150) );
  INV_X1 U7442 ( .A(n9150), .ZN(n7284) );
  XNOR2_X2 U7443 ( .A(n6283), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6922) );
  INV_X1 U7444 ( .A(n7096), .ZN(n6889) );
  NAND2_X1 U7445 ( .A1(n9150), .A2(n6889), .ZN(n8724) );
  NAND2_X1 U7446 ( .A1(n8725), .A2(n8724), .ZN(n7098) );
  NAND2_X1 U7447 ( .A1(n7095), .A2(n8722), .ZN(n6285) );
  NAND2_X1 U7448 ( .A1(n6285), .A2(n8725), .ZN(n7280) );
  NAND2_X1 U7449 ( .A1(n6601), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6291) );
  OR2_X1 U7450 ( .A1(n6436), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6290) );
  INV_X1 U7451 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6286) );
  OR2_X1 U7452 ( .A1(n8645), .A2(n6286), .ZN(n6289) );
  INV_X1 U7453 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6287) );
  OR2_X1 U7454 ( .A1(n8649), .A2(n6287), .ZN(n6288) );
  NAND2_X1 U7455 ( .A1(n6292), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U7456 ( .A1(n6293), .A2(n6294), .ZN(n6320) );
  NAND2_X1 U7457 ( .A1(n6320), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6296) );
  INV_X1 U7458 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U7459 ( .A1(n6296), .A2(n6295), .ZN(n6306) );
  OR2_X1 U7460 ( .A1(n6296), .A2(n6295), .ZN(n6297) );
  NAND2_X1 U7461 ( .A1(n6484), .A2(n6919), .ZN(n6298) );
  OR2_X1 U7462 ( .A1(n7384), .A2(n9017), .ZN(n8748) );
  NAND2_X1 U7463 ( .A1(n7384), .A2(n9017), .ZN(n8732) );
  NAND2_X1 U7464 ( .A1(n7280), .A2(n8663), .ZN(n7389) );
  NAND2_X1 U7465 ( .A1(n7389), .A2(n8732), .ZN(n6310) );
  NAND2_X1 U7466 ( .A1(n6601), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6304) );
  INV_X1 U7467 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7133) );
  OR2_X1 U7468 ( .A1(n8645), .A2(n7133), .ZN(n6303) );
  INV_X2 U7469 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10466) );
  NAND2_X1 U7470 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6300) );
  AND2_X1 U7471 ( .A1(n6312), .A2(n6300), .ZN(n9083) );
  OR2_X1 U7472 ( .A1(n6436), .A2(n9083), .ZN(n6302) );
  INV_X1 U7473 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7123) );
  OR2_X1 U7474 ( .A1(n8649), .A2(n7123), .ZN(n6301) );
  NAND4_X1 U7475 ( .A1(n6304), .A2(n6303), .A3(n6302), .A4(n6301), .ZN(n9148)
         );
  NAND2_X1 U7476 ( .A1(n8643), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6309) );
  NAND2_X1 U7477 ( .A1(n6306), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6307) );
  NAND2_X1 U7478 ( .A1(n6484), .A2(n7134), .ZN(n6308) );
  OAI211_X1 U7479 ( .C1(n6780), .C2(n6319), .A(n6309), .B(n6308), .ZN(n9082)
         );
  NAND2_X1 U7480 ( .A1(n7484), .A2(n9082), .ZN(n8745) );
  INV_X1 U7481 ( .A(n9082), .ZN(n7476) );
  NAND2_X1 U7482 ( .A1(n9148), .A2(n7476), .ZN(n8734) );
  NAND2_X1 U7483 ( .A1(n6310), .A2(n7388), .ZN(n7387) );
  NAND2_X1 U7484 ( .A1(n6601), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6318) );
  INV_X1 U7485 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7490) );
  OR2_X1 U7486 ( .A1(n8645), .A2(n7490), .ZN(n6317) );
  NAND2_X1 U7487 ( .A1(n6312), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6313) );
  AND2_X1 U7488 ( .A1(n6331), .A2(n6313), .ZN(n7208) );
  OR2_X1 U7489 ( .A1(n6436), .A2(n7208), .ZN(n6316) );
  INV_X1 U7490 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6314) );
  OR2_X1 U7491 ( .A1(n8649), .A2(n6314), .ZN(n6315) );
  NAND4_X1 U7492 ( .A1(n6318), .A2(n6317), .A3(n6316), .A4(n6315), .ZN(n9147)
         );
  INV_X4 U7493 ( .A(n6319), .ZN(n8656) );
  NAND2_X1 U7494 ( .A1(n6777), .A2(n8656), .ZN(n6325) );
  INV_X1 U7495 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U7496 ( .A1(n6326), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6321) );
  XNOR2_X1 U7497 ( .A(n6322), .B(n6321), .ZN(n7224) );
  OAI22_X1 U7498 ( .A1(n6305), .A2(n6778), .B1(n6766), .B2(n7224), .ZN(n6323)
         );
  INV_X1 U7499 ( .A(n6323), .ZN(n6324) );
  NAND2_X1 U7500 ( .A1(n6325), .A2(n6324), .ZN(n7492) );
  NAND2_X1 U7501 ( .A1(n7775), .A2(n7492), .ZN(n8746) );
  INV_X1 U7502 ( .A(n7492), .ZN(n7550) );
  NAND2_X1 U7503 ( .A1(n7550), .A2(n9147), .ZN(n8733) );
  NAND2_X1 U7504 ( .A1(n6788), .A2(n8656), .ZN(n6329) );
  INV_X1 U7505 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6791) );
  OAI22_X1 U7506 ( .A1(n6305), .A2(n6791), .B1(n6766), .B2(n7349), .ZN(n6327)
         );
  INV_X1 U7507 ( .A(n6327), .ZN(n6328) );
  NAND2_X1 U7508 ( .A1(n6329), .A2(n6328), .ZN(n7293) );
  NAND2_X1 U7509 ( .A1(n6601), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6337) );
  INV_X1 U7510 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6330) );
  OR2_X1 U7511 ( .A1(n8645), .A2(n6330), .ZN(n6336) );
  NAND2_X1 U7512 ( .A1(n6331), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6332) );
  AND2_X1 U7513 ( .A1(n6349), .A2(n6332), .ZN(n7872) );
  INV_X1 U7514 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6333) );
  OR2_X1 U7515 ( .A1(n8649), .A2(n6333), .ZN(n6334) );
  NAND2_X1 U7516 ( .A1(n7873), .A2(n9146), .ZN(n8736) );
  NAND2_X1 U7517 ( .A1(n7483), .A2(n7293), .ZN(n8751) );
  NAND2_X1 U7518 ( .A1(n6792), .A2(n8656), .ZN(n6345) );
  INV_X1 U7519 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6795) );
  INV_X1 U7520 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6368) );
  NAND2_X1 U7521 ( .A1(n6338), .A2(n6368), .ZN(n6339) );
  NAND2_X1 U7522 ( .A1(n6339), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6341) );
  INV_X1 U7523 ( .A(n6341), .ZN(n6340) );
  NAND2_X1 U7524 ( .A1(n6340), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n6342) );
  INV_X1 U7525 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6369) );
  NAND2_X1 U7526 ( .A1(n6341), .A2(n6369), .ZN(n6355) );
  INV_X1 U7527 ( .A(n7537), .ZN(n7528) );
  OAI22_X1 U7528 ( .A1(n6305), .A2(n6795), .B1(n6766), .B2(n7528), .ZN(n6343)
         );
  INV_X1 U7529 ( .A(n6343), .ZN(n6344) );
  NAND2_X1 U7530 ( .A1(n6601), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6354) );
  INV_X1 U7531 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7813) );
  OR2_X1 U7532 ( .A1(n8645), .A2(n7813), .ZN(n6353) );
  INV_X1 U7533 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6346) );
  OR2_X1 U7534 ( .A1(n8649), .A2(n6346), .ZN(n6352) );
  INV_X1 U7535 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6347) );
  NAND2_X1 U7536 ( .A1(n6349), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6350) );
  AND2_X1 U7537 ( .A1(n6360), .A2(n6350), .ZN(n7514) );
  OR2_X1 U7538 ( .A1(n6436), .A2(n7514), .ZN(n6351) );
  NAND4_X1 U7539 ( .A1(n6354), .A2(n6353), .A3(n6352), .A4(n6351), .ZN(n9145)
         );
  XNOR2_X1 U7540 ( .A(n8705), .B(n8704), .ZN(n7795) );
  NAND2_X1 U7541 ( .A1(n7794), .A2(n8740), .ZN(n7793) );
  OR2_X1 U7542 ( .A1(n8705), .A2(n8704), .ZN(n8755) );
  NAND2_X1 U7543 ( .A1(n7793), .A2(n8755), .ZN(n7982) );
  INV_X1 U7544 ( .A(n7982), .ZN(n6366) );
  NAND2_X1 U7545 ( .A1(n6796), .A2(n8656), .ZN(n6359) );
  NAND2_X1 U7546 ( .A1(n6355), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6356) );
  INV_X1 U7547 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6367) );
  XNOR2_X1 U7548 ( .A(n6356), .B(n6367), .ZN(n7630) );
  OAI22_X1 U7549 ( .A1(n6305), .A2(n6799), .B1(n6766), .B2(n7630), .ZN(n6357)
         );
  INV_X1 U7550 ( .A(n6357), .ZN(n6358) );
  NAND2_X1 U7551 ( .A1(n6601), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6365) );
  INV_X1 U7552 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8002) );
  OR2_X1 U7553 ( .A1(n8645), .A2(n8002), .ZN(n6364) );
  NAND2_X1 U7554 ( .A1(n6360), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6361) );
  AND2_X1 U7555 ( .A1(n6380), .A2(n6361), .ZN(n7609) );
  OR2_X1 U7556 ( .A1(n6436), .A2(n7609), .ZN(n6363) );
  INV_X1 U7557 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7527) );
  OR2_X1 U7558 ( .A1(n8649), .A2(n7527), .ZN(n6362) );
  NAND4_X1 U7559 ( .A1(n6365), .A2(n6364), .A3(n6363), .A4(n6362), .ZN(n9144)
         );
  NAND2_X1 U7560 ( .A1(n8004), .A2(n7673), .ZN(n8707) );
  NAND2_X1 U7561 ( .A1(n6808), .A2(n8656), .ZN(n6375) );
  AND3_X1 U7562 ( .A1(n6369), .A2(n6368), .A3(n6367), .ZN(n6370) );
  NAND2_X1 U7563 ( .A1(n6371), .A2(n6370), .ZN(n6386) );
  NAND2_X1 U7564 ( .A1(n6386), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6372) );
  XNOR2_X1 U7565 ( .A(n6372), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7749) );
  INV_X1 U7566 ( .A(n7749), .ZN(n7740) );
  OAI22_X1 U7567 ( .A1(n6305), .A2(n6809), .B1(n6766), .B2(n7740), .ZN(n6373)
         );
  INV_X1 U7568 ( .A(n6373), .ZN(n6374) );
  NAND2_X1 U7569 ( .A1(n6601), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6385) );
  INV_X1 U7570 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6376) );
  OR2_X1 U7571 ( .A1(n8645), .A2(n6376), .ZN(n6384) );
  INV_X1 U7572 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6377) );
  OR2_X1 U7573 ( .A1(n8649), .A2(n6377), .ZN(n6383) );
  INV_X1 U7574 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6378) );
  NAND2_X1 U7575 ( .A1(n6380), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6381) );
  AND2_X1 U7576 ( .A1(n6392), .A2(n6381), .ZN(n7670) );
  OR2_X1 U7577 ( .A1(n6436), .A2(n7670), .ZN(n6382) );
  NAND4_X1 U7578 ( .A1(n6385), .A2(n6384), .A3(n6383), .A4(n6382), .ZN(n9143)
         );
  NAND2_X1 U7579 ( .A1(n8760), .A2(n8708), .ZN(n8671) );
  NAND2_X1 U7580 ( .A1(n6806), .A2(n8656), .ZN(n6391) );
  NAND2_X1 U7581 ( .A1(n6398), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6388) );
  INV_X1 U7582 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6387) );
  XNOR2_X1 U7583 ( .A(n6388), .B(n6387), .ZN(n7938) );
  OAI22_X1 U7584 ( .A1(n6305), .A2(n6813), .B1(n6766), .B2(n7938), .ZN(n6389)
         );
  INV_X1 U7585 ( .A(n6389), .ZN(n6390) );
  NAND2_X1 U7586 ( .A1(n6601), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6397) );
  INV_X1 U7587 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8015) );
  OR2_X1 U7588 ( .A1(n8645), .A2(n8015), .ZN(n6396) );
  NAND2_X1 U7589 ( .A1(n6392), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6393) );
  AND2_X1 U7590 ( .A1(n6402), .A2(n6393), .ZN(n8014) );
  OR2_X1 U7591 ( .A1(n6436), .A2(n8014), .ZN(n6395) );
  INV_X1 U7592 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7739) );
  OR2_X1 U7593 ( .A1(n8649), .A2(n7739), .ZN(n6394) );
  NAND2_X1 U7594 ( .A1(n8144), .A2(n8057), .ZN(n8762) );
  NAND2_X1 U7595 ( .A1(n6831), .A2(n8656), .ZN(n6400) );
  OAI21_X1 U7596 ( .B1(n6398), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6424) );
  XNOR2_X1 U7597 ( .A(n6424), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10675) );
  AOI22_X1 U7598 ( .A1(n8643), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6484), .B2(
        n10675), .ZN(n6399) );
  NAND2_X1 U7599 ( .A1(n6400), .A2(n6399), .ZN(n8060) );
  NAND2_X1 U7600 ( .A1(n6601), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6408) );
  INV_X1 U7601 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6401) );
  OR2_X1 U7602 ( .A1(n8645), .A2(n6401), .ZN(n6407) );
  NAND2_X1 U7603 ( .A1(n6402), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6403) );
  AND2_X1 U7604 ( .A1(n6417), .A2(n6403), .ZN(n8058) );
  OR2_X1 U7605 ( .A1(n6436), .A2(n8058), .ZN(n6406) );
  INV_X1 U7606 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6404) );
  OR2_X1 U7607 ( .A1(n8649), .A2(n6404), .ZN(n6405) );
  NAND4_X1 U7608 ( .A1(n6408), .A2(n6407), .A3(n6406), .A4(n6405), .ZN(n9141)
         );
  OR2_X1 U7609 ( .A1(n8060), .A2(n8021), .ZN(n8765) );
  NAND2_X1 U7610 ( .A1(n8060), .A2(n8021), .ZN(n8763) );
  NAND2_X1 U7611 ( .A1(n8054), .A2(n8675), .ZN(n6409) );
  NAND2_X1 U7612 ( .A1(n6893), .A2(n8656), .ZN(n6415) );
  INV_X1 U7613 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6894) );
  NAND2_X1 U7614 ( .A1(n6424), .A2(n6410), .ZN(n6411) );
  NAND2_X1 U7615 ( .A1(n6411), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6412) );
  XNOR2_X1 U7616 ( .A(n6412), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7941) );
  INV_X1 U7617 ( .A(n7941), .ZN(n8154) );
  OAI22_X1 U7618 ( .A1(n6305), .A2(n6894), .B1(n6766), .B2(n8154), .ZN(n6413)
         );
  INV_X1 U7619 ( .A(n6413), .ZN(n6414) );
  NAND2_X1 U7620 ( .A1(n6601), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6423) );
  INV_X1 U7621 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8134) );
  OR2_X1 U7622 ( .A1(n8645), .A2(n8134), .ZN(n6422) );
  INV_X1 U7623 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10545) );
  NAND2_X1 U7624 ( .A1(n6417), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6418) );
  AND2_X1 U7625 ( .A1(n6434), .A2(n6418), .ZN(n8133) );
  OR2_X1 U7626 ( .A1(n6436), .A2(n8133), .ZN(n6421) );
  INV_X1 U7627 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6419) );
  OR2_X1 U7628 ( .A1(n8649), .A2(n6419), .ZN(n6420) );
  NAND4_X1 U7629 ( .A1(n6423), .A2(n6422), .A3(n6421), .A4(n6420), .ZN(n9140)
         );
  INV_X1 U7630 ( .A(n9140), .ZN(n9470) );
  NAND2_X1 U7631 ( .A1(n8768), .A2(n9470), .ZN(n8769) );
  NAND2_X1 U7632 ( .A1(n6898), .A2(n8656), .ZN(n6429) );
  INV_X1 U7633 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6985) );
  NOR2_X1 U7634 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n6425) );
  OAI21_X1 U7635 ( .B1(n6425), .B2(n9613), .A(n6424), .ZN(n6441) );
  INV_X1 U7636 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6426) );
  XNOR2_X1 U7637 ( .A(n6441), .B(n6426), .ZN(n9167) );
  INV_X1 U7638 ( .A(n9167), .ZN(n9158) );
  OAI22_X1 U7639 ( .A1(n6305), .A2(n6985), .B1(n9158), .B2(n6766), .ZN(n6427)
         );
  INV_X1 U7640 ( .A(n6427), .ZN(n6428) );
  NAND2_X1 U7641 ( .A1(n6601), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6440) );
  INV_X1 U7642 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6430) );
  OR2_X1 U7643 ( .A1(n8645), .A2(n6430), .ZN(n6439) );
  INV_X1 U7644 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6431) );
  OR2_X1 U7645 ( .A1(n8649), .A2(n6431), .ZN(n6438) );
  INV_X1 U7646 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6432) );
  NAND2_X1 U7647 ( .A1(n6434), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6435) );
  AND2_X1 U7648 ( .A1(n6459), .A2(n6435), .ZN(n9474) );
  OR2_X1 U7649 ( .A1(n6436), .A2(n9474), .ZN(n6437) );
  OR2_X1 U7650 ( .A1(n9567), .A2(n8239), .ZN(n8775) );
  NAND2_X1 U7651 ( .A1(n6986), .A2(n8656), .ZN(n6444) );
  OR2_X1 U7652 ( .A1(n6441), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U7653 ( .A1(n6442), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6454) );
  XNOR2_X1 U7654 ( .A(n6454), .B(P2_IR_REG_14__SCAN_IN), .ZN(n9170) );
  AOI22_X1 U7655 ( .A1(n8643), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6484), .B2(
        n9170), .ZN(n6443) );
  NAND2_X1 U7656 ( .A1(n6601), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6449) );
  INV_X1 U7657 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9171) );
  OR2_X1 U7658 ( .A1(n8645), .A2(n9171), .ZN(n6448) );
  XNOR2_X1 U7659 ( .A(n6459), .B(n10542), .ZN(n10839) );
  OR2_X1 U7660 ( .A1(n6436), .A2(n10839), .ZN(n6447) );
  INV_X1 U7661 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6445) );
  OR2_X1 U7662 ( .A1(n8649), .A2(n6445), .ZN(n6446) );
  NAND4_X1 U7663 ( .A1(n6449), .A2(n6448), .A3(n6447), .A4(n6446), .ZN(n9139)
         );
  NAND2_X1 U7664 ( .A1(n8780), .A2(n9139), .ZN(n8791) );
  OR2_X1 U7665 ( .A1(n8780), .A2(n9139), .ZN(n6450) );
  INV_X1 U7666 ( .A(n9139), .ZN(n9472) );
  OR2_X1 U7667 ( .A1(n8780), .A2(n9472), .ZN(n6451) );
  NAND2_X1 U7668 ( .A1(n6452), .A2(n6451), .ZN(n9454) );
  NAND2_X1 U7669 ( .A1(n7072), .A2(n8656), .ZN(n6457) );
  NAND2_X1 U7670 ( .A1(n6454), .A2(n6453), .ZN(n6455) );
  NAND2_X1 U7671 ( .A1(n6455), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6468) );
  XNOR2_X1 U7672 ( .A(n6468), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9213) );
  AOI22_X1 U7673 ( .A1(n6484), .A2(n9213), .B1(n8643), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6456) );
  INV_X1 U7674 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8272) );
  OAI21_X1 U7675 ( .B1(n8272), .B2(n6460), .A(n6475), .ZN(n9459) );
  NAND2_X1 U7676 ( .A1(n6458), .A2(n9459), .ZN(n6466) );
  INV_X1 U7677 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9461) );
  OR2_X1 U7678 ( .A1(n8645), .A2(n9461), .ZN(n6465) );
  INV_X1 U7679 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6461) );
  OR2_X1 U7680 ( .A1(n8649), .A2(n6461), .ZN(n6464) );
  INV_X1 U7681 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n6462) );
  OR2_X1 U7682 ( .A1(n8647), .A2(n6462), .ZN(n6463) );
  NAND4_X1 U7683 ( .A1(n6466), .A2(n6465), .A3(n6464), .A4(n6463), .ZN(n9551)
         );
  INV_X1 U7684 ( .A(n9551), .ZN(n10576) );
  NAND2_X1 U7685 ( .A1(n9545), .A2(n10576), .ZN(n8784) );
  NAND2_X1 U7686 ( .A1(n7318), .A2(n8656), .ZN(n6474) );
  INV_X1 U7687 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U7688 ( .A1(n6468), .A2(n6467), .ZN(n6469) );
  NAND2_X1 U7689 ( .A1(n6469), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U7690 ( .A1(n6471), .A2(n6470), .ZN(n6482) );
  OR2_X1 U7691 ( .A1(n6471), .A2(n6470), .ZN(n6472) );
  AND2_X1 U7692 ( .A1(n6482), .A2(n6472), .ZN(n9207) );
  AOI22_X1 U7693 ( .A1(n9207), .A2(n6484), .B1(n8643), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n6473) );
  AND2_X1 U7694 ( .A1(n6475), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6476) );
  OR2_X1 U7695 ( .A1(n6476), .A2(n6490), .ZN(n9442) );
  NAND2_X1 U7696 ( .A1(n9442), .A2(n6458), .ZN(n6480) );
  INV_X1 U7697 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9444) );
  OR2_X1 U7698 ( .A1(n8645), .A2(n9444), .ZN(n6479) );
  NAND2_X1 U7699 ( .A1(n6601), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6478) );
  INV_X1 U7700 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9202) );
  OR2_X1 U7701 ( .A1(n8649), .A2(n9202), .ZN(n6477) );
  NAND4_X1 U7702 ( .A1(n6480), .A2(n6479), .A3(n6478), .A4(n6477), .ZN(n9428)
         );
  INV_X1 U7703 ( .A(n9428), .ZN(n9458) );
  NAND2_X1 U7704 ( .A1(n9538), .A2(n9458), .ZN(n8794) );
  NAND2_X1 U7705 ( .A1(n8795), .A2(n8794), .ZN(n9446) );
  INV_X1 U7706 ( .A(n8784), .ZN(n9447) );
  NOR2_X1 U7707 ( .A1(n9446), .A2(n9447), .ZN(n6481) );
  NAND2_X1 U7708 ( .A1(n7365), .A2(n8656), .ZN(n6486) );
  NAND2_X1 U7709 ( .A1(n6482), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6483) );
  XNOR2_X1 U7710 ( .A(n6483), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9246) );
  AOI22_X1 U7711 ( .A1(n9246), .A2(n6484), .B1(n8643), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n6485) );
  INV_X1 U7712 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n6487) );
  OR2_X1 U7713 ( .A1(n8647), .A2(n6487), .ZN(n6489) );
  INV_X1 U7714 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9432) );
  OR2_X1 U7715 ( .A1(n8645), .A2(n9432), .ZN(n6488) );
  AND2_X1 U7716 ( .A1(n6489), .A2(n6488), .ZN(n6494) );
  INV_X1 U7717 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10457) );
  OR2_X1 U7718 ( .A1(n6490), .A2(n10457), .ZN(n6491) );
  NAND2_X1 U7719 ( .A1(n6502), .A2(n6491), .ZN(n9430) );
  NAND2_X1 U7720 ( .A1(n9430), .A2(n6458), .ZN(n6493) );
  INV_X1 U7721 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9226) );
  OR2_X1 U7722 ( .A1(n8649), .A2(n9226), .ZN(n6492) );
  XNOR2_X1 U7723 ( .A(n9534), .B(n9060), .ZN(n6639) );
  INV_X1 U7724 ( .A(n6639), .ZN(n9434) );
  OR2_X1 U7725 ( .A1(n9534), .A2(n9060), .ZN(n6495) );
  NAND2_X1 U7726 ( .A1(n7469), .A2(n8656), .ZN(n6501) );
  NAND2_X1 U7727 ( .A1(n6496), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6498) );
  INV_X1 U7728 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6497) );
  XNOR2_X1 U7729 ( .A(n6498), .B(n6497), .ZN(n10705) );
  OAI22_X1 U7730 ( .A1(n6305), .A2(n7472), .B1(n6766), .B2(n10705), .ZN(n6499)
         );
  INV_X1 U7731 ( .A(n6499), .ZN(n6500) );
  NAND2_X1 U7732 ( .A1(n6502), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U7733 ( .A1(n6512), .A2(n6503), .ZN(n9417) );
  NAND2_X1 U7734 ( .A1(n9417), .A2(n6458), .ZN(n6508) );
  INV_X1 U7735 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9257) );
  NAND2_X1 U7736 ( .A1(n6621), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6505) );
  NAND2_X1 U7737 ( .A1(n6601), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6504) );
  OAI211_X1 U7738 ( .C1(n9257), .C2(n8649), .A(n6505), .B(n6504), .ZN(n6506)
         );
  INV_X1 U7739 ( .A(n6506), .ZN(n6507) );
  NAND2_X1 U7740 ( .A1(n6508), .A2(n6507), .ZN(n9427) );
  INV_X1 U7741 ( .A(n9427), .ZN(n9406) );
  NAND2_X1 U7742 ( .A1(n9530), .A2(n9406), .ZN(n8808) );
  NAND2_X1 U7743 ( .A1(n7599), .A2(n8656), .ZN(n6511) );
  OAI22_X1 U7744 ( .A1(n6305), .A2(n7600), .B1(n6766), .B2(n8696), .ZN(n6509)
         );
  INV_X1 U7745 ( .A(n6509), .ZN(n6510) );
  AND2_X1 U7746 ( .A1(n6512), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6513) );
  OR2_X1 U7747 ( .A1(n6513), .A2(n6522), .ZN(n9408) );
  NAND2_X1 U7748 ( .A1(n9408), .A2(n6458), .ZN(n6519) );
  INV_X1 U7749 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9410) );
  INV_X1 U7750 ( .A(n8649), .ZN(n6514) );
  NAND2_X1 U7751 ( .A1(n6514), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6516) );
  NAND2_X1 U7752 ( .A1(n6601), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6515) );
  OAI211_X1 U7753 ( .C1(n8645), .C2(n9410), .A(n6516), .B(n6515), .ZN(n6517)
         );
  INV_X1 U7754 ( .A(n6517), .ZN(n6518) );
  NAND2_X1 U7755 ( .A1(n9523), .A2(n9113), .ZN(n8811) );
  NAND2_X1 U7756 ( .A1(n8810), .A2(n8811), .ZN(n8607) );
  NAND2_X1 U7757 ( .A1(n9399), .A2(n8810), .ZN(n9383) );
  NAND2_X1 U7758 ( .A1(n7695), .A2(n8656), .ZN(n6521) );
  NAND2_X1 U7759 ( .A1(n8643), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6520) );
  NAND2_X2 U7760 ( .A1(n6521), .A2(n6520), .ZN(n9519) );
  INV_X1 U7761 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9093) );
  NOR2_X1 U7762 ( .A1(n6522), .A2(n9093), .ZN(n6523) );
  OR2_X1 U7763 ( .A1(n6532), .A2(n6523), .ZN(n9384) );
  NAND2_X1 U7764 ( .A1(n9384), .A2(n6458), .ZN(n6529) );
  INV_X1 U7765 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U7766 ( .A1(n6601), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6525) );
  NAND2_X1 U7767 ( .A1(n6621), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6524) );
  OAI211_X1 U7768 ( .C1(n6526), .C2(n8649), .A(n6525), .B(n6524), .ZN(n6527)
         );
  INV_X1 U7769 ( .A(n6527), .ZN(n6528) );
  NAND2_X1 U7770 ( .A1(n9519), .A2(n9407), .ZN(n8816) );
  NAND2_X1 U7771 ( .A1(n9383), .A2(n9388), .ZN(n9382) );
  NAND2_X1 U7772 ( .A1(n9382), .A2(n8815), .ZN(n9376) );
  NAND2_X1 U7773 ( .A1(n7790), .A2(n8656), .ZN(n6531) );
  NAND2_X1 U7774 ( .A1(n8643), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6530) );
  INV_X1 U7775 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10544) );
  OR2_X1 U7776 ( .A1(n6532), .A2(n10544), .ZN(n6533) );
  NAND2_X1 U7777 ( .A1(n6542), .A2(n6533), .ZN(n9374) );
  NAND2_X1 U7778 ( .A1(n9374), .A2(n6458), .ZN(n6538) );
  INV_X1 U7779 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9517) );
  NAND2_X1 U7780 ( .A1(n6601), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6535) );
  NAND2_X1 U7781 ( .A1(n6621), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6534) );
  OAI211_X1 U7782 ( .C1(n9517), .C2(n8649), .A(n6535), .B(n6534), .ZN(n6536)
         );
  INV_X1 U7783 ( .A(n6536), .ZN(n6537) );
  NAND2_X1 U7784 ( .A1(n6538), .A2(n6537), .ZN(n9391) );
  NAND2_X1 U7785 ( .A1(n9375), .A2(n9391), .ZN(n8701) );
  INV_X1 U7786 ( .A(n9391), .ZN(n9095) );
  OR2_X1 U7787 ( .A1(n9375), .A2(n9095), .ZN(n6539) );
  NAND2_X1 U7788 ( .A1(n9515), .A2(n6539), .ZN(n9356) );
  NAND2_X1 U7789 ( .A1(n7879), .A2(n8656), .ZN(n6541) );
  NAND2_X1 U7790 ( .A1(n8643), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6540) );
  NAND2_X1 U7791 ( .A1(n6542), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6543) );
  NAND2_X1 U7792 ( .A1(n6551), .A2(n6543), .ZN(n9358) );
  NAND2_X1 U7793 ( .A1(n9358), .A2(n6458), .ZN(n6548) );
  INV_X1 U7794 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U7795 ( .A1(n6621), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6545) );
  NAND2_X1 U7796 ( .A1(n6601), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6544) );
  OAI211_X1 U7797 ( .C1(n8649), .C2(n9511), .A(n6545), .B(n6544), .ZN(n6546)
         );
  INV_X1 U7798 ( .A(n6546), .ZN(n6547) );
  NAND2_X1 U7799 ( .A1(n6548), .A2(n6547), .ZN(n9338) );
  OR2_X1 U7800 ( .A1(n9101), .A2(n9373), .ZN(n8824) );
  NAND2_X2 U7801 ( .A1(n9357), .A2(n8824), .ZN(n9341) );
  NAND2_X1 U7802 ( .A1(n7909), .A2(n8656), .ZN(n6550) );
  NAND2_X1 U7803 ( .A1(n8643), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U7804 ( .A1(n6551), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U7805 ( .A1(n6561), .A2(n6552), .ZN(n9342) );
  NAND2_X1 U7806 ( .A1(n9342), .A2(n6458), .ZN(n6558) );
  INV_X1 U7807 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n6555) );
  NAND2_X1 U7808 ( .A1(n6601), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U7809 ( .A1(n6621), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6553) );
  OAI211_X1 U7810 ( .C1(n6555), .C2(n8649), .A(n6554), .B(n6553), .ZN(n6556)
         );
  INV_X1 U7811 ( .A(n6556), .ZN(n6557) );
  NOR2_X1 U7812 ( .A1(n9503), .A2(n9330), .ZN(n8828) );
  NAND2_X1 U7813 ( .A1(n9503), .A2(n9330), .ZN(n8662) );
  NAND2_X1 U7814 ( .A1(n8033), .A2(n8656), .ZN(n6560) );
  NAND2_X1 U7815 ( .A1(n8643), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6559) );
  AND2_X1 U7816 ( .A1(n6561), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6562) );
  OR2_X1 U7817 ( .A1(n6562), .A2(n6569), .ZN(n9332) );
  INV_X1 U7818 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9501) );
  NAND2_X1 U7819 ( .A1(n6601), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6564) );
  NAND2_X1 U7820 ( .A1(n6621), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6563) );
  OAI211_X1 U7821 ( .C1(n9501), .C2(n8649), .A(n6564), .B(n6563), .ZN(n6565)
         );
  XNOR2_X1 U7822 ( .A(n8698), .B(n9316), .ZN(n9326) );
  NAND2_X1 U7823 ( .A1(n8051), .A2(n8656), .ZN(n6567) );
  NAND2_X1 U7824 ( .A1(n8643), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6566) );
  INV_X1 U7825 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6568) );
  OR2_X1 U7826 ( .A1(n6569), .A2(n6568), .ZN(n6570) );
  NAND2_X1 U7827 ( .A1(n6578), .A2(n6570), .ZN(n9320) );
  NAND2_X1 U7828 ( .A1(n9320), .A2(n6458), .ZN(n6575) );
  INV_X1 U7829 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9497) );
  NAND2_X1 U7830 ( .A1(n6621), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6572) );
  NAND2_X1 U7831 ( .A1(n6601), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6571) );
  OAI211_X1 U7832 ( .C1(n8649), .C2(n9497), .A(n6572), .B(n6571), .ZN(n6573)
         );
  INV_X1 U7833 ( .A(n6573), .ZN(n6574) );
  NAND2_X1 U7834 ( .A1(n9318), .A2(n9329), .ZN(n8661) );
  NAND2_X1 U7835 ( .A1(n8643), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6576) );
  NAND2_X1 U7836 ( .A1(n6578), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6579) );
  NAND2_X1 U7837 ( .A1(n6598), .A2(n6579), .ZN(n9309) );
  NAND2_X1 U7838 ( .A1(n9309), .A2(n6458), .ZN(n6584) );
  INV_X1 U7839 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9493) );
  NAND2_X1 U7840 ( .A1(n6621), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6581) );
  NAND2_X1 U7841 ( .A1(n6601), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6580) );
  OAI211_X1 U7842 ( .C1(n9493), .C2(n8649), .A(n6581), .B(n6580), .ZN(n6582)
         );
  INV_X1 U7843 ( .A(n6582), .ZN(n6583) );
  NAND2_X1 U7844 ( .A1(n8993), .A2(n8656), .ZN(n6586) );
  NAND2_X1 U7845 ( .A1(n8643), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6585) );
  NAND2_X1 U7846 ( .A1(n6601), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6594) );
  INV_X1 U7847 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n9289) );
  OR2_X1 U7848 ( .A1(n8645), .A2(n9289), .ZN(n6593) );
  INV_X1 U7849 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6587) );
  NAND2_X1 U7850 ( .A1(n6587), .A2(n6588), .ZN(n8588) );
  INV_X1 U7851 ( .A(n6588), .ZN(n6599) );
  NAND2_X1 U7852 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(n6599), .ZN(n6589) );
  OR2_X1 U7853 ( .A1(n6436), .A2(n9288), .ZN(n6592) );
  INV_X1 U7854 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6590) );
  OR2_X1 U7855 ( .A1(n8649), .A2(n6590), .ZN(n6591) );
  NAND2_X2 U7856 ( .A1(n6608), .A2(n6611), .ZN(n9285) );
  INV_X1 U7857 ( .A(n9285), .ZN(n6595) );
  AOI22_X1 U7858 ( .A1(n6610), .A2(n6595), .B1(n8836), .B2(n6611), .ZN(n6609)
         );
  NAND2_X1 U7859 ( .A1(n8264), .A2(n8656), .ZN(n6597) );
  NAND2_X1 U7860 ( .A1(n8643), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U7861 ( .A1(n6598), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6600) );
  NAND2_X1 U7862 ( .A1(n6600), .A2(n6599), .ZN(n9298) );
  NAND2_X1 U7863 ( .A1(n9298), .A2(n6458), .ZN(n6606) );
  INV_X1 U7864 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9489) );
  NAND2_X1 U7865 ( .A1(n6621), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U7866 ( .A1(n6601), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6602) );
  OAI211_X1 U7867 ( .C1(n9489), .C2(n8649), .A(n6603), .B(n6602), .ZN(n6604)
         );
  INV_X1 U7868 ( .A(n6604), .ZN(n6605) );
  INV_X1 U7869 ( .A(n8660), .ZN(n8839) );
  NAND2_X1 U7870 ( .A1(n6611), .A2(n8839), .ZN(n6607) );
  OAI211_X1 U7871 ( .C1(n6609), .C2(n8840), .A(n6608), .B(n6607), .ZN(n6627)
         );
  INV_X1 U7872 ( .A(n6614), .ZN(n6615) );
  NAND2_X1 U7873 ( .A1(n6615), .A2(n10491), .ZN(n6616) );
  INV_X1 U7874 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n6618) );
  INV_X1 U7875 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10351) );
  MUX2_X1 U7876 ( .A(n6618), .B(n10351), .S(n8328), .Z(n8279) );
  NAND2_X1 U7877 ( .A1(n9619), .A2(n8656), .ZN(n6620) );
  NAND2_X1 U7878 ( .A1(n8643), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6619) );
  NAND2_X1 U7879 ( .A1(n6621), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6624) );
  INV_X1 U7880 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6760) );
  OR2_X1 U7881 ( .A1(n8649), .A2(n6760), .ZN(n6623) );
  INV_X1 U7882 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6711) );
  OR2_X1 U7883 ( .A1(n8647), .A2(n6711), .ZN(n6622) );
  NAND4_X1 U7884 ( .A1(n8653), .A2(n6624), .A3(n6623), .A4(n6622), .ZN(n9282)
         );
  INV_X1 U7885 ( .A(n9282), .ZN(n6625) );
  NAND2_X1 U7886 ( .A1(n6712), .A2(n6625), .ZN(n8688) );
  NOR2_X1 U7887 ( .A1(n8302), .A2(n7194), .ZN(n7076) );
  NOR2_X1 U7888 ( .A1(n9151), .A2(n7359), .ZN(n7099) );
  NOR2_X1 U7889 ( .A1(n7282), .A2(n7384), .ZN(n6631) );
  INV_X1 U7890 ( .A(n7282), .ZN(n6630) );
  OAI22_X1 U7891 ( .A1(n6631), .A2(n9017), .B1(n6630), .B2(n9149), .ZN(n7383)
         );
  INV_X1 U7892 ( .A(n8705), .ZN(n7844) );
  NAND2_X1 U7893 ( .A1(n8144), .A2(n9142), .ZN(n8008) );
  INV_X1 U7894 ( .A(n8060), .ZN(n8063) );
  NAND2_X1 U7895 ( .A1(n8768), .A2(n9140), .ZN(n6634) );
  INV_X1 U7896 ( .A(n9467), .ZN(n6636) );
  INV_X1 U7897 ( .A(n8239), .ZN(n9554) );
  NAND2_X1 U7898 ( .A1(n9550), .A2(n9549), .ZN(n9548) );
  NAND2_X1 U7899 ( .A1(n9538), .A2(n9428), .ZN(n6637) );
  INV_X1 U7900 ( .A(n9060), .ZN(n9440) );
  NAND2_X1 U7901 ( .A1(n9534), .A2(n9440), .ZN(n6640) );
  INV_X1 U7902 ( .A(n9530), .ZN(n9115) );
  NOR2_X1 U7903 ( .A1(n9115), .A2(n9406), .ZN(n9400) );
  INV_X1 U7904 ( .A(n9113), .ZN(n9415) );
  AND2_X1 U7905 ( .A1(n9523), .A2(n9415), .ZN(n6643) );
  OR2_X1 U7906 ( .A1(n9400), .A2(n6643), .ZN(n9385) );
  INV_X1 U7907 ( .A(n9519), .ZN(n9100) );
  NAND2_X1 U7908 ( .A1(n9100), .A2(n9407), .ZN(n9369) );
  NAND2_X1 U7909 ( .A1(n9115), .A2(n9406), .ZN(n9401) );
  AND2_X1 U7910 ( .A1(n5033), .A2(n9401), .ZN(n6642) );
  OR2_X1 U7911 ( .A1(n6643), .A2(n6642), .ZN(n9386) );
  AND2_X1 U7912 ( .A1(n9369), .A2(n9367), .ZN(n6644) );
  NAND2_X1 U7913 ( .A1(n9503), .A2(n9353), .ZN(n6647) );
  NOR2_X1 U7914 ( .A1(n9503), .A2(n9353), .ZN(n6646) );
  NAND2_X1 U7915 ( .A1(n5510), .A2(n9316), .ZN(n6648) );
  NAND2_X1 U7916 ( .A1(n9327), .A2(n6648), .ZN(n6650) );
  NAND2_X1 U7917 ( .A1(n8698), .A2(n5509), .ZN(n6649) );
  NOR2_X1 U7918 ( .A1(n9589), .A2(n9329), .ZN(n6652) );
  NAND2_X1 U7919 ( .A1(n9589), .A2(n9329), .ZN(n6651) );
  NOR2_X1 U7920 ( .A1(n9581), .A2(n9305), .ZN(n6654) );
  NAND2_X1 U7921 ( .A1(n9581), .A2(n9305), .ZN(n6653) );
  INV_X1 U7922 ( .A(n9295), .ZN(n9136) );
  NOR2_X1 U7923 ( .A1(n9483), .A2(n9136), .ZN(n6655) );
  INV_X1 U7924 ( .A(n9483), .ZN(n9287) );
  XNOR2_X1 U7925 ( .A(n6656), .B(n8686), .ZN(n6659) );
  OR2_X1 U7926 ( .A1(n8712), .A2(n7696), .ZN(n6658) );
  AND2_X1 U7927 ( .A1(n8867), .A2(n9266), .ZN(n6697) );
  INV_X1 U7928 ( .A(n6697), .ZN(n6657) );
  NAND2_X1 U7929 ( .A1(n6658), .A2(n6657), .ZN(n9547) );
  NAND2_X1 U7930 ( .A1(n6659), .A2(n9547), .ZN(n6668) );
  OAI21_X1 U7931 ( .B1(n8864), .B2(n4946), .A(n6766), .ZN(n6861) );
  NOR2_X2 U7932 ( .A1(n6861), .A2(n8842), .ZN(n9553) );
  NAND2_X1 U7933 ( .A1(n6861), .A2(n8849), .ZN(n9473) );
  AND2_X1 U7934 ( .A1(n6766), .A2(P2_B_REG_SCAN_IN), .ZN(n6660) );
  NOR2_X1 U7935 ( .A1(n9473), .A2(n6660), .ZN(n9274) );
  INV_X1 U7936 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6661) );
  OR2_X1 U7937 ( .A1(n8647), .A2(n6661), .ZN(n6666) );
  INV_X1 U7938 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6662) );
  OR2_X1 U7939 ( .A1(n8645), .A2(n6662), .ZN(n6665) );
  INV_X1 U7940 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6663) );
  OR2_X1 U7941 ( .A1(n8649), .A2(n6663), .ZN(n6664) );
  NAND4_X1 U7942 ( .A1(n8653), .A2(n6666), .A3(n6665), .A4(n6664), .ZN(n9135)
         );
  AOI22_X1 U7943 ( .A1(n9136), .A2(n9553), .B1(n9274), .B2(n9135), .ZN(n6667)
         );
  NAND2_X1 U7944 ( .A1(n7696), .A2(n9266), .ZN(n7371) );
  OR2_X1 U7945 ( .A1(n7371), .A2(n8867), .ZN(n8141) );
  NOR2_X1 U7946 ( .A1(n8594), .A2(n8141), .ZN(n6669) );
  INV_X1 U7947 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6670) );
  NAND2_X1 U7948 ( .A1(n6709), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6672) );
  INV_X1 U7949 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6671) );
  XNOR2_X1 U7950 ( .A(n6703), .B(P2_B_REG_SCAN_IN), .ZN(n6676) );
  INV_X1 U7951 ( .A(n6709), .ZN(n6673) );
  NAND2_X1 U7952 ( .A1(n6673), .A2(n6671), .ZN(n6677) );
  NAND2_X1 U7953 ( .A1(n6677), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6675) );
  INV_X1 U7954 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6674) );
  XNOR2_X1 U7955 ( .A(n6675), .B(n6674), .ZN(n6702) );
  NAND2_X1 U7956 ( .A1(n6676), .A2(n6702), .ZN(n6679) );
  OAI21_X2 U7957 ( .B1(n6677), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6678) );
  XNOR2_X2 U7958 ( .A(n6678), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6704) );
  INV_X1 U7959 ( .A(n6704), .ZN(n6683) );
  NAND2_X1 U7960 ( .A1(n6683), .A2(n6703), .ZN(n6680) );
  OR2_X1 U7961 ( .A1(n6682), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6685) );
  NAND2_X1 U7962 ( .A1(n6683), .A2(n6702), .ZN(n6684) );
  AND2_X1 U7963 ( .A1(n7182), .A2(n9612), .ZN(n6752) );
  NOR2_X1 U7964 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6689) );
  NOR4_X1 U7965 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6688) );
  NOR4_X1 U7966 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6687) );
  NOR4_X1 U7967 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6686) );
  NAND4_X1 U7968 ( .A1(n6689), .A2(n6688), .A3(n6687), .A4(n6686), .ZN(n6695)
         );
  NOR4_X1 U7969 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6693) );
  NOR4_X1 U7970 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6692) );
  NOR4_X1 U7971 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6691) );
  NOR4_X1 U7972 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6690) );
  NAND4_X1 U7973 ( .A1(n6693), .A2(n6692), .A3(n6691), .A4(n6690), .ZN(n6694)
         );
  NOR2_X1 U7974 ( .A1(n6695), .A2(n6694), .ZN(n6696) );
  OR2_X1 U7975 ( .A1(n6682), .A2(n6696), .ZN(n6750) );
  NAND2_X1 U7976 ( .A1(n6752), .A2(n6750), .ZN(n6872) );
  INV_X1 U7977 ( .A(n7696), .ZN(n8862) );
  AND3_X1 U7978 ( .A1(n8712), .A2(n8862), .A3(n6697), .ZN(n6848) );
  INV_X1 U7979 ( .A(n6848), .ZN(n6870) );
  AND2_X1 U7980 ( .A1(n6870), .A2(n7188), .ZN(n6701) );
  INV_X1 U7981 ( .A(n9612), .ZN(n6756) );
  NAND3_X1 U7982 ( .A1(n6681), .A2(n6756), .A3(n6750), .ZN(n6855) );
  INV_X1 U7983 ( .A(n6855), .ZN(n6699) );
  NAND2_X1 U7984 ( .A1(n8842), .A2(n9559), .ZN(n6871) );
  OR2_X1 U7985 ( .A1(n6871), .A2(n6848), .ZN(n6698) );
  INV_X1 U7986 ( .A(n7371), .ZN(n8859) );
  OR2_X1 U7987 ( .A1(n9559), .A2(n8859), .ZN(n10840) );
  NAND2_X1 U7988 ( .A1(n6698), .A2(n10840), .ZN(n6846) );
  NAND2_X1 U7989 ( .A1(n6699), .A2(n6846), .ZN(n6700) );
  OAI21_X1 U7990 ( .B1(n6872), .B2(n6701), .A(n6700), .ZN(n6713) );
  INV_X1 U7991 ( .A(n6702), .ZN(n8052) );
  INV_X1 U7992 ( .A(n6703), .ZN(n8034) );
  AND2_X1 U7993 ( .A1(n8052), .A2(n8034), .ZN(n6705) );
  NAND2_X1 U7994 ( .A1(n6705), .A2(n6704), .ZN(n6910) );
  INV_X1 U7995 ( .A(n6706), .ZN(n6707) );
  NAND2_X1 U7996 ( .A1(n6707), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6708) );
  MUX2_X1 U7997 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6708), .S(
        P2_IR_REG_23__SCAN_IN), .Z(n6710) );
  NAND2_X1 U7998 ( .A1(n6710), .A2(n6709), .ZN(n6909) );
  AND2_X1 U7999 ( .A1(n6909), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6768) );
  NAND2_X1 U8000 ( .A1(n6910), .A2(n6768), .ZN(n9611) );
  INV_X1 U8001 ( .A(n9611), .ZN(n6873) );
  AND2_X2 U8002 ( .A1(n6713), .A2(n6873), .ZN(n10852) );
  NOR2_X1 U8003 ( .A1(n10852), .A2(n6711), .ZN(n6715) );
  NOR2_X1 U8004 ( .A1(n9611), .A2(n9559), .ZN(n6857) );
  NAND2_X1 U8005 ( .A1(n6713), .A2(n6857), .ZN(n9606) );
  NOR2_X1 U8006 ( .A1(n6715), .A2(n6714), .ZN(n6716) );
  NOR2_X1 U8007 ( .A1(n9983), .A2(n9792), .ZN(n6717) );
  NAND2_X1 U8008 ( .A1(n9619), .A2(n8333), .ZN(n6720) );
  OR2_X1 U8009 ( .A1(n8287), .A2(n10351), .ZN(n6719) );
  NAND2_X1 U8010 ( .A1(n6734), .A2(n9979), .ZN(n8503) );
  XNOR2_X1 U8011 ( .A(n6722), .B(n6721), .ZN(n9966) );
  AND2_X1 U8012 ( .A1(n6723), .A2(n8502), .ZN(n6724) );
  INV_X1 U8013 ( .A(P1_B_REG_SCAN_IN), .ZN(n6725) );
  NOR2_X1 U8014 ( .A1(n8304), .A2(n6725), .ZN(n6726) );
  OR2_X1 U8015 ( .A1(n10794), .A2(n6726), .ZN(n8298) );
  NAND2_X1 U8016 ( .A1(n8292), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6731) );
  INV_X1 U8017 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9960) );
  OR2_X1 U8018 ( .A1(n6727), .A2(n9960), .ZN(n6730) );
  INV_X1 U8019 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n6728) );
  OR2_X1 U8020 ( .A1(n8294), .A2(n6728), .ZN(n6729) );
  AND3_X1 U8021 ( .A1(n6731), .A2(n6730), .A3(n6729), .ZN(n8439) );
  OAI22_X1 U8022 ( .A1(n8298), .A2(n8439), .B1(n10205), .B2(n10796), .ZN(n6732) );
  INV_X1 U8023 ( .A(n6735), .ZN(n6736) );
  OAI211_X1 U8024 ( .C1(n6747), .C2(n6736), .A(n10782), .B(n8289), .ZN(n9969)
         );
  INV_X1 U8025 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6738) );
  NOR2_X1 U8026 ( .A1(n10834), .A2(n6738), .ZN(n6739) );
  NOR2_X1 U8027 ( .A1(n6737), .A2(n6739), .ZN(n6740) );
  OAI21_X1 U8028 ( .B1(n6749), .B2(n6207), .A(n6740), .ZN(P1_U3519) );
  AND2_X1 U8029 ( .A1(n6741), .A2(n7014), .ZN(n6743) );
  AND2_X2 U8030 ( .A1(n6743), .A2(n6742), .ZN(n10831) );
  NAND2_X1 U8031 ( .A1(n10831), .A2(n10283), .ZN(n10298) );
  NAND2_X1 U8032 ( .A1(n6873), .A2(n6750), .ZN(n6751) );
  NOR2_X1 U8033 ( .A1(n6752), .A2(n6751), .ZN(n7186) );
  OAI21_X1 U8034 ( .B1(n8693), .B2(n8141), .A(n7182), .ZN(n6757) );
  OR2_X1 U8035 ( .A1(n8842), .A2(n8860), .ZN(n6847) );
  INV_X1 U8036 ( .A(n6753), .ZN(n6754) );
  OR2_X1 U8037 ( .A1(n6754), .A2(n7696), .ZN(n6755) );
  NAND2_X1 U8038 ( .A1(n8842), .A2(n6755), .ZN(n7178) );
  NAND2_X1 U8039 ( .A1(n6847), .A2(n7178), .ZN(n7180) );
  AOI22_X1 U8040 ( .A1(n6757), .A2(n7180), .B1(n6756), .B2(n7178), .ZN(n6758)
         );
  AND2_X2 U8041 ( .A1(n7186), .A2(n6758), .ZN(n9561) );
  OR2_X1 U8042 ( .A1(n9570), .A2(n9559), .ZN(n9529) );
  INV_X1 U8043 ( .A(n6762), .ZN(n6763) );
  NAND2_X1 U8044 ( .A1(n6764), .A2(n6763), .ZN(P2_U3488) );
  NAND2_X1 U8045 ( .A1(n6910), .A2(n8842), .ZN(n6765) );
  NAND2_X1 U8046 ( .A1(n6765), .A2(n6909), .ZN(n6912) );
  NAND2_X1 U8047 ( .A1(n6912), .A2(n6766), .ZN(n6767) );
  NAND2_X1 U8048 ( .A1(n6767), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8049 ( .A(n6768), .ZN(n6801) );
  OR2_X1 U8050 ( .A1(n6910), .A2(n6801), .ZN(n10574) );
  INV_X2 U8051 ( .A(n10574), .ZN(P2_U3893) );
  NOR2_X1 U8052 ( .A1(n7028), .A2(P1_U3086), .ZN(n6769) );
  NAND2_X1 U8053 ( .A1(n7910), .A2(n6769), .ZN(n7071) );
  NOR2_X1 U8054 ( .A1(n8328), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10345) );
  INV_X1 U8055 ( .A(n10345), .ZN(n10350) );
  OAI222_X1 U8056 ( .A1(n6953), .A2(P1_U3086), .B1(n10354), .B2(n6775), .C1(
        n6770), .C2(n10350), .ZN(P1_U3352) );
  INV_X1 U8057 ( .A(n9623), .ZN(n7792) );
  INV_X1 U8058 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6772) );
  OAI222_X1 U8059 ( .A1(n7792), .A2(n6772), .B1(n9625), .B2(n6783), .C1(
        P2_U3151), .C2(n5359), .ZN(P2_U3294) );
  INV_X1 U8060 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6773) );
  OAI222_X1 U8061 ( .A1(n7792), .A2(n6773), .B1(n9625), .B2(n6782), .C1(
        P2_U3151), .C2(n7122), .ZN(P2_U3293) );
  INV_X1 U8062 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6774) );
  INV_X1 U8063 ( .A(n7134), .ZN(n7167) );
  OAI222_X1 U8064 ( .A1(n7792), .A2(n6774), .B1(n9625), .B2(n6780), .C1(
        P2_U3151), .C2(n7167), .ZN(P2_U3291) );
  INV_X1 U8065 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6776) );
  OAI222_X1 U8066 ( .A1(n7792), .A2(n6776), .B1(n9625), .B2(n6775), .C1(
        P2_U3151), .C2(n7126), .ZN(P2_U3292) );
  INV_X1 U8067 ( .A(n6777), .ZN(n6786) );
  OAI222_X1 U8068 ( .A1(n7792), .A2(n6778), .B1(n9625), .B2(n6786), .C1(
        P2_U3151), .C2(n7224), .ZN(P2_U3290) );
  OAI222_X1 U8069 ( .A1(n9852), .A2(P1_U3086), .B1(n10354), .B2(n6780), .C1(
        n6779), .C2(n10350), .ZN(P1_U3351) );
  OAI222_X1 U8070 ( .A1(n6951), .A2(P1_U3086), .B1(n10354), .B2(n6782), .C1(
        n6781), .C2(n10350), .ZN(P1_U3353) );
  OAI222_X1 U8071 ( .A1(n10350), .A2(n6784), .B1(n10354), .B2(n6783), .C1(
        n6949), .C2(P1_U3086), .ZN(P1_U3354) );
  INV_X1 U8072 ( .A(n9872), .ZN(n6787) );
  OAI222_X1 U8073 ( .A1(n6787), .A2(P1_U3086), .B1(n10354), .B2(n6786), .C1(
        n6785), .C2(n10350), .ZN(P1_U3350) );
  INV_X1 U8074 ( .A(n6788), .ZN(n6790) );
  AOI22_X1 U8075 ( .A1(n9887), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n10345), .ZN(n6789) );
  OAI21_X1 U8076 ( .B1(n6790), .B2(n10354), .A(n6789), .ZN(P1_U3349) );
  OAI222_X1 U8077 ( .A1(n7792), .A2(n6791), .B1(n9625), .B2(n6790), .C1(
        P2_U3151), .C2(n7349), .ZN(P2_U3289) );
  INV_X1 U8078 ( .A(n6792), .ZN(n6794) );
  AOI22_X1 U8079 ( .A1(n6978), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10345), .ZN(n6793) );
  OAI21_X1 U8080 ( .B1(n6794), .B2(n10354), .A(n6793), .ZN(P1_U3348) );
  OAI222_X1 U8081 ( .A1(n7792), .A2(n6795), .B1(n9625), .B2(n6794), .C1(
        P2_U3151), .C2(n7528), .ZN(P2_U3288) );
  INV_X1 U8082 ( .A(n6796), .ZN(n6798) );
  AOI22_X1 U8083 ( .A1(n9903), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10345), .ZN(n6797) );
  OAI21_X1 U8084 ( .B1(n6798), .B2(n10354), .A(n6797), .ZN(P1_U3347) );
  OAI222_X1 U8085 ( .A1(n7792), .A2(n6799), .B1(n9625), .B2(n6798), .C1(
        P2_U3151), .C2(n7630), .ZN(P2_U3287) );
  INV_X1 U8086 ( .A(n6682), .ZN(n6800) );
  INV_X1 U8087 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6803) );
  NOR3_X1 U8088 ( .A1(n6704), .A2(n6801), .A3(n8034), .ZN(n6802) );
  AOI21_X1 U8089 ( .B1(n8278), .B2(n6803), .A(n6802), .ZN(P2_U3376) );
  INV_X1 U8090 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6805) );
  NAND2_X1 U8091 ( .A1(n7014), .A2(n7023), .ZN(n6804) );
  OAI21_X1 U8092 ( .B1(n7023), .B2(n6805), .A(n6804), .ZN(P1_U3439) );
  INV_X1 U8093 ( .A(n6806), .ZN(n6812) );
  AOI22_X1 U8094 ( .A1(n7309), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10345), .ZN(n6807) );
  OAI21_X1 U8095 ( .B1(n6812), .B2(n10354), .A(n6807), .ZN(P1_U3345) );
  INV_X1 U8096 ( .A(n6808), .ZN(n6811) );
  OAI222_X1 U8097 ( .A1(n7792), .A2(n6809), .B1(n9625), .B2(n6811), .C1(n7740), 
        .C2(P2_U3151), .ZN(P2_U3286) );
  INV_X1 U8098 ( .A(n7086), .ZN(n6965) );
  OAI222_X1 U8099 ( .A1(P1_U3086), .A2(n6965), .B1(n10354), .B2(n6811), .C1(
        n6810), .C2(n10350), .ZN(P1_U3346) );
  OAI222_X1 U8100 ( .A1(n7792), .A2(n6813), .B1(n9625), .B2(n6812), .C1(n7938), 
        .C2(P2_U3151), .ZN(P2_U3285) );
  INV_X1 U8101 ( .A(n7028), .ZN(n6999) );
  NAND2_X1 U8102 ( .A1(n7910), .A2(n6999), .ZN(n6814) );
  NAND2_X1 U8103 ( .A1(n6814), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6818) );
  INV_X1 U8104 ( .A(n6818), .ZN(n6817) );
  NAND2_X1 U8105 ( .A1(n7016), .A2(n7910), .ZN(n6816) );
  NAND2_X1 U8106 ( .A1(n6816), .A2(n6815), .ZN(n6819) );
  AND2_X1 U8107 ( .A1(n6817), .A2(n6819), .ZN(n9950) );
  INV_X1 U8108 ( .A(n9950), .ZN(n9920) );
  INV_X1 U8109 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6825) );
  OR2_X1 U8110 ( .A1(n6819), .A2(n6818), .ZN(n6963) );
  INV_X1 U8111 ( .A(n6963), .ZN(n6823) );
  INV_X1 U8112 ( .A(n8304), .ZN(n6962) );
  NOR2_X1 U8113 ( .A1(n8995), .A2(n6962), .ZN(n9824) );
  INV_X1 U8114 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10739) );
  OR2_X1 U8115 ( .A1(n8995), .A2(n8304), .ZN(n8323) );
  INV_X1 U8116 ( .A(n8323), .ZN(n6820) );
  AOI22_X1 U8117 ( .A1(n9824), .A2(P1_REG1_REG_0__SCAN_IN), .B1(n6820), .B2(
        P1_REG2_REG_0__SCAN_IN), .ZN(n6821) );
  XNOR2_X1 U8118 ( .A(n6821), .B(P1_IR_REG_0__SCAN_IN), .ZN(n6822) );
  AOI22_X1 U8119 ( .A1(n6823), .A2(n6822), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n6824) );
  OAI21_X1 U8120 ( .B1(n9920), .B2(n6825), .A(n6824), .ZN(P1_U3243) );
  NOR2_X1 U8121 ( .A1(n9950), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8122 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6830) );
  NAND2_X1 U8123 ( .A1(n7023), .A2(n6826), .ZN(n10356) );
  INV_X1 U8124 ( .A(n10356), .ZN(n6828) );
  OAI21_X1 U8125 ( .B1(n6828), .B2(P1_D_REG_1__SCAN_IN), .A(n6827), .ZN(n6829)
         );
  OAI21_X1 U8126 ( .B1(n7023), .B2(n6830), .A(n6829), .ZN(P1_U3440) );
  INV_X1 U8127 ( .A(n6831), .ZN(n6834) );
  AOI22_X1 U8128 ( .A1(n7430), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10345), .ZN(n6832) );
  OAI21_X1 U8129 ( .B1(n6834), .B2(n10354), .A(n6832), .ZN(P1_U3344) );
  AOI22_X1 U8130 ( .A1(n10675), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n9623), .ZN(n6833) );
  OAI21_X1 U8131 ( .B1(n6834), .B2(n9625), .A(n6833), .ZN(P2_U3284) );
  NAND2_X1 U8132 ( .A1(P1_U3973), .A2(n5056), .ZN(n6835) );
  OAI21_X1 U8133 ( .B1(P1_U3973), .B2(n6270), .A(n6835), .ZN(P1_U3554) );
  INV_X1 U8134 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7791) );
  NAND2_X1 U8135 ( .A1(n10249), .A2(P1_U3973), .ZN(n6836) );
  OAI21_X1 U8136 ( .B1(n7791), .B2(P1_U3973), .A(n6836), .ZN(P1_U3575) );
  NAND2_X1 U8137 ( .A1(n10236), .A2(P1_U3973), .ZN(n6837) );
  OAI21_X1 U8138 ( .B1(P1_U3973), .B2(n6015), .A(n6837), .ZN(P1_U3577) );
  NAND2_X1 U8139 ( .A1(n8140), .A2(n8141), .ZN(n9525) );
  OR2_X1 U8140 ( .A1(n6838), .A2(n8302), .ZN(n8718) );
  NAND2_X1 U8141 ( .A1(n8718), .A2(n8713), .ZN(n7187) );
  OAI21_X1 U8142 ( .B1(n9547), .B2(n9525), .A(n7187), .ZN(n6841) );
  NOR2_X1 U8143 ( .A1(n6839), .A2(n9473), .ZN(n7190) );
  INV_X1 U8144 ( .A(n7190), .ZN(n6840) );
  OAI211_X1 U8145 ( .C1(n9559), .C2(n7194), .A(n6841), .B(n6840), .ZN(n6843)
         );
  NAND2_X1 U8146 ( .A1(n6843), .A2(n9561), .ZN(n6842) );
  OAI21_X1 U8147 ( .B1(n9561), .B2(n6264), .A(n6842), .ZN(P2_U3459) );
  INV_X1 U8148 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6845) );
  NAND2_X1 U8149 ( .A1(n6843), .A2(n10852), .ZN(n6844) );
  OAI21_X1 U8150 ( .B1(n10852), .B2(n6845), .A(n6844), .ZN(P2_U3390) );
  NAND2_X1 U8151 ( .A1(n6872), .A2(n6846), .ZN(n6850) );
  AND2_X1 U8152 ( .A1(n6847), .A2(n6909), .ZN(n6849) );
  NAND2_X1 U8153 ( .A1(n6855), .A2(n6848), .ZN(n6874) );
  NAND4_X1 U8154 ( .A1(n6850), .A2(n6849), .A3(n6910), .A4(n6874), .ZN(n6851)
         );
  NAND2_X1 U8155 ( .A1(n6851), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6853) );
  NOR2_X1 U8156 ( .A1(n9611), .A2(n7188), .ZN(n6854) );
  NAND2_X1 U8157 ( .A1(n6855), .A2(n6854), .ZN(n6852) );
  NAND2_X1 U8158 ( .A1(n6853), .A2(n6852), .ZN(n9125) );
  NOR2_X1 U8159 ( .A1(n9125), .A2(P2_U3151), .ZN(n6902) );
  INV_X1 U8160 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10674) );
  INV_X1 U8161 ( .A(n6854), .ZN(n8866) );
  NOR2_X1 U8162 ( .A1(n6855), .A2(n8866), .ZN(n6860) );
  INV_X1 U8163 ( .A(n6872), .ZN(n6856) );
  NAND2_X1 U8164 ( .A1(n6856), .A2(n6857), .ZN(n6858) );
  NAND2_X1 U8165 ( .A1(n6858), .A2(n10838), .ZN(n9131) );
  INV_X1 U8166 ( .A(n6860), .ZN(n6862) );
  OAI22_X1 U8167 ( .A1(n9114), .A2(n6859), .B1(n8302), .B2(n9094), .ZN(n6863)
         );
  AOI21_X1 U8168 ( .B1(n9081), .B2(n9150), .A(n6863), .ZN(n6879) );
  AND2_X1 U8169 ( .A1(n8712), .A2(n7371), .ZN(n6864) );
  NAND2_X1 U8170 ( .A1(n8693), .A2(n7696), .ZN(n6866) );
  NAND2_X2 U8171 ( .A1(n6867), .A2(n6866), .ZN(n8600) );
  XNOR2_X1 U8172 ( .A(n6880), .B(n9151), .ZN(n6868) );
  OAI21_X1 U8173 ( .B1(n6869), .B2(n6868), .A(n4959), .ZN(n6877) );
  OAI21_X1 U8174 ( .B1(n6872), .B2(n6871), .A(n6870), .ZN(n6876) );
  AND2_X1 U8175 ( .A1(n6874), .A2(n6873), .ZN(n6875) );
  NAND2_X1 U8176 ( .A1(n6876), .A2(n6875), .ZN(n9133) );
  INV_X1 U8177 ( .A(n9133), .ZN(n9091) );
  NAND2_X1 U8178 ( .A1(n6877), .A2(n9091), .ZN(n6878) );
  OAI211_X1 U8179 ( .C1(n6902), .C2(n10674), .A(n6879), .B(n6878), .ZN(
        P2_U3162) );
  INV_X1 U8180 ( .A(n4959), .ZN(n6882) );
  NAND2_X1 U8181 ( .A1(n6880), .A2(n6839), .ZN(n6883) );
  INV_X1 U8182 ( .A(n6883), .ZN(n6881) );
  XNOR2_X1 U8183 ( .A(n7198), .B(n9150), .ZN(n6885) );
  NOR3_X1 U8184 ( .A1(n6882), .A2(n6881), .A3(n6885), .ZN(n6888) );
  NAND2_X1 U8185 ( .A1(n6884), .A2(n6883), .ZN(n6886) );
  NAND2_X1 U8186 ( .A1(n6886), .A2(n6885), .ZN(n7200) );
  INV_X1 U8187 ( .A(n7200), .ZN(n6887) );
  OAI21_X1 U8188 ( .B1(n6888), .B2(n6887), .A(n9091), .ZN(n6892) );
  OAI22_X1 U8189 ( .A1(n9114), .A2(n6889), .B1(n6839), .B2(n9094), .ZN(n6890)
         );
  AOI21_X1 U8190 ( .B1(n9081), .B2(n9149), .A(n6890), .ZN(n6891) );
  OAI211_X1 U8191 ( .C1(n6275), .C2(n6902), .A(n6892), .B(n6891), .ZN(P2_U3177) );
  INV_X1 U8192 ( .A(n6893), .ZN(n6896) );
  OAI222_X1 U8193 ( .A1(n7792), .A2(n6894), .B1(n9625), .B2(n6896), .C1(n8154), 
        .C2(P2_U3151), .ZN(P2_U3283) );
  INV_X1 U8194 ( .A(n7621), .ZN(n7428) );
  INV_X1 U8195 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6895) );
  OAI222_X1 U8196 ( .A1(P1_U3086), .A2(n7428), .B1(n10354), .B2(n6896), .C1(
        n6895), .C2(n10350), .ZN(P1_U3343) );
  INV_X1 U8197 ( .A(n9407), .ZN(n9037) );
  NAND2_X1 U8198 ( .A1(n9037), .A2(P2_U3893), .ZN(n6897) );
  OAI21_X1 U8199 ( .B1(P2_U3893), .B2(n7652), .A(n6897), .ZN(P2_U3511) );
  INV_X1 U8200 ( .A(n6898), .ZN(n6984) );
  AOI22_X1 U8201 ( .A1(n7823), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10345), .ZN(n6899) );
  OAI21_X1 U8202 ( .B1(n6984), .B2(n10354), .A(n6899), .ZN(P1_U3342) );
  INV_X1 U8203 ( .A(n9081), .ZN(n9129) );
  OAI22_X1 U8204 ( .A1(n9114), .A2(n7194), .B1(n9129), .B2(n6839), .ZN(n6900)
         );
  AOI21_X1 U8205 ( .B1(n9091), .B2(n7187), .A(n6900), .ZN(n6901) );
  OAI21_X1 U8206 ( .B1(n6902), .B2(n7193), .A(n6901), .ZN(P2_U3172) );
  NOR2_X1 U8207 ( .A1(n4947), .A2(P2_U3151), .ZN(n8265) );
  AND2_X1 U8208 ( .A1(n6912), .A2(n8265), .ZN(n6903) );
  MUX2_X1 U8209 ( .A(n6903), .B(P2_U3893), .S(n5093), .Z(n10676) );
  INV_X1 U8210 ( .A(n10676), .ZN(n10706) );
  MUX2_X1 U8211 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n4946), .Z(n6905) );
  MUX2_X1 U8212 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n9256), .Z(n6904) );
  XNOR2_X1 U8213 ( .A(n10655), .B(n6904), .ZN(n10659) );
  MUX2_X1 U8214 ( .A(n6263), .B(n6264), .S(n4947), .Z(n7036) );
  NAND2_X1 U8215 ( .A1(n7036), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10658) );
  AND2_X1 U8216 ( .A1(n10659), .A2(n10658), .ZN(n10656) );
  AOI21_X1 U8217 ( .B1(n6904), .B2(n5359), .A(n10656), .ZN(n7106) );
  XOR2_X1 U8218 ( .A(n6922), .B(n6905), .Z(n7107) );
  NOR2_X1 U8219 ( .A1(n7106), .A2(n7107), .ZN(n7105) );
  AOI21_X1 U8220 ( .B1(n6905), .B2(n7122), .A(n7105), .ZN(n6907) );
  MUX2_X1 U8221 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n4946), .Z(n7127) );
  XNOR2_X1 U8222 ( .A(n7127), .B(n6919), .ZN(n6906) );
  NAND2_X1 U8223 ( .A1(n6907), .A2(n6906), .ZN(n7125) );
  OAI21_X1 U8224 ( .B1(n6907), .B2(n6906), .A(n7125), .ZN(n6908) );
  AND2_X1 U8225 ( .A1(P2_U3893), .A2(n8864), .ZN(n10690) );
  NAND2_X1 U8226 ( .A1(n6908), .A2(n10690), .ZN(n6936) );
  INV_X1 U8227 ( .A(n6909), .ZN(n7890) );
  NOR2_X1 U8228 ( .A1(n6910), .A2(n7890), .ZN(n6911) );
  OR2_X1 U8229 ( .A1(P2_U3150), .A2(n6911), .ZN(n9263) );
  INV_X1 U8230 ( .A(n9263), .ZN(n10698) );
  NOR2_X1 U8231 ( .A1(n8864), .A2(P2_U3151), .ZN(n9622) );
  NAND2_X1 U8232 ( .A1(n6912), .A2(n9622), .ZN(n7035) );
  INV_X1 U8233 ( .A(n4946), .ZN(n8865) );
  OR2_X1 U8234 ( .A1(n7035), .A2(n8865), .ZN(n10713) );
  NAND2_X1 U8235 ( .A1(n6924), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6913) );
  NAND2_X1 U8236 ( .A1(n10655), .A2(n6913), .ZN(n6914) );
  NAND2_X1 U8237 ( .A1(n6293), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6915) );
  NAND2_X1 U8238 ( .A1(n6914), .A2(n6915), .ZN(n10660) );
  NOR2_X1 U8239 ( .A1(n10660), .A2(n6250), .ZN(n10663) );
  INV_X1 U8240 ( .A(n6915), .ZN(n6916) );
  NOR2_X1 U8241 ( .A1(n10663), .A2(n6916), .ZN(n7114) );
  OAI21_X1 U8242 ( .B1(n6922), .B2(n6917), .A(n6918), .ZN(n7113) );
  NOR2_X1 U8243 ( .A1(n7114), .A2(n7113), .ZN(n7112) );
  AOI21_X1 U8244 ( .B1(n6287), .B2(n6920), .A(n7156), .ZN(n6921) );
  NOR2_X1 U8245 ( .A1(n10713), .A2(n6921), .ZN(n6934) );
  OR2_X1 U8246 ( .A1(n7035), .A2(n4947), .ZN(n10682) );
  INV_X1 U8247 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6923) );
  MUX2_X1 U8248 ( .A(n6923), .B(P2_REG2_REG_2__SCAN_IN), .S(n6922), .Z(n7111)
         );
  NAND2_X1 U8249 ( .A1(n6924), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6925) );
  NAND2_X1 U8250 ( .A1(n10655), .A2(n6925), .ZN(n6926) );
  NAND2_X1 U8251 ( .A1(n6293), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6927) );
  NAND2_X1 U8252 ( .A1(n6926), .A2(n6927), .ZN(n10670) );
  OR2_X1 U8253 ( .A1(n10670), .A2(n6246), .ZN(n10668) );
  NAND2_X1 U8254 ( .A1(n10668), .A2(n6927), .ZN(n7110) );
  NAND2_X1 U8255 ( .A1(n7122), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6928) );
  INV_X1 U8256 ( .A(n7153), .ZN(n6929) );
  AOI21_X1 U8257 ( .B1(n6286), .B2(n6930), .A(n6929), .ZN(n6932) );
  NOR2_X1 U8258 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10466), .ZN(n9016) );
  INV_X1 U8259 ( .A(n9016), .ZN(n6931) );
  OAI21_X1 U8260 ( .B1(n10682), .B2(n6932), .A(n6931), .ZN(n6933) );
  AOI211_X1 U8261 ( .C1(n10698), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6934), .B(
        n6933), .ZN(n6935) );
  OAI211_X1 U8262 ( .C1(n10706), .C2(n7126), .A(n6936), .B(n6935), .ZN(
        P2_U3185) );
  XNOR2_X1 U8263 ( .A(n7086), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n6948) );
  XNOR2_X1 U8264 ( .A(n6951), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n9831) );
  XNOR2_X1 U8265 ( .A(n6949), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9813) );
  AND2_X1 U8266 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9812) );
  NAND2_X1 U8267 ( .A1(n9813), .A2(n9812), .ZN(n9811) );
  INV_X1 U8268 ( .A(n6949), .ZN(n9814) );
  NAND2_X1 U8269 ( .A1(n9814), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6937) );
  NAND2_X1 U8270 ( .A1(n9811), .A2(n6937), .ZN(n9830) );
  NAND2_X1 U8271 ( .A1(n9831), .A2(n9830), .ZN(n9829) );
  INV_X1 U8272 ( .A(n6951), .ZN(n9828) );
  NAND2_X1 U8273 ( .A1(n9828), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6938) );
  NAND2_X1 U8274 ( .A1(n9829), .A2(n6938), .ZN(n9844) );
  XNOR2_X1 U8275 ( .A(n6953), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9845) );
  NAND2_X1 U8276 ( .A1(n9844), .A2(n9845), .ZN(n9843) );
  INV_X1 U8277 ( .A(n6953), .ZN(n9842) );
  NAND2_X1 U8278 ( .A1(n9842), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6939) );
  NAND2_X1 U8279 ( .A1(n9843), .A2(n6939), .ZN(n9859) );
  MUX2_X1 U8280 ( .A(n5777), .B(P1_REG2_REG_4__SCAN_IN), .S(n9852), .Z(n9860)
         );
  NAND2_X1 U8281 ( .A1(n9859), .A2(n9860), .ZN(n9858) );
  INV_X1 U8282 ( .A(n9852), .ZN(n6956) );
  NAND2_X1 U8283 ( .A1(n6956), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6940) );
  NAND2_X1 U8284 ( .A1(n9858), .A2(n6940), .ZN(n9874) );
  INV_X1 U8285 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6941) );
  XNOR2_X1 U8286 ( .A(n9872), .B(n6941), .ZN(n9875) );
  NAND2_X1 U8287 ( .A1(n9874), .A2(n9875), .ZN(n9873) );
  NAND2_X1 U8288 ( .A1(n9872), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6942) );
  NAND2_X1 U8289 ( .A1(n9873), .A2(n6942), .ZN(n9889) );
  MUX2_X1 U8290 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7856), .S(n9887), .Z(n9890)
         );
  NAND2_X1 U8291 ( .A1(n9889), .A2(n9890), .ZN(n9888) );
  NAND2_X1 U8292 ( .A1(n9887), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6943) );
  NAND2_X1 U8293 ( .A1(n9888), .A2(n6943), .ZN(n6973) );
  XNOR2_X1 U8294 ( .A(n6978), .B(n7579), .ZN(n6974) );
  AND2_X1 U8295 ( .A1(n6973), .A2(n6974), .ZN(n6975) );
  AND2_X1 U8296 ( .A1(n6978), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6944) );
  XNOR2_X1 U8297 ( .A(n9903), .B(n7861), .ZN(n9907) );
  NAND2_X1 U8298 ( .A1(n9906), .A2(n9907), .ZN(n9904) );
  NAND2_X1 U8299 ( .A1(n9903), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6945) );
  NAND2_X1 U8300 ( .A1(n9904), .A2(n6945), .ZN(n6947) );
  INV_X1 U8301 ( .A(n7081), .ZN(n6946) );
  AOI21_X1 U8302 ( .B1(n6948), .B2(n6947), .A(n6946), .ZN(n6969) );
  OR2_X1 U8303 ( .A1(n6963), .A2(n8323), .ZN(n9953) );
  XNOR2_X1 U8304 ( .A(n6949), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9810) );
  NAND3_X1 U8305 ( .A1(n9810), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9808) );
  OAI21_X1 U8306 ( .B1(n6950), .B2(n6949), .A(n9808), .ZN(n9833) );
  XNOR2_X1 U8307 ( .A(n6951), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9834) );
  NAND2_X1 U8308 ( .A1(n9833), .A2(n9834), .ZN(n9832) );
  OAI21_X1 U8309 ( .B1(n6952), .B2(n6951), .A(n9832), .ZN(n9847) );
  XNOR2_X1 U8310 ( .A(n6953), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9848) );
  NAND2_X1 U8311 ( .A1(n9847), .A2(n9848), .ZN(n9846) );
  OAI21_X1 U8312 ( .B1(n6954), .B2(n6953), .A(n9846), .ZN(n9856) );
  MUX2_X1 U8313 ( .A(n5778), .B(P1_REG1_REG_4__SCAN_IN), .S(n9852), .Z(n9857)
         );
  NAND2_X1 U8314 ( .A1(n9856), .A2(n9857), .ZN(n9855) );
  INV_X1 U8315 ( .A(n9855), .ZN(n6955) );
  AOI21_X1 U8316 ( .B1(n6956), .B2(P1_REG1_REG_4__SCAN_IN), .A(n6955), .ZN(
        n9867) );
  XNOR2_X1 U8317 ( .A(n9872), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9866) );
  NOR2_X1 U8318 ( .A1(n9867), .A2(n9866), .ZN(n9865) );
  AOI21_X1 U8319 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n9872), .A(n9865), .ZN(
        n9881) );
  MUX2_X1 U8320 ( .A(n6957), .B(P1_REG1_REG_6__SCAN_IN), .S(n9887), .Z(n9880)
         );
  NOR2_X1 U8321 ( .A1(n9881), .A2(n9880), .ZN(n9879) );
  AOI21_X1 U8322 ( .B1(n9887), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9879), .ZN(
        n6972) );
  XNOR2_X1 U8323 ( .A(n6978), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n6971) );
  NOR2_X1 U8324 ( .A1(n6972), .A2(n6971), .ZN(n6970) );
  AOI21_X1 U8325 ( .B1(n6978), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6970), .ZN(
        n9897) );
  MUX2_X1 U8326 ( .A(n6958), .B(P1_REG1_REG_8__SCAN_IN), .S(n9903), .Z(n9896)
         );
  NOR2_X1 U8327 ( .A1(n9897), .A2(n9896), .ZN(n9894) );
  AOI21_X1 U8328 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9903), .A(n9894), .ZN(
        n6961) );
  MUX2_X1 U8329 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n6959), .S(n7086), .Z(n6960)
         );
  NAND2_X1 U8330 ( .A1(n6961), .A2(n6960), .ZN(n7085) );
  OAI21_X1 U8331 ( .B1(n6961), .B2(n6960), .A(n7085), .ZN(n6967) );
  NOR2_X1 U8332 ( .A1(n6963), .A2(n6962), .ZN(n9944) );
  OR2_X1 U8333 ( .A1(n6963), .A2(n9819), .ZN(n9947) );
  AND2_X1 U8334 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7786) );
  AOI21_X1 U8335 ( .B1(n9950), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7786), .ZN(
        n6964) );
  OAI21_X1 U8336 ( .B1(n9947), .B2(n6965), .A(n6964), .ZN(n6966) );
  AOI21_X1 U8337 ( .B1(n6967), .B2(n9944), .A(n6966), .ZN(n6968) );
  OAI21_X1 U8338 ( .B1(n6969), .B2(n9953), .A(n6968), .ZN(P1_U3252) );
  INV_X1 U8339 ( .A(n9944), .ZN(n9895) );
  AOI211_X1 U8340 ( .C1(n6972), .C2(n6971), .A(n9895), .B(n6970), .ZN(n6983)
         );
  INV_X1 U8341 ( .A(n6973), .ZN(n6977) );
  INV_X1 U8342 ( .A(n6974), .ZN(n6976) );
  AOI211_X1 U8343 ( .C1(n6977), .C2(n6976), .A(n6975), .B(n9953), .ZN(n6982)
         );
  INV_X1 U8344 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6980) );
  INV_X1 U8345 ( .A(n9947), .ZN(n9930) );
  NAND2_X1 U8346 ( .A1(n9930), .A2(n6978), .ZN(n6979) );
  NAND2_X1 U8347 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8309) );
  OAI211_X1 U8348 ( .C1(n6980), .C2(n9920), .A(n6979), .B(n8309), .ZN(n6981)
         );
  OR3_X1 U8349 ( .A1(n6983), .A2(n6982), .A3(n6981), .ZN(P1_U3250) );
  OAI222_X1 U8350 ( .A1(n6985), .A2(n7792), .B1(P2_U3151), .B2(n9158), .C1(
        n9625), .C2(n6984), .ZN(P2_U3282) );
  INV_X1 U8351 ( .A(n6986), .ZN(n6988) );
  AOI22_X1 U8352 ( .A1(n8074), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10345), .ZN(n6987) );
  OAI21_X1 U8353 ( .B1(n6988), .B2(n10354), .A(n6987), .ZN(P1_U3341) );
  INV_X1 U8354 ( .A(n9170), .ZN(n9191) );
  OAI222_X1 U8355 ( .A1(n7792), .A2(n6989), .B1(n9625), .B2(n6988), .C1(
        P2_U3151), .C2(n9191), .ZN(P2_U3281) );
  NAND2_X1 U8356 ( .A1(n7574), .A2(n8577), .ZN(n6990) );
  NAND2_X1 U8357 ( .A1(n6995), .A2(n6990), .ZN(n6991) );
  NAND2_X1 U8358 ( .A1(n7254), .A2(n9807), .ZN(n6994) );
  AND2_X4 U8359 ( .A1(n6992), .A2(n7028), .ZN(n8916) );
  NAND2_X1 U8360 ( .A1(n8916), .A2(n10193), .ZN(n6993) );
  NAND2_X1 U8361 ( .A1(n6994), .A2(n6993), .ZN(n7255) );
  NAND2_X1 U8362 ( .A1(n7269), .A2(n10722), .ZN(n6997) );
  NAND2_X1 U8363 ( .A1(n10194), .A2(n8916), .ZN(n6996) );
  NAND2_X1 U8364 ( .A1(n6999), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n7000) );
  OAI211_X1 U8365 ( .C1(n8903), .C2(n8449), .A(n7001), .B(n7000), .ZN(n8318)
         );
  NAND2_X1 U8366 ( .A1(n8319), .A2(n8318), .ZN(n8317) );
  OR2_X1 U8367 ( .A1(n7002), .A2(n8963), .ZN(n7003) );
  NAND2_X1 U8368 ( .A1(n7269), .A2(n10193), .ZN(n7005) );
  NAND2_X1 U8369 ( .A1(n9807), .A2(n8916), .ZN(n7004) );
  NAND2_X1 U8370 ( .A1(n7005), .A2(n7004), .ZN(n7007) );
  INV_X2 U8371 ( .A(n8975), .ZN(n8883) );
  XNOR2_X1 U8372 ( .A(n7007), .B(n8883), .ZN(n7009) );
  INV_X1 U8373 ( .A(n7009), .ZN(n7010) );
  NAND2_X1 U8374 ( .A1(n7011), .A2(n7010), .ZN(n7257) );
  NAND2_X1 U8375 ( .A1(n7256), .A2(n7257), .ZN(n7012) );
  XOR2_X1 U8376 ( .A(n7255), .B(n7012), .Z(n7034) );
  NAND3_X1 U8377 ( .A1(n7014), .A2(n7571), .A3(n7013), .ZN(n7027) );
  INV_X1 U8378 ( .A(n7027), .ZN(n7015) );
  NAND2_X1 U8379 ( .A1(n7015), .A2(n7023), .ZN(n7025) );
  INV_X1 U8380 ( .A(n7025), .ZN(n7018) );
  INV_X1 U8381 ( .A(n10283), .ZN(n10824) );
  INV_X1 U8382 ( .A(n7016), .ZN(n8511) );
  AND2_X1 U8383 ( .A1(n10824), .A2(n8511), .ZN(n7017) );
  NAND2_X1 U8384 ( .A1(n7018), .A2(n7017), .ZN(n9788) );
  OR2_X1 U8385 ( .A1(n7020), .A2(n7019), .ZN(n8324) );
  NOR2_X1 U8386 ( .A1(n7027), .A2(n8324), .ZN(n7021) );
  NAND2_X1 U8387 ( .A1(n7021), .A2(n8995), .ZN(n9779) );
  NAND2_X1 U8388 ( .A1(n7021), .A2(n9819), .ZN(n9783) );
  INV_X1 U8389 ( .A(n9783), .ZN(n9767) );
  AOI22_X1 U8390 ( .A1(n9768), .A2(n9806), .B1(n9767), .B2(n5056), .ZN(n7033)
         );
  OR2_X1 U8391 ( .A1(n7022), .A2(n8576), .ZN(n7577) );
  NAND2_X1 U8392 ( .A1(n8515), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7650) );
  NAND2_X1 U8393 ( .A1(n10283), .A2(n7650), .ZN(n7026) );
  NAND2_X1 U8394 ( .A1(n7027), .A2(n7026), .ZN(n7031) );
  AND3_X1 U8395 ( .A1(n7029), .A2(n7910), .A3(n7028), .ZN(n7030) );
  NAND2_X1 U8396 ( .A1(n7031), .A2(n7030), .ZN(n7273) );
  OR2_X1 U8397 ( .A1(n7273), .A2(P1_U3086), .ZN(n8320) );
  AOI22_X1 U8398 ( .A1(n4944), .A2(n10193), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n8320), .ZN(n7032) );
  OAI211_X1 U8399 ( .C1(n7034), .C2(n9788), .A(n7033), .B(n7032), .ZN(P1_U3222) );
  INV_X1 U8400 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n7041) );
  INV_X1 U8401 ( .A(n10690), .ZN(n10695) );
  NAND2_X1 U8402 ( .A1(n10695), .A2(n7035), .ZN(n7038) );
  OAI21_X1 U8403 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n7036), .A(n10658), .ZN(
        n7037) );
  AOI22_X1 U8404 ( .A1(n7038), .A2(n7037), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n7040) );
  NAND2_X1 U8405 ( .A1(n10676), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7039) );
  OAI211_X1 U8406 ( .C1(n9263), .C2(n7041), .A(n7040), .B(n7039), .ZN(P2_U3182) );
  OAI21_X1 U8407 ( .B1(n7043), .B2(n8453), .A(n7042), .ZN(n7767) );
  INV_X1 U8408 ( .A(n10782), .ZN(n10174) );
  AOI211_X1 U8409 ( .C1(n7276), .C2(n7704), .A(n10174), .B(n7044), .ZN(n7762)
         );
  XNOR2_X1 U8410 ( .A(n8453), .B(n7045), .ZN(n7046) );
  INV_X1 U8411 ( .A(n10162), .ZN(n10791) );
  OAI222_X1 U8412 ( .A1(n10796), .A2(n10186), .B1(n10794), .B2(n7415), .C1(
        n7046), .C2(n10791), .ZN(n7761) );
  AOI211_X1 U8413 ( .C1(n5053), .C2(n7767), .A(n7762), .B(n7761), .ZN(n7241)
         );
  OAI22_X1 U8414 ( .A1(n10340), .A2(n7765), .B1(n10834), .B2(n5772), .ZN(n7047) );
  INV_X1 U8415 ( .A(n7047), .ZN(n7048) );
  OAI21_X1 U8416 ( .B1(n7241), .B2(n6207), .A(n7048), .ZN(P1_U3462) );
  XNOR2_X1 U8417 ( .A(n7049), .B(n8454), .ZN(n7662) );
  OAI21_X1 U8418 ( .B1(n7051), .B2(n8454), .A(n7050), .ZN(n7660) );
  NAND2_X1 U8419 ( .A1(n7052), .A2(n10782), .ZN(n7053) );
  NOR2_X1 U8420 ( .A1(n7687), .A2(n7053), .ZN(n7653) );
  OAI22_X1 U8421 ( .A1(n7657), .A2(n10796), .B1(n9726), .B2(n10794), .ZN(n7054) );
  AOI211_X1 U8422 ( .C1(n7660), .C2(n10828), .A(n7653), .B(n7054), .ZN(n7055)
         );
  OAI21_X1 U8423 ( .B1(n10791), .B2(n7662), .A(n7055), .ZN(n7246) );
  INV_X1 U8424 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7056) );
  OAI22_X1 U8425 ( .A1(n10340), .A2(n5290), .B1(n10834), .B2(n7056), .ZN(n7057) );
  AOI21_X1 U8426 ( .B1(n7246), .B2(n10834), .A(n7057), .ZN(n7058) );
  INV_X1 U8427 ( .A(n7058), .ZN(P1_U3465) );
  OAI21_X1 U8428 ( .B1(n7064), .B2(n7060), .A(n7059), .ZN(n10188) );
  AOI22_X1 U8429 ( .A1(n10268), .A2(n9806), .B1(n10267), .B2(n5056), .ZN(n7063) );
  NAND2_X1 U8430 ( .A1(n10193), .A2(n10722), .ZN(n7061) );
  NAND2_X1 U8431 ( .A1(n10782), .A2(n7061), .ZN(n7062) );
  OR2_X1 U8432 ( .A1(n7062), .A2(n7705), .ZN(n10183) );
  NAND2_X1 U8433 ( .A1(n7063), .A2(n10183), .ZN(n7067) );
  INV_X1 U8434 ( .A(n8450), .ZN(n7065) );
  XNOR2_X1 U8435 ( .A(n7065), .B(n7064), .ZN(n7066) );
  AND2_X1 U8436 ( .A1(n7066), .A2(n10162), .ZN(n10196) );
  AOI211_X1 U8437 ( .C1(n5053), .C2(n10188), .A(n7067), .B(n10196), .ZN(n7250)
         );
  OAI22_X1 U8438 ( .A1(n10340), .A2(n8520), .B1(n10834), .B2(n5722), .ZN(n7068) );
  INV_X1 U8439 ( .A(n7068), .ZN(n7069) );
  OAI21_X1 U8440 ( .B1(n7250), .B2(n6207), .A(n7069), .ZN(P1_U3456) );
  NAND2_X1 U8441 ( .A1(n7071), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7070) );
  OAI21_X1 U8442 ( .B1(n7071), .B2(n9979), .A(n7070), .ZN(P1_U3583) );
  INV_X1 U8443 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7073) );
  INV_X1 U8444 ( .A(n7072), .ZN(n7074) );
  INV_X1 U8445 ( .A(n9213), .ZN(n9206) );
  OAI222_X1 U8446 ( .A1(n7792), .A2(n7073), .B1(n9625), .B2(n7074), .C1(n9206), 
        .C2(P2_U3151), .ZN(P2_U3280) );
  INV_X1 U8447 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10575) );
  OAI222_X1 U8448 ( .A1(P1_U3086), .A2(n8173), .B1(n10354), .B2(n7074), .C1(
        n10575), .C2(n10350), .ZN(P1_U3340) );
  OAI21_X1 U8449 ( .B1(n6274), .B2(n6273), .A(n7075), .ZN(n7362) );
  NOR2_X1 U8450 ( .A1(n6859), .A2(n9559), .ZN(n7078) );
  INV_X1 U8451 ( .A(n9547), .ZN(n9468) );
  AOI21_X1 U8452 ( .B1(n7076), .B2(n6274), .A(n7100), .ZN(n7077) );
  OAI222_X1 U8453 ( .A1(n9473), .A2(n7284), .B1(n9471), .B2(n8302), .C1(n9468), 
        .C2(n7077), .ZN(n7357) );
  AOI211_X1 U8454 ( .C1(n9525), .C2(n7362), .A(n7078), .B(n7357), .ZN(n10741)
         );
  OR2_X1 U8455 ( .A1(n10741), .A2(n9570), .ZN(n7079) );
  OAI21_X1 U8456 ( .B1(n9561), .B2(n6250), .A(n7079), .ZN(P2_U3460) );
  OR2_X1 U8457 ( .A1(n7086), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7080) );
  MUX2_X1 U8458 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n7590), .S(n7309), .Z(n7082)
         );
  INV_X1 U8459 ( .A(n9953), .ZN(n9905) );
  OAI21_X1 U8460 ( .B1(n7083), .B2(n7082), .A(n9905), .ZN(n7094) );
  MUX2_X1 U8461 ( .A(n7084), .B(P1_REG1_REG_10__SCAN_IN), .S(n7309), .Z(n7088)
         );
  OAI21_X1 U8462 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n7086), .A(n7085), .ZN(
        n7087) );
  NOR2_X1 U8463 ( .A1(n7087), .A2(n7088), .ZN(n7304) );
  AOI211_X1 U8464 ( .C1(n7088), .C2(n7087), .A(n9895), .B(n7304), .ZN(n7089)
         );
  INV_X1 U8465 ( .A(n7089), .ZN(n7093) );
  INV_X1 U8466 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7090) );
  NAND2_X1 U8467 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n7964) );
  OAI21_X1 U8468 ( .B1(n9920), .B2(n7090), .A(n7964), .ZN(n7091) );
  AOI21_X1 U8469 ( .B1(n7309), .B2(n9930), .A(n7091), .ZN(n7092) );
  OAI211_X1 U8470 ( .C1(n7308), .C2(n7094), .A(n7093), .B(n7092), .ZN(P1_U3253) );
  XNOR2_X1 U8471 ( .A(n8722), .B(n7095), .ZN(n7373) );
  INV_X1 U8472 ( .A(n9559), .ZN(n9568) );
  AND2_X1 U8473 ( .A1(n7096), .A2(n9568), .ZN(n7372) );
  INV_X1 U8474 ( .A(n7097), .ZN(n7102) );
  NOR3_X1 U8475 ( .A1(n7100), .A2(n7099), .A3(n7098), .ZN(n7101) );
  NOR2_X1 U8476 ( .A1(n7102), .A2(n7101), .ZN(n7103) );
  OAI222_X1 U8477 ( .A1(n9473), .A2(n7384), .B1(n9471), .B2(n6839), .C1(n9468), 
        .C2(n7103), .ZN(n7369) );
  AOI211_X1 U8478 ( .C1(n7373), .C2(n9525), .A(n7372), .B(n7369), .ZN(n10748)
         );
  NAND2_X1 U8479 ( .A1(n9570), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7104) );
  OAI21_X1 U8480 ( .B1(n10748), .B2(n9570), .A(n7104), .ZN(P2_U3461) );
  AOI211_X1 U8481 ( .C1(n7107), .C2(n7106), .A(n10695), .B(n7105), .ZN(n7108)
         );
  INV_X1 U8482 ( .A(n7108), .ZN(n7121) );
  INV_X1 U8483 ( .A(n10682), .ZN(n10710) );
  OAI21_X1 U8484 ( .B1(n7111), .B2(n7110), .A(n7109), .ZN(n7119) );
  NOR2_X1 U8485 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6275), .ZN(n7118) );
  INV_X1 U8486 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7116) );
  AOI21_X1 U8487 ( .B1(n7114), .B2(n7113), .A(n7112), .ZN(n7115) );
  OAI22_X1 U8488 ( .A1(n9263), .A2(n7116), .B1(n10713), .B2(n7115), .ZN(n7117)
         );
  AOI211_X1 U8489 ( .C1(n10710), .C2(n7119), .A(n7118), .B(n7117), .ZN(n7120)
         );
  OAI211_X1 U8490 ( .C1(n10706), .C2(n7122), .A(n7121), .B(n7120), .ZN(
        P2_U3184) );
  MUX2_X1 U8491 ( .A(n7123), .B(P2_REG1_REG_4__SCAN_IN), .S(n7134), .Z(n7157)
         );
  OAI21_X1 U8492 ( .B1(n7134), .B2(n7123), .A(n7160), .ZN(n7219) );
  XNOR2_X1 U8493 ( .A(n7219), .B(n7224), .ZN(n7124) );
  AOI21_X1 U8494 ( .B1(n6314), .B2(n7124), .A(n7220), .ZN(n7145) );
  MUX2_X1 U8495 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n4947), .Z(n7216) );
  XNOR2_X1 U8496 ( .A(n7216), .B(n7224), .ZN(n7130) );
  MUX2_X1 U8497 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n4946), .Z(n7128) );
  OAI21_X1 U8498 ( .B1(n7127), .B2(n7126), .A(n7125), .ZN(n7147) );
  XOR2_X1 U8499 ( .A(n7134), .B(n7128), .Z(n7148) );
  NOR2_X1 U8500 ( .A1(n7147), .A2(n7148), .ZN(n7146) );
  AOI21_X1 U8501 ( .B1(n7128), .B2(n7167), .A(n7146), .ZN(n7129) );
  NOR2_X1 U8502 ( .A1(n7129), .A2(n7130), .ZN(n7215) );
  AOI211_X1 U8503 ( .C1(n7130), .C2(n7129), .A(n10695), .B(n7215), .ZN(n7131)
         );
  INV_X1 U8504 ( .A(n7131), .ZN(n7144) );
  NAND2_X1 U8505 ( .A1(n7153), .A2(n7151), .ZN(n7132) );
  MUX2_X1 U8506 ( .A(n7133), .B(P2_REG2_REG_4__SCAN_IN), .S(n7134), .Z(n7150)
         );
  NAND2_X1 U8507 ( .A1(n7132), .A2(n7150), .ZN(n7155) );
  OR2_X1 U8508 ( .A1(n7134), .A2(n7133), .ZN(n7135) );
  NAND2_X1 U8509 ( .A1(n7155), .A2(n7135), .ZN(n7225) );
  INV_X1 U8510 ( .A(n7224), .ZN(n7137) );
  OAI21_X1 U8511 ( .B1(n7136), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7227), .ZN(
        n7142) );
  INV_X1 U8512 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7140) );
  NAND2_X1 U8513 ( .A1(n10676), .A2(n7137), .ZN(n7139) );
  INV_X1 U8514 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10459) );
  NOR2_X1 U8515 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10459), .ZN(n7210) );
  INV_X1 U8516 ( .A(n7210), .ZN(n7138) );
  OAI211_X1 U8517 ( .C1(n9263), .C2(n7140), .A(n7139), .B(n7138), .ZN(n7141)
         );
  AOI21_X1 U8518 ( .B1(n10710), .B2(n7142), .A(n7141), .ZN(n7143) );
  OAI211_X1 U8519 ( .C1(n7145), .C2(n10713), .A(n7144), .B(n7143), .ZN(
        P2_U3187) );
  AOI211_X1 U8520 ( .C1(n7148), .C2(n7147), .A(n10695), .B(n7146), .ZN(n7149)
         );
  INV_X1 U8521 ( .A(n7149), .ZN(n7166) );
  INV_X1 U8522 ( .A(n7150), .ZN(n7152) );
  NAND3_X1 U8523 ( .A1(n7153), .A2(n7152), .A3(n7151), .ZN(n7154) );
  AOI21_X1 U8524 ( .B1(n7155), .B2(n7154), .A(n10682), .ZN(n7164) );
  OR3_X1 U8525 ( .A1(n7158), .A2(n7157), .A3(n7156), .ZN(n7159) );
  AOI21_X1 U8526 ( .B1(n7160), .B2(n7159), .A(n10713), .ZN(n7163) );
  INV_X1 U8527 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7161) );
  NOR2_X1 U8528 ( .A1(n9263), .A2(n7161), .ZN(n7162) );
  AND2_X1 U8529 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3151), .ZN(n9080) );
  NOR4_X1 U8530 ( .A1(n7164), .A2(n7163), .A3(n7162), .A4(n9080), .ZN(n7165)
         );
  OAI211_X1 U8531 ( .C1(n10706), .C2(n7167), .A(n7166), .B(n7165), .ZN(
        P2_U3186) );
  NAND2_X1 U8532 ( .A1(n9353), .A2(P2_U3893), .ZN(n7168) );
  OAI21_X1 U8533 ( .B1(P2_U3893), .B2(n7912), .A(n7168), .ZN(P2_U3514) );
  OAI21_X1 U8534 ( .B1(n7170), .B2(n8353), .A(n7169), .ZN(n7855) );
  NAND2_X1 U8535 ( .A1(n7855), .A2(n5053), .ZN(n7174) );
  AOI22_X1 U8536 ( .A1(n10267), .A2(n9803), .B1(n10268), .B2(n9801), .ZN(n7173) );
  INV_X1 U8537 ( .A(n8353), .ZN(n8366) );
  XNOR2_X1 U8538 ( .A(n7171), .B(n8366), .ZN(n7172) );
  NAND2_X1 U8539 ( .A1(n7172), .A2(n10162), .ZN(n7857) );
  OAI211_X1 U8540 ( .C1(n7685), .C2(n5824), .A(n10782), .B(n7326), .ZN(n7853)
         );
  NAND4_X1 U8541 ( .A1(n7174), .A2(n7173), .A3(n7857), .A4(n7853), .ZN(n7243)
         );
  INV_X1 U8542 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7175) );
  OAI22_X1 U8543 ( .A1(n10340), .A2(n5824), .B1(n10834), .B2(n7175), .ZN(n7176) );
  AOI21_X1 U8544 ( .B1(n7243), .B2(n10834), .A(n7176), .ZN(n7177) );
  INV_X1 U8545 ( .A(n7177), .ZN(P1_U3471) );
  INV_X1 U8546 ( .A(n7178), .ZN(n7179) );
  NAND2_X1 U8547 ( .A1(n9612), .A2(n7179), .ZN(n7184) );
  INV_X1 U8548 ( .A(n7180), .ZN(n7181) );
  NAND2_X1 U8549 ( .A1(n7182), .A2(n7181), .ZN(n7183) );
  NAND2_X1 U8550 ( .A1(n7184), .A2(n7183), .ZN(n7185) );
  NAND2_X1 U8551 ( .A1(n7186), .A2(n7185), .ZN(n7192) );
  INV_X1 U8552 ( .A(n7187), .ZN(n8664) );
  INV_X1 U8553 ( .A(n7188), .ZN(n7189) );
  NOR3_X1 U8554 ( .A1(n8664), .A2(n9568), .A3(n7189), .ZN(n7191) );
  OAI21_X1 U8555 ( .B1(n7191), .B2(n7190), .A(n10846), .ZN(n7197) );
  OR2_X1 U8556 ( .A1(n7192), .A2(n10840), .ZN(n9360) );
  OAI22_X1 U8557 ( .A1(n9360), .A2(n7194), .B1(n7193), .B2(n10838), .ZN(n7195)
         );
  INV_X1 U8558 ( .A(n7195), .ZN(n7196) );
  OAI211_X1 U8559 ( .C1(n6263), .C2(n10846), .A(n7197), .B(n7196), .ZN(
        P2_U3233) );
  NAND2_X1 U8560 ( .A1(n7198), .A2(n7284), .ZN(n7199) );
  NAND2_X1 U8561 ( .A1(n7200), .A2(n7199), .ZN(n9012) );
  INV_X1 U8562 ( .A(n9012), .ZN(n7202) );
  XNOR2_X1 U8563 ( .A(n8600), .B(n9017), .ZN(n7203) );
  XNOR2_X1 U8564 ( .A(n7203), .B(n7384), .ZN(n9013) );
  INV_X1 U8565 ( .A(n9013), .ZN(n7201) );
  INV_X1 U8566 ( .A(n7203), .ZN(n7204) );
  NAND2_X1 U8567 ( .A1(n7204), .A2(n9149), .ZN(n7205) );
  XNOR2_X1 U8568 ( .A(n8600), .B(n9082), .ZN(n7206) );
  XNOR2_X1 U8569 ( .A(n7206), .B(n9148), .ZN(n9078) );
  NAND2_X1 U8570 ( .A1(n7206), .A2(n7484), .ZN(n7207) );
  XNOR2_X1 U8571 ( .A(n8635), .B(n7492), .ZN(n7289) );
  XNOR2_X1 U8572 ( .A(n7289), .B(n9147), .ZN(n7287) );
  XOR2_X1 U8573 ( .A(n7288), .B(n7287), .Z(n7214) );
  INV_X1 U8574 ( .A(n7208), .ZN(n7491) );
  NOR2_X1 U8575 ( .A1(n9094), .A2(n7484), .ZN(n7209) );
  AOI211_X1 U8576 ( .C1(n9081), .C2(n9146), .A(n7210), .B(n7209), .ZN(n7211)
         );
  OAI21_X1 U8577 ( .B1(n7550), .B2(n9114), .A(n7211), .ZN(n7212) );
  AOI21_X1 U8578 ( .B1(n7491), .B2(n9125), .A(n7212), .ZN(n7213) );
  OAI21_X1 U8579 ( .B1(n7214), .B2(n9133), .A(n7213), .ZN(P2_U3167) );
  AOI21_X1 U8580 ( .B1(n7216), .B2(n7224), .A(n7215), .ZN(n7218) );
  MUX2_X1 U8581 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n4947), .Z(n7338) );
  XNOR2_X1 U8582 ( .A(n7338), .B(n4948), .ZN(n7217) );
  NAND2_X1 U8583 ( .A1(n7218), .A2(n7217), .ZN(n7337) );
  OAI21_X1 U8584 ( .B1(n7218), .B2(n7217), .A(n7337), .ZN(n7237) );
  AOI22_X1 U8585 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(n4948), .B1(n7349), .B2(
        n6333), .ZN(n7221) );
  AOI21_X1 U8586 ( .B1(n7222), .B2(n7221), .A(n7348), .ZN(n7223) );
  NOR2_X1 U8587 ( .A1(n7223), .A2(n10713), .ZN(n7236) );
  NAND2_X1 U8588 ( .A1(n7225), .A2(n7224), .ZN(n7226) );
  AOI21_X1 U8589 ( .B1(n7229), .B2(n7228), .A(n7342), .ZN(n7230) );
  OR2_X1 U8590 ( .A1(n7230), .A2(n10682), .ZN(n7234) );
  NAND2_X1 U8591 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3151), .ZN(n7298) );
  NAND2_X1 U8592 ( .A1(n10676), .A2(n4948), .ZN(n7233) );
  NAND2_X1 U8593 ( .A1(n10698), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7232) );
  NAND4_X1 U8594 ( .A1(n7234), .A2(n7298), .A3(n7233), .A4(n7232), .ZN(n7235)
         );
  AOI211_X1 U8595 ( .C1(n7237), .C2(n10690), .A(n7236), .B(n7235), .ZN(n7238)
         );
  INV_X1 U8596 ( .A(n7238), .ZN(P2_U3188) );
  OAI22_X1 U8597 ( .A1(n10298), .A2(n7765), .B1(n10831), .B2(n6954), .ZN(n7239) );
  INV_X1 U8598 ( .A(n7239), .ZN(n7240) );
  OAI21_X1 U8599 ( .B1(n7241), .B2(n10830), .A(n7240), .ZN(P1_U3525) );
  OAI22_X1 U8600 ( .A1(n10298), .A2(n5824), .B1(n10831), .B2(n6957), .ZN(n7242) );
  AOI21_X1 U8601 ( .B1(n7243), .B2(n10831), .A(n7242), .ZN(n7244) );
  INV_X1 U8602 ( .A(n7244), .ZN(P1_U3528) );
  OAI22_X1 U8603 ( .A1(n10298), .A2(n5290), .B1(n10831), .B2(n5778), .ZN(n7245) );
  AOI21_X1 U8604 ( .B1(n7246), .B2(n10831), .A(n7245), .ZN(n7247) );
  INV_X1 U8605 ( .A(n7247), .ZN(P1_U3526) );
  OAI22_X1 U8606 ( .A1(n10298), .A2(n8520), .B1(n10831), .B2(n6950), .ZN(n7248) );
  INV_X1 U8607 ( .A(n7248), .ZN(n7249) );
  OAI21_X1 U8608 ( .B1(n7250), .B2(n10830), .A(n7249), .ZN(P1_U3523) );
  NAND2_X1 U8609 ( .A1(n7269), .A2(n7706), .ZN(n7252) );
  NAND2_X1 U8610 ( .A1(n5063), .A2(n8916), .ZN(n7251) );
  XNOR2_X1 U8611 ( .A(n7253), .B(n8883), .ZN(n7266) );
  AOI22_X1 U8612 ( .A1(n7254), .A2(n9806), .B1(n8916), .B2(n7706), .ZN(n7265)
         );
  NAND2_X1 U8613 ( .A1(n7256), .A2(n7255), .ZN(n7258) );
  INV_X1 U8614 ( .A(n7268), .ZN(n7260) );
  AOI21_X1 U8615 ( .B1(n7261), .B2(n7259), .A(n7260), .ZN(n7264) );
  AOI22_X1 U8616 ( .A1(n9768), .A2(n9805), .B1(n9767), .B2(n9807), .ZN(n7263)
         );
  AOI22_X1 U8617 ( .A1(n4944), .A2(n7706), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n8320), .ZN(n7262) );
  OAI211_X1 U8618 ( .C1(n7264), .C2(n9788), .A(n7263), .B(n7262), .ZN(P1_U3237) );
  NAND2_X1 U8619 ( .A1(n7266), .A2(n7265), .ZN(n7267) );
  NAND2_X1 U8620 ( .A1(n7269), .A2(n7276), .ZN(n7271) );
  NAND2_X1 U8621 ( .A1(n9805), .A2(n8916), .ZN(n7270) );
  AOI22_X1 U8622 ( .A1(n7254), .A2(n9805), .B1(n8916), .B2(n7276), .ZN(n7396)
         );
  XNOR2_X1 U8623 ( .A(n7395), .B(n7396), .ZN(n7399) );
  XOR2_X1 U8624 ( .A(n7399), .B(n7400), .Z(n7279) );
  NAND2_X1 U8625 ( .A1(n7273), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9781) );
  INV_X1 U8626 ( .A(n9781), .ZN(n9769) );
  INV_X1 U8627 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7274) );
  AOI22_X1 U8628 ( .A1(n9768), .A2(n9804), .B1(n9769), .B2(n7274), .ZN(n7278)
         );
  NOR2_X1 U8629 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7274), .ZN(n9838) );
  NOR2_X1 U8630 ( .A1(n9783), .A2(n10186), .ZN(n7275) );
  AOI211_X1 U8631 ( .C1(n7276), .C2(n4944), .A(n9838), .B(n7275), .ZN(n7277)
         );
  OAI211_X1 U8632 ( .C1(n7279), .C2(n9788), .A(n7278), .B(n7277), .ZN(P1_U3218) );
  OAI21_X1 U8633 ( .B1(n7280), .B2(n8663), .A(n7389), .ZN(n7379) );
  INV_X1 U8634 ( .A(n9017), .ZN(n7281) );
  NOR2_X1 U8635 ( .A1(n7281), .A2(n9559), .ZN(n7285) );
  XNOR2_X1 U8636 ( .A(n7282), .B(n8663), .ZN(n7283) );
  OAI222_X1 U8637 ( .A1(n9473), .A2(n7484), .B1(n9471), .B2(n7284), .C1(n9468), 
        .C2(n7283), .ZN(n7376) );
  AOI211_X1 U8638 ( .C1(n9525), .C2(n7379), .A(n7285), .B(n7376), .ZN(n10750)
         );
  OR2_X1 U8639 ( .A1(n10750), .A2(n9570), .ZN(n7286) );
  OAI21_X1 U8640 ( .B1(n9561), .B2(n6287), .A(n7286), .ZN(P2_U3462) );
  NAND2_X1 U8641 ( .A1(n7288), .A2(n7287), .ZN(n7291) );
  NAND2_X1 U8642 ( .A1(n7289), .A2(n7775), .ZN(n7290) );
  XNOR2_X1 U8643 ( .A(n7293), .B(n8630), .ZN(n7509) );
  XNOR2_X1 U8644 ( .A(n7509), .B(n9146), .ZN(n7295) );
  AOI21_X1 U8645 ( .B1(n7294), .B2(n7295), .A(n9133), .ZN(n7297) );
  INV_X1 U8646 ( .A(n7295), .ZN(n7296) );
  NAND2_X1 U8647 ( .A1(n7297), .A2(n7511), .ZN(n7303) );
  INV_X1 U8648 ( .A(n7872), .ZN(n7301) );
  NAND2_X1 U8649 ( .A1(n9081), .A2(n9145), .ZN(n7299) );
  OAI211_X1 U8650 ( .C1(n7775), .C2(n9094), .A(n7299), .B(n7298), .ZN(n7300)
         );
  AOI21_X1 U8651 ( .B1(n7301), .B2(n9125), .A(n7300), .ZN(n7302) );
  OAI211_X1 U8652 ( .C1(n7873), .C2(n9114), .A(n7303), .B(n7302), .ZN(P2_U3179) );
  AOI21_X1 U8653 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n7309), .A(n7304), .ZN(
        n7307) );
  MUX2_X1 U8654 ( .A(n7305), .B(P1_REG1_REG_11__SCAN_IN), .S(n7430), .Z(n7306)
         );
  NOR2_X1 U8655 ( .A1(n7307), .A2(n7306), .ZN(n7429) );
  AOI211_X1 U8656 ( .C1(n7307), .C2(n7306), .A(n7429), .B(n9895), .ZN(n7317)
         );
  AOI21_X1 U8657 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n7309), .A(n7308), .ZN(
        n7312) );
  NAND2_X1 U8658 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7430), .ZN(n7310) );
  OAI21_X1 U8659 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7430), .A(n7310), .ZN(
        n7311) );
  NOR2_X1 U8660 ( .A1(n7312), .A2(n7311), .ZN(n7422) );
  AOI211_X1 U8661 ( .C1(n7312), .C2(n7311), .A(n7422), .B(n9953), .ZN(n7316)
         );
  INV_X1 U8662 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7314) );
  NAND2_X1 U8663 ( .A1(n9930), .A2(n7430), .ZN(n7313) );
  NAND2_X1 U8664 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n8096) );
  OAI211_X1 U8665 ( .C1(n7314), .C2(n9920), .A(n7313), .B(n8096), .ZN(n7315)
         );
  OR3_X1 U8666 ( .A1(n7317), .A2(n7316), .A3(n7315), .ZN(P1_U3254) );
  INV_X1 U8667 ( .A(n8232), .ZN(n8172) );
  INV_X1 U8668 ( .A(n7318), .ZN(n7320) );
  OAI222_X1 U8669 ( .A1(n8172), .A2(P1_U3086), .B1(n10354), .B2(n7320), .C1(
        n7319), .C2(n10350), .ZN(P1_U3339) );
  INV_X1 U8670 ( .A(n9207), .ZN(n9233) );
  OAI222_X1 U8671 ( .A1(n7792), .A2(n7321), .B1(n9625), .B2(n7320), .C1(
        P2_U3151), .C2(n9233), .ZN(P2_U3279) );
  OAI21_X1 U8672 ( .B1(n7323), .B2(n8358), .A(n7322), .ZN(n7576) );
  NAND2_X1 U8673 ( .A1(n7324), .A2(n8354), .ZN(n7325) );
  NOR2_X1 U8674 ( .A1(n7325), .A2(n8358), .ZN(n7460) );
  AOI21_X1 U8675 ( .B1(n8358), .B2(n7325), .A(n7460), .ZN(n7587) );
  AOI22_X1 U8676 ( .A1(n10267), .A2(n9802), .B1(n10268), .B2(n9800), .ZN(n7328) );
  INV_X1 U8677 ( .A(n7326), .ZN(n7327) );
  INV_X1 U8678 ( .A(n8313), .ZN(n7333) );
  OAI211_X1 U8679 ( .C1(n7327), .C2(n7333), .A(n10782), .B(n7462), .ZN(n7582)
         );
  OAI211_X1 U8680 ( .C1(n7587), .C2(n10791), .A(n7328), .B(n7582), .ZN(n7329)
         );
  AOI21_X1 U8681 ( .B1(n5053), .B2(n7576), .A(n7329), .ZN(n7336) );
  OAI22_X1 U8682 ( .A1(n10298), .A2(n7333), .B1(n10831), .B2(n5836), .ZN(n7330) );
  INV_X1 U8683 ( .A(n7330), .ZN(n7331) );
  OAI21_X1 U8684 ( .B1(n7336), .B2(n10830), .A(n7331), .ZN(P1_U3529) );
  INV_X1 U8685 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7332) );
  OAI22_X1 U8686 ( .A1(n10340), .A2(n7333), .B1(n10834), .B2(n7332), .ZN(n7334) );
  INV_X1 U8687 ( .A(n7334), .ZN(n7335) );
  OAI21_X1 U8688 ( .B1(n7336), .B2(n6207), .A(n7335), .ZN(P1_U3474) );
  OAI21_X1 U8689 ( .B1(n7338), .B2(n7349), .A(n7337), .ZN(n7340) );
  MUX2_X1 U8690 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n4947), .Z(n7529) );
  XNOR2_X1 U8691 ( .A(n7529), .B(n7537), .ZN(n7339) );
  NAND2_X1 U8692 ( .A1(n7340), .A2(n7339), .ZN(n7530) );
  OAI21_X1 U8693 ( .B1(n7340), .B2(n7339), .A(n7530), .ZN(n7341) );
  NAND2_X1 U8694 ( .A1(n7341), .A2(n10690), .ZN(n7356) );
  INV_X1 U8695 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7347) );
  AOI21_X1 U8696 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n7349), .A(n7342), .ZN(
        n7536) );
  AND2_X1 U8697 ( .A1(n7343), .A2(n7813), .ZN(n7344) );
  OAI21_X1 U8698 ( .B1(n7538), .B2(n7344), .A(n10710), .ZN(n7346) );
  NOR2_X1 U8699 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6347), .ZN(n7515) );
  INV_X1 U8700 ( .A(n7515), .ZN(n7345) );
  OAI211_X1 U8701 ( .C1(n9263), .C2(n7347), .A(n7346), .B(n7345), .ZN(n7354)
         );
  NAND2_X1 U8702 ( .A1(n7349), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7350) );
  AOI21_X1 U8703 ( .B1(n6346), .B2(n7351), .A(n7523), .ZN(n7352) );
  NOR2_X1 U8704 ( .A1(n7352), .A2(n10713), .ZN(n7353) );
  AOI211_X1 U8705 ( .C1(n10676), .C2(n7537), .A(n7354), .B(n7353), .ZN(n7355)
         );
  NAND2_X1 U8706 ( .A1(n7356), .A2(n7355), .ZN(P2_U3189) );
  INV_X1 U8707 ( .A(n7357), .ZN(n7364) );
  NOR2_X1 U8708 ( .A1(n8712), .A2(n7371), .ZN(n7482) );
  INV_X1 U8709 ( .A(n7482), .ZN(n7358) );
  NAND2_X1 U8710 ( .A1(n8140), .A2(n7358), .ZN(n10844) );
  INV_X1 U8711 ( .A(n10838), .ZN(n10770) );
  AOI22_X1 U8712 ( .A1(n10768), .A2(n7359), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n10770), .ZN(n7360) );
  OAI21_X1 U8713 ( .B1(n6246), .B2(n10846), .A(n7360), .ZN(n7361) );
  AOI21_X1 U8714 ( .B1(n9377), .B2(n7362), .A(n7361), .ZN(n7363) );
  OAI21_X1 U8715 ( .B1(n7364), .B2(n4949), .A(n7363), .ZN(P2_U3232) );
  INV_X1 U8716 ( .A(n7365), .ZN(n7367) );
  OAI222_X1 U8717 ( .A1(n7792), .A2(n7366), .B1(n9625), .B2(n7367), .C1(n5210), 
        .C2(P2_U3151), .ZN(P2_U3278) );
  INV_X1 U8718 ( .A(n9922), .ZN(n9911) );
  OAI222_X1 U8719 ( .A1(n10350), .A2(n7368), .B1(n10354), .B2(n7367), .C1(
        P1_U3086), .C2(n9911), .ZN(P1_U3338) );
  NOR2_X1 U8720 ( .A1(n10838), .A2(n6275), .ZN(n7370) );
  AOI211_X1 U8721 ( .C1(n7372), .C2(n7371), .A(n7370), .B(n7369), .ZN(n7375)
         );
  AOI22_X1 U8722 ( .A1(n7373), .A2(n9377), .B1(n4949), .B2(
        P2_REG2_REG_2__SCAN_IN), .ZN(n7374) );
  OAI21_X1 U8723 ( .B1(n7375), .B2(n4949), .A(n7374), .ZN(P2_U3231) );
  INV_X1 U8724 ( .A(n7376), .ZN(n7381) );
  AOI22_X1 U8725 ( .A1(n10768), .A2(n9017), .B1(n10770), .B2(n10466), .ZN(
        n7377) );
  OAI21_X1 U8726 ( .B1(n6286), .B2(n10846), .A(n7377), .ZN(n7378) );
  AOI21_X1 U8727 ( .B1(n7379), .B2(n9377), .A(n7378), .ZN(n7380) );
  OAI21_X1 U8728 ( .B1(n7381), .B2(n4949), .A(n7380), .ZN(P2_U3230) );
  AOI211_X1 U8729 ( .C1(n7388), .C2(n7383), .A(n9468), .B(n7382), .ZN(n7386)
         );
  OAI22_X1 U8730 ( .A1(n7775), .A2(n9473), .B1(n7384), .B2(n9471), .ZN(n7385)
         );
  OR2_X1 U8731 ( .A1(n7386), .A2(n7385), .ZN(n7477) );
  INV_X1 U8732 ( .A(n7477), .ZN(n7394) );
  INV_X1 U8733 ( .A(n7388), .ZN(n8729) );
  NAND3_X1 U8734 ( .A1(n7389), .A2(n8729), .A3(n8732), .ZN(n7390) );
  NAND2_X1 U8735 ( .A1(n7387), .A2(n7390), .ZN(n7479) );
  NOR2_X1 U8736 ( .A1(n10846), .A2(n7133), .ZN(n7392) );
  OAI22_X1 U8737 ( .A1(n9360), .A2(n7476), .B1(n9083), .B2(n10838), .ZN(n7391)
         );
  AOI211_X1 U8738 ( .C1(n7479), .C2(n9377), .A(n7392), .B(n7391), .ZN(n7393)
         );
  OAI21_X1 U8739 ( .B1(n7394), .B2(n4949), .A(n7393), .ZN(P2_U3229) );
  INV_X1 U8740 ( .A(n7395), .ZN(n7397) );
  AND2_X1 U8741 ( .A1(n7397), .A2(n7396), .ZN(n7398) );
  NAND2_X1 U8742 ( .A1(n8977), .A2(n9728), .ZN(n7402) );
  NAND2_X1 U8743 ( .A1(n9804), .A2(n8916), .ZN(n7401) );
  NAND2_X1 U8744 ( .A1(n7402), .A2(n7401), .ZN(n7403) );
  XNOR2_X1 U8745 ( .A(n7403), .B(n8963), .ZN(n7404) );
  AOI22_X1 U8746 ( .A1(n7254), .A2(n9804), .B1(n8916), .B2(n9728), .ZN(n7405)
         );
  XNOR2_X1 U8747 ( .A(n7404), .B(n7405), .ZN(n9722) );
  INV_X1 U8748 ( .A(n7404), .ZN(n7406) );
  OR2_X1 U8749 ( .A1(n7406), .A2(n7405), .ZN(n7407) );
  NAND2_X1 U8750 ( .A1(n8977), .A2(n7689), .ZN(n7409) );
  NAND2_X1 U8751 ( .A1(n9803), .A2(n8965), .ZN(n7408) );
  NAND2_X1 U8752 ( .A1(n7409), .A2(n7408), .ZN(n7410) );
  XNOR2_X1 U8753 ( .A(n7410), .B(n8963), .ZN(n7412) );
  NAND2_X1 U8754 ( .A1(n7439), .A2(n7438), .ZN(n7413) );
  AOI22_X1 U8755 ( .A1(n7254), .A2(n9803), .B1(n7689), .B2(n8965), .ZN(n7437)
         );
  XNOR2_X1 U8756 ( .A(n7413), .B(n7437), .ZN(n7420) );
  INV_X1 U8757 ( .A(n7414), .ZN(n7688) );
  AOI22_X1 U8758 ( .A1(n9768), .A2(n9802), .B1(n9769), .B2(n7688), .ZN(n7419)
         );
  NAND2_X1 U8759 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9869) );
  INV_X1 U8760 ( .A(n9869), .ZN(n7417) );
  NOR2_X1 U8761 ( .A1(n9783), .A2(n7415), .ZN(n7416) );
  AOI211_X1 U8762 ( .C1(n7689), .C2(n4944), .A(n7417), .B(n7416), .ZN(n7418)
         );
  OAI211_X1 U8763 ( .C1(n7420), .C2(n9788), .A(n7419), .B(n7418), .ZN(P1_U3227) );
  NOR2_X1 U8764 ( .A1(n7621), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7421) );
  AOI21_X1 U8765 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7621), .A(n7421), .ZN(
        n7424) );
  AOI21_X1 U8766 ( .B1(n7430), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7422), .ZN(
        n7423) );
  NAND2_X1 U8767 ( .A1(n7424), .A2(n7423), .ZN(n7616) );
  OAI21_X1 U8768 ( .B1(n7424), .B2(n7423), .A(n7616), .ZN(n7425) );
  INV_X1 U8769 ( .A(n7425), .ZN(n7436) );
  NOR2_X1 U8770 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7426), .ZN(n8197) );
  NOR2_X1 U8771 ( .A1(n9947), .A2(n7428), .ZN(n7427) );
  AOI211_X1 U8772 ( .C1(n9950), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n8197), .B(
        n7427), .ZN(n7435) );
  AOI22_X1 U8773 ( .A1(n7621), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n5699), .B2(
        n7428), .ZN(n7432) );
  AOI21_X1 U8774 ( .B1(n7430), .B2(P1_REG1_REG_11__SCAN_IN), .A(n7429), .ZN(
        n7431) );
  NAND2_X1 U8775 ( .A1(n7432), .A2(n7431), .ZN(n7620) );
  OAI21_X1 U8776 ( .B1(n7432), .B2(n7431), .A(n7620), .ZN(n7433) );
  NAND2_X1 U8777 ( .A1(n7433), .A2(n9944), .ZN(n7434) );
  OAI211_X1 U8778 ( .C1(n7436), .C2(n9953), .A(n7435), .B(n7434), .ZN(P1_U3255) );
  NAND2_X1 U8779 ( .A1(n8977), .A2(n7851), .ZN(n7441) );
  NAND2_X1 U8780 ( .A1(n9802), .A2(n8916), .ZN(n7440) );
  NAND2_X1 U8781 ( .A1(n7441), .A2(n7440), .ZN(n7442) );
  XNOR2_X1 U8782 ( .A(n7442), .B(n8883), .ZN(n7445) );
  NAND2_X1 U8783 ( .A1(n7851), .A2(n8965), .ZN(n7444) );
  NAND2_X1 U8784 ( .A1(n7254), .A2(n9802), .ZN(n7443) );
  AND2_X1 U8785 ( .A1(n7444), .A2(n7443), .ZN(n7446) );
  AND2_X1 U8786 ( .A1(n7445), .A2(n7446), .ZN(n7712) );
  INV_X1 U8787 ( .A(n7712), .ZN(n7449) );
  INV_X1 U8788 ( .A(n7445), .ZN(n7448) );
  INV_X1 U8789 ( .A(n7446), .ZN(n7447) );
  NAND2_X1 U8790 ( .A1(n7448), .A2(n7447), .ZN(n7711) );
  NAND2_X1 U8791 ( .A1(n7449), .A2(n7711), .ZN(n7450) );
  XNOR2_X1 U8792 ( .A(n7713), .B(n7450), .ZN(n7456) );
  INV_X1 U8793 ( .A(n7848), .ZN(n7451) );
  AOI22_X1 U8794 ( .A1(n9768), .A2(n9801), .B1(n9769), .B2(n7451), .ZN(n7455)
         );
  NOR2_X1 U8795 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7452), .ZN(n9883) );
  NOR2_X1 U8796 ( .A1(n9783), .A2(n9726), .ZN(n7453) );
  AOI211_X1 U8797 ( .C1(n7851), .C2(n4944), .A(n9883), .B(n7453), .ZN(n7454)
         );
  OAI211_X1 U8798 ( .C1(n7456), .C2(n9788), .A(n7455), .B(n7454), .ZN(P1_U3239) );
  INV_X1 U8799 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7468) );
  OAI21_X1 U8800 ( .B1(n7458), .B2(n8359), .A(n7457), .ZN(n7869) );
  NAND2_X1 U8801 ( .A1(n7869), .A2(n5053), .ZN(n7465) );
  AOI22_X1 U8802 ( .A1(n10267), .A2(n9801), .B1(n10268), .B2(n9799), .ZN(n7464) );
  INV_X1 U8803 ( .A(n8360), .ZN(n7459) );
  NOR2_X1 U8804 ( .A1(n7460), .A2(n7459), .ZN(n7498) );
  XNOR2_X1 U8805 ( .A(n7498), .B(n8359), .ZN(n7461) );
  NAND2_X1 U8806 ( .A1(n7461), .A2(n10162), .ZN(n7871) );
  AOI21_X1 U8807 ( .B1(n7462), .B2(n8374), .A(n10174), .ZN(n7463) );
  NAND2_X1 U8808 ( .A1(n7463), .A2(n7501), .ZN(n7867) );
  NAND4_X1 U8809 ( .A1(n7465), .A2(n7464), .A3(n7871), .A4(n7867), .ZN(n7473)
         );
  NAND2_X1 U8810 ( .A1(n7473), .A2(n10834), .ZN(n7467) );
  NAND2_X1 U8811 ( .A1(n6205), .A2(n8374), .ZN(n7466) );
  OAI211_X1 U8812 ( .C1(n10834), .C2(n7468), .A(n7467), .B(n7466), .ZN(
        P1_U3477) );
  INV_X1 U8813 ( .A(n7469), .ZN(n7471) );
  INV_X1 U8814 ( .A(n9929), .ZN(n9915) );
  OAI222_X1 U8815 ( .A1(n10350), .A2(n7470), .B1(n10354), .B2(n7471), .C1(
        P1_U3086), .C2(n9915), .ZN(P1_U3337) );
  OAI222_X1 U8816 ( .A1(n7792), .A2(n7472), .B1(n9625), .B2(n7471), .C1(n10705), .C2(P2_U3151), .ZN(P2_U3277) );
  NAND2_X1 U8817 ( .A1(n7473), .A2(n10831), .ZN(n7475) );
  INV_X1 U8818 ( .A(n10298), .ZN(n7919) );
  NAND2_X1 U8819 ( .A1(n7919), .A2(n8374), .ZN(n7474) );
  OAI211_X1 U8820 ( .C1(n10831), .C2(n6958), .A(n7475), .B(n7474), .ZN(
        P1_U3530) );
  NOR2_X1 U8821 ( .A1(n7476), .A2(n9559), .ZN(n7478) );
  AOI211_X1 U8822 ( .C1(n9525), .C2(n7479), .A(n7478), .B(n7477), .ZN(n10752)
         );
  OR2_X1 U8823 ( .A1(n10752), .A2(n9570), .ZN(n7480) );
  OAI21_X1 U8824 ( .B1(n9561), .B2(n7123), .A(n7480), .ZN(P2_U3463) );
  OAI21_X1 U8825 ( .B1(n7481), .B2(n8665), .A(n7771), .ZN(n7553) );
  INV_X1 U8826 ( .A(n7553), .ZN(n7495) );
  NAND2_X1 U8827 ( .A1(n10846), .A2(n7482), .ZN(n8593) );
  XNOR2_X1 U8828 ( .A(n5050), .B(n8665), .ZN(n7488) );
  INV_X1 U8829 ( .A(n8140), .ZN(n7486) );
  OAI22_X1 U8830 ( .A1(n7484), .A2(n9471), .B1(n7483), .B2(n9473), .ZN(n7485)
         );
  AOI21_X1 U8831 ( .B1(n7553), .B2(n7486), .A(n7485), .ZN(n7487) );
  OAI21_X1 U8832 ( .B1(n7488), .B2(n9468), .A(n7487), .ZN(n7551) );
  INV_X1 U8833 ( .A(n7551), .ZN(n7489) );
  MUX2_X1 U8834 ( .A(n7490), .B(n7489), .S(n10846), .Z(n7494) );
  AOI22_X1 U8835 ( .A1(n10768), .A2(n7492), .B1(n10770), .B2(n7491), .ZN(n7493) );
  OAI211_X1 U8836 ( .C1(n7495), .C2(n8593), .A(n7494), .B(n7493), .ZN(P2_U3228) );
  OAI21_X1 U8837 ( .B1(n7497), .B2(n7499), .A(n7496), .ZN(n7808) );
  OAI21_X1 U8838 ( .B1(n7498), .B2(n8359), .A(n8369), .ZN(n7500) );
  INV_X1 U8839 ( .A(n7499), .ZN(n8372) );
  XNOR2_X1 U8840 ( .A(n7500), .B(n8372), .ZN(n7800) );
  NAND2_X1 U8841 ( .A1(n7800), .A2(n10162), .ZN(n7503) );
  AOI211_X1 U8842 ( .C1(n7807), .C2(n7501), .A(n10174), .B(n7560), .ZN(n7502)
         );
  AOI21_X1 U8843 ( .B1(n10268), .B2(n9798), .A(n7502), .ZN(n7804) );
  OAI211_X1 U8844 ( .C1(n8373), .C2(n10796), .A(n7503), .B(n7804), .ZN(n7504)
         );
  AOI21_X1 U8845 ( .B1(n5053), .B2(n7808), .A(n7504), .ZN(n7508) );
  AOI22_X1 U8846 ( .A1(n7919), .A2(n7807), .B1(n10830), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7505) );
  OAI21_X1 U8847 ( .B1(n7508), .B2(n10830), .A(n7505), .ZN(P1_U3531) );
  OAI22_X1 U8848 ( .A1(n10340), .A2(n5295), .B1(n10834), .B2(n5863), .ZN(n7506) );
  INV_X1 U8849 ( .A(n7506), .ZN(n7507) );
  OAI21_X1 U8850 ( .B1(n7508), .B2(n6207), .A(n7507), .ZN(P1_U3480) );
  NAND2_X1 U8851 ( .A1(n7509), .A2(n9146), .ZN(n7510) );
  XNOR2_X1 U8852 ( .A(n8705), .B(n8635), .ZN(n7603) );
  XNOR2_X1 U8853 ( .A(n7603), .B(n9145), .ZN(n7513) );
  OAI21_X1 U8854 ( .B1(n7512), .B2(n7513), .A(n7605), .ZN(n7520) );
  NOR2_X1 U8855 ( .A1(n9114), .A2(n7844), .ZN(n7519) );
  INV_X1 U8856 ( .A(n7514), .ZN(n7814) );
  NAND2_X1 U8857 ( .A1(n9125), .A2(n7814), .ZN(n7517) );
  INV_X1 U8858 ( .A(n9094), .ZN(n9126) );
  AOI21_X1 U8859 ( .B1(n9126), .B2(n9146), .A(n7515), .ZN(n7516) );
  OAI211_X1 U8860 ( .C1(n7673), .C2(n9129), .A(n7517), .B(n7516), .ZN(n7518)
         );
  AOI211_X1 U8861 ( .C1(n7520), .C2(n9091), .A(n7519), .B(n7518), .ZN(n7521)
         );
  INV_X1 U8862 ( .A(n7521), .ZN(P2_U3153) );
  NOR2_X1 U8863 ( .A1(n7537), .A2(n7522), .ZN(n7524) );
  NAND2_X1 U8864 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7630), .ZN(n7640) );
  OAI21_X1 U8865 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7630), .A(n7640), .ZN(
        n7525) );
  AOI21_X1 U8866 ( .B1(n7526), .B2(n7525), .A(n7642), .ZN(n7548) );
  MUX2_X1 U8867 ( .A(n8002), .B(n7527), .S(n4946), .Z(n7632) );
  XNOR2_X1 U8868 ( .A(n7632), .B(n7630), .ZN(n7533) );
  OR2_X1 U8869 ( .A1(n7529), .A2(n7528), .ZN(n7531) );
  NAND2_X1 U8870 ( .A1(n7531), .A2(n7530), .ZN(n7532) );
  NAND2_X1 U8871 ( .A1(n7533), .A2(n7532), .ZN(n7633) );
  OAI21_X1 U8872 ( .B1(n7533), .B2(n7532), .A(n7633), .ZN(n7546) );
  INV_X1 U8873 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7535) );
  NAND2_X1 U8874 ( .A1(n10676), .A2(n5073), .ZN(n7534) );
  NAND2_X1 U8875 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7610) );
  OAI211_X1 U8876 ( .C1(n9263), .C2(n7535), .A(n7534), .B(n7610), .ZN(n7545)
         );
  NOR2_X1 U8877 ( .A1(n7537), .A2(n7536), .ZN(n7539) );
  NAND2_X1 U8878 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7630), .ZN(n7540) );
  OAI21_X1 U8879 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7630), .A(n7540), .ZN(
        n7541) );
  NOR2_X1 U8880 ( .A1(n7542), .A2(n7541), .ZN(n7629) );
  AOI21_X1 U8881 ( .B1(n7542), .B2(n7541), .A(n7629), .ZN(n7543) );
  NOR2_X1 U8882 ( .A1(n7543), .A2(n10682), .ZN(n7544) );
  AOI211_X1 U8883 ( .C1(n10690), .C2(n7546), .A(n7545), .B(n7544), .ZN(n7547)
         );
  OAI21_X1 U8884 ( .B1(n7548), .B2(n10713), .A(n7547), .ZN(P2_U3190) );
  INV_X1 U8885 ( .A(n9305), .ZN(n9283) );
  NAND2_X1 U8886 ( .A1(n9283), .A2(P2_U3893), .ZN(n7549) );
  OAI21_X1 U8887 ( .B1(P2_U3893), .B2(n6097), .A(n7549), .ZN(P2_U3518) );
  INV_X1 U8888 ( .A(n8141), .ZN(n7554) );
  NOR2_X1 U8889 ( .A1(n7550), .A2(n9559), .ZN(n7552) );
  AOI211_X1 U8890 ( .C1(n7554), .C2(n7553), .A(n7552), .B(n7551), .ZN(n10754)
         );
  OR2_X1 U8891 ( .A1(n10754), .A2(n9570), .ZN(n7555) );
  OAI21_X1 U8892 ( .B1(n9561), .B2(n6314), .A(n7555), .ZN(P2_U3464) );
  OAI21_X1 U8893 ( .B1(n7557), .B2(n8460), .A(n7556), .ZN(n7589) );
  NAND3_X1 U8894 ( .A1(n7558), .A2(n8460), .A3(n8536), .ZN(n7559) );
  NAND2_X1 U8895 ( .A1(n10790), .A2(n7559), .ZN(n7588) );
  NAND2_X1 U8896 ( .A1(n7588), .A2(n10162), .ZN(n7563) );
  AOI22_X1 U8897 ( .A1(n10267), .A2(n9799), .B1(n10268), .B2(n9797), .ZN(n7562) );
  OAI21_X1 U8898 ( .B1(n7560), .B2(n7567), .A(n10782), .ZN(n7561) );
  OR2_X1 U8899 ( .A1(n10784), .A2(n7561), .ZN(n7593) );
  NAND3_X1 U8900 ( .A1(n7563), .A2(n7562), .A3(n7593), .ZN(n7564) );
  AOI21_X1 U8901 ( .B1(n7589), .B2(n5053), .A(n7564), .ZN(n7570) );
  AOI22_X1 U8902 ( .A1(n7919), .A2(n7969), .B1(n10830), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7565) );
  OAI21_X1 U8903 ( .B1(n7570), .B2(n10830), .A(n7565), .ZN(P1_U3532) );
  INV_X1 U8904 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7566) );
  OAI22_X1 U8905 ( .A1(n7567), .A2(n10340), .B1(n10834), .B2(n7566), .ZN(n7568) );
  INV_X1 U8906 ( .A(n7568), .ZN(n7569) );
  OAI21_X1 U8907 ( .B1(n7570), .B2(n6207), .A(n7569), .ZN(P1_U3483) );
  NAND2_X1 U8908 ( .A1(n7572), .A2(n7571), .ZN(n7573) );
  NAND2_X1 U8909 ( .A1(n10732), .A2(n10162), .ZN(n10160) );
  OR2_X1 U8910 ( .A1(n7574), .A2(n9946), .ZN(n10811) );
  NAND2_X1 U8911 ( .A1(n10786), .A2(n10811), .ZN(n7575) );
  NAND2_X1 U8912 ( .A1(n7576), .A2(n10189), .ZN(n7586) );
  INV_X1 U8913 ( .A(n7577), .ZN(n7578) );
  NAND2_X1 U8914 ( .A1(n10732), .A2(n10268), .ZN(n10185) );
  AND2_X1 U8915 ( .A1(n10732), .A2(n10267), .ZN(n10195) );
  OAI22_X1 U8916 ( .A1(n10732), .A2(n7579), .B1(n8310), .B2(n10729), .ZN(n7580) );
  AOI21_X1 U8917 ( .B1(n10195), .B2(n9802), .A(n7580), .ZN(n7581) );
  OAI21_X1 U8918 ( .B1(n8373), .B2(n10185), .A(n7581), .ZN(n7584) );
  NAND2_X1 U8919 ( .A1(n10732), .A2(n9946), .ZN(n10184) );
  NOR2_X1 U8920 ( .A1(n7582), .A2(n10184), .ZN(n7583) );
  AOI211_X1 U8921 ( .C1(n10809), .C2(n8313), .A(n7584), .B(n7583), .ZN(n7585)
         );
  OAI211_X1 U8922 ( .C1(n7587), .C2(n10160), .A(n7586), .B(n7585), .ZN(
        P1_U3286) );
  INV_X1 U8923 ( .A(n7588), .ZN(n7598) );
  NAND2_X1 U8924 ( .A1(n7589), .A2(n10189), .ZN(n7597) );
  INV_X1 U8925 ( .A(n10195), .ZN(n10156) );
  INV_X1 U8926 ( .A(n10185), .ZN(n10153) );
  OAI22_X1 U8927 ( .A1(n10732), .A2(n7590), .B1(n7965), .B2(n10729), .ZN(n7591) );
  AOI21_X1 U8928 ( .B1(n10153), .B2(n9797), .A(n7591), .ZN(n7592) );
  OAI21_X1 U8929 ( .B1(n7966), .B2(n10156), .A(n7592), .ZN(n7595) );
  NOR2_X1 U8930 ( .A1(n7593), .A2(n10184), .ZN(n7594) );
  AOI211_X1 U8931 ( .C1(n10809), .C2(n7969), .A(n7595), .B(n7594), .ZN(n7596)
         );
  OAI211_X1 U8932 ( .C1(n7598), .C2(n10160), .A(n7597), .B(n7596), .ZN(
        P1_U3283) );
  INV_X1 U8933 ( .A(n7599), .ZN(n7602) );
  OAI222_X1 U8934 ( .A1(n7792), .A2(n7600), .B1(n9625), .B2(n7602), .C1(n8696), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OAI222_X1 U8935 ( .A1(n9946), .A2(P1_U3086), .B1(n10354), .B2(n7602), .C1(
        n7601), .C2(n10350), .ZN(P1_U3336) );
  INV_X1 U8936 ( .A(n8004), .ZN(n7615) );
  INV_X1 U8937 ( .A(n7605), .ZN(n7604) );
  XNOR2_X1 U8938 ( .A(n8004), .B(n8635), .ZN(n7663) );
  XNOR2_X1 U8939 ( .A(n7663), .B(n9144), .ZN(n7606) );
  NOR3_X1 U8940 ( .A1(n7604), .A2(n5052), .A3(n7606), .ZN(n7608) );
  INV_X1 U8941 ( .A(n7665), .ZN(n7607) );
  OAI21_X1 U8942 ( .B1(n7608), .B2(n7607), .A(n9091), .ZN(n7614) );
  INV_X1 U8943 ( .A(n7609), .ZN(n8003) );
  NAND2_X1 U8944 ( .A1(n9081), .A2(n9143), .ZN(n7611) );
  OAI211_X1 U8945 ( .C1(n8704), .C2(n9094), .A(n7611), .B(n7610), .ZN(n7612)
         );
  AOI21_X1 U8946 ( .B1(n8003), .B2(n9125), .A(n7612), .ZN(n7613) );
  OAI211_X1 U8947 ( .C1(n7615), .C2(n9114), .A(n7614), .B(n7613), .ZN(P2_U3161) );
  OAI21_X1 U8948 ( .B1(n7621), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7616), .ZN(
        n7619) );
  NAND2_X1 U8949 ( .A1(n7823), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7617) );
  OAI21_X1 U8950 ( .B1(n7823), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7617), .ZN(
        n7618) );
  NOR2_X1 U8951 ( .A1(n7618), .A2(n7619), .ZN(n7822) );
  AOI211_X1 U8952 ( .C1(n7619), .C2(n7618), .A(n7822), .B(n9953), .ZN(n7628)
         );
  OAI21_X1 U8953 ( .B1(n7621), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7620), .ZN(
        n7623) );
  XNOR2_X1 U8954 ( .A(n7823), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n7622) );
  NOR2_X1 U8955 ( .A1(n7623), .A2(n7622), .ZN(n7818) );
  AOI211_X1 U8956 ( .C1(n7623), .C2(n7622), .A(n7818), .B(n9895), .ZN(n7627)
         );
  INV_X1 U8957 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7625) );
  NAND2_X1 U8958 ( .A1(n9930), .A2(n7823), .ZN(n7624) );
  NAND2_X1 U8959 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8221) );
  OAI211_X1 U8960 ( .C1(n7625), .C2(n9920), .A(n7624), .B(n8221), .ZN(n7626)
         );
  OR3_X1 U8961 ( .A1(n7628), .A2(n7627), .A3(n7626), .ZN(P1_U3256) );
  XNOR2_X1 U8962 ( .A(n7748), .B(n7749), .ZN(n7631) );
  AOI21_X1 U8963 ( .B1(n7631), .B2(n6376), .A(n7750), .ZN(n7649) );
  MUX2_X1 U8964 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n4947), .Z(n7741) );
  XNOR2_X1 U8965 ( .A(n7741), .B(n7749), .ZN(n7636) );
  NAND2_X1 U8966 ( .A1(n5073), .A2(n7632), .ZN(n7634) );
  NAND2_X1 U8967 ( .A1(n7634), .A2(n7633), .ZN(n7635) );
  NAND2_X1 U8968 ( .A1(n7636), .A2(n7635), .ZN(n7742) );
  OAI21_X1 U8969 ( .B1(n7636), .B2(n7635), .A(n7742), .ZN(n7647) );
  INV_X1 U8970 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7639) );
  NAND2_X1 U8971 ( .A1(n10676), .A2(n7749), .ZN(n7638) );
  NOR2_X1 U8972 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6378), .ZN(n7671) );
  INV_X1 U8973 ( .A(n7671), .ZN(n7637) );
  OAI211_X1 U8974 ( .C1(n7639), .C2(n9263), .A(n7638), .B(n7637), .ZN(n7646)
         );
  INV_X1 U8975 ( .A(n7640), .ZN(n7641) );
  AOI21_X1 U8976 ( .B1(n6377), .B2(n7643), .A(n7734), .ZN(n7644) );
  NOR2_X1 U8977 ( .A1(n7644), .A2(n10713), .ZN(n7645) );
  AOI211_X1 U8978 ( .C1(n10690), .C2(n7647), .A(n7646), .B(n7645), .ZN(n7648)
         );
  OAI21_X1 U8979 ( .B1(n7649), .B2(n10682), .A(n7648), .ZN(P2_U3191) );
  NAND2_X1 U8980 ( .A1(n7695), .A2(n10343), .ZN(n7651) );
  OAI211_X1 U8981 ( .C1(n7652), .C2(n10350), .A(n7651), .B(n7650), .ZN(
        P1_U3335) );
  INV_X1 U8982 ( .A(n7653), .ZN(n7654) );
  OAI22_X1 U8983 ( .A1(n7654), .A2(n10184), .B1(n10185), .B2(n9726), .ZN(n7659) );
  OAI22_X1 U8984 ( .A1(n10732), .A2(n5777), .B1(n9724), .B2(n10729), .ZN(n7655) );
  AOI21_X1 U8985 ( .B1(n10809), .B2(n9728), .A(n7655), .ZN(n7656) );
  OAI21_X1 U8986 ( .B1(n7657), .B2(n10156), .A(n7656), .ZN(n7658) );
  AOI211_X1 U8987 ( .C1(n10189), .C2(n7660), .A(n7659), .B(n7658), .ZN(n7661)
         );
  OAI21_X1 U8988 ( .B1(n10160), .B2(n7662), .A(n7661), .ZN(P1_U3289) );
  INV_X1 U8989 ( .A(n10769), .ZN(n7677) );
  NAND2_X1 U8990 ( .A1(n7663), .A2(n7673), .ZN(n7664) );
  XNOR2_X1 U8991 ( .A(n10769), .B(n8630), .ZN(n7881) );
  XNOR2_X1 U8992 ( .A(n7881), .B(n9143), .ZN(n7667) );
  AOI21_X1 U8993 ( .B1(n7666), .B2(n7667), .A(n9133), .ZN(n7669) );
  INV_X1 U8994 ( .A(n7667), .ZN(n7668) );
  NAND2_X1 U8995 ( .A1(n7669), .A2(n7883), .ZN(n7676) );
  INV_X1 U8996 ( .A(n7670), .ZN(n10771) );
  AOI21_X1 U8997 ( .B1(n9081), .B2(n9142), .A(n7671), .ZN(n7672) );
  OAI21_X1 U8998 ( .B1(n7673), .B2(n9094), .A(n7672), .ZN(n7674) );
  AOI21_X1 U8999 ( .B1(n10771), .B2(n9125), .A(n7674), .ZN(n7675) );
  OAI211_X1 U9000 ( .C1(n7677), .C2(n9114), .A(n7676), .B(n7675), .ZN(P2_U3171) );
  INV_X2 U9001 ( .A(n10732), .ZN(n10820) );
  NAND2_X1 U9002 ( .A1(n7678), .A2(n8344), .ZN(n7679) );
  XNOR2_X1 U9003 ( .A(n7679), .B(n8455), .ZN(n7680) );
  NAND2_X1 U9004 ( .A1(n7680), .A2(n10162), .ZN(n7682) );
  AOI22_X1 U9005 ( .A1(n10267), .A2(n9804), .B1(n10268), .B2(n9802), .ZN(n7681) );
  NAND2_X1 U9006 ( .A1(n7682), .A2(n7681), .ZN(n10757) );
  INV_X1 U9007 ( .A(n10757), .ZN(n7694) );
  OAI21_X1 U9008 ( .B1(n7684), .B2(n8455), .A(n7683), .ZN(n10759) );
  INV_X1 U9009 ( .A(n7685), .ZN(n7686) );
  OAI211_X1 U9010 ( .C1(n10756), .C2(n7687), .A(n7686), .B(n10782), .ZN(n10755) );
  INV_X1 U9011 ( .A(n10729), .ZN(n10807) );
  AOI22_X1 U9012 ( .A1(n10820), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7688), .B2(
        n10807), .ZN(n7691) );
  NAND2_X1 U9013 ( .A1(n10809), .A2(n7689), .ZN(n7690) );
  OAI211_X1 U9014 ( .C1(n10755), .C2(n10184), .A(n7691), .B(n7690), .ZN(n7692)
         );
  AOI21_X1 U9015 ( .B1(n10759), .B2(n10189), .A(n7692), .ZN(n7693) );
  OAI21_X1 U9016 ( .B1(n10820), .B2(n7694), .A(n7693), .ZN(P1_U3288) );
  INV_X1 U9017 ( .A(n7695), .ZN(n7697) );
  OAI222_X1 U9018 ( .A1(n7792), .A2(n7698), .B1(n9625), .B2(n7697), .C1(n7696), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  XNOR2_X1 U9019 ( .A(n8523), .B(n8452), .ZN(n7699) );
  NAND2_X1 U9020 ( .A1(n7699), .A2(n10162), .ZN(n7701) );
  AOI22_X1 U9021 ( .A1(n10268), .A2(n9805), .B1(n10267), .B2(n9807), .ZN(n7700) );
  NAND2_X1 U9022 ( .A1(n7701), .A2(n7700), .ZN(n10744) );
  AOI21_X1 U9023 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n10807), .A(n10744), .ZN(
        n7710) );
  OAI21_X1 U9024 ( .B1(n7703), .B2(n8342), .A(n7702), .ZN(n10746) );
  OAI211_X1 U9025 ( .C1(n7705), .C2(n10743), .A(n7704), .B(n10782), .ZN(n10742) );
  AOI22_X1 U9026 ( .A1(n10809), .A2(n7706), .B1(n10820), .B2(
        P1_REG2_REG_2__SCAN_IN), .ZN(n7707) );
  OAI21_X1 U9027 ( .B1(n10184), .B2(n10742), .A(n7707), .ZN(n7708) );
  AOI21_X1 U9028 ( .B1(n10189), .B2(n10746), .A(n7708), .ZN(n7709) );
  OAI21_X1 U9029 ( .B1(n10820), .B2(n7710), .A(n7709), .ZN(P1_U3291) );
  NAND2_X1 U9030 ( .A1(n8313), .A2(n8965), .ZN(n7715) );
  NAND2_X1 U9031 ( .A1(n7254), .A2(n9801), .ZN(n7714) );
  NAND2_X1 U9032 ( .A1(n7715), .A2(n7714), .ZN(n8306) );
  NAND2_X1 U9033 ( .A1(n8313), .A2(n8977), .ZN(n7717) );
  NAND2_X1 U9034 ( .A1(n9801), .A2(n8916), .ZN(n7716) );
  NAND2_X1 U9035 ( .A1(n7717), .A2(n7716), .ZN(n7718) );
  XNOR2_X1 U9036 ( .A(n7718), .B(n8963), .ZN(n8305) );
  NAND2_X1 U9037 ( .A1(n8308), .A2(n8306), .ZN(n7719) );
  NAND2_X1 U9038 ( .A1(n7720), .A2(n7719), .ZN(n7780) );
  NAND2_X1 U9039 ( .A1(n8374), .A2(n8965), .ZN(n7722) );
  NAND2_X1 U9040 ( .A1(n7254), .A2(n9800), .ZN(n7721) );
  NAND2_X1 U9041 ( .A1(n7722), .A2(n7721), .ZN(n7778) );
  NAND2_X1 U9042 ( .A1(n8374), .A2(n8977), .ZN(n7724) );
  NAND2_X1 U9043 ( .A1(n9800), .A2(n8965), .ZN(n7723) );
  NAND2_X1 U9044 ( .A1(n7724), .A2(n7723), .ZN(n7725) );
  XNOR2_X1 U9045 ( .A(n7725), .B(n8963), .ZN(n7779) );
  XOR2_X1 U9046 ( .A(n7778), .B(n7779), .Z(n7726) );
  XNOR2_X1 U9047 ( .A(n7727), .B(n7726), .ZN(n7732) );
  NOR2_X1 U9048 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7728), .ZN(n9899) );
  OAI22_X1 U9049 ( .A1(n9779), .A2(n7966), .B1(n9781), .B2(n7860), .ZN(n7729)
         );
  AOI211_X1 U9050 ( .C1(n9767), .C2(n9801), .A(n9899), .B(n7729), .ZN(n7731)
         );
  NAND2_X1 U9051 ( .A1(n4944), .A2(n8374), .ZN(n7730) );
  OAI211_X1 U9052 ( .C1(n7732), .C2(n9788), .A(n7731), .B(n7730), .ZN(P1_U3221) );
  NOR2_X1 U9053 ( .A1(n7749), .A2(n7733), .ZN(n7735) );
  NAND2_X1 U9054 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7938), .ZN(n7736) );
  OAI21_X1 U9055 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7938), .A(n7736), .ZN(
        n7737) );
  AOI21_X1 U9056 ( .B1(n7738), .B2(n7737), .A(n7922), .ZN(n7760) );
  MUX2_X1 U9057 ( .A(n8015), .B(n7739), .S(n4946), .Z(n7928) );
  XNOR2_X1 U9058 ( .A(n7928), .B(n7938), .ZN(n7745) );
  OR2_X1 U9059 ( .A1(n7741), .A2(n7740), .ZN(n7743) );
  NAND2_X1 U9060 ( .A1(n7743), .A2(n7742), .ZN(n7744) );
  NAND2_X1 U9061 ( .A1(n7745), .A2(n7744), .ZN(n7930) );
  OAI21_X1 U9062 ( .B1(n7745), .B2(n7744), .A(n7930), .ZN(n7758) );
  INV_X1 U9063 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7747) );
  INV_X1 U9064 ( .A(n7938), .ZN(n7929) );
  NAND2_X1 U9065 ( .A1(n10676), .A2(n7929), .ZN(n7746) );
  NAND2_X1 U9066 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7884) );
  OAI211_X1 U9067 ( .C1(n9263), .C2(n7747), .A(n7746), .B(n7884), .ZN(n7757)
         );
  NOR2_X1 U9068 ( .A1(n7749), .A2(n7748), .ZN(n7751) );
  NAND2_X1 U9069 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7938), .ZN(n7752) );
  OAI21_X1 U9070 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7938), .A(n7752), .ZN(
        n7753) );
  AOI21_X1 U9071 ( .B1(n7754), .B2(n7753), .A(n7937), .ZN(n7755) );
  NOR2_X1 U9072 ( .A1(n7755), .A2(n10682), .ZN(n7756) );
  AOI211_X1 U9073 ( .C1(n10690), .C2(n7758), .A(n7757), .B(n7756), .ZN(n7759)
         );
  OAI21_X1 U9074 ( .B1(n7760), .B2(n10713), .A(n7759), .ZN(P2_U3192) );
  INV_X1 U9075 ( .A(n7761), .ZN(n7769) );
  INV_X1 U9076 ( .A(n10809), .ZN(n10178) );
  NAND2_X1 U9077 ( .A1(n7762), .A2(n10814), .ZN(n7764) );
  AOI22_X1 U9078 ( .A1(n10820), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10807), .B2(
        n7274), .ZN(n7763) );
  OAI211_X1 U9079 ( .C1(n10178), .C2(n7765), .A(n7764), .B(n7763), .ZN(n7766)
         );
  AOI21_X1 U9080 ( .B1(n10189), .B2(n7767), .A(n7766), .ZN(n7768) );
  OAI21_X1 U9081 ( .B1(n10820), .B2(n7769), .A(n7768), .ZN(P1_U3290) );
  NAND3_X1 U9082 ( .A1(n7771), .A2(n5467), .A3(n8746), .ZN(n7772) );
  NAND2_X1 U9083 ( .A1(n7770), .A2(n7772), .ZN(n7877) );
  NOR2_X1 U9084 ( .A1(n7873), .A2(n9559), .ZN(n7776) );
  XNOR2_X1 U9085 ( .A(n7773), .B(n8668), .ZN(n7774) );
  OAI222_X1 U9086 ( .A1(n9473), .A2(n8704), .B1(n9471), .B2(n7775), .C1(n7774), 
        .C2(n9468), .ZN(n7874) );
  AOI211_X1 U9087 ( .C1(n9525), .C2(n7877), .A(n7776), .B(n7874), .ZN(n10762)
         );
  OR2_X1 U9088 ( .A1(n10762), .A2(n9570), .ZN(n7777) );
  OAI21_X1 U9089 ( .B1(n9561), .B2(n6333), .A(n7777), .ZN(P2_U3465) );
  NAND2_X1 U9090 ( .A1(n7807), .A2(n8977), .ZN(n7782) );
  NAND2_X1 U9091 ( .A1(n9799), .A2(n8965), .ZN(n7781) );
  NAND2_X1 U9092 ( .A1(n7782), .A2(n7781), .ZN(n7783) );
  XNOR2_X1 U9093 ( .A(n7783), .B(n8883), .ZN(n7954) );
  NOR2_X1 U9094 ( .A1(n7966), .A2(n8902), .ZN(n7784) );
  AOI21_X1 U9095 ( .B1(n7807), .B2(n8965), .A(n7784), .ZN(n7953) );
  XNOR2_X1 U9096 ( .A(n7954), .B(n7953), .ZN(n7951) );
  XOR2_X1 U9097 ( .A(n7952), .B(n7951), .Z(n7789) );
  OAI22_X1 U9098 ( .A1(n9783), .A2(n8373), .B1(n9781), .B2(n7801), .ZN(n7785)
         );
  AOI211_X1 U9099 ( .C1(n9768), .C2(n9798), .A(n7786), .B(n7785), .ZN(n7788)
         );
  NAND2_X1 U9100 ( .A1(n4944), .A2(n7807), .ZN(n7787) );
  OAI211_X1 U9101 ( .C1(n7789), .C2(n9788), .A(n7788), .B(n7787), .ZN(P1_U3231) );
  INV_X1 U9102 ( .A(n7790), .ZN(n7842) );
  OAI222_X1 U9103 ( .A1(n9625), .A2(n7842), .B1(n7792), .B2(n7791), .C1(n8712), 
        .C2(P2_U3151), .ZN(P2_U3274) );
  INV_X1 U9104 ( .A(n9525), .ZN(n9563) );
  INV_X1 U9105 ( .A(n7795), .ZN(n8740) );
  OAI21_X1 U9106 ( .B1(n7794), .B2(n8740), .A(n7793), .ZN(n7817) );
  XNOR2_X1 U9107 ( .A(n7796), .B(n7795), .ZN(n7797) );
  INV_X1 U9108 ( .A(n9473), .ZN(n9552) );
  AOI222_X1 U9109 ( .A1(n9547), .A2(n7797), .B1(n9144), .B2(n9552), .C1(n9146), 
        .C2(n9553), .ZN(n7812) );
  OAI21_X1 U9110 ( .B1(n9563), .B2(n7817), .A(n7812), .ZN(n7846) );
  INV_X1 U9111 ( .A(n7846), .ZN(n7799) );
  INV_X1 U9112 ( .A(n9529), .ZN(n7997) );
  AOI22_X1 U9113 ( .A1(n7997), .A2(n8705), .B1(n9570), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n7798) );
  OAI21_X1 U9114 ( .B1(n7799), .B2(n9570), .A(n7798), .ZN(P2_U3466) );
  INV_X1 U9115 ( .A(n7800), .ZN(n7811) );
  INV_X1 U9116 ( .A(n7801), .ZN(n7802) );
  AOI22_X1 U9117 ( .A1(n10820), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7802), .B2(
        n10807), .ZN(n7803) );
  OAI21_X1 U9118 ( .B1(n10156), .B2(n8373), .A(n7803), .ZN(n7806) );
  NOR2_X1 U9119 ( .A1(n7804), .A2(n10184), .ZN(n7805) );
  AOI211_X1 U9120 ( .C1(n10809), .C2(n7807), .A(n7806), .B(n7805), .ZN(n7810)
         );
  NAND2_X1 U9121 ( .A1(n7808), .A2(n10189), .ZN(n7809) );
  OAI211_X1 U9122 ( .C1(n7811), .C2(n10160), .A(n7810), .B(n7809), .ZN(
        P1_U3284) );
  MUX2_X1 U9123 ( .A(n7813), .B(n7812), .S(n10846), .Z(n7816) );
  AOI22_X1 U9124 ( .A1(n10768), .A2(n8705), .B1(n10770), .B2(n7814), .ZN(n7815) );
  OAI211_X1 U9125 ( .C1(n9479), .C2(n7817), .A(n7816), .B(n7815), .ZN(P2_U3226) );
  AOI21_X1 U9126 ( .B1(n7823), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7818), .ZN(
        n7820) );
  XNOR2_X1 U9127 ( .A(n8074), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n7819) );
  NOR2_X1 U9128 ( .A1(n7819), .A2(n7820), .ZN(n8071) );
  AOI211_X1 U9129 ( .C1(n7820), .C2(n7819), .A(n8071), .B(n9895), .ZN(n7830)
         );
  NOR2_X1 U9130 ( .A1(n8074), .A2(n8042), .ZN(n7821) );
  AOI21_X1 U9131 ( .B1(n8074), .B2(n8042), .A(n7821), .ZN(n7825) );
  AOI21_X1 U9132 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n7823), .A(n7822), .ZN(
        n7824) );
  NOR2_X1 U9133 ( .A1(n7825), .A2(n7824), .ZN(n8073) );
  AOI211_X1 U9134 ( .C1(n7825), .C2(n7824), .A(n8073), .B(n9953), .ZN(n7829)
         );
  INV_X1 U9135 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7827) );
  NAND2_X1 U9136 ( .A1(n9930), .A2(n8074), .ZN(n7826) );
  NAND2_X1 U9137 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9644) );
  OAI211_X1 U9138 ( .C1(n7827), .C2(n9920), .A(n7826), .B(n9644), .ZN(n7828)
         );
  OR3_X1 U9139 ( .A1(n7830), .A2(n7829), .A3(n7828), .ZN(P1_U3257) );
  XNOR2_X1 U9140 ( .A(n7831), .B(n8463), .ZN(n10829) );
  INV_X1 U9141 ( .A(n10829), .ZN(n7840) );
  INV_X1 U9142 ( .A(n10189), .ZN(n10098) );
  NAND3_X1 U9143 ( .A1(n5237), .A2(n10787), .A3(n8386), .ZN(n7832) );
  NAND3_X1 U9144 ( .A1(n7893), .A2(n10162), .A3(n7832), .ZN(n7834) );
  AOI22_X1 U9145 ( .A1(n10267), .A2(n9797), .B1(n10268), .B2(n9795), .ZN(n7833) );
  NAND2_X1 U9146 ( .A1(n7834), .A2(n7833), .ZN(n10827) );
  OAI211_X1 U9147 ( .C1(n10781), .C2(n10825), .A(n10782), .B(n7899), .ZN(
        n10823) );
  OAI22_X1 U9148 ( .A1(n10732), .A2(n7835), .B1(n8194), .B2(n10729), .ZN(n7836) );
  AOI21_X1 U9149 ( .B1(n8188), .B2(n10809), .A(n7836), .ZN(n7837) );
  OAI21_X1 U9150 ( .B1(n10823), .B2(n10184), .A(n7837), .ZN(n7838) );
  AOI21_X1 U9151 ( .B1(n10732), .B2(n10827), .A(n7838), .ZN(n7839) );
  OAI21_X1 U9152 ( .B1(n7840), .B2(n10098), .A(n7839), .ZN(P1_U3281) );
  OAI222_X1 U9153 ( .A1(P1_U3086), .A2(n8519), .B1(n10354), .B2(n7842), .C1(
        n7841), .C2(n10350), .ZN(P1_U3334) );
  INV_X1 U9154 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7843) );
  OAI22_X1 U9155 ( .A1(n9606), .A2(n7844), .B1(n10852), .B2(n7843), .ZN(n7845)
         );
  AOI21_X1 U9156 ( .B1(n7846), .B2(n10852), .A(n7845), .ZN(n7847) );
  INV_X1 U9157 ( .A(n7847), .ZN(P2_U3411) );
  OAI22_X1 U9158 ( .A1(n10185), .A2(n7864), .B1(n10729), .B2(n7848), .ZN(n7850) );
  NOR2_X1 U9159 ( .A1(n10156), .A2(n9726), .ZN(n7849) );
  AOI211_X1 U9160 ( .C1(n10809), .C2(n7851), .A(n7850), .B(n7849), .ZN(n7852)
         );
  OAI21_X1 U9161 ( .B1(n10184), .B2(n7853), .A(n7852), .ZN(n7854) );
  AOI21_X1 U9162 ( .B1(n10189), .B2(n7855), .A(n7854), .ZN(n7859) );
  MUX2_X1 U9163 ( .A(n7857), .B(n7856), .S(n10820), .Z(n7858) );
  NAND2_X1 U9164 ( .A1(n7859), .A2(n7858), .ZN(P1_U3287) );
  OAI22_X1 U9165 ( .A1(n10732), .A2(n7861), .B1(n7860), .B2(n10729), .ZN(n7862) );
  AOI21_X1 U9166 ( .B1(n10153), .B2(n9799), .A(n7862), .ZN(n7863) );
  OAI21_X1 U9167 ( .B1(n7864), .B2(n10156), .A(n7863), .ZN(n7865) );
  AOI21_X1 U9168 ( .B1(n10809), .B2(n8374), .A(n7865), .ZN(n7866) );
  OAI21_X1 U9169 ( .B1(n10184), .B2(n7867), .A(n7866), .ZN(n7868) );
  AOI21_X1 U9170 ( .B1(n7869), .B2(n10189), .A(n7868), .ZN(n7870) );
  OAI21_X1 U9171 ( .B1(n10820), .B2(n7871), .A(n7870), .ZN(P1_U3285) );
  OAI22_X1 U9172 ( .A1(n9360), .A2(n7873), .B1(n7872), .B2(n10838), .ZN(n7876)
         );
  MUX2_X1 U9173 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7874), .S(n10846), .Z(n7875)
         );
  AOI211_X1 U9174 ( .C1(n9377), .C2(n7877), .A(n7876), .B(n7875), .ZN(n7878)
         );
  INV_X1 U9175 ( .A(n7878), .ZN(P2_U3227) );
  INV_X1 U9176 ( .A(n7879), .ZN(n8989) );
  AOI22_X1 U9177 ( .A1(n8867), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n9623), .ZN(n7880) );
  OAI21_X1 U9178 ( .B1(n8989), .B2(n9625), .A(n7880), .ZN(P2_U3273) );
  NAND2_X1 U9179 ( .A1(n7881), .A2(n9143), .ZN(n7882) );
  XNOR2_X1 U9180 ( .A(n8144), .B(n8635), .ZN(n7973) );
  XNOR2_X1 U9181 ( .A(n7972), .B(n9142), .ZN(n7889) );
  INV_X1 U9182 ( .A(n9125), .ZN(n9006) );
  OAI21_X1 U9183 ( .B1(n9094), .B2(n8013), .A(n7884), .ZN(n7885) );
  AOI21_X1 U9184 ( .B1(n9081), .B2(n9141), .A(n7885), .ZN(n7886) );
  OAI21_X1 U9185 ( .B1(n9006), .B2(n8014), .A(n7886), .ZN(n7887) );
  AOI21_X1 U9186 ( .B1(n8144), .B2(n9131), .A(n7887), .ZN(n7888) );
  OAI21_X1 U9187 ( .B1(n7889), .B2(n9133), .A(n7888), .ZN(P2_U3157) );
  INV_X1 U9188 ( .A(n7909), .ZN(n7892) );
  NAND2_X1 U9189 ( .A1(n9623), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7891) );
  NAND2_X1 U9190 ( .A1(n7890), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8870) );
  OAI211_X1 U9191 ( .C1(n7892), .C2(n9625), .A(n7891), .B(n8870), .ZN(P2_U3272) );
  INV_X1 U9192 ( .A(n8464), .ZN(n7895) );
  NAND2_X1 U9193 ( .A1(n7893), .A2(n8391), .ZN(n7894) );
  NAND2_X1 U9194 ( .A1(n7895), .A2(n7894), .ZN(n7897) );
  AND2_X1 U9195 ( .A1(n7897), .A2(n7896), .ZN(n7915) );
  XNOR2_X1 U9196 ( .A(n7898), .B(n8464), .ZN(n7917) );
  NAND2_X1 U9197 ( .A1(n7917), .A2(n10189), .ZN(n7908) );
  AOI21_X1 U9198 ( .B1(n7899), .B2(n8213), .A(n10174), .ZN(n7900) );
  NAND2_X1 U9199 ( .A1(n7900), .A2(n8043), .ZN(n7913) );
  INV_X1 U9200 ( .A(n7913), .ZN(n7906) );
  NAND2_X1 U9201 ( .A1(n8213), .A2(n10809), .ZN(n7904) );
  INV_X1 U9202 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7901) );
  OAI22_X1 U9203 ( .A1(n10732), .A2(n7901), .B1(n8222), .B2(n10729), .ZN(n7902) );
  AOI21_X1 U9204 ( .B1(n10153), .B2(n9794), .A(n7902), .ZN(n7903) );
  OAI211_X1 U9205 ( .C1(n10795), .C2(n10156), .A(n7904), .B(n7903), .ZN(n7905)
         );
  AOI21_X1 U9206 ( .B1(n7906), .B2(n10814), .A(n7905), .ZN(n7907) );
  OAI211_X1 U9207 ( .C1(n7915), .C2(n10160), .A(n7908), .B(n7907), .ZN(
        P1_U3280) );
  NAND2_X1 U9208 ( .A1(n7909), .A2(n10343), .ZN(n7911) );
  OR2_X1 U9209 ( .A1(n7910), .A2(P1_U3086), .ZN(n8579) );
  OAI211_X1 U9210 ( .C1(n7912), .C2(n10350), .A(n7911), .B(n8579), .ZN(
        P1_U3332) );
  AOI22_X1 U9211 ( .A1(n10267), .A2(n9796), .B1(n10268), .B2(n9794), .ZN(n7914) );
  OAI211_X1 U9212 ( .C1(n7915), .C2(n10791), .A(n7914), .B(n7913), .ZN(n7916)
         );
  AOI21_X1 U9213 ( .B1(n7917), .B2(n5053), .A(n7916), .ZN(n7921) );
  AOI22_X1 U9214 ( .A1(n8213), .A2(n6205), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n6207), .ZN(n7918) );
  OAI21_X1 U9215 ( .B1(n7921), .B2(n6207), .A(n7918), .ZN(P1_U3492) );
  AOI22_X1 U9216 ( .A1(n8213), .A2(n7919), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n10830), .ZN(n7920) );
  OAI21_X1 U9217 ( .B1(n7921), .B2(n10830), .A(n7920), .ZN(P1_U3535) );
  XNOR2_X1 U9218 ( .A(n10675), .B(n7923), .ZN(n10685) );
  AOI22_X1 U9219 ( .A1(n7941), .A2(P2_REG1_REG_12__SCAN_IN), .B1(n6419), .B2(
        n8154), .ZN(n7924) );
  AOI21_X1 U9220 ( .B1(n7925), .B2(n7924), .A(n8146), .ZN(n7950) );
  MUX2_X1 U9221 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n4946), .Z(n8148) );
  XNOR2_X1 U9222 ( .A(n8148), .B(n7941), .ZN(n7934) );
  MUX2_X1 U9223 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n4947), .Z(n7927) );
  INV_X1 U9224 ( .A(n7927), .ZN(n7926) );
  NAND2_X1 U9225 ( .A1(n10675), .A2(n7926), .ZN(n7932) );
  XNOR2_X1 U9226 ( .A(n7927), .B(n10675), .ZN(n10679) );
  NAND2_X1 U9227 ( .A1(n7929), .A2(n7928), .ZN(n7931) );
  NAND2_X1 U9228 ( .A1(n7931), .A2(n7930), .ZN(n10678) );
  NAND2_X1 U9229 ( .A1(n10679), .A2(n10678), .ZN(n10677) );
  NAND2_X1 U9230 ( .A1(n7932), .A2(n10677), .ZN(n7933) );
  NAND2_X1 U9231 ( .A1(n7934), .A2(n7933), .ZN(n8149) );
  OAI21_X1 U9232 ( .B1(n7934), .B2(n7933), .A(n8149), .ZN(n7948) );
  INV_X1 U9233 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7936) );
  NAND2_X1 U9234 ( .A1(n10676), .A2(n7941), .ZN(n7935) );
  OR2_X1 U9235 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10545), .ZN(n8028) );
  OAI211_X1 U9236 ( .C1(n7936), .C2(n9263), .A(n7935), .B(n8028), .ZN(n7947)
         );
  NOR2_X1 U9237 ( .A1(n10675), .A2(n7939), .ZN(n7940) );
  XNOR2_X1 U9238 ( .A(n10675), .B(n7939), .ZN(n10681) );
  NOR2_X1 U9239 ( .A1(n6401), .A2(n10681), .ZN(n10680) );
  MUX2_X1 U9240 ( .A(n8134), .B(P2_REG2_REG_12__SCAN_IN), .S(n7941), .Z(n7942)
         );
  INV_X1 U9241 ( .A(n7942), .ZN(n7943) );
  NOR2_X1 U9242 ( .A1(n7944), .A2(n7943), .ZN(n8153) );
  AOI21_X1 U9243 ( .B1(n7944), .B2(n7943), .A(n8153), .ZN(n7945) );
  NOR2_X1 U9244 ( .A1(n7945), .A2(n10682), .ZN(n7946) );
  AOI211_X1 U9245 ( .C1(n10690), .C2(n7948), .A(n7947), .B(n7946), .ZN(n7949)
         );
  OAI21_X1 U9246 ( .B1(n7950), .B2(n10713), .A(n7949), .ZN(P2_U3194) );
  INV_X1 U9247 ( .A(n7961), .ZN(n7959) );
  NAND2_X1 U9248 ( .A1(n7969), .A2(n8977), .ZN(n7956) );
  NAND2_X1 U9249 ( .A1(n9798), .A2(n8965), .ZN(n7955) );
  NAND2_X1 U9250 ( .A1(n7956), .A2(n7955), .ZN(n7957) );
  XNOR2_X1 U9251 ( .A(n7957), .B(n8883), .ZN(n7960) );
  NAND2_X1 U9252 ( .A1(n7959), .A2(n7958), .ZN(n8083) );
  NAND2_X1 U9253 ( .A1(n7961), .A2(n7960), .ZN(n8084) );
  NAND2_X1 U9254 ( .A1(n8083), .A2(n8084), .ZN(n7963) );
  NOR2_X1 U9255 ( .A1(n10797), .A2(n8902), .ZN(n7962) );
  AOI21_X1 U9256 ( .B1(n7969), .B2(n8965), .A(n7962), .ZN(n8082) );
  XNOR2_X1 U9257 ( .A(n7963), .B(n8082), .ZN(n7971) );
  OAI21_X1 U9258 ( .B1(n9779), .B2(n8195), .A(n7964), .ZN(n7968) );
  OAI22_X1 U9259 ( .A1(n9783), .A2(n7966), .B1(n9781), .B2(n7965), .ZN(n7967)
         );
  AOI211_X1 U9260 ( .C1(n7969), .C2(n4944), .A(n7968), .B(n7967), .ZN(n7970)
         );
  OAI21_X1 U9261 ( .B1(n7971), .B2(n9788), .A(n7970), .ZN(P1_U3217) );
  NAND2_X1 U9262 ( .A1(n7974), .A2(n7973), .ZN(n7975) );
  XNOR2_X1 U9263 ( .A(n8060), .B(n8635), .ZN(n8022) );
  XNOR2_X1 U9264 ( .A(n8022), .B(n9141), .ZN(n8019) );
  XOR2_X1 U9265 ( .A(n8020), .B(n8019), .Z(n7981) );
  INV_X1 U9266 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10693) );
  OAI22_X1 U9267 ( .A1(n9094), .A2(n8057), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10693), .ZN(n7977) );
  AOI21_X1 U9268 ( .B1(n9081), .B2(n9140), .A(n7977), .ZN(n7978) );
  OAI21_X1 U9269 ( .B1(n9006), .B2(n8058), .A(n7978), .ZN(n7979) );
  AOI21_X1 U9270 ( .B1(n8060), .B2(n9131), .A(n7979), .ZN(n7980) );
  OAI21_X1 U9271 ( .B1(n7981), .B2(n9133), .A(n7980), .ZN(P2_U3176) );
  XNOR2_X1 U9272 ( .A(n7982), .B(n8669), .ZN(n8007) );
  NOR2_X1 U9273 ( .A1(n8007), .A2(n9563), .ZN(n7985) );
  XOR2_X1 U9274 ( .A(n8669), .B(n7983), .Z(n7984) );
  OAI222_X1 U9275 ( .A1(n9473), .A2(n8013), .B1(n9471), .B2(n8704), .C1(n9468), 
        .C2(n7984), .ZN(n8000) );
  AOI211_X1 U9276 ( .C1(n9568), .C2(n8004), .A(n7985), .B(n8000), .ZN(n10764)
         );
  OR2_X1 U9277 ( .A1(n10764), .A2(n9570), .ZN(n7986) );
  OAI21_X1 U9278 ( .B1(n9561), .B2(n7527), .A(n7986), .ZN(P2_U3467) );
  INV_X1 U9279 ( .A(n8671), .ZN(n7988) );
  OAI21_X1 U9280 ( .B1(n7989), .B2(n7988), .A(n7987), .ZN(n10766) );
  XNOR2_X1 U9281 ( .A(n7990), .B(n8671), .ZN(n7991) );
  AOI222_X1 U9282 ( .A1(n9547), .A2(n7991), .B1(n9142), .B2(n9552), .C1(n9144), 
        .C2(n9553), .ZN(n10765) );
  OAI21_X1 U9283 ( .B1(n9563), .B2(n10766), .A(n10765), .ZN(n7992) );
  INV_X1 U9284 ( .A(n7992), .ZN(n7999) );
  INV_X1 U9285 ( .A(n9606), .ZN(n7995) );
  INV_X1 U9286 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7993) );
  NOR2_X1 U9287 ( .A1(n10852), .A2(n7993), .ZN(n7994) );
  AOI21_X1 U9288 ( .B1(n7995), .B2(n10769), .A(n7994), .ZN(n7996) );
  OAI21_X1 U9289 ( .B1(n7999), .B2(n10850), .A(n7996), .ZN(P2_U3417) );
  AOI22_X1 U9290 ( .A1(n10769), .A2(n7997), .B1(n9570), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n7998) );
  OAI21_X1 U9291 ( .B1(n7999), .B2(n9570), .A(n7998), .ZN(P2_U3468) );
  INV_X1 U9292 ( .A(n8000), .ZN(n8001) );
  MUX2_X1 U9293 ( .A(n8002), .B(n8001), .S(n10846), .Z(n8006) );
  AOI22_X1 U9294 ( .A1(n10768), .A2(n8004), .B1(n10770), .B2(n8003), .ZN(n8005) );
  OAI211_X1 U9295 ( .C1(n8007), .C2(n9479), .A(n8006), .B(n8005), .ZN(P2_U3225) );
  NAND2_X1 U9296 ( .A1(n8009), .A2(n8008), .ZN(n8673) );
  XNOR2_X1 U9297 ( .A(n8010), .B(n8673), .ZN(n8139) );
  XNOR2_X1 U9298 ( .A(n8011), .B(n8673), .ZN(n8012) );
  OAI222_X1 U9299 ( .A1(n9471), .A2(n8013), .B1(n9473), .B2(n8021), .C1(n8012), 
        .C2(n9468), .ZN(n8142) );
  NAND2_X1 U9300 ( .A1(n8142), .A2(n10846), .ZN(n8018) );
  OAI22_X1 U9301 ( .A1(n10846), .A2(n8015), .B1(n8014), .B2(n10838), .ZN(n8016) );
  AOI21_X1 U9302 ( .B1(n8144), .B2(n10768), .A(n8016), .ZN(n8017) );
  OAI211_X1 U9303 ( .C1(n8139), .C2(n9479), .A(n8018), .B(n8017), .ZN(P2_U3223) );
  INV_X1 U9304 ( .A(n8768), .ZN(n8256) );
  NAND2_X1 U9305 ( .A1(n8022), .A2(n8021), .ZN(n8023) );
  XNOR2_X1 U9306 ( .A(n8768), .B(n8630), .ZN(n8101) );
  XNOR2_X1 U9307 ( .A(n8101), .B(n9140), .ZN(n8025) );
  AOI21_X1 U9308 ( .B1(n8024), .B2(n8025), .A(n9133), .ZN(n8027) );
  INV_X1 U9309 ( .A(n8025), .ZN(n8026) );
  NAND2_X1 U9310 ( .A1(n8027), .A2(n8103), .ZN(n8032) );
  OAI21_X1 U9311 ( .B1(n9129), .B2(n8239), .A(n8028), .ZN(n8030) );
  NOR2_X1 U9312 ( .A1(n9006), .A2(n8133), .ZN(n8029) );
  AOI211_X1 U9313 ( .C1(n9126), .C2(n9141), .A(n8030), .B(n8029), .ZN(n8031)
         );
  OAI211_X1 U9314 ( .C1(n8256), .C2(n9114), .A(n8032), .B(n8031), .ZN(P2_U3164) );
  INV_X1 U9315 ( .A(n8033), .ZN(n8069) );
  AOI22_X1 U9316 ( .A1(n8034), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n9623), .ZN(n8035) );
  OAI21_X1 U9317 ( .B1(n8069), .B2(n9625), .A(n8035), .ZN(P2_U3271) );
  NAND2_X1 U9318 ( .A1(n8036), .A2(n8466), .ZN(n8037) );
  NAND3_X1 U9319 ( .A1(n8119), .A2(n10162), .A3(n8037), .ZN(n8039) );
  AOI22_X1 U9320 ( .A1(n10267), .A2(n9795), .B1(n10268), .B2(n10165), .ZN(
        n8038) );
  NAND2_X1 U9321 ( .A1(n8039), .A2(n8038), .ZN(n8203) );
  INV_X1 U9322 ( .A(n8203), .ZN(n8050) );
  NOR2_X1 U9323 ( .A1(n8040), .A2(n8466), .ZN(n8200) );
  INV_X1 U9324 ( .A(n8200), .ZN(n8041) );
  NAND3_X1 U9325 ( .A1(n8041), .A2(n10189), .A3(n8204), .ZN(n8049) );
  OAI22_X1 U9326 ( .A1(n10732), .A2(n8042), .B1(n9645), .B2(n10729), .ZN(n8047) );
  INV_X1 U9327 ( .A(n8043), .ZN(n8045) );
  INV_X1 U9328 ( .A(n8044), .ZN(n8115) );
  OAI211_X1 U9329 ( .C1(n8877), .C2(n8045), .A(n8115), .B(n10782), .ZN(n8201)
         );
  NOR2_X1 U9330 ( .A1(n8201), .A2(n10184), .ZN(n8046) );
  AOI211_X1 U9331 ( .C1(n10809), .C2(n9649), .A(n8047), .B(n8046), .ZN(n8048)
         );
  OAI211_X1 U9332 ( .C1(n10820), .C2(n8050), .A(n8049), .B(n8048), .ZN(
        P1_U3279) );
  INV_X1 U9333 ( .A(n8051), .ZN(n8111) );
  AOI22_X1 U9334 ( .A1(n8052), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n9623), .ZN(n8053) );
  OAI21_X1 U9335 ( .B1(n8111), .B2(n9625), .A(n8053), .ZN(P2_U3270) );
  XOR2_X1 U9336 ( .A(n8675), .B(n8054), .Z(n8064) );
  XNOR2_X1 U9337 ( .A(n8055), .B(n8675), .ZN(n8056) );
  OAI222_X1 U9338 ( .A1(n9473), .A2(n9470), .B1(n9471), .B2(n8057), .C1(n9468), 
        .C2(n8056), .ZN(n8066) );
  NAND2_X1 U9339 ( .A1(n8066), .A2(n10846), .ZN(n8062) );
  OAI22_X1 U9340 ( .A1(n10846), .A2(n6401), .B1(n8058), .B2(n10838), .ZN(n8059) );
  AOI21_X1 U9341 ( .B1(n8060), .B2(n10768), .A(n8059), .ZN(n8061) );
  OAI211_X1 U9342 ( .C1(n8064), .C2(n9479), .A(n8062), .B(n8061), .ZN(P2_U3222) );
  OAI22_X1 U9343 ( .A1(n8064), .A2(n9563), .B1(n8063), .B2(n9559), .ZN(n8065)
         );
  NOR2_X1 U9344 ( .A1(n8066), .A2(n8065), .ZN(n10777) );
  NAND2_X1 U9345 ( .A1(n9570), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8067) );
  OAI21_X1 U9346 ( .B1(n10777), .B2(n9570), .A(n8067), .ZN(P2_U3470) );
  OAI222_X1 U9347 ( .A1(P1_U3086), .A2(n8070), .B1(n10354), .B2(n8069), .C1(
        n8068), .C2(n10350), .ZN(P1_U3331) );
  AOI21_X1 U9348 ( .B1(n8074), .B2(P1_REG1_REG_14__SCAN_IN), .A(n8071), .ZN(
        n8166) );
  XNOR2_X1 U9349 ( .A(n8166), .B(n8173), .ZN(n8072) );
  NOR2_X1 U9350 ( .A1(n10296), .A2(n8072), .ZN(n8167) );
  AOI211_X1 U9351 ( .C1(n8072), .C2(n10296), .A(n8167), .B(n9895), .ZN(n8081)
         );
  AOI21_X1 U9352 ( .B1(n8074), .B2(P1_REG2_REG_14__SCAN_IN), .A(n8073), .ZN(
        n8174) );
  XNOR2_X1 U9353 ( .A(n8174), .B(n8173), .ZN(n8075) );
  NOR2_X1 U9354 ( .A1(n8116), .A2(n8075), .ZN(n8175) );
  AOI211_X1 U9355 ( .C1(n8075), .C2(n8116), .A(n8175), .B(n9953), .ZN(n8080)
         );
  INV_X1 U9356 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n8078) );
  NAND2_X1 U9357 ( .A1(n9930), .A2(n8076), .ZN(n8077) );
  NAND2_X1 U9358 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9778) );
  OAI211_X1 U9359 ( .C1(n8078), .C2(n9920), .A(n8077), .B(n9778), .ZN(n8079)
         );
  OR3_X1 U9360 ( .A1(n8081), .A2(n8080), .A3(n8079), .ZN(P1_U3258) );
  INV_X1 U9361 ( .A(n4944), .ZN(n9737) );
  NAND2_X1 U9362 ( .A1(n8083), .A2(n8082), .ZN(n8085) );
  NAND2_X1 U9363 ( .A1(n10810), .A2(n8977), .ZN(n8087) );
  NAND2_X1 U9364 ( .A1(n9797), .A2(n8965), .ZN(n8086) );
  NAND2_X1 U9365 ( .A1(n8087), .A2(n8086), .ZN(n8088) );
  XNOR2_X1 U9366 ( .A(n8088), .B(n8963), .ZN(n8092) );
  NAND2_X1 U9367 ( .A1(n10810), .A2(n8965), .ZN(n8090) );
  NAND2_X1 U9368 ( .A1(n7254), .A2(n9797), .ZN(n8089) );
  NAND2_X1 U9369 ( .A1(n8090), .A2(n8089), .ZN(n8091) );
  NOR2_X1 U9370 ( .A1(n8092), .A2(n8091), .ZN(n8094) );
  INV_X1 U9371 ( .A(n9788), .ZN(n9764) );
  OAI21_X1 U9372 ( .B1(n8094), .B2(n8190), .A(n8093), .ZN(n8095) );
  OAI211_X1 U9373 ( .C1(n5403), .C2(n8190), .A(n9764), .B(n8095), .ZN(n8100)
         );
  INV_X1 U9374 ( .A(n8096), .ZN(n8098) );
  OAI22_X1 U9375 ( .A1(n9783), .A2(n10797), .B1(n9781), .B2(n10806), .ZN(n8097) );
  AOI211_X1 U9376 ( .C1(n9768), .C2(n9796), .A(n8098), .B(n8097), .ZN(n8099)
         );
  OAI211_X1 U9377 ( .C1(n10785), .C2(n9737), .A(n8100), .B(n8099), .ZN(
        P1_U3236) );
  NAND2_X1 U9378 ( .A1(n8101), .A2(n9140), .ZN(n8102) );
  XNOR2_X1 U9379 ( .A(n9567), .B(n8635), .ZN(n8242) );
  XNOR2_X1 U9380 ( .A(n8242), .B(n9554), .ZN(n8104) );
  XNOR2_X1 U9381 ( .A(n8241), .B(n8104), .ZN(n8109) );
  NAND2_X1 U9382 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8156) );
  OAI21_X1 U9383 ( .B1(n9129), .B2(n9472), .A(n8156), .ZN(n8105) );
  AOI21_X1 U9384 ( .B1(n9126), .B2(n9140), .A(n8105), .ZN(n8106) );
  OAI21_X1 U9385 ( .B1(n9474), .B2(n9006), .A(n8106), .ZN(n8107) );
  AOI21_X1 U9386 ( .B1(n9567), .B2(n9131), .A(n8107), .ZN(n8108) );
  OAI21_X1 U9387 ( .B1(n8109), .B2(n9133), .A(n8108), .ZN(P2_U3174) );
  OAI222_X1 U9388 ( .A1(P1_U3086), .A2(n8112), .B1(n10354), .B2(n8111), .C1(
        n8110), .C2(n10350), .ZN(P1_U3330) );
  OAI21_X1 U9389 ( .B1(n8114), .B2(n8467), .A(n8113), .ZN(n10292) );
  AOI211_X1 U9390 ( .C1(n9786), .C2(n8115), .A(n10174), .B(n10171), .ZN(n10294) );
  NOR2_X1 U9391 ( .A1(n10341), .A2(n10178), .ZN(n8118) );
  OAI22_X1 U9392 ( .A1(n10732), .A2(n8116), .B1(n9780), .B2(n10729), .ZN(n8117) );
  AOI211_X1 U9393 ( .C1(n10294), .C2(n10814), .A(n8118), .B(n8117), .ZN(n8125)
         );
  NAND3_X1 U9394 ( .A1(n8119), .A2(n8397), .A3(n8467), .ZN(n8120) );
  NAND3_X1 U9395 ( .A1(n8121), .A2(n10162), .A3(n8120), .ZN(n8123) );
  AOI22_X1 U9396 ( .A1(n10267), .A2(n9794), .B1(n10268), .B2(n9793), .ZN(n8122) );
  NAND2_X1 U9397 ( .A1(n8123), .A2(n8122), .ZN(n10293) );
  NAND2_X1 U9398 ( .A1(n10293), .A2(n10732), .ZN(n8124) );
  OAI211_X1 U9399 ( .C1(n10292), .C2(n10098), .A(n8125), .B(n8124), .ZN(
        P1_U3278) );
  INV_X1 U9400 ( .A(n8126), .ZN(n8128) );
  OAI211_X1 U9401 ( .C1(n8128), .C2(n5460), .A(n8127), .B(n9547), .ZN(n8130)
         );
  AOI22_X1 U9402 ( .A1(n9554), .A2(n9552), .B1(n9553), .B2(n9141), .ZN(n8129)
         );
  NAND2_X1 U9403 ( .A1(n8130), .A2(n8129), .ZN(n8257) );
  INV_X1 U9404 ( .A(n8257), .ZN(n8138) );
  OAI21_X1 U9405 ( .B1(n8132), .B2(n8767), .A(n8131), .ZN(n8259) );
  NOR2_X1 U9406 ( .A1(n8256), .A2(n9360), .ZN(n8136) );
  OAI22_X1 U9407 ( .A1(n10846), .A2(n8134), .B1(n8133), .B2(n10838), .ZN(n8135) );
  AOI211_X1 U9408 ( .C1(n8259), .C2(n9377), .A(n8136), .B(n8135), .ZN(n8137)
         );
  OAI21_X1 U9409 ( .B1(n8138), .B2(n4949), .A(n8137), .ZN(P2_U3221) );
  AOI21_X1 U9410 ( .B1(n8141), .B2(n8140), .A(n8139), .ZN(n8143) );
  AOI211_X1 U9411 ( .C1(n9568), .C2(n8144), .A(n8143), .B(n8142), .ZN(n10775)
         );
  OR2_X1 U9412 ( .A1(n10775), .A2(n9570), .ZN(n8145) );
  OAI21_X1 U9413 ( .B1(n9561), .B2(n7739), .A(n8145), .ZN(P2_U3469) );
  AOI21_X1 U9414 ( .B1(n6431), .B2(n8147), .A(n9153), .ZN(n8165) );
  MUX2_X1 U9415 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n4947), .Z(n9157) );
  XNOR2_X1 U9416 ( .A(n9157), .B(n9167), .ZN(n8152) );
  OR2_X1 U9417 ( .A1(n8148), .A2(n8154), .ZN(n8150) );
  NAND2_X1 U9418 ( .A1(n8150), .A2(n8149), .ZN(n8151) );
  NAND2_X1 U9419 ( .A1(n8152), .A2(n8151), .ZN(n9159) );
  OAI21_X1 U9420 ( .B1(n8152), .B2(n8151), .A(n9159), .ZN(n8163) );
  INV_X1 U9421 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8161) );
  AOI21_X1 U9422 ( .B1(n8155), .B2(n6430), .A(n9168), .ZN(n8157) );
  OAI21_X1 U9423 ( .B1(n10682), .B2(n8157), .A(n8156), .ZN(n8158) );
  INV_X1 U9424 ( .A(n8158), .ZN(n8160) );
  NAND2_X1 U9425 ( .A1(n10676), .A2(n9167), .ZN(n8159) );
  OAI211_X1 U9426 ( .C1(n8161), .C2(n9263), .A(n8160), .B(n8159), .ZN(n8162)
         );
  AOI21_X1 U9427 ( .B1(n10690), .B2(n8163), .A(n8162), .ZN(n8164) );
  OAI21_X1 U9428 ( .B1(n8165), .B2(n10713), .A(n8164), .ZN(P2_U3195) );
  NOR2_X1 U9429 ( .A1(n8166), .A2(n8173), .ZN(n8168) );
  NOR2_X1 U9430 ( .A1(n8168), .A2(n8167), .ZN(n8170) );
  AOI22_X1 U9431 ( .A1(n8232), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n10290), .B2(
        n8172), .ZN(n8169) );
  NAND2_X1 U9432 ( .A1(n8169), .A2(n8170), .ZN(n8230) );
  OAI21_X1 U9433 ( .B1(n8170), .B2(n8169), .A(n8230), .ZN(n8182) );
  AND2_X1 U9434 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9697) );
  AOI21_X1 U9435 ( .B1(n9950), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n9697), .ZN(
        n8171) );
  OAI21_X1 U9436 ( .B1(n9947), .B2(n8172), .A(n8171), .ZN(n8181) );
  NOR2_X1 U9437 ( .A1(n8174), .A2(n8173), .ZN(n8176) );
  NOR2_X1 U9438 ( .A1(n8176), .A2(n8175), .ZN(n8179) );
  NAND2_X1 U9439 ( .A1(n8232), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8177) );
  OAI21_X1 U9440 ( .B1(n8232), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8177), .ZN(
        n8178) );
  NOR2_X1 U9441 ( .A1(n8179), .A2(n8178), .ZN(n8231) );
  AOI211_X1 U9442 ( .C1(n8179), .C2(n8178), .A(n8231), .B(n9953), .ZN(n8180)
         );
  AOI211_X1 U9443 ( .C1(n9944), .C2(n8182), .A(n8181), .B(n8180), .ZN(n8183)
         );
  INV_X1 U9444 ( .A(n8183), .ZN(P1_U3259) );
  NAND2_X1 U9445 ( .A1(n8188), .A2(n8977), .ZN(n8185) );
  NAND2_X1 U9446 ( .A1(n9796), .A2(n8965), .ZN(n8184) );
  NAND2_X1 U9447 ( .A1(n8185), .A2(n8184), .ZN(n8186) );
  XNOR2_X1 U9448 ( .A(n8186), .B(n8883), .ZN(n8214) );
  NOR2_X1 U9449 ( .A1(n10795), .A2(n8902), .ZN(n8187) );
  AOI21_X1 U9450 ( .B1(n8188), .B2(n8965), .A(n8187), .ZN(n8215) );
  XNOR2_X1 U9451 ( .A(n8214), .B(n8215), .ZN(n8189) );
  OAI21_X1 U9452 ( .B1(n8191), .B2(n8190), .A(n8189), .ZN(n8192) );
  INV_X1 U9453 ( .A(n8192), .ZN(n8193) );
  OAI21_X1 U9454 ( .B1(n5039), .B2(n8193), .A(n9764), .ZN(n8199) );
  OAI22_X1 U9455 ( .A1(n9783), .A2(n8195), .B1(n9781), .B2(n8194), .ZN(n8196)
         );
  AOI211_X1 U9456 ( .C1(n9768), .C2(n9795), .A(n8197), .B(n8196), .ZN(n8198)
         );
  OAI211_X1 U9457 ( .C1(n10825), .C2(n9737), .A(n8199), .B(n8198), .ZN(
        P1_U3224) );
  INV_X1 U9458 ( .A(n10828), .ZN(n10735) );
  NOR2_X1 U9459 ( .A1(n8200), .A2(n10735), .ZN(n8205) );
  OAI21_X1 U9460 ( .B1(n8877), .B2(n10824), .A(n8201), .ZN(n8202) );
  AOI211_X1 U9461 ( .C1(n8205), .C2(n8204), .A(n8203), .B(n8202), .ZN(n8208)
         );
  NAND2_X1 U9462 ( .A1(n6207), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8206) );
  OAI21_X1 U9463 ( .B1(n8208), .B2(n6207), .A(n8206), .ZN(P1_U3495) );
  NAND2_X1 U9464 ( .A1(n10830), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8207) );
  OAI21_X1 U9465 ( .B1(n8208), .B2(n10830), .A(n8207), .ZN(P1_U3536) );
  NAND2_X1 U9466 ( .A1(n8213), .A2(n8977), .ZN(n8210) );
  NAND2_X1 U9467 ( .A1(n9795), .A2(n8965), .ZN(n8209) );
  NAND2_X1 U9468 ( .A1(n8210), .A2(n8209), .ZN(n8211) );
  XNOR2_X1 U9469 ( .A(n8211), .B(n8883), .ZN(n8872) );
  NOR2_X1 U9470 ( .A1(n9646), .A2(n8902), .ZN(n8212) );
  AOI21_X1 U9471 ( .B1(n8213), .B2(n8965), .A(n8212), .ZN(n8873) );
  XNOR2_X1 U9472 ( .A(n8872), .B(n8873), .ZN(n8218) );
  INV_X1 U9473 ( .A(n8214), .ZN(n8217) );
  INV_X1 U9474 ( .A(n8215), .ZN(n8216) );
  NOR2_X1 U9475 ( .A1(n8217), .A2(n8216), .ZN(n8219) );
  OAI21_X1 U9476 ( .B1(n5039), .B2(n8219), .A(n8218), .ZN(n8220) );
  NAND3_X1 U9477 ( .A1(n5045), .A2(n9764), .A3(n8220), .ZN(n8226) );
  INV_X1 U9478 ( .A(n8221), .ZN(n8224) );
  OAI22_X1 U9479 ( .A1(n9779), .A2(n9782), .B1(n9781), .B2(n8222), .ZN(n8223)
         );
  AOI211_X1 U9480 ( .C1(n9767), .C2(n9796), .A(n8224), .B(n8223), .ZN(n8225)
         );
  OAI211_X1 U9481 ( .C1(n8227), .C2(n9737), .A(n8226), .B(n8225), .ZN(P1_U3234) );
  INV_X1 U9482 ( .A(n8228), .ZN(n8262) );
  AOI22_X1 U9483 ( .A1(n6704), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n9623), .ZN(n8229) );
  OAI21_X1 U9484 ( .B1(n8262), .B2(n9625), .A(n8229), .ZN(P2_U3269) );
  OAI21_X1 U9485 ( .B1(n8232), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8230), .ZN(
        n9914) );
  XOR2_X1 U9486 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9922), .Z(n9913) );
  XNOR2_X1 U9487 ( .A(n9914), .B(n9913), .ZN(n8237) );
  XNOR2_X1 U9488 ( .A(n9922), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n9924) );
  AOI21_X1 U9489 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n8232), .A(n8231), .ZN(
        n9921) );
  XNOR2_X1 U9490 ( .A(n9924), .B(n9921), .ZN(n8233) );
  NOR2_X1 U9491 ( .A1(n9953), .A2(n8233), .ZN(n8236) );
  NAND2_X1 U9492 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9706) );
  NAND2_X1 U9493 ( .A1(n9950), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n8234) );
  OAI211_X1 U9494 ( .C1(n9947), .C2(n9911), .A(n9706), .B(n8234), .ZN(n8235)
         );
  AOI211_X1 U9495 ( .C1(n8237), .C2(n9944), .A(n8236), .B(n8235), .ZN(n8238)
         );
  INV_X1 U9496 ( .A(n8238), .ZN(P1_U3260) );
  XNOR2_X1 U9497 ( .A(n8780), .B(n8630), .ZN(n8267) );
  XNOR2_X1 U9498 ( .A(n8267), .B(n9139), .ZN(n8250) );
  NAND2_X1 U9499 ( .A1(n8242), .A2(n8239), .ZN(n8240) );
  NAND2_X1 U9500 ( .A1(n8241), .A2(n8240), .ZN(n8245) );
  INV_X1 U9501 ( .A(n8242), .ZN(n8243) );
  NAND2_X1 U9502 ( .A1(n8243), .A2(n9554), .ZN(n8244) );
  NAND2_X1 U9503 ( .A1(n8245), .A2(n8244), .ZN(n8249) );
  INV_X1 U9504 ( .A(n8249), .ZN(n8247) );
  INV_X1 U9505 ( .A(n8270), .ZN(n8248) );
  AOI21_X1 U9506 ( .B1(n8250), .B2(n8249), .A(n8248), .ZN(n8255) );
  INV_X1 U9507 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10542) );
  OR2_X1 U9508 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10542), .ZN(n9163) );
  OAI21_X1 U9509 ( .B1(n9129), .B2(n10576), .A(n9163), .ZN(n8251) );
  AOI21_X1 U9510 ( .B1(n9126), .B2(n9554), .A(n8251), .ZN(n8252) );
  OAI21_X1 U9511 ( .B1(n9006), .B2(n10839), .A(n8252), .ZN(n8253) );
  AOI21_X1 U9512 ( .B1(n8780), .B2(n9131), .A(n8253), .ZN(n8254) );
  OAI21_X1 U9513 ( .B1(n8255), .B2(n9133), .A(n8254), .ZN(P2_U3155) );
  NOR2_X1 U9514 ( .A1(n8256), .A2(n9559), .ZN(n8258) );
  AOI211_X1 U9515 ( .C1(n9525), .C2(n8259), .A(n8258), .B(n8257), .ZN(n10822)
         );
  OR2_X1 U9516 ( .A1(n10822), .A2(n9570), .ZN(n8260) );
  OAI21_X1 U9517 ( .B1(n9561), .B2(n6419), .A(n8260), .ZN(P2_U3471) );
  OAI222_X1 U9518 ( .A1(n8263), .A2(P1_U3086), .B1(n10354), .B2(n8262), .C1(
        n8261), .C2(n10350), .ZN(P1_U3329) );
  INV_X1 U9519 ( .A(n8264), .ZN(n8303) );
  AOI21_X1 U9520 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n9623), .A(n8265), .ZN(
        n8266) );
  OAI21_X1 U9521 ( .B1(n8303), .B2(n9625), .A(n8266), .ZN(P2_U3268) );
  INV_X1 U9522 ( .A(n9545), .ZN(n8277) );
  INV_X1 U9523 ( .A(n8267), .ZN(n8268) );
  NAND2_X1 U9524 ( .A1(n8268), .A2(n9472), .ZN(n8269) );
  XNOR2_X1 U9525 ( .A(n9545), .B(n8635), .ZN(n8595) );
  XNOR2_X1 U9526 ( .A(n8595), .B(n9551), .ZN(n8271) );
  OAI211_X1 U9527 ( .C1(n5048), .C2(n8271), .A(n8598), .B(n9091), .ZN(n8276)
         );
  NOR2_X1 U9528 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8272), .ZN(n9184) );
  AOI21_X1 U9529 ( .B1(n9081), .B2(n9428), .A(n9184), .ZN(n8273) );
  OAI21_X1 U9530 ( .B1(n9472), .B2(n9094), .A(n8273), .ZN(n8274) );
  AOI21_X1 U9531 ( .B1(n9459), .B2(n9125), .A(n8274), .ZN(n8275) );
  OAI211_X1 U9532 ( .C1(n8277), .C2(n9114), .A(n8276), .B(n8275), .ZN(P2_U3181) );
  AND2_X1 U9533 ( .A1(n8278), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U9534 ( .A1(n8278), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U9535 ( .A1(n8278), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U9536 ( .A1(n8278), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U9537 ( .A1(n8278), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U9538 ( .A1(n8278), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U9539 ( .A1(n8278), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U9540 ( .A1(n8278), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U9541 ( .A1(n8278), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U9542 ( .A1(n8278), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U9543 ( .A1(n8278), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U9544 ( .A1(n8278), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U9545 ( .A1(n8278), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U9546 ( .A1(n8278), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U9547 ( .A1(n8278), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U9548 ( .A1(n8278), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U9549 ( .A1(n8278), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U9550 ( .A1(n8278), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U9551 ( .A1(n8278), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U9552 ( .A1(n8278), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U9553 ( .A1(n8278), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U9554 ( .A1(n8278), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U9555 ( .A1(n8278), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U9556 ( .A1(n8278), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U9557 ( .A1(n8278), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U9558 ( .A1(n8278), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U9559 ( .A1(n8278), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U9560 ( .A1(n8278), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U9561 ( .A1(n8278), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U9562 ( .A1(n8278), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  INV_X1 U9563 ( .A(SI_29_), .ZN(n10487) );
  INV_X1 U9564 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8283) );
  INV_X1 U9565 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8992) );
  MUX2_X1 U9566 ( .A(n8283), .B(n8992), .S(n8328), .Z(n8284) );
  INV_X1 U9567 ( .A(SI_30_), .ZN(n10484) );
  NAND2_X1 U9568 ( .A1(n8284), .A2(n10484), .ZN(n8325) );
  INV_X1 U9569 ( .A(n8284), .ZN(n8285) );
  NAND2_X1 U9570 ( .A1(n8285), .A2(SI_30_), .ZN(n8286) );
  NAND2_X1 U9571 ( .A1(n8325), .A2(n8286), .ZN(n8326) );
  OR2_X1 U9572 ( .A1(n8287), .A2(n8992), .ZN(n8288) );
  NAND2_X1 U9573 ( .A1(n10306), .A2(n8290), .ZN(n9955) );
  OR2_X1 U9574 ( .A1(n8290), .A2(n10306), .ZN(n8291) );
  NAND3_X1 U9575 ( .A1(n9955), .A2(n8291), .A3(n10782), .ZN(n9965) );
  NAND2_X1 U9576 ( .A1(n8292), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8297) );
  INV_X1 U9577 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8293) );
  OR2_X1 U9578 ( .A1(n6727), .A2(n8293), .ZN(n8296) );
  INV_X1 U9579 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10300) );
  OR2_X1 U9580 ( .A1(n8294), .A2(n10300), .ZN(n8295) );
  AND3_X1 U9581 ( .A1(n8297), .A2(n8296), .A3(n8295), .ZN(n8440) );
  NOR2_X1 U9582 ( .A1(n8298), .A2(n8440), .ZN(n10201) );
  INV_X1 U9583 ( .A(n10201), .ZN(n9957) );
  NAND2_X1 U9584 ( .A1(n9965), .A2(n9957), .ZN(n10303) );
  MUX2_X1 U9585 ( .A(n10303), .B(P1_REG1_REG_30__SCAN_IN), .S(n10830), .Z(
        n8299) );
  INV_X1 U9586 ( .A(n8299), .ZN(n8300) );
  OAI21_X1 U9587 ( .B1(n10306), .B2(n10298), .A(n8300), .ZN(P1_U3552) );
  NAND2_X1 U9588 ( .A1(n10574), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8301) );
  OAI21_X1 U9589 ( .B1(n8302), .B2(n10574), .A(n8301), .ZN(P2_U3491) );
  OAI222_X1 U9590 ( .A1(n8304), .A2(P1_U3086), .B1(n10354), .B2(n8303), .C1(
        n10350), .C2(n6097), .ZN(P1_U3328) );
  XOR2_X1 U9591 ( .A(n8306), .B(n8305), .Z(n8307) );
  XNOR2_X1 U9592 ( .A(n8308), .B(n8307), .ZN(n8316) );
  INV_X1 U9593 ( .A(n8309), .ZN(n8312) );
  OAI22_X1 U9594 ( .A1(n9779), .A2(n8373), .B1(n9781), .B2(n8310), .ZN(n8311)
         );
  AOI211_X1 U9595 ( .C1(n9767), .C2(n9802), .A(n8312), .B(n8311), .ZN(n8315)
         );
  NAND2_X1 U9596 ( .A1(n4944), .A2(n8313), .ZN(n8314) );
  OAI211_X1 U9597 ( .C1(n8316), .C2(n9788), .A(n8315), .B(n8314), .ZN(P1_U3213) );
  OAI21_X1 U9598 ( .B1(n8319), .B2(n8318), .A(n8317), .ZN(n9821) );
  AOI22_X1 U9599 ( .A1(n4944), .A2(n10722), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n8320), .ZN(n8322) );
  NAND2_X1 U9600 ( .A1(n9768), .A2(n9807), .ZN(n8321) );
  OAI211_X1 U9601 ( .C1(n9788), .C2(n9821), .A(n8322), .B(n8321), .ZN(P1_U3232) );
  NOR2_X1 U9602 ( .A1(n8324), .A2(n8323), .ZN(n8586) );
  OAI21_X1 U9603 ( .B1(n8579), .B2(n8481), .A(P1_B_REG_SCAN_IN), .ZN(n8585) );
  MUX2_X1 U9604 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n8328), .Z(n8329) );
  XOR2_X1 U9605 ( .A(n8329), .B(SI_31_), .Z(n8330) );
  INV_X1 U9606 ( .A(n8440), .ZN(n9790) );
  NAND2_X1 U9607 ( .A1(n10302), .A2(n9790), .ZN(n8574) );
  INV_X1 U9608 ( .A(n8574), .ZN(n8507) );
  MUX2_X1 U9609 ( .A(n8499), .B(n8502), .S(n8442), .Z(n8437) );
  INV_X1 U9610 ( .A(n8483), .ZN(n8429) );
  INV_X1 U9611 ( .A(n8421), .ZN(n10051) );
  AND2_X1 U9612 ( .A1(n9793), .A2(n8442), .ZN(n8336) );
  OAI21_X1 U9613 ( .B1(n8442), .B2(n9793), .A(n10176), .ZN(n8335) );
  OAI21_X1 U9614 ( .B1(n8336), .B2(n10176), .A(n8335), .ZN(n8404) );
  AND2_X1 U9615 ( .A1(n8522), .A2(n8528), .ZN(n8338) );
  NAND2_X1 U9616 ( .A1(n8344), .A2(n8341), .ZN(n8337) );
  AOI21_X1 U9617 ( .B1(n8339), .B2(n8338), .A(n8337), .ZN(n8347) );
  AND2_X1 U9618 ( .A1(n8341), .A2(n8340), .ZN(n8527) );
  OAI21_X1 U9619 ( .B1(n8523), .B2(n8342), .A(n8527), .ZN(n8343) );
  NAND2_X1 U9620 ( .A1(n8343), .A2(n8528), .ZN(n8345) );
  AOI21_X1 U9621 ( .B1(n8345), .B2(n8344), .A(n8350), .ZN(n8346) );
  INV_X1 U9622 ( .A(n8442), .ZN(n8445) );
  MUX2_X1 U9623 ( .A(n8347), .B(n8346), .S(n8445), .Z(n8349) );
  INV_X1 U9624 ( .A(n8455), .ZN(n8348) );
  NAND2_X1 U9625 ( .A1(n8349), .A2(n8348), .ZN(n8368) );
  NAND2_X1 U9626 ( .A1(n8350), .A2(n8365), .ZN(n8352) );
  NAND2_X1 U9627 ( .A1(n8352), .A2(n8351), .ZN(n8531) );
  NOR2_X1 U9628 ( .A1(n8531), .A2(n8353), .ZN(n8356) );
  INV_X1 U9629 ( .A(n8354), .ZN(n8355) );
  AOI21_X1 U9630 ( .B1(n8368), .B2(n8356), .A(n8355), .ZN(n8357) );
  MUX2_X1 U9631 ( .A(n8361), .B(n8360), .S(n8442), .Z(n8362) );
  NAND2_X1 U9632 ( .A1(n8363), .A2(n8362), .ZN(n8364) );
  INV_X1 U9633 ( .A(n8364), .ZN(n8367) );
  NAND4_X1 U9634 ( .A1(n8368), .A2(n8367), .A3(n8366), .A4(n8365), .ZN(n8370)
         );
  NAND3_X1 U9635 ( .A1(n8370), .A2(n10789), .A3(n8369), .ZN(n8371) );
  INV_X1 U9636 ( .A(n8375), .ZN(n8376) );
  NAND2_X1 U9637 ( .A1(n10789), .A2(n8376), .ZN(n8377) );
  AND2_X1 U9638 ( .A1(n8377), .A2(n8540), .ZN(n8382) );
  NAND2_X1 U9639 ( .A1(n8385), .A2(n10789), .ZN(n8539) );
  INV_X1 U9640 ( .A(n8378), .ZN(n8379) );
  AND2_X1 U9641 ( .A1(n8540), .A2(n8379), .ZN(n8380) );
  NOR2_X1 U9642 ( .A1(n8539), .A2(n8380), .ZN(n8381) );
  MUX2_X1 U9643 ( .A(n8382), .B(n8381), .S(n8442), .Z(n8383) );
  NAND2_X1 U9644 ( .A1(n8384), .A2(n8383), .ZN(n8390) );
  NAND2_X1 U9645 ( .A1(n8392), .A2(n8385), .ZN(n8387) );
  NAND2_X1 U9646 ( .A1(n8391), .A2(n8386), .ZN(n8542) );
  MUX2_X1 U9647 ( .A(n8387), .B(n8542), .S(n8442), .Z(n8388) );
  INV_X1 U9648 ( .A(n8388), .ZN(n8389) );
  NAND2_X1 U9649 ( .A1(n8390), .A2(n8389), .ZN(n8395) );
  NAND2_X1 U9650 ( .A1(n9649), .A2(n9782), .ZN(n8396) );
  AND2_X1 U9651 ( .A1(n8393), .A2(n8392), .ZN(n8544) );
  INV_X1 U9652 ( .A(n8545), .ZN(n8394) );
  AOI21_X1 U9653 ( .B1(n8395), .B2(n8544), .A(n8394), .ZN(n8399) );
  INV_X1 U9654 ( .A(n8396), .ZN(n8398) );
  AND2_X1 U9655 ( .A1(n8518), .A2(n8397), .ZN(n8546) );
  OAI21_X1 U9656 ( .B1(n8399), .B2(n8398), .A(n8546), .ZN(n8401) );
  NAND4_X1 U9657 ( .A1(n8401), .A2(n8442), .A3(n8400), .A4(n8549), .ZN(n8402)
         );
  NAND4_X1 U9658 ( .A1(n10147), .A2(n8404), .A3(n8403), .A4(n8402), .ZN(n8409)
         );
  NAND2_X1 U9659 ( .A1(n8409), .A2(n8405), .ZN(n8406) );
  AND2_X1 U9660 ( .A1(n8408), .A2(n8407), .ZN(n8555) );
  NAND2_X1 U9661 ( .A1(n8409), .A2(n8555), .ZN(n8410) );
  INV_X1 U9662 ( .A(n8415), .ZN(n8556) );
  AND2_X1 U9663 ( .A1(n8418), .A2(n8411), .ZN(n8559) );
  OAI211_X1 U9664 ( .C1(n8414), .C2(n10084), .A(n8422), .B(n8413), .ZN(n8420)
         );
  NAND3_X1 U9665 ( .A1(n8416), .A2(n8415), .A3(n10082), .ZN(n8417) );
  AOI21_X1 U9666 ( .B1(n8418), .B2(n8417), .A(n10084), .ZN(n8419) );
  NAND2_X1 U9667 ( .A1(n8424), .A2(n8421), .ZN(n8486) );
  NAND2_X1 U9668 ( .A1(n8487), .A2(n8422), .ZN(n8491) );
  MUX2_X1 U9669 ( .A(n8486), .B(n8491), .S(n8442), .Z(n8423) );
  INV_X1 U9670 ( .A(n8472), .ZN(n10040) );
  INV_X1 U9671 ( .A(n8424), .ZN(n8425) );
  NAND3_X1 U9672 ( .A1(n8426), .A2(n8488), .A3(n8483), .ZN(n8427) );
  NAND2_X1 U9673 ( .A1(n8427), .A2(n9995), .ZN(n8428) );
  INV_X1 U9674 ( .A(n8487), .ZN(n8430) );
  OAI211_X1 U9675 ( .C1(n8431), .C2(n8430), .A(n10026), .B(n8484), .ZN(n8432)
         );
  NAND4_X1 U9676 ( .A1(n8432), .A2(n8445), .A3(n10007), .A4(n8495), .ZN(n8433)
         );
  NAND2_X1 U9677 ( .A1(n8433), .A2(n9996), .ZN(n8436) );
  MUX2_X1 U9678 ( .A(n8501), .B(n8564), .S(n8442), .Z(n8434) );
  MUX2_X1 U9679 ( .A(n8503), .B(n8438), .S(n8442), .Z(n8441) );
  OAI21_X1 U9680 ( .B1(n10306), .B2(n9790), .A(n8567), .ZN(n8508) );
  INV_X1 U9681 ( .A(n8439), .ZN(n9791) );
  NOR2_X1 U9682 ( .A1(n8571), .A2(n8440), .ZN(n8482) );
  OAI21_X1 U9683 ( .B1(n8444), .B2(n8443), .A(n8574), .ZN(n8446) );
  AOI211_X1 U9684 ( .C1(n6137), .C2(n8507), .A(n8481), .B(n8447), .ZN(n8583)
         );
  NAND2_X1 U9685 ( .A1(n8571), .A2(n8567), .ZN(n8477) );
  XNOR2_X1 U9686 ( .A(n10143), .B(n10279), .ZN(n10131) );
  INV_X1 U9687 ( .A(n10779), .ZN(n10788) );
  INV_X1 U9688 ( .A(n8448), .ZN(n8459) );
  AND2_X1 U9689 ( .A1(n8449), .A2(n5056), .ZN(n8521) );
  NOR2_X1 U9690 ( .A1(n8450), .A2(n8521), .ZN(n10734) );
  NAND4_X1 U9691 ( .A1(n10734), .A2(n8452), .A3(n8519), .A4(n8451), .ZN(n8456)
         );
  NOR4_X1 U9692 ( .A1(n8456), .A2(n8455), .A3(n8454), .A4(n8453), .ZN(n8458)
         );
  NAND4_X1 U9693 ( .A1(n8535), .A2(n8459), .A3(n8458), .A4(n8457), .ZN(n8461)
         );
  NOR2_X1 U9694 ( .A1(n8461), .A2(n8460), .ZN(n8462) );
  NAND4_X1 U9695 ( .A1(n8464), .A2(n8463), .A3(n10788), .A4(n8462), .ZN(n8465)
         );
  NOR3_X1 U9696 ( .A1(n8467), .A2(n8466), .A3(n8465), .ZN(n8468) );
  NAND3_X1 U9697 ( .A1(n10147), .A2(n10169), .A3(n8468), .ZN(n8469) );
  NOR4_X1 U9698 ( .A1(n10101), .A2(n10113), .A3(n10131), .A4(n8469), .ZN(n8470) );
  NAND4_X1 U9699 ( .A1(n10054), .A2(n5167), .A3(n10063), .A4(n8470), .ZN(n8471) );
  NOR2_X1 U9700 ( .A1(n8472), .A2(n8471), .ZN(n8473) );
  NAND4_X1 U9701 ( .A1(n9996), .A2(n10026), .A3(n10007), .A4(n8473), .ZN(n8474) );
  OAI211_X1 U9702 ( .C1(n8481), .C2(n8519), .A(n8480), .B(n6137), .ZN(n8517)
         );
  INV_X1 U9703 ( .A(n8482), .ZN(n8510) );
  NAND2_X1 U9704 ( .A1(n8499), .A2(n8483), .ZN(n8570) );
  INV_X1 U9705 ( .A(n8484), .ZN(n8485) );
  AOI21_X1 U9706 ( .B1(n8487), .B2(n8486), .A(n8485), .ZN(n8490) );
  INV_X1 U9707 ( .A(n8494), .ZN(n8489) );
  OAI21_X1 U9708 ( .B1(n8490), .B2(n8489), .A(n8488), .ZN(n8563) );
  INV_X1 U9709 ( .A(n8491), .ZN(n8493) );
  AND3_X1 U9710 ( .A1(n8494), .A2(n8493), .A3(n8492), .ZN(n8496) );
  OAI211_X1 U9711 ( .C1(n8563), .C2(n8496), .A(n9995), .B(n8495), .ZN(n8565)
         );
  NOR2_X1 U9712 ( .A1(n8563), .A2(n8497), .ZN(n8498) );
  OAI21_X1 U9713 ( .B1(n8565), .B2(n8498), .A(n8564), .ZN(n8506) );
  INV_X1 U9714 ( .A(n8499), .ZN(n8500) );
  AOI21_X1 U9715 ( .B1(n8502), .B2(n8501), .A(n8500), .ZN(n8505) );
  INV_X1 U9716 ( .A(n8503), .ZN(n8504) );
  NOR2_X1 U9717 ( .A1(n8505), .A2(n8504), .ZN(n8568) );
  OAI21_X1 U9718 ( .B1(n8570), .B2(n8506), .A(n8568), .ZN(n8509) );
  AOI211_X1 U9719 ( .C1(n8510), .C2(n8509), .A(n8508), .B(n8507), .ZN(n8512)
         );
  NOR3_X1 U9720 ( .A1(n8512), .A2(n8573), .A3(n8511), .ZN(n8514) );
  OAI21_X1 U9721 ( .B1(n8514), .B2(n8513), .A(n9946), .ZN(n8516) );
  INV_X1 U9722 ( .A(n8518), .ZN(n8551) );
  AOI21_X1 U9723 ( .B1(n8520), .B2(n9807), .A(n8519), .ZN(n8526) );
  INV_X1 U9724 ( .A(n8521), .ZN(n8525) );
  INV_X1 U9725 ( .A(n8522), .ZN(n8524) );
  AOI211_X1 U9726 ( .C1(n8526), .C2(n8525), .A(n8524), .B(n8523), .ZN(n8530)
         );
  INV_X1 U9727 ( .A(n8527), .ZN(n8529) );
  OAI21_X1 U9728 ( .B1(n8530), .B2(n8529), .A(n8528), .ZN(n8534) );
  AOI211_X1 U9729 ( .C1(n8534), .C2(n8533), .A(n8532), .B(n8531), .ZN(n8538)
         );
  INV_X1 U9730 ( .A(n8535), .ZN(n8537) );
  OAI21_X1 U9731 ( .B1(n8538), .B2(n8537), .A(n8536), .ZN(n8541) );
  AOI21_X1 U9732 ( .B1(n8541), .B2(n8540), .A(n8539), .ZN(n8543) );
  NOR2_X1 U9733 ( .A1(n8543), .A2(n8542), .ZN(n8548) );
  INV_X1 U9734 ( .A(n8544), .ZN(n8547) );
  OAI211_X1 U9735 ( .C1(n8548), .C2(n8547), .A(n8546), .B(n8545), .ZN(n8550)
         );
  OAI211_X1 U9736 ( .C1(n5042), .C2(n8551), .A(n8550), .B(n8549), .ZN(n8552)
         );
  NAND3_X1 U9737 ( .A1(n10128), .A2(n8553), .A3(n8552), .ZN(n8554) );
  NAND2_X1 U9738 ( .A1(n8555), .A2(n8554), .ZN(n8557) );
  AOI21_X1 U9739 ( .B1(n8558), .B2(n8557), .A(n8556), .ZN(n8561) );
  INV_X1 U9740 ( .A(n8559), .ZN(n8560) );
  NOR4_X1 U9741 ( .A1(n8563), .A2(n8562), .A3(n8561), .A4(n8560), .ZN(n8566)
         );
  OAI21_X1 U9742 ( .B1(n8566), .B2(n8565), .A(n8564), .ZN(n8569) );
  OAI211_X1 U9743 ( .C1(n8570), .C2(n8569), .A(n8568), .B(n8567), .ZN(n8572)
         );
  NAND2_X1 U9744 ( .A1(n8572), .A2(n8571), .ZN(n8575) );
  AND2_X1 U9745 ( .A1(n6137), .A2(n8576), .ZN(n10724) );
  NOR2_X1 U9746 ( .A1(n8580), .A2(n8577), .ZN(n8578) );
  AOI211_X1 U9747 ( .C1(n8580), .C2(n10724), .A(n8579), .B(n8578), .ZN(n8581)
         );
  OAI21_X1 U9748 ( .B1(n8583), .B2(n8582), .A(n8581), .ZN(n8584) );
  OAI21_X1 U9749 ( .B1(n8586), .B2(n8585), .A(n8584), .ZN(P1_U3242) );
  NAND2_X1 U9750 ( .A1(n8587), .A2(n10846), .ZN(n8592) );
  NOR2_X1 U9751 ( .A1(n10838), .A2(n8588), .ZN(n9273) );
  NOR2_X1 U9752 ( .A1(n8589), .A2(n9360), .ZN(n8590) );
  AOI211_X1 U9753 ( .C1(n4949), .C2(P2_REG2_REG_29__SCAN_IN), .A(n9273), .B(
        n8590), .ZN(n8591) );
  OAI211_X1 U9754 ( .C1(n8594), .C2(n8593), .A(n8592), .B(n8591), .ZN(P2_U3204) );
  INV_X1 U9755 ( .A(n8595), .ZN(n8596) );
  NAND2_X1 U9756 ( .A1(n8596), .A2(n9551), .ZN(n8597) );
  XNOR2_X1 U9757 ( .A(n9538), .B(n8630), .ZN(n9051) );
  AND2_X1 U9758 ( .A1(n9051), .A2(n9428), .ZN(n8599) );
  XNOR2_X1 U9759 ( .A(n9534), .B(n8635), .ZN(n9061) );
  AND2_X1 U9760 ( .A1(n9061), .A2(n9060), .ZN(n8603) );
  INV_X1 U9761 ( .A(n9061), .ZN(n8601) );
  NAND2_X1 U9762 ( .A1(n8601), .A2(n9440), .ZN(n8602) );
  OAI21_X1 U9763 ( .B1(n9059), .B2(n8603), .A(n8602), .ZN(n9110) );
  XNOR2_X1 U9764 ( .A(n9530), .B(n8635), .ZN(n8604) );
  XNOR2_X1 U9765 ( .A(n8604), .B(n9427), .ZN(n9111) );
  INV_X1 U9766 ( .A(n8604), .ZN(n8605) );
  AOI21_X2 U9767 ( .B1(n9110), .B2(n9111), .A(n8606), .ZN(n9023) );
  XNOR2_X1 U9768 ( .A(n8607), .B(n8630), .ZN(n9022) );
  NAND2_X1 U9769 ( .A1(n9023), .A2(n9022), .ZN(n8610) );
  XNOR2_X1 U9770 ( .A(n9519), .B(n8635), .ZN(n8611) );
  NAND2_X1 U9771 ( .A1(n8611), .A2(n9407), .ZN(n9030) );
  INV_X1 U9772 ( .A(n8611), .ZN(n8612) );
  NAND2_X1 U9773 ( .A1(n8612), .A2(n9037), .ZN(n8613) );
  XNOR2_X1 U9774 ( .A(n9375), .B(n8635), .ZN(n8615) );
  XNOR2_X1 U9775 ( .A(n8615), .B(n9391), .ZN(n9031) );
  NAND2_X1 U9776 ( .A1(n8615), .A2(n9095), .ZN(n8616) );
  XNOR2_X1 U9777 ( .A(n9101), .B(n8630), .ZN(n8618) );
  XNOR2_X1 U9778 ( .A(n8618), .B(n9338), .ZN(n9102) );
  INV_X1 U9779 ( .A(n9102), .ZN(n8617) );
  NAND2_X1 U9780 ( .A1(n8618), .A2(n9338), .ZN(n8619) );
  XNOR2_X1 U9781 ( .A(n9503), .B(n8630), .ZN(n8620) );
  INV_X1 U9782 ( .A(n8623), .ZN(n9069) );
  XNOR2_X1 U9783 ( .A(n8698), .B(n8635), .ZN(n8624) );
  NAND2_X1 U9784 ( .A1(n8624), .A2(n9316), .ZN(n8627) );
  INV_X1 U9785 ( .A(n8624), .ZN(n8625) );
  NAND2_X1 U9786 ( .A1(n8625), .A2(n5509), .ZN(n8626) );
  NAND2_X1 U9787 ( .A1(n8627), .A2(n8626), .ZN(n9068) );
  INV_X1 U9788 ( .A(n8627), .ZN(n9044) );
  XNOR2_X1 U9789 ( .A(n9318), .B(n8635), .ZN(n8628) );
  XNOR2_X1 U9790 ( .A(n8628), .B(n9138), .ZN(n9043) );
  XNOR2_X1 U9791 ( .A(n9308), .B(n8630), .ZN(n8631) );
  NOR2_X1 U9792 ( .A1(n8631), .A2(n9137), .ZN(n9120) );
  NAND2_X1 U9793 ( .A1(n8631), .A2(n9137), .ZN(n9121) );
  XNOR2_X1 U9794 ( .A(n8632), .B(n8635), .ZN(n8633) );
  NOR2_X1 U9795 ( .A1(n8633), .A2(n9305), .ZN(n8634) );
  AOI21_X1 U9796 ( .B1(n9305), .B2(n8633), .A(n8634), .ZN(n8997) );
  XOR2_X1 U9797 ( .A(n8635), .B(n9285), .Z(n8636) );
  AOI22_X1 U9798 ( .A1(n9081), .A2(n9282), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8639) );
  INV_X1 U9799 ( .A(n9288), .ZN(n8637) );
  NAND2_X1 U9800 ( .A1(n9125), .A2(n8637), .ZN(n8638) );
  OAI211_X1 U9801 ( .C1(n9305), .C2(n9094), .A(n8639), .B(n8638), .ZN(n8640)
         );
  AOI21_X1 U9802 ( .B1(n9483), .B2(n9131), .A(n8640), .ZN(n8641) );
  OAI21_X1 U9803 ( .B1(n8642), .B2(n9133), .A(n8641), .ZN(P2_U3160) );
  INV_X1 U9804 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8644) );
  OR2_X1 U9805 ( .A1(n8645), .A2(n8644), .ZN(n8652) );
  INV_X1 U9806 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8646) );
  OR2_X1 U9807 ( .A1(n8647), .A2(n8646), .ZN(n8651) );
  INV_X1 U9808 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8648) );
  OR2_X1 U9809 ( .A1(n8649), .A2(n8648), .ZN(n8650) );
  NAND4_X1 U9810 ( .A1(n8653), .A2(n8652), .A3(n8651), .A4(n8650), .ZN(n9275)
         );
  NOR2_X1 U9811 ( .A1(n9573), .A2(n9275), .ZN(n8855) );
  INV_X1 U9812 ( .A(n9573), .ZN(n8655) );
  INV_X1 U9813 ( .A(n9275), .ZN(n8654) );
  NAND2_X1 U9814 ( .A1(n8990), .A2(n8656), .ZN(n8658) );
  NAND2_X1 U9815 ( .A1(n8643), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8657) );
  INV_X1 U9816 ( .A(n9135), .ZN(n8659) );
  INV_X1 U9817 ( .A(n8689), .ZN(n8854) );
  INV_X1 U9818 ( .A(n8661), .ZN(n8831) );
  OR2_X1 U9819 ( .A1(n8828), .A2(n5505), .ZN(n9340) );
  NAND4_X1 U9820 ( .A1(n8722), .A2(n8664), .A3(n8663), .A4(n6274), .ZN(n8667)
         );
  INV_X1 U9821 ( .A(n8665), .ZN(n8666) );
  NOR3_X1 U9822 ( .A1(n8667), .A2(n8666), .A3(n8729), .ZN(n8670) );
  NAND4_X1 U9823 ( .A1(n8670), .A2(n8669), .A3(n8668), .A4(n8740), .ZN(n8672)
         );
  NOR2_X1 U9824 ( .A1(n8672), .A2(n8671), .ZN(n8674) );
  NAND3_X1 U9825 ( .A1(n8675), .A2(n8674), .A3(n8673), .ZN(n8676) );
  NOR2_X1 U9826 ( .A1(n9466), .A2(n8676), .ZN(n8677) );
  NAND3_X1 U9827 ( .A1(n9557), .A2(n8677), .A3(n8767), .ZN(n8678) );
  NOR2_X1 U9828 ( .A1(n8678), .A2(n9455), .ZN(n8679) );
  AND4_X1 U9829 ( .A1(n9421), .A2(n5349), .A3(n8679), .A4(n9434), .ZN(n8680)
         );
  NAND4_X1 U9830 ( .A1(n4982), .A2(n9403), .A3(n9388), .A4(n8680), .ZN(n8681)
         );
  OR3_X1 U9831 ( .A1(n9340), .A2(n9352), .A3(n8681), .ZN(n8682) );
  NOR2_X1 U9832 ( .A1(n9321), .A2(n8682), .ZN(n8683) );
  INV_X1 U9833 ( .A(n9326), .ZN(n9333) );
  NAND4_X1 U9834 ( .A1(n9296), .A2(n9306), .A3(n8683), .A4(n9333), .ZN(n8684)
         );
  NOR2_X1 U9835 ( .A1(n8684), .A2(n9285), .ZN(n8685) );
  NAND4_X1 U9836 ( .A1(n8853), .A2(n8686), .A3(n8854), .A4(n8685), .ZN(n8687)
         );
  NOR3_X1 U9837 ( .A1(n8855), .A2(n8856), .A3(n8687), .ZN(n8695) );
  INV_X1 U9838 ( .A(n8688), .ZN(n8851) );
  OAI21_X1 U9839 ( .B1(n9278), .B2(n9275), .A(n9573), .ZN(n8692) );
  AOI21_X1 U9840 ( .B1(n8853), .B2(n9275), .A(n9573), .ZN(n8691) );
  MUX2_X1 U9841 ( .A(n8695), .B(n8694), .S(n8693), .Z(n8697) );
  XNOR2_X1 U9842 ( .A(n8697), .B(n8696), .ZN(n8863) );
  NOR3_X1 U9843 ( .A1(n8698), .A2(n9316), .A3(n8842), .ZN(n8700) );
  NOR3_X1 U9844 ( .A1(n5510), .A2(n8849), .A3(n5509), .ZN(n8699) );
  NOR3_X1 U9845 ( .A1(n9321), .A2(n8700), .A3(n8699), .ZN(n8835) );
  INV_X1 U9846 ( .A(n8701), .ZN(n8823) );
  MUX2_X1 U9847 ( .A(n9391), .B(n9375), .S(n8849), .Z(n8819) );
  INV_X1 U9848 ( .A(n8819), .ZN(n8822) );
  INV_X1 U9849 ( .A(n8702), .ZN(n8820) );
  INV_X1 U9850 ( .A(n8760), .ZN(n8703) );
  NAND2_X1 U9851 ( .A1(n8705), .A2(n8704), .ZN(n8706) );
  AND2_X1 U9852 ( .A1(n8707), .A2(n8706), .ZN(n8709) );
  OAI211_X1 U9853 ( .C1(n8711), .C2(n8709), .A(n8708), .B(n8762), .ZN(n8710)
         );
  NAND2_X1 U9854 ( .A1(n8710), .A2(n8849), .ZN(n8743) );
  INV_X1 U9855 ( .A(n8711), .ZN(n8758) );
  NAND2_X1 U9856 ( .A1(n8713), .A2(n8712), .ZN(n8714) );
  NAND3_X1 U9857 ( .A1(n8718), .A2(n8714), .A3(n8717), .ZN(n8715) );
  NAND2_X1 U9858 ( .A1(n8715), .A2(n8716), .ZN(n8721) );
  INV_X1 U9859 ( .A(n8716), .ZN(n8719) );
  OAI21_X1 U9860 ( .B1(n8719), .B2(n8718), .A(n8717), .ZN(n8720) );
  MUX2_X1 U9861 ( .A(n8721), .B(n8720), .S(n8849), .Z(n8723) );
  NAND2_X1 U9862 ( .A1(n8723), .A2(n8722), .ZN(n8731) );
  NAND2_X1 U9863 ( .A1(n8748), .A2(n8724), .ZN(n8727) );
  NAND2_X1 U9864 ( .A1(n8732), .A2(n8725), .ZN(n8726) );
  MUX2_X1 U9865 ( .A(n8727), .B(n8726), .S(n8842), .Z(n8728) );
  INV_X1 U9866 ( .A(n8728), .ZN(n8730) );
  AOI21_X1 U9867 ( .B1(n8731), .B2(n8730), .A(n8729), .ZN(n8749) );
  NAND2_X1 U9868 ( .A1(n8749), .A2(n8732), .ZN(n8735) );
  AND2_X1 U9869 ( .A1(n8736), .A2(n8733), .ZN(n8750) );
  NAND3_X1 U9870 ( .A1(n8735), .A2(n8750), .A3(n8734), .ZN(n8739) );
  NAND2_X1 U9871 ( .A1(n8751), .A2(n8746), .ZN(n8737) );
  AOI21_X1 U9872 ( .B1(n8737), .B2(n8736), .A(n8842), .ZN(n8738) );
  NAND2_X1 U9873 ( .A1(n8739), .A2(n8738), .ZN(n8741) );
  NAND3_X1 U9874 ( .A1(n8758), .A2(n8741), .A3(n8740), .ZN(n8742) );
  NAND2_X1 U9875 ( .A1(n8743), .A2(n8742), .ZN(n8752) );
  NAND3_X1 U9876 ( .A1(n8752), .A2(n8765), .A3(n4987), .ZN(n8744) );
  NAND2_X1 U9877 ( .A1(n8744), .A2(n8763), .ZN(n8766) );
  NAND2_X1 U9878 ( .A1(n8746), .A2(n8745), .ZN(n8747) );
  AOI21_X1 U9879 ( .B1(n8749), .B2(n8748), .A(n8747), .ZN(n8754) );
  INV_X1 U9880 ( .A(n8750), .ZN(n8753) );
  OAI211_X1 U9881 ( .C1(n8754), .C2(n8753), .A(n8752), .B(n8751), .ZN(n8761)
         );
  NAND2_X1 U9882 ( .A1(n8756), .A2(n8755), .ZN(n8757) );
  NAND2_X1 U9883 ( .A1(n8758), .A2(n8757), .ZN(n8759) );
  NAND4_X1 U9884 ( .A1(n8761), .A2(n8760), .A3(n4987), .A4(n8759), .ZN(n8764)
         );
  NOR2_X1 U9885 ( .A1(n8768), .A2(n9470), .ZN(n8770) );
  MUX2_X1 U9886 ( .A(n8770), .B(n5463), .S(n8849), .Z(n8771) );
  NOR2_X1 U9887 ( .A1(n9466), .A2(n8771), .ZN(n8772) );
  NAND2_X1 U9888 ( .A1(n8773), .A2(n8772), .ZN(n8779) );
  NAND2_X1 U9889 ( .A1(n8774), .A2(n8842), .ZN(n8777) );
  OR2_X1 U9890 ( .A1(n8775), .A2(n8842), .ZN(n8776) );
  AND2_X1 U9891 ( .A1(n8777), .A2(n8776), .ZN(n8778) );
  NAND2_X1 U9892 ( .A1(n8779), .A2(n8778), .ZN(n8790) );
  NAND2_X1 U9893 ( .A1(n8790), .A2(n9557), .ZN(n8783) );
  INV_X1 U9894 ( .A(n8780), .ZN(n10841) );
  AND2_X1 U9895 ( .A1(n8784), .A2(n10841), .ZN(n8782) );
  INV_X1 U9896 ( .A(n8786), .ZN(n8781) );
  AOI21_X1 U9897 ( .B1(n8783), .B2(n8782), .A(n8781), .ZN(n8789) );
  NAND2_X1 U9898 ( .A1(n8783), .A2(n9472), .ZN(n8785) );
  NAND2_X1 U9899 ( .A1(n8785), .A2(n8784), .ZN(n8787) );
  NAND2_X1 U9900 ( .A1(n8787), .A2(n8786), .ZN(n8788) );
  MUX2_X1 U9901 ( .A(n8789), .B(n8788), .S(n8849), .Z(n8799) );
  INV_X1 U9902 ( .A(n8790), .ZN(n8793) );
  NOR2_X1 U9903 ( .A1(n9455), .A2(n8791), .ZN(n8792) );
  AOI21_X1 U9904 ( .B1(n8793), .B2(n8792), .A(n9446), .ZN(n8798) );
  MUX2_X1 U9905 ( .A(n8795), .B(n8794), .S(n8842), .Z(n8796) );
  INV_X1 U9906 ( .A(n8796), .ZN(n8797) );
  INV_X1 U9907 ( .A(n9534), .ZN(n8800) );
  MUX2_X1 U9908 ( .A(n9060), .B(n8800), .S(n8842), .Z(n8805) );
  NAND2_X1 U9909 ( .A1(n8808), .A2(n8800), .ZN(n8802) );
  NAND2_X1 U9910 ( .A1(n8807), .A2(n9060), .ZN(n8801) );
  MUX2_X1 U9911 ( .A(n8802), .B(n8801), .S(n8842), .Z(n8803) );
  AOI21_X1 U9912 ( .B1(n8804), .B2(n8805), .A(n8803), .ZN(n8814) );
  INV_X1 U9913 ( .A(n8805), .ZN(n8806) );
  MUX2_X1 U9914 ( .A(n8808), .B(n8807), .S(n8849), .Z(n8809) );
  MUX2_X1 U9915 ( .A(n8811), .B(n8810), .S(n8842), .Z(n8812) );
  OAI211_X1 U9916 ( .C1(n8814), .C2(n8813), .A(n9388), .B(n8812), .ZN(n8818)
         );
  MUX2_X1 U9917 ( .A(n8816), .B(n8815), .S(n8849), .Z(n8817) );
  OAI211_X1 U9918 ( .C1(n8820), .C2(n8819), .A(n8818), .B(n8817), .ZN(n8821)
         );
  OAI211_X1 U9919 ( .C1(n8823), .C2(n8822), .A(n9355), .B(n8821), .ZN(n8827)
         );
  NAND2_X1 U9920 ( .A1(n9101), .A2(n9373), .ZN(n8825) );
  MUX2_X1 U9921 ( .A(n8825), .B(n8824), .S(n8849), .Z(n8826) );
  AOI21_X1 U9922 ( .B1(n8827), .B2(n8826), .A(n9340), .ZN(n8830) );
  MUX2_X1 U9923 ( .A(n8828), .B(n5505), .S(n8842), .Z(n8829) );
  MUX2_X1 U9924 ( .A(n8832), .B(n8831), .S(n8849), .Z(n8834) );
  MUX2_X1 U9925 ( .A(n8837), .B(n8836), .S(n8849), .Z(n8838) );
  MUX2_X1 U9926 ( .A(n8840), .B(n8839), .S(n8842), .Z(n8841) );
  INV_X1 U9927 ( .A(n8845), .ZN(n8848) );
  MUX2_X1 U9928 ( .A(n9136), .B(n9483), .S(n8842), .Z(n8847) );
  INV_X1 U9929 ( .A(n8847), .ZN(n8844) );
  MUX2_X1 U9930 ( .A(n9136), .B(n9483), .S(n8849), .Z(n8843) );
  OAI21_X1 U9931 ( .B1(n8845), .B2(n8844), .A(n8843), .ZN(n8846) );
  OAI21_X1 U9932 ( .B1(n8848), .B2(n8847), .A(n8846), .ZN(n8850) );
  INV_X1 U9933 ( .A(n8855), .ZN(n8857) );
  MUX2_X1 U9934 ( .A(n8860), .B(n8859), .S(n8858), .Z(n8861) );
  AOI21_X1 U9935 ( .B1(n8863), .B2(n8862), .A(n8861), .ZN(n8871) );
  NOR3_X1 U9936 ( .A1(n8866), .A2(n8865), .A3(n8864), .ZN(n8869) );
  OAI21_X1 U9937 ( .B1(n8870), .B2(n8867), .A(P2_B_REG_SCAN_IN), .ZN(n8868) );
  OAI22_X1 U9938 ( .A1(n8871), .A2(n8870), .B1(n8869), .B2(n8868), .ZN(
        P2_U3296) );
  INV_X1 U9939 ( .A(n8872), .ZN(n8875) );
  INV_X1 U9940 ( .A(n8873), .ZN(n8874) );
  AOI22_X1 U9941 ( .A1(n9649), .A2(n8977), .B1(n8916), .B2(n9794), .ZN(n8876)
         );
  XNOR2_X1 U9942 ( .A(n8876), .B(n8963), .ZN(n8878) );
  OAI22_X1 U9943 ( .A1(n8877), .A2(n8903), .B1(n9782), .B2(n8902), .ZN(n9642)
         );
  NAND2_X1 U9944 ( .A1(n8879), .A2(n8878), .ZN(n9639) );
  AOI22_X1 U9945 ( .A1(n9786), .A2(n8916), .B1(n7254), .B2(n10165), .ZN(n9774)
         );
  AOI22_X1 U9946 ( .A1(n9786), .A2(n8977), .B1(n8916), .B2(n10165), .ZN(n8880)
         );
  XNOR2_X1 U9947 ( .A(n8880), .B(n8963), .ZN(n9775) );
  NAND2_X1 U9948 ( .A1(n10176), .A2(n8977), .ZN(n8882) );
  NAND2_X1 U9949 ( .A1(n9793), .A2(n8965), .ZN(n8881) );
  NAND2_X1 U9950 ( .A1(n8882), .A2(n8881), .ZN(n8884) );
  XNOR2_X1 U9951 ( .A(n8884), .B(n8883), .ZN(n8887) );
  INV_X1 U9952 ( .A(n8887), .ZN(n8889) );
  NOR2_X1 U9953 ( .A1(n10278), .A2(n8902), .ZN(n8885) );
  AOI21_X1 U9954 ( .B1(n10176), .B2(n8965), .A(n8885), .ZN(n8886) );
  INV_X1 U9955 ( .A(n8886), .ZN(n8888) );
  AOI21_X1 U9956 ( .B1(n8889), .B2(n8888), .A(n8890), .ZN(n9693) );
  INV_X1 U9957 ( .A(n8890), .ZN(n8891) );
  NAND2_X1 U9958 ( .A1(n10282), .A2(n8977), .ZN(n8893) );
  NAND2_X1 U9959 ( .A1(n10266), .A2(n8965), .ZN(n8892) );
  NAND2_X1 U9960 ( .A1(n8893), .A2(n8892), .ZN(n8894) );
  XNOR2_X1 U9961 ( .A(n8894), .B(n8963), .ZN(n8897) );
  NAND2_X1 U9962 ( .A1(n10282), .A2(n8965), .ZN(n8896) );
  NAND2_X1 U9963 ( .A1(n7254), .A2(n10266), .ZN(n8895) );
  NAND2_X1 U9964 ( .A1(n8896), .A2(n8895), .ZN(n8898) );
  NAND2_X1 U9965 ( .A1(n8897), .A2(n8898), .ZN(n9702) );
  INV_X1 U9966 ( .A(n8897), .ZN(n8900) );
  INV_X1 U9967 ( .A(n8898), .ZN(n8899) );
  NAND2_X1 U9968 ( .A1(n8900), .A2(n8899), .ZN(n9704) );
  NAND2_X1 U9969 ( .A1(n9700), .A2(n9704), .ZN(n8905) );
  AOI22_X1 U9970 ( .A1(n10143), .A2(n8977), .B1(n8916), .B2(n10257), .ZN(n8901) );
  XNOR2_X1 U9971 ( .A(n8901), .B(n8963), .ZN(n8904) );
  NAND2_X1 U9972 ( .A1(n8905), .A2(n8904), .ZN(n9751) );
  OAI22_X1 U9973 ( .A1(n10331), .A2(n8903), .B1(n10279), .B2(n8902), .ZN(n9754) );
  NAND2_X1 U9974 ( .A1(n10125), .A2(n8977), .ZN(n8907) );
  NAND2_X1 U9975 ( .A1(n10269), .A2(n8965), .ZN(n8906) );
  NAND2_X1 U9976 ( .A1(n8907), .A2(n8906), .ZN(n8908) );
  XNOR2_X1 U9977 ( .A(n8908), .B(n8975), .ZN(n8911) );
  AOI22_X1 U9978 ( .A1(n10125), .A2(n8916), .B1(n7254), .B2(n10269), .ZN(n8909) );
  XNOR2_X1 U9979 ( .A(n8911), .B(n8909), .ZN(n9668) );
  INV_X1 U9980 ( .A(n8909), .ZN(n8910) );
  NAND2_X1 U9981 ( .A1(n9666), .A2(n8912), .ZN(n9733) );
  NAND2_X1 U9982 ( .A1(n10110), .A2(n8977), .ZN(n8914) );
  NAND2_X1 U9983 ( .A1(n10258), .A2(n8965), .ZN(n8913) );
  NAND2_X1 U9984 ( .A1(n8914), .A2(n8913), .ZN(n8915) );
  XNOR2_X1 U9985 ( .A(n8915), .B(n8963), .ZN(n8919) );
  AOI22_X1 U9986 ( .A1(n10110), .A2(n8916), .B1(n7254), .B2(n10258), .ZN(n8917) );
  XNOR2_X1 U9987 ( .A(n8919), .B(n8917), .ZN(n9734) );
  INV_X1 U9988 ( .A(n8917), .ZN(n8918) );
  AOI22_X1 U9989 ( .A1(n10091), .A2(n8977), .B1(n8916), .B2(n10249), .ZN(n8921) );
  XNOR2_X1 U9990 ( .A(n8921), .B(n8975), .ZN(n8922) );
  AOI22_X1 U9991 ( .A1(n10091), .A2(n8916), .B1(n7254), .B2(n10249), .ZN(n8923) );
  XNOR2_X1 U9992 ( .A(n8922), .B(n8923), .ZN(n9673) );
  INV_X1 U9993 ( .A(n8922), .ZN(n8925) );
  INV_X1 U9994 ( .A(n8923), .ZN(n8924) );
  AOI22_X1 U9995 ( .A1(n10232), .A2(n8977), .B1(n8916), .B2(n10236), .ZN(n8926) );
  XOR2_X1 U9996 ( .A(n8963), .B(n8926), .Z(n9656) );
  NAND2_X1 U9997 ( .A1(n10232), .A2(n8965), .ZN(n8928) );
  NAND2_X1 U9998 ( .A1(n10236), .A2(n7254), .ZN(n8927) );
  NAND2_X1 U9999 ( .A1(n8928), .A2(n8927), .ZN(n9655) );
  NAND2_X1 U10000 ( .A1(n10077), .A2(n8965), .ZN(n8930) );
  NAND2_X1 U10001 ( .A1(n10086), .A2(n7254), .ZN(n8929) );
  NAND2_X1 U10002 ( .A1(n8930), .A2(n8929), .ZN(n9744) );
  NAND2_X1 U10003 ( .A1(n10077), .A2(n8977), .ZN(n8932) );
  NAND2_X1 U10004 ( .A1(n10086), .A2(n8965), .ZN(n8931) );
  NAND2_X1 U10005 ( .A1(n8932), .A2(n8931), .ZN(n8933) );
  XNOR2_X1 U10006 ( .A(n8933), .B(n8975), .ZN(n9652) );
  AOI22_X1 U10007 ( .A1(n9656), .A2(n9655), .B1(n9744), .B2(n9652), .ZN(n8934)
         );
  INV_X1 U10008 ( .A(n9656), .ZN(n8937) );
  OAI21_X1 U10009 ( .B1(n9652), .B2(n9744), .A(n9655), .ZN(n8936) );
  NOR3_X1 U10010 ( .A1(n9652), .A2(n9655), .A3(n9744), .ZN(n8935) );
  AOI21_X1 U10011 ( .B1(n8937), .B2(n8936), .A(n8935), .ZN(n8938) );
  NAND2_X1 U10012 ( .A1(n8939), .A2(n8938), .ZN(n9711) );
  NAND2_X1 U10013 ( .A1(n10227), .A2(n8977), .ZN(n8941) );
  NAND2_X1 U10014 ( .A1(n10056), .A2(n8965), .ZN(n8940) );
  NAND2_X1 U10015 ( .A1(n8941), .A2(n8940), .ZN(n8942) );
  XNOR2_X1 U10016 ( .A(n8942), .B(n8975), .ZN(n8945) );
  NAND2_X1 U10017 ( .A1(n10227), .A2(n8965), .ZN(n8944) );
  NAND2_X1 U10018 ( .A1(n10056), .A2(n7254), .ZN(n8943) );
  NAND2_X1 U10019 ( .A1(n8944), .A2(n8943), .ZN(n8946) );
  NAND2_X1 U10020 ( .A1(n8945), .A2(n8946), .ZN(n9712) );
  NAND2_X1 U10021 ( .A1(n9711), .A2(n9712), .ZN(n8949) );
  INV_X1 U10022 ( .A(n8945), .ZN(n8948) );
  INV_X1 U10023 ( .A(n8946), .ZN(n8947) );
  NAND2_X1 U10024 ( .A1(n8948), .A2(n8947), .ZN(n9713) );
  NAND2_X1 U10025 ( .A1(n8949), .A2(n9713), .ZN(n9682) );
  NAND2_X1 U10026 ( .A1(n10220), .A2(n8977), .ZN(n8951) );
  NAND2_X1 U10027 ( .A1(n10005), .A2(n8965), .ZN(n8950) );
  NAND2_X1 U10028 ( .A1(n8951), .A2(n8950), .ZN(n8952) );
  XNOR2_X1 U10029 ( .A(n8952), .B(n8963), .ZN(n8957) );
  AOI22_X1 U10030 ( .A1(n10220), .A2(n8916), .B1(n7254), .B2(n10005), .ZN(
        n8958) );
  XNOR2_X1 U10031 ( .A(n8957), .B(n8958), .ZN(n9684) );
  NAND2_X1 U10032 ( .A1(n9682), .A2(n9684), .ZN(n9683) );
  NAND2_X1 U10033 ( .A1(n10214), .A2(n8977), .ZN(n8954) );
  NAND2_X1 U10034 ( .A1(n10028), .A2(n8965), .ZN(n8953) );
  NAND2_X1 U10035 ( .A1(n8954), .A2(n8953), .ZN(n8955) );
  XNOR2_X1 U10036 ( .A(n8955), .B(n8975), .ZN(n8972) );
  AND2_X1 U10037 ( .A1(n10028), .A2(n7254), .ZN(n8956) );
  AOI21_X1 U10038 ( .B1(n10214), .B2(n8916), .A(n8956), .ZN(n8970) );
  XNOR2_X1 U10039 ( .A(n8972), .B(n8970), .ZN(n9765) );
  INV_X1 U10040 ( .A(n8957), .ZN(n8959) );
  NAND2_X1 U10041 ( .A1(n8959), .A2(n8958), .ZN(n9762) );
  NAND2_X1 U10042 ( .A1(n9990), .A2(n8977), .ZN(n8962) );
  NAND2_X1 U10043 ( .A1(n10004), .A2(n8965), .ZN(n8961) );
  NAND2_X1 U10044 ( .A1(n8962), .A2(n8961), .ZN(n8964) );
  XNOR2_X1 U10045 ( .A(n8964), .B(n8963), .ZN(n8969) );
  NAND2_X1 U10046 ( .A1(n9990), .A2(n8965), .ZN(n8967) );
  NAND2_X1 U10047 ( .A1(n7254), .A2(n10004), .ZN(n8966) );
  NAND2_X1 U10048 ( .A1(n8967), .A2(n8966), .ZN(n8968) );
  NOR2_X1 U10049 ( .A1(n8969), .A2(n8968), .ZN(n8973) );
  AOI21_X1 U10050 ( .B1(n8969), .B2(n8968), .A(n8973), .ZN(n9630) );
  INV_X1 U10051 ( .A(n8970), .ZN(n8971) );
  NAND2_X1 U10052 ( .A1(n8972), .A2(n8971), .ZN(n9631) );
  INV_X1 U10053 ( .A(n8973), .ZN(n8974) );
  AOI22_X1 U10054 ( .A1(n9983), .A2(n8916), .B1(n7254), .B2(n9792), .ZN(n8976)
         );
  XNOR2_X1 U10055 ( .A(n8976), .B(n8975), .ZN(n8979) );
  AOI22_X1 U10056 ( .A1(n9983), .A2(n8977), .B1(n8916), .B2(n9792), .ZN(n8978)
         );
  XNOR2_X1 U10057 ( .A(n8979), .B(n8978), .ZN(n8980) );
  XNOR2_X1 U10058 ( .A(n8981), .B(n8980), .ZN(n8987) );
  OAI22_X1 U10059 ( .A1(n9783), .A2(n8983), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8982), .ZN(n8985) );
  OAI22_X1 U10060 ( .A1(n9779), .A2(n9979), .B1(n9781), .B2(n9976), .ZN(n8984)
         );
  AOI211_X1 U10061 ( .C1(n9983), .C2(n4944), .A(n8985), .B(n8984), .ZN(n8986)
         );
  OAI21_X1 U10062 ( .B1(n8987), .B2(n9788), .A(n8986), .ZN(P1_U3220) );
  OAI222_X1 U10063 ( .A1(n6135), .A2(P1_U3086), .B1(n10354), .B2(n8989), .C1(
        n8988), .C2(n10350), .ZN(P1_U3333) );
  INV_X1 U10064 ( .A(n8990), .ZN(n9618) );
  OAI222_X1 U10065 ( .A1(n10350), .A2(n8992), .B1(n10354), .B2(n9618), .C1(
        P1_U3086), .C2(n8991), .ZN(P1_U3325) );
  INV_X1 U10066 ( .A(n8993), .ZN(n9626) );
  OAI222_X1 U10067 ( .A1(P1_U3086), .A2(n8995), .B1(n10354), .B2(n9626), .C1(
        n8994), .C2(n10350), .ZN(P1_U3327) );
  INV_X1 U10068 ( .A(n9298), .ZN(n9000) );
  AOI22_X1 U10069 ( .A1(n9081), .A2(n9136), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8999) );
  OAI21_X1 U10070 ( .B1(n9000), .B2(n9006), .A(n8999), .ZN(n9001) );
  AOI21_X1 U10071 ( .B1(n9126), .B2(n9137), .A(n9001), .ZN(n9002) );
  INV_X1 U10072 ( .A(n9503), .ZN(n9011) );
  OAI21_X1 U10073 ( .B1(n9330), .B2(n4964), .A(n9070), .ZN(n9004) );
  NAND2_X1 U10074 ( .A1(n9004), .A2(n9091), .ZN(n9010) );
  INV_X1 U10075 ( .A(n9342), .ZN(n9007) );
  AOI22_X1 U10076 ( .A1(n9338), .A2(n9126), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n9005) );
  OAI21_X1 U10077 ( .B1(n9007), .B2(n9006), .A(n9005), .ZN(n9008) );
  AOI21_X1 U10078 ( .B1(n5509), .B2(n9081), .A(n9008), .ZN(n9009) );
  OAI211_X1 U10079 ( .C1(n9011), .C2(n9114), .A(n9010), .B(n9009), .ZN(
        P2_U3156) );
  AOI21_X1 U10080 ( .B1(n9012), .B2(n9013), .A(n9133), .ZN(n9015) );
  NAND2_X1 U10081 ( .A1(n9015), .A2(n9014), .ZN(n9021) );
  AOI21_X1 U10082 ( .B1(n9126), .B2(n9150), .A(n9016), .ZN(n9020) );
  AOI22_X1 U10083 ( .A1(n9017), .A2(n9131), .B1(n9081), .B2(n9148), .ZN(n9019)
         );
  NAND2_X1 U10084 ( .A1(n9125), .A2(n10466), .ZN(n9018) );
  NAND4_X1 U10085 ( .A1(n9021), .A2(n9020), .A3(n9019), .A4(n9018), .ZN(
        P2_U3158) );
  XOR2_X1 U10086 ( .A(n9023), .B(n9022), .Z(n9028) );
  INV_X1 U10087 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10468) );
  NOR2_X1 U10088 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10468), .ZN(n9265) );
  AOI21_X1 U10089 ( .B1(n9037), .B2(n9081), .A(n9265), .ZN(n9025) );
  NAND2_X1 U10090 ( .A1(n9125), .A2(n9408), .ZN(n9024) );
  OAI211_X1 U10091 ( .C1(n9406), .C2(n9094), .A(n9025), .B(n9024), .ZN(n9026)
         );
  AOI21_X1 U10092 ( .B1(n9523), .B2(n9131), .A(n9026), .ZN(n9027) );
  OAI21_X1 U10093 ( .B1(n9028), .B2(n9133), .A(n9027), .ZN(P2_U3159) );
  INV_X1 U10094 ( .A(n9375), .ZN(n9601) );
  INV_X1 U10095 ( .A(n4952), .ZN(n9033) );
  INV_X1 U10096 ( .A(n9030), .ZN(n9032) );
  NOR3_X1 U10097 ( .A1(n9033), .A2(n9032), .A3(n9031), .ZN(n9036) );
  INV_X1 U10098 ( .A(n9034), .ZN(n9035) );
  OAI21_X1 U10099 ( .B1(n9036), .B2(n9035), .A(n9091), .ZN(n9041) );
  AOI22_X1 U10100 ( .A1(n9037), .A2(n9126), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n9038) );
  OAI21_X1 U10101 ( .B1(n9373), .B2(n9129), .A(n9038), .ZN(n9039) );
  AOI21_X1 U10102 ( .B1(n9374), .B2(n9125), .A(n9039), .ZN(n9040) );
  OAI211_X1 U10103 ( .C1(n9601), .C2(n9114), .A(n9041), .B(n9040), .ZN(
        P2_U3163) );
  INV_X1 U10104 ( .A(n9042), .ZN(n9046) );
  NOR3_X1 U10105 ( .A1(n9072), .A2(n9044), .A3(n9043), .ZN(n9045) );
  OAI21_X1 U10106 ( .B1(n9046), .B2(n9045), .A(n9091), .ZN(n9050) );
  AOI22_X1 U10107 ( .A1(n9320), .A2(n9125), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n9047) );
  OAI21_X1 U10108 ( .B1(n9316), .B2(n9094), .A(n9047), .ZN(n9048) );
  AOI21_X1 U10109 ( .B1(n9081), .B2(n9137), .A(n9048), .ZN(n9049) );
  OAI211_X1 U10110 ( .C1(n9589), .C2(n9114), .A(n9050), .B(n9049), .ZN(
        P2_U3165) );
  XNOR2_X1 U10111 ( .A(n9051), .B(n9458), .ZN(n9052) );
  XNOR2_X1 U10112 ( .A(n9053), .B(n9052), .ZN(n9058) );
  NAND2_X1 U10113 ( .A1(n9081), .A2(n9440), .ZN(n9054) );
  NAND2_X1 U10114 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3151), .ZN(n9211) );
  OAI211_X1 U10115 ( .C1(n10576), .C2(n9094), .A(n9054), .B(n9211), .ZN(n9055)
         );
  AOI21_X1 U10116 ( .B1(n9442), .B2(n9125), .A(n9055), .ZN(n9057) );
  NAND2_X1 U10117 ( .A1(n9538), .A2(n9131), .ZN(n9056) );
  OAI211_X1 U10118 ( .C1(n9058), .C2(n9133), .A(n9057), .B(n9056), .ZN(
        P2_U3166) );
  XNOR2_X1 U10119 ( .A(n9061), .B(n9060), .ZN(n9062) );
  XNOR2_X1 U10120 ( .A(n9059), .B(n9062), .ZN(n9067) );
  NAND2_X1 U10121 ( .A1(n9125), .A2(n9430), .ZN(n9064) );
  NOR2_X1 U10122 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10457), .ZN(n9238) );
  AOI21_X1 U10123 ( .B1(n9126), .B2(n9428), .A(n9238), .ZN(n9063) );
  OAI211_X1 U10124 ( .C1(n9406), .C2(n9129), .A(n9064), .B(n9063), .ZN(n9065)
         );
  AOI21_X1 U10125 ( .B1(n9534), .B2(n9131), .A(n9065), .ZN(n9066) );
  OAI21_X1 U10126 ( .B1(n9067), .B2(n9133), .A(n9066), .ZN(P2_U3168) );
  AND3_X1 U10127 ( .A1(n9070), .A2(n9069), .A3(n9068), .ZN(n9071) );
  OAI21_X1 U10128 ( .B1(n9072), .B2(n9071), .A(n9091), .ZN(n9076) );
  INV_X1 U10129 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10460) );
  OAI22_X1 U10130 ( .A1(n9330), .A2(n9094), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10460), .ZN(n9074) );
  NOR2_X1 U10131 ( .A1(n9329), .A2(n9129), .ZN(n9073) );
  AOI211_X1 U10132 ( .C1(n9332), .C2(n9125), .A(n9074), .B(n9073), .ZN(n9075)
         );
  OAI211_X1 U10133 ( .C1(n5510), .C2(n9114), .A(n9076), .B(n9075), .ZN(
        P2_U3169) );
  NAND2_X1 U10134 ( .A1(n9079), .A2(n9091), .ZN(n9088) );
  AOI21_X1 U10135 ( .B1(n9081), .B2(n9147), .A(n9080), .ZN(n9087) );
  AOI22_X1 U10136 ( .A1(n9082), .A2(n9131), .B1(n9126), .B2(n9149), .ZN(n9086)
         );
  INV_X1 U10137 ( .A(n9083), .ZN(n9084) );
  NAND2_X1 U10138 ( .A1(n9125), .A2(n9084), .ZN(n9085) );
  NAND4_X1 U10139 ( .A1(n9088), .A2(n9087), .A3(n9086), .A4(n9085), .ZN(
        P2_U3170) );
  OAI21_X1 U10140 ( .B1(n9090), .B2(n9089), .A(n4952), .ZN(n9092) );
  NAND2_X1 U10141 ( .A1(n9092), .A2(n9091), .ZN(n9099) );
  OAI22_X1 U10142 ( .A1(n9113), .A2(n9094), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9093), .ZN(n9097) );
  NOR2_X1 U10143 ( .A1(n9095), .A2(n9129), .ZN(n9096) );
  AOI211_X1 U10144 ( .C1(n9384), .C2(n9125), .A(n9097), .B(n9096), .ZN(n9098)
         );
  OAI211_X1 U10145 ( .C1(n9100), .C2(n9114), .A(n9099), .B(n9098), .ZN(
        P2_U3173) );
  INV_X1 U10146 ( .A(n9101), .ZN(n9597) );
  AOI21_X1 U10147 ( .B1(n9103), .B2(n9102), .A(n9133), .ZN(n9105) );
  NAND2_X1 U10148 ( .A1(n9105), .A2(n9104), .ZN(n9109) );
  AOI22_X1 U10149 ( .A1(n9391), .A2(n9126), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n9106) );
  OAI21_X1 U10150 ( .B1(n9330), .B2(n9129), .A(n9106), .ZN(n9107) );
  AOI21_X1 U10151 ( .B1(n9358), .B2(n9125), .A(n9107), .ZN(n9108) );
  OAI211_X1 U10152 ( .C1(n9597), .C2(n9114), .A(n9109), .B(n9108), .ZN(
        P2_U3175) );
  XNOR2_X1 U10153 ( .A(n9110), .B(n9111), .ZN(n9119) );
  NAND2_X1 U10154 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3151), .ZN(n10717)
         );
  NAND2_X1 U10155 ( .A1(n9126), .A2(n9440), .ZN(n9112) );
  OAI211_X1 U10156 ( .C1(n9113), .C2(n9129), .A(n10717), .B(n9112), .ZN(n9117)
         );
  NOR2_X1 U10157 ( .A1(n9115), .A2(n9114), .ZN(n9116) );
  AOI211_X1 U10158 ( .C1(n9417), .C2(n9125), .A(n9117), .B(n9116), .ZN(n9118)
         );
  OAI21_X1 U10159 ( .B1(n9119), .B2(n9133), .A(n9118), .ZN(P2_U3178) );
  INV_X1 U10160 ( .A(n9120), .ZN(n9122) );
  NAND2_X1 U10161 ( .A1(n9122), .A2(n9121), .ZN(n9123) );
  XNOR2_X1 U10162 ( .A(n9124), .B(n9123), .ZN(n9134) );
  AOI22_X1 U10163 ( .A1(n9309), .A2(n9125), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n9128) );
  NAND2_X1 U10164 ( .A1(n9138), .A2(n9126), .ZN(n9127) );
  OAI211_X1 U10165 ( .C1(n9305), .C2(n9129), .A(n9128), .B(n9127), .ZN(n9130)
         );
  AOI21_X1 U10166 ( .B1(n9308), .B2(n9131), .A(n9130), .ZN(n9132) );
  OAI21_X1 U10167 ( .B1(n9134), .B2(n9133), .A(n9132), .ZN(P2_U3180) );
  MUX2_X1 U10168 ( .A(n9275), .B(P2_DATAO_REG_31__SCAN_IN), .S(n10574), .Z(
        P2_U3522) );
  MUX2_X1 U10169 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n9135), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10170 ( .A(n9282), .B(P2_DATAO_REG_29__SCAN_IN), .S(n10574), .Z(
        P2_U3520) );
  MUX2_X1 U10171 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n9136), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10172 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n9137), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10173 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9138), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10174 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n5509), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10175 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9338), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10176 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9391), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10177 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9415), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10178 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9427), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10179 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9440), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10180 ( .A(n9428), .B(P2_DATAO_REG_16__SCAN_IN), .S(n10574), .Z(
        P2_U3507) );
  MUX2_X1 U10181 ( .A(n9139), .B(P2_DATAO_REG_14__SCAN_IN), .S(n10574), .Z(
        P2_U3505) );
  MUX2_X1 U10182 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n9554), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10183 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n9140), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U10184 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n9141), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10185 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n9142), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10186 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n9143), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10187 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n9144), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U10188 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n9145), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U10189 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n9146), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U10190 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n9147), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U10191 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n9148), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10192 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n9149), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U10193 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n9150), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U10194 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n9151), .S(P2_U3893), .Z(
        P2_U3492) );
  NOR2_X1 U10195 ( .A1(n9167), .A2(n9152), .ZN(n9154) );
  AOI22_X1 U10196 ( .A1(n9170), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n6445), .B2(
        n9191), .ZN(n9155) );
  AOI21_X1 U10197 ( .B1(n9156), .B2(n9155), .A(n9180), .ZN(n9178) );
  MUX2_X1 U10198 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n4947), .Z(n9185) );
  XNOR2_X1 U10199 ( .A(n9185), .B(n9170), .ZN(n9162) );
  OR2_X1 U10200 ( .A1(n9158), .A2(n9157), .ZN(n9160) );
  NAND2_X1 U10201 ( .A1(n9160), .A2(n9159), .ZN(n9161) );
  NAND2_X1 U10202 ( .A1(n9162), .A2(n9161), .ZN(n9186) );
  OAI21_X1 U10203 ( .B1(n9162), .B2(n9161), .A(n9186), .ZN(n9176) );
  INV_X1 U10204 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9165) );
  NAND2_X1 U10205 ( .A1(n10676), .A2(n9170), .ZN(n9164) );
  OAI211_X1 U10206 ( .C1(n9165), .C2(n9263), .A(n9164), .B(n9163), .ZN(n9175)
         );
  NOR2_X1 U10207 ( .A1(n9167), .A2(n9166), .ZN(n9169) );
  MUX2_X1 U10208 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n9171), .S(n9170), .Z(n9172) );
  AOI21_X1 U10209 ( .B1(n4997), .B2(n9172), .A(n9190), .ZN(n9173) );
  NOR2_X1 U10210 ( .A1(n9173), .A2(n10682), .ZN(n9174) );
  AOI211_X1 U10211 ( .C1(n10690), .C2(n9176), .A(n9175), .B(n9174), .ZN(n9177)
         );
  OAI21_X1 U10212 ( .B1(n9178), .B2(n10713), .A(n9177), .ZN(P2_U3196) );
  NOR2_X1 U10213 ( .A1(n9170), .A2(n6445), .ZN(n9179) );
  AOI21_X1 U10214 ( .B1(n6461), .B2(n9181), .A(n9201), .ZN(n9198) );
  INV_X1 U10215 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9182) );
  NOR2_X1 U10216 ( .A1(n9263), .A2(n9182), .ZN(n9183) );
  AOI211_X1 U10217 ( .C1(n10676), .C2(n9213), .A(n9184), .B(n9183), .ZN(n9197)
         );
  MUX2_X1 U10218 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n4946), .Z(n9205) );
  XNOR2_X1 U10219 ( .A(n9213), .B(n9205), .ZN(n9189) );
  OR2_X1 U10220 ( .A1(n9185), .A2(n9191), .ZN(n9187) );
  NAND2_X1 U10221 ( .A1(n9187), .A2(n9186), .ZN(n9188) );
  NAND2_X1 U10222 ( .A1(n9189), .A2(n9188), .ZN(n9204) );
  OAI21_X1 U10223 ( .B1(n9189), .B2(n9188), .A(n9204), .ZN(n9195) );
  AOI21_X1 U10224 ( .B1(n9192), .B2(n9461), .A(n9214), .ZN(n9193) );
  NOR2_X1 U10225 ( .A1(n9193), .A2(n10682), .ZN(n9194) );
  AOI21_X1 U10226 ( .B1(n10690), .B2(n9195), .A(n9194), .ZN(n9196) );
  OAI211_X1 U10227 ( .C1(n9198), .C2(n10713), .A(n9197), .B(n9196), .ZN(
        P2_U3197) );
  NOR2_X1 U10228 ( .A1(n9213), .A2(n9199), .ZN(n9200) );
  AOI22_X1 U10229 ( .A1(n9207), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n9202), .B2(
        n9233), .ZN(n9203) );
  AOI21_X1 U10230 ( .B1(n4998), .B2(n9203), .A(n9224), .ZN(n9223) );
  OAI21_X1 U10231 ( .B1(n9206), .B2(n9205), .A(n9204), .ZN(n9209) );
  MUX2_X1 U10232 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n4947), .Z(n9227) );
  XNOR2_X1 U10233 ( .A(n9207), .B(n9227), .ZN(n9208) );
  NAND2_X1 U10234 ( .A1(n9208), .A2(n9209), .ZN(n9228) );
  OAI21_X1 U10235 ( .B1(n9209), .B2(n9208), .A(n9228), .ZN(n9221) );
  NAND2_X1 U10236 ( .A1(n10698), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n9210) );
  OAI211_X1 U10237 ( .C1(n10706), .C2(n9233), .A(n9211), .B(n9210), .ZN(n9220)
         );
  NOR2_X1 U10238 ( .A1(n9213), .A2(n9212), .ZN(n9215) );
  NAND2_X1 U10239 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n9233), .ZN(n9216) );
  OAI21_X1 U10240 ( .B1(n9233), .B2(P2_REG2_REG_16__SCAN_IN), .A(n9216), .ZN(
        n9217) );
  AOI21_X1 U10241 ( .B1(n4999), .B2(n9217), .A(n9232), .ZN(n9218) );
  NOR2_X1 U10242 ( .A1(n9218), .A2(n10682), .ZN(n9219) );
  AOI211_X1 U10243 ( .C1(n10690), .C2(n9221), .A(n9220), .B(n9219), .ZN(n9222)
         );
  OAI21_X1 U10244 ( .B1(n9223), .B2(n10713), .A(n9222), .ZN(P2_U3198) );
  AOI21_X1 U10245 ( .B1(n9226), .B2(n9225), .A(n9247), .ZN(n9244) );
  MUX2_X1 U10246 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n4946), .Z(n9255) );
  XNOR2_X1 U10247 ( .A(n9246), .B(n9255), .ZN(n9231) );
  OR2_X1 U10248 ( .A1(n9227), .A2(n9233), .ZN(n9229) );
  NAND2_X1 U10249 ( .A1(n9229), .A2(n9228), .ZN(n9230) );
  NAND2_X1 U10250 ( .A1(n9231), .A2(n9230), .ZN(n9254) );
  OAI21_X1 U10251 ( .B1(n9231), .B2(n9230), .A(n9254), .ZN(n9242) );
  AOI21_X1 U10252 ( .B1(n9235), .B2(n9432), .A(n10699), .ZN(n9240) );
  INV_X1 U10253 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9236) );
  NOR2_X1 U10254 ( .A1(n9263), .A2(n9236), .ZN(n9237) );
  AOI211_X1 U10255 ( .C1(n10676), .C2(n9246), .A(n9238), .B(n9237), .ZN(n9239)
         );
  OAI21_X1 U10256 ( .B1(n9240), .B2(n10682), .A(n9239), .ZN(n9241) );
  AOI21_X1 U10257 ( .B1(n10690), .B2(n9242), .A(n9241), .ZN(n9243) );
  OAI21_X1 U10258 ( .B1(n9244), .B2(n10713), .A(n9243), .ZN(P2_U3199) );
  NAND2_X1 U10259 ( .A1(n10705), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9249) );
  OAI21_X1 U10260 ( .B1(n10705), .B2(P2_REG1_REG_18__SCAN_IN), .A(n9249), .ZN(
        n10711) );
  INV_X1 U10261 ( .A(n9249), .ZN(n9250) );
  NOR2_X1 U10262 ( .A1(n10715), .A2(n9250), .ZN(n9251) );
  XNOR2_X1 U10263 ( .A(n9266), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9252) );
  XNOR2_X1 U10264 ( .A(n9251), .B(n9252), .ZN(n9272) );
  MUX2_X1 U10265 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n9410), .S(n9266), .Z(n9262) );
  INV_X1 U10266 ( .A(n9252), .ZN(n9253) );
  MUX2_X1 U10267 ( .A(n9262), .B(n9253), .S(n4946), .Z(n9261) );
  OAI21_X1 U10268 ( .B1(n5210), .B2(n9255), .A(n9254), .ZN(n9259) );
  INV_X1 U10269 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9419) );
  MUX2_X1 U10270 ( .A(n9419), .B(n9257), .S(n4947), .Z(n9258) );
  NAND2_X1 U10271 ( .A1(n9259), .A2(n9258), .ZN(n10703) );
  NOR2_X1 U10272 ( .A1(n9259), .A2(n9258), .ZN(n10694) );
  AOI21_X1 U10273 ( .B1(n10705), .B2(n10703), .A(n10694), .ZN(n9260) );
  XOR2_X1 U10274 ( .A(n9261), .B(n9260), .Z(n9270) );
  XOR2_X1 U10275 ( .A(P2_REG2_REG_18__SCAN_IN), .B(n10705), .Z(n10701) );
  NOR2_X1 U10276 ( .A1(n9263), .A2(n5345), .ZN(n9264) );
  AOI211_X1 U10277 ( .C1(n10676), .C2(n9266), .A(n9265), .B(n9264), .ZN(n9267)
         );
  OAI21_X1 U10278 ( .B1(n9268), .B2(n10682), .A(n9267), .ZN(n9269) );
  AOI21_X1 U10279 ( .B1(n9270), .B2(n10690), .A(n9269), .ZN(n9271) );
  OAI21_X1 U10280 ( .B1(n9272), .B2(n10713), .A(n9271), .ZN(P2_U3201) );
  NOR2_X1 U10281 ( .A1(n4949), .A2(n9273), .ZN(n9276) );
  NAND2_X1 U10282 ( .A1(n9275), .A2(n9274), .ZN(n9571) );
  NAND2_X1 U10283 ( .A1(n9276), .A2(n9571), .ZN(n9279) );
  OAI21_X1 U10284 ( .B1(n10846), .B2(P2_REG2_REG_31__SCAN_IN), .A(n9279), .ZN(
        n9277) );
  OAI21_X1 U10285 ( .B1(n9573), .B2(n9360), .A(n9277), .ZN(P2_U3202) );
  OAI21_X1 U10286 ( .B1(n10846), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9279), .ZN(
        n9280) );
  OAI21_X1 U10287 ( .B1(n9576), .B2(n9360), .A(n9280), .ZN(P2_U3203) );
  XNOR2_X1 U10288 ( .A(n9281), .B(n9285), .ZN(n9284) );
  XNOR2_X1 U10289 ( .A(n9286), .B(n9285), .ZN(n9484) );
  NOR2_X1 U10290 ( .A1(n9287), .A2(n9360), .ZN(n9291) );
  OAI22_X1 U10291 ( .A1(n10846), .A2(n9289), .B1(n9288), .B2(n10838), .ZN(
        n9290) );
  AOI211_X1 U10292 ( .C1(n9484), .C2(n9377), .A(n9291), .B(n9290), .ZN(n9292)
         );
  OAI21_X1 U10293 ( .B1(n9486), .B2(n4949), .A(n9292), .ZN(P2_U3205) );
  OAI222_X1 U10294 ( .A1(n9471), .A2(n9317), .B1(n9473), .B2(n9295), .C1(n9294), .C2(n9468), .ZN(n9487) );
  INV_X1 U10295 ( .A(n9487), .ZN(n9302) );
  XNOR2_X1 U10296 ( .A(n9297), .B(n9296), .ZN(n9488) );
  AOI22_X1 U10297 ( .A1(n9298), .A2(n10770), .B1(n4949), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n9299) );
  OAI21_X1 U10298 ( .B1(n9581), .B2(n9360), .A(n9299), .ZN(n9300) );
  AOI21_X1 U10299 ( .B1(n9488), .B2(n9377), .A(n9300), .ZN(n9301) );
  OAI21_X1 U10300 ( .B1(n9302), .B2(n4949), .A(n9301), .ZN(P2_U3206) );
  XNOR2_X1 U10301 ( .A(n9303), .B(n9306), .ZN(n9304) );
  OAI222_X1 U10302 ( .A1(n9473), .A2(n9305), .B1(n9471), .B2(n9329), .C1(n9468), .C2(n9304), .ZN(n9491) );
  INV_X1 U10303 ( .A(n9491), .ZN(n9313) );
  XNOR2_X1 U10304 ( .A(n9307), .B(n9306), .ZN(n9492) );
  INV_X1 U10305 ( .A(n9308), .ZN(n9585) );
  AOI22_X1 U10306 ( .A1(n9309), .A2(n10770), .B1(n4949), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n9310) );
  OAI21_X1 U10307 ( .B1(n9585), .B2(n9360), .A(n9310), .ZN(n9311) );
  AOI21_X1 U10308 ( .B1(n9492), .B2(n9377), .A(n9311), .ZN(n9312) );
  OAI21_X1 U10309 ( .B1(n9313), .B2(n4949), .A(n9312), .ZN(P2_U3207) );
  INV_X1 U10310 ( .A(n10840), .ZN(n9319) );
  XNOR2_X1 U10311 ( .A(n9314), .B(n9321), .ZN(n9315) );
  OAI222_X1 U10312 ( .A1(n9473), .A2(n9317), .B1(n9471), .B2(n9316), .C1(n9315), .C2(n9468), .ZN(n9495) );
  AOI21_X1 U10313 ( .B1(n9319), .B2(n9318), .A(n9495), .ZN(n9325) );
  AOI22_X1 U10314 ( .A1(n9320), .A2(n10770), .B1(n4949), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n9324) );
  XNOR2_X1 U10315 ( .A(n9322), .B(n9321), .ZN(n9496) );
  NAND2_X1 U10316 ( .A1(n9496), .A2(n9377), .ZN(n9323) );
  OAI211_X1 U10317 ( .C1(n9325), .C2(n4949), .A(n9324), .B(n9323), .ZN(
        P2_U3208) );
  NOR2_X1 U10318 ( .A1(n5510), .A2(n10840), .ZN(n9331) );
  XNOR2_X1 U10319 ( .A(n9327), .B(n9326), .ZN(n9328) );
  OAI222_X1 U10320 ( .A1(n9471), .A2(n9330), .B1(n9473), .B2(n9329), .C1(n9328), .C2(n9468), .ZN(n9499) );
  AOI211_X1 U10321 ( .C1(n10770), .C2(n9332), .A(n9331), .B(n9499), .ZN(n9336)
         );
  XNOR2_X1 U10322 ( .A(n9334), .B(n9333), .ZN(n9500) );
  AOI22_X1 U10323 ( .A1(n9500), .A2(n9377), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n4949), .ZN(n9335) );
  OAI21_X1 U10324 ( .B1(n9336), .B2(n4949), .A(n9335), .ZN(P2_U3209) );
  XNOR2_X1 U10325 ( .A(n9337), .B(n9340), .ZN(n9339) );
  AOI222_X1 U10326 ( .A1(n9547), .A2(n9339), .B1(n5509), .B2(n9552), .C1(n9338), .C2(n9553), .ZN(n9506) );
  XNOR2_X1 U10327 ( .A(n9341), .B(n9340), .ZN(n9504) );
  NAND2_X1 U10328 ( .A1(n9503), .A2(n10768), .ZN(n9344) );
  AOI22_X1 U10329 ( .A1(n9342), .A2(n10770), .B1(n4949), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n9343) );
  NAND2_X1 U10330 ( .A1(n9344), .A2(n9343), .ZN(n9345) );
  AOI21_X1 U10331 ( .B1(n9504), .B2(n9377), .A(n9345), .ZN(n9346) );
  OAI21_X1 U10332 ( .B1(n9506), .B2(n4949), .A(n9346), .ZN(P2_U3210) );
  OR2_X1 U10333 ( .A1(n9347), .A2(n9348), .ZN(n9365) );
  NAND2_X1 U10334 ( .A1(n9365), .A2(n9349), .ZN(n9351) );
  OAI21_X1 U10335 ( .B1(n9352), .B2(n9351), .A(n9350), .ZN(n9354) );
  AOI222_X1 U10336 ( .A1(n9547), .A2(n9354), .B1(n9391), .B2(n9553), .C1(n9353), .C2(n9552), .ZN(n9508) );
  NOR2_X1 U10337 ( .A1(n9356), .A2(n9355), .ZN(n9507) );
  NOR2_X1 U10338 ( .A1(n9507), .A2(n9479), .ZN(n9362) );
  AOI22_X1 U10339 ( .A1(n9358), .A2(n10770), .B1(n4949), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n9359) );
  OAI21_X1 U10340 ( .B1(n9597), .B2(n9360), .A(n9359), .ZN(n9361) );
  AOI21_X1 U10341 ( .B1(n9362), .B2(n9357), .A(n9361), .ZN(n9363) );
  OAI21_X1 U10342 ( .B1(n9508), .B2(n4949), .A(n9363), .ZN(P2_U3211) );
  AND2_X1 U10343 ( .A1(n9365), .A2(n9364), .ZN(n9371) );
  OR2_X1 U10344 ( .A1(n9347), .A2(n9366), .ZN(n9368) );
  NAND3_X1 U10345 ( .A1(n9389), .A2(n4982), .A3(n9369), .ZN(n9370) );
  OAI222_X1 U10346 ( .A1(n9473), .A2(n9373), .B1(n9471), .B2(n9407), .C1(n9468), .C2(n9372), .ZN(n9514) );
  AOI21_X1 U10347 ( .B1(n10770), .B2(n9374), .A(n9514), .ZN(n9381) );
  AOI22_X1 U10348 ( .A1(n9375), .A2(n10768), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n4949), .ZN(n9380) );
  NOR2_X1 U10349 ( .A1(n9376), .A2(n4982), .ZN(n9513) );
  INV_X1 U10350 ( .A(n9513), .ZN(n9378) );
  NAND3_X1 U10351 ( .A1(n9378), .A2(n9377), .A3(n9515), .ZN(n9379) );
  OAI211_X1 U10352 ( .C1(n9381), .C2(n4949), .A(n9380), .B(n9379), .ZN(
        P2_U3212) );
  OAI21_X1 U10353 ( .B1(n9383), .B2(n9388), .A(n9382), .ZN(n9522) );
  INV_X1 U10354 ( .A(n9384), .ZN(n9393) );
  OR2_X1 U10355 ( .A1(n9347), .A2(n9385), .ZN(n9387) );
  INV_X1 U10356 ( .A(n9388), .ZN(n9390) );
  OAI21_X1 U10357 ( .B1(n5554), .B2(n9390), .A(n9389), .ZN(n9392) );
  AOI222_X1 U10358 ( .A1(n9547), .A2(n9392), .B1(n9391), .B2(n9552), .C1(n9415), .C2(n9553), .ZN(n9521) );
  OAI21_X1 U10359 ( .B1(n9393), .B2(n10838), .A(n9521), .ZN(n9394) );
  NAND2_X1 U10360 ( .A1(n9394), .A2(n10846), .ZN(n9396) );
  AOI22_X1 U10361 ( .A1(n9519), .A2(n10768), .B1(P2_REG2_REG_20__SCAN_IN), 
        .B2(n4949), .ZN(n9395) );
  OAI211_X1 U10362 ( .C1(n9522), .C2(n9479), .A(n9396), .B(n9395), .ZN(
        P2_U3213) );
  OR2_X1 U10363 ( .A1(n9397), .A2(n9403), .ZN(n9398) );
  AND2_X1 U10364 ( .A1(n9399), .A2(n9398), .ZN(n9526) );
  INV_X1 U10365 ( .A(n9526), .ZN(n9414) );
  OR2_X1 U10366 ( .A1(n9347), .A2(n9400), .ZN(n9402) );
  NAND2_X1 U10367 ( .A1(n9402), .A2(n9401), .ZN(n9404) );
  XNOR2_X1 U10368 ( .A(n9404), .B(n9403), .ZN(n9405) );
  OAI222_X1 U10369 ( .A1(n9473), .A2(n9407), .B1(n9471), .B2(n9406), .C1(n9468), .C2(n9405), .ZN(n9524) );
  NAND2_X1 U10370 ( .A1(n9524), .A2(n10846), .ZN(n9413) );
  INV_X1 U10371 ( .A(n9408), .ZN(n9409) );
  OAI22_X1 U10372 ( .A1(n10846), .A2(n9410), .B1(n9409), .B2(n10838), .ZN(
        n9411) );
  AOI21_X1 U10373 ( .B1(n9523), .B2(n10768), .A(n9411), .ZN(n9412) );
  OAI211_X1 U10374 ( .C1(n9414), .C2(n9479), .A(n9413), .B(n9412), .ZN(
        P2_U3214) );
  XNOR2_X1 U10375 ( .A(n9347), .B(n9421), .ZN(n9416) );
  AOI222_X1 U10376 ( .A1(n9547), .A2(n9416), .B1(n9415), .B2(n9552), .C1(n9440), .C2(n9553), .ZN(n9532) );
  INV_X1 U10377 ( .A(n9417), .ZN(n9418) );
  OAI22_X1 U10378 ( .A1(n10846), .A2(n9419), .B1(n9418), .B2(n10838), .ZN(
        n9424) );
  OAI21_X1 U10379 ( .B1(n9422), .B2(n9421), .A(n9420), .ZN(n9533) );
  NOR2_X1 U10380 ( .A1(n9533), .A2(n9479), .ZN(n9423) );
  AOI211_X1 U10381 ( .C1(n10768), .C2(n9530), .A(n9424), .B(n9423), .ZN(n9425)
         );
  OAI21_X1 U10382 ( .B1(n9532), .B2(n4949), .A(n9425), .ZN(P2_U3215) );
  XNOR2_X1 U10383 ( .A(n9426), .B(n9434), .ZN(n9429) );
  AOI222_X1 U10384 ( .A1(n9547), .A2(n9429), .B1(n9428), .B2(n9553), .C1(n9427), .C2(n9552), .ZN(n9536) );
  INV_X1 U10385 ( .A(n9430), .ZN(n9431) );
  OAI22_X1 U10386 ( .A1(n10846), .A2(n9432), .B1(n9431), .B2(n10838), .ZN(
        n9437) );
  OAI21_X1 U10387 ( .B1(n9435), .B2(n9434), .A(n9433), .ZN(n9537) );
  NOR2_X1 U10388 ( .A1(n9537), .A2(n9479), .ZN(n9436) );
  AOI211_X1 U10389 ( .C1(n10768), .C2(n9534), .A(n9437), .B(n9436), .ZN(n9438)
         );
  OAI21_X1 U10390 ( .B1(n9536), .B2(n4949), .A(n9438), .ZN(P2_U3216) );
  XNOR2_X1 U10391 ( .A(n9439), .B(n5349), .ZN(n9441) );
  AOI222_X1 U10392 ( .A1(n9547), .A2(n9441), .B1(n9440), .B2(n9552), .C1(n9551), .C2(n9553), .ZN(n9540) );
  INV_X1 U10393 ( .A(n9442), .ZN(n9443) );
  OAI22_X1 U10394 ( .A1(n10846), .A2(n9444), .B1(n9443), .B2(n10838), .ZN(
        n9451) );
  INV_X1 U10395 ( .A(n9445), .ZN(n9453) );
  OAI21_X1 U10396 ( .B1(n9453), .B2(n9447), .A(n9446), .ZN(n9449) );
  NAND2_X1 U10397 ( .A1(n9449), .A2(n9448), .ZN(n9541) );
  NOR2_X1 U10398 ( .A1(n9541), .A2(n9479), .ZN(n9450) );
  AOI211_X1 U10399 ( .C1(n10768), .C2(n9538), .A(n9451), .B(n9450), .ZN(n9452)
         );
  OAI21_X1 U10400 ( .B1(n9540), .B2(n4949), .A(n9452), .ZN(P2_U3217) );
  AOI21_X1 U10401 ( .B1(n9455), .B2(n9454), .A(n9453), .ZN(n9542) );
  XNOR2_X1 U10402 ( .A(n9456), .B(n9455), .ZN(n9457) );
  OAI222_X1 U10403 ( .A1(n9473), .A2(n9458), .B1(n9471), .B2(n9472), .C1(n9457), .C2(n9468), .ZN(n9543) );
  NAND2_X1 U10404 ( .A1(n9543), .A2(n10846), .ZN(n9464) );
  INV_X1 U10405 ( .A(n9459), .ZN(n9460) );
  OAI22_X1 U10406 ( .A1(n10846), .A2(n9461), .B1(n9460), .B2(n10838), .ZN(
        n9462) );
  AOI21_X1 U10407 ( .B1(n9545), .B2(n10768), .A(n9462), .ZN(n9463) );
  OAI211_X1 U10408 ( .C1(n9542), .C2(n9479), .A(n9464), .B(n9463), .ZN(
        P2_U3218) );
  XNOR2_X1 U10409 ( .A(n9465), .B(n9466), .ZN(n9564) );
  XNOR2_X1 U10410 ( .A(n9467), .B(n9466), .ZN(n9469) );
  OAI222_X1 U10411 ( .A1(n9473), .A2(n9472), .B1(n9471), .B2(n9470), .C1(n9469), .C2(n9468), .ZN(n9565) );
  INV_X1 U10412 ( .A(n9567), .ZN(n9475) );
  OAI22_X1 U10413 ( .A1(n9475), .A2(n10840), .B1(n9474), .B2(n10838), .ZN(
        n9476) );
  OAI21_X1 U10414 ( .B1(n9565), .B2(n9476), .A(n10846), .ZN(n9478) );
  NAND2_X1 U10415 ( .A1(n4949), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9477) );
  OAI211_X1 U10416 ( .C1(n9564), .C2(n9479), .A(n9478), .B(n9477), .ZN(
        P2_U3220) );
  NOR2_X1 U10417 ( .A1(n9570), .A2(n9571), .ZN(n9481) );
  AOI21_X1 U10418 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n9570), .A(n9481), .ZN(
        n9480) );
  OAI21_X1 U10419 ( .B1(n9573), .B2(n9529), .A(n9480), .ZN(P2_U3490) );
  AOI21_X1 U10420 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n9570), .A(n9481), .ZN(
        n9482) );
  OAI21_X1 U10421 ( .B1(n9576), .B2(n9529), .A(n9482), .ZN(P2_U3489) );
  AOI22_X1 U10422 ( .A1(n9484), .A2(n9525), .B1(n9568), .B2(n9483), .ZN(n9485)
         );
  MUX2_X1 U10423 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9577), .S(n9561), .Z(
        P2_U3487) );
  AOI21_X1 U10424 ( .B1(n9525), .B2(n9488), .A(n9487), .ZN(n9578) );
  MUX2_X1 U10425 ( .A(n9489), .B(n9578), .S(n9561), .Z(n9490) );
  OAI21_X1 U10426 ( .B1(n9581), .B2(n9529), .A(n9490), .ZN(P2_U3486) );
  AOI21_X1 U10427 ( .B1(n9492), .B2(n9525), .A(n9491), .ZN(n9582) );
  MUX2_X1 U10428 ( .A(n9493), .B(n9582), .S(n9561), .Z(n9494) );
  OAI21_X1 U10429 ( .B1(n9585), .B2(n9529), .A(n9494), .ZN(P2_U3485) );
  AOI21_X1 U10430 ( .B1(n9525), .B2(n9496), .A(n9495), .ZN(n9586) );
  MUX2_X1 U10431 ( .A(n9497), .B(n9586), .S(n9561), .Z(n9498) );
  OAI21_X1 U10432 ( .B1(n9589), .B2(n9529), .A(n9498), .ZN(P2_U3484) );
  AOI21_X1 U10433 ( .B1(n9525), .B2(n9500), .A(n9499), .ZN(n9590) );
  MUX2_X1 U10434 ( .A(n9501), .B(n9590), .S(n9561), .Z(n9502) );
  OAI21_X1 U10435 ( .B1(n5510), .B2(n9529), .A(n9502), .ZN(P2_U3483) );
  AOI22_X1 U10436 ( .A1(n9504), .A2(n9525), .B1(n9568), .B2(n9503), .ZN(n9505)
         );
  NAND2_X1 U10437 ( .A1(n9506), .A2(n9505), .ZN(n9593) );
  MUX2_X1 U10438 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9593), .S(n9561), .Z(
        P2_U3482) );
  NOR2_X1 U10439 ( .A1(n9507), .A2(n9563), .ZN(n9510) );
  INV_X1 U10440 ( .A(n9508), .ZN(n9509) );
  AOI21_X1 U10441 ( .B1(n9510), .B2(n9357), .A(n9509), .ZN(n9594) );
  MUX2_X1 U10442 ( .A(n9511), .B(n9594), .S(n9561), .Z(n9512) );
  OAI21_X1 U10443 ( .B1(n9597), .B2(n9529), .A(n9512), .ZN(P2_U3481) );
  NOR2_X1 U10444 ( .A1(n9513), .A2(n9563), .ZN(n9516) );
  AOI21_X1 U10445 ( .B1(n9516), .B2(n9515), .A(n9514), .ZN(n9598) );
  MUX2_X1 U10446 ( .A(n9517), .B(n9598), .S(n9561), .Z(n9518) );
  OAI21_X1 U10447 ( .B1(n9601), .B2(n9529), .A(n9518), .ZN(P2_U3480) );
  NAND2_X1 U10448 ( .A1(n9519), .A2(n9568), .ZN(n9520) );
  OAI211_X1 U10449 ( .C1(n9563), .C2(n9522), .A(n9521), .B(n9520), .ZN(n9602)
         );
  MUX2_X1 U10450 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9602), .S(n9561), .Z(
        P2_U3479) );
  INV_X1 U10451 ( .A(n9523), .ZN(n9607) );
  INV_X1 U10452 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9527) );
  AOI21_X1 U10453 ( .B1(n9526), .B2(n9525), .A(n9524), .ZN(n9603) );
  MUX2_X1 U10454 ( .A(n9527), .B(n9603), .S(n9561), .Z(n9528) );
  OAI21_X1 U10455 ( .B1(n9607), .B2(n9529), .A(n9528), .ZN(P2_U3478) );
  NAND2_X1 U10456 ( .A1(n9530), .A2(n9568), .ZN(n9531) );
  OAI211_X1 U10457 ( .C1(n9563), .C2(n9533), .A(n9532), .B(n9531), .ZN(n9608)
         );
  MUX2_X1 U10458 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9608), .S(n9561), .Z(
        P2_U3477) );
  NAND2_X1 U10459 ( .A1(n9534), .A2(n9568), .ZN(n9535) );
  OAI211_X1 U10460 ( .C1(n9563), .C2(n9537), .A(n9536), .B(n9535), .ZN(n9609)
         );
  MUX2_X1 U10461 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9609), .S(n9561), .Z(
        P2_U3476) );
  NAND2_X1 U10462 ( .A1(n9538), .A2(n9568), .ZN(n9539) );
  OAI211_X1 U10463 ( .C1(n9563), .C2(n9541), .A(n9540), .B(n9539), .ZN(n9610)
         );
  MUX2_X1 U10464 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9610), .S(n9561), .Z(
        P2_U3475) );
  NOR2_X1 U10465 ( .A1(n9542), .A2(n9563), .ZN(n9544) );
  AOI211_X1 U10466 ( .C1(n9568), .C2(n9545), .A(n9544), .B(n9543), .ZN(n10851)
         );
  NAND2_X1 U10467 ( .A1(n9570), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n9546) );
  OAI21_X1 U10468 ( .B1(n10851), .B2(n9570), .A(n9546), .ZN(P2_U3474) );
  OAI211_X1 U10469 ( .C1(n9550), .C2(n9549), .A(n9548), .B(n9547), .ZN(n9556)
         );
  AOI22_X1 U10470 ( .A1(n9554), .A2(n9553), .B1(n9552), .B2(n9551), .ZN(n9555)
         );
  NAND2_X1 U10471 ( .A1(n9556), .A2(n9555), .ZN(n10842) );
  XNOR2_X1 U10472 ( .A(n9558), .B(n9557), .ZN(n10837) );
  OAI22_X1 U10473 ( .A1(n10837), .A2(n9563), .B1(n10841), .B2(n9559), .ZN(
        n9560) );
  NOR2_X1 U10474 ( .A1(n10842), .A2(n9560), .ZN(n10849) );
  OR2_X1 U10475 ( .A1(n9561), .A2(n6445), .ZN(n9562) );
  OAI21_X1 U10476 ( .B1(n10849), .B2(n9570), .A(n9562), .ZN(P2_U3473) );
  NOR2_X1 U10477 ( .A1(n9564), .A2(n9563), .ZN(n9566) );
  AOI211_X1 U10478 ( .C1(n9568), .C2(n9567), .A(n9566), .B(n9565), .ZN(n10836)
         );
  NAND2_X1 U10479 ( .A1(n9570), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9569) );
  OAI21_X1 U10480 ( .B1(n10836), .B2(n9570), .A(n9569), .ZN(P2_U3472) );
  NOR2_X1 U10481 ( .A1(n10850), .A2(n9571), .ZN(n9574) );
  AOI21_X1 U10482 ( .B1(P2_REG0_REG_31__SCAN_IN), .B2(n10850), .A(n9574), .ZN(
        n9572) );
  OAI21_X1 U10483 ( .B1(n9573), .B2(n9606), .A(n9572), .ZN(P2_U3458) );
  AOI21_X1 U10484 ( .B1(P2_REG0_REG_30__SCAN_IN), .B2(n10850), .A(n9574), .ZN(
        n9575) );
  OAI21_X1 U10485 ( .B1(n9576), .B2(n9606), .A(n9575), .ZN(P2_U3457) );
  MUX2_X1 U10486 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9577), .S(n10852), .Z(
        P2_U3455) );
  INV_X1 U10487 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9579) );
  MUX2_X1 U10488 ( .A(n9579), .B(n9578), .S(n10852), .Z(n9580) );
  OAI21_X1 U10489 ( .B1(n9581), .B2(n9606), .A(n9580), .ZN(P2_U3454) );
  INV_X1 U10490 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9583) );
  MUX2_X1 U10491 ( .A(n9583), .B(n9582), .S(n10852), .Z(n9584) );
  OAI21_X1 U10492 ( .B1(n9585), .B2(n9606), .A(n9584), .ZN(P2_U3453) );
  INV_X1 U10493 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9587) );
  MUX2_X1 U10494 ( .A(n9587), .B(n9586), .S(n10852), .Z(n9588) );
  OAI21_X1 U10495 ( .B1(n9589), .B2(n9606), .A(n9588), .ZN(P2_U3452) );
  INV_X1 U10496 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9591) );
  MUX2_X1 U10497 ( .A(n9591), .B(n9590), .S(n10852), .Z(n9592) );
  OAI21_X1 U10498 ( .B1(n5510), .B2(n9606), .A(n9592), .ZN(P2_U3451) );
  MUX2_X1 U10499 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9593), .S(n10852), .Z(
        P2_U3450) );
  INV_X1 U10500 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9595) );
  MUX2_X1 U10501 ( .A(n9595), .B(n9594), .S(n10852), .Z(n9596) );
  OAI21_X1 U10502 ( .B1(n9597), .B2(n9606), .A(n9596), .ZN(P2_U3449) );
  INV_X1 U10503 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9599) );
  MUX2_X1 U10504 ( .A(n9599), .B(n9598), .S(n10852), .Z(n9600) );
  OAI21_X1 U10505 ( .B1(n9601), .B2(n9606), .A(n9600), .ZN(P2_U3448) );
  MUX2_X1 U10506 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9602), .S(n10852), .Z(
        P2_U3447) );
  INV_X1 U10507 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9604) );
  MUX2_X1 U10508 ( .A(n9604), .B(n9603), .S(n10852), .Z(n9605) );
  OAI21_X1 U10509 ( .B1(n9607), .B2(n9606), .A(n9605), .ZN(P2_U3446) );
  MUX2_X1 U10510 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9608), .S(n10852), .Z(
        P2_U3444) );
  MUX2_X1 U10511 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9609), .S(n10852), .Z(
        P2_U3441) );
  MUX2_X1 U10512 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9610), .S(n10852), .Z(
        P2_U3438) );
  MUX2_X1 U10513 ( .A(n9612), .B(P2_D_REG_1__SCAN_IN), .S(n9611), .Z(P2_U3377)
         );
  INV_X1 U10514 ( .A(n10344), .ZN(n9616) );
  NOR4_X1 U10515 ( .A1(n6240), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9613), .A4(
        P2_U3151), .ZN(n9614) );
  AOI21_X1 U10516 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n9623), .A(n9614), .ZN(
        n9615) );
  OAI21_X1 U10517 ( .B1(n9616), .B2(n9625), .A(n9615), .ZN(P2_U3264) );
  AOI22_X1 U10518 ( .A1(n6242), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9623), .ZN(n9617) );
  OAI21_X1 U10519 ( .B1(n9618), .B2(n9625), .A(n9617), .ZN(P2_U3265) );
  INV_X1 U10520 ( .A(n9619), .ZN(n10353) );
  AOI22_X1 U10521 ( .A1(n9620), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9623), .ZN(n9621) );
  OAI21_X1 U10522 ( .B1(n10353), .B2(n9625), .A(n9621), .ZN(P2_U3266) );
  AOI21_X1 U10523 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n9623), .A(n9622), .ZN(
        n9624) );
  OAI21_X1 U10524 ( .B1(n9626), .B2(n9625), .A(n9624), .ZN(P2_U3267) );
  INV_X1 U10525 ( .A(n9627), .ZN(n9628) );
  MUX2_X1 U10526 ( .A(n9628), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10527 ( .A(n9629), .ZN(n9633) );
  AOI21_X1 U10528 ( .B1(n9763), .B2(n9631), .A(n9630), .ZN(n9632) );
  OAI21_X1 U10529 ( .B1(n9633), .B2(n9632), .A(n9764), .ZN(n9638) );
  OAI22_X1 U10530 ( .A1(n9779), .A2(n10205), .B1(n9781), .B2(n9991), .ZN(n9636) );
  NOR2_X1 U10531 ( .A1(n9634), .A2(n9783), .ZN(n9635) );
  AOI211_X1 U10532 ( .C1(P1_REG3_REG_27__SCAN_IN), .C2(P1_U3086), .A(n9636), 
        .B(n9635), .ZN(n9637) );
  OAI211_X1 U10533 ( .C1(n10206), .C2(n9737), .A(n9638), .B(n9637), .ZN(
        P1_U3214) );
  INV_X1 U10534 ( .A(n9639), .ZN(n9640) );
  NOR2_X1 U10535 ( .A1(n9641), .A2(n9640), .ZN(n9643) );
  XNOR2_X1 U10536 ( .A(n9643), .B(n9642), .ZN(n9651) );
  OAI21_X1 U10537 ( .B1(n9779), .B2(n9695), .A(n9644), .ZN(n9648) );
  OAI22_X1 U10538 ( .A1(n9783), .A2(n9646), .B1(n9781), .B2(n9645), .ZN(n9647)
         );
  AOI211_X1 U10539 ( .C1(n9649), .C2(n4944), .A(n9648), .B(n9647), .ZN(n9650)
         );
  OAI21_X1 U10540 ( .B1(n9651), .B2(n9788), .A(n9650), .ZN(P1_U3215) );
  INV_X1 U10541 ( .A(n9652), .ZN(n9653) );
  NAND2_X1 U10542 ( .A1(n9654), .A2(n9653), .ZN(n9741) );
  AOI21_X1 U10543 ( .B1(n9744), .B2(n9741), .A(n9743), .ZN(n9658) );
  XNOR2_X1 U10544 ( .A(n9656), .B(n9655), .ZN(n9657) );
  XNOR2_X1 U10545 ( .A(n9658), .B(n9657), .ZN(n9665) );
  OAI22_X1 U10546 ( .A1(n9660), .A2(n9779), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9659), .ZN(n9663) );
  INV_X1 U10547 ( .A(n10048), .ZN(n9661) );
  OAI22_X1 U10548 ( .A1(n9783), .A2(n9677), .B1(n9781), .B2(n9661), .ZN(n9662)
         );
  AOI211_X1 U10549 ( .C1(n10232), .C2(n4944), .A(n9663), .B(n9662), .ZN(n9664)
         );
  OAI21_X1 U10550 ( .B1(n9665), .B2(n9788), .A(n9664), .ZN(P1_U3216) );
  OAI21_X1 U10551 ( .B1(n9668), .B2(n9667), .A(n9666), .ZN(n9669) );
  NAND2_X1 U10552 ( .A1(n9669), .A2(n9764), .ZN(n9672) );
  AND2_X1 U10553 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9949) );
  OAI22_X1 U10554 ( .A1(n9783), .A2(n10279), .B1(n9781), .B2(n10117), .ZN(
        n9670) );
  AOI211_X1 U10555 ( .C1(n9768), .C2(n10258), .A(n9949), .B(n9670), .ZN(n9671)
         );
  OAI211_X1 U10556 ( .C1(n10327), .C2(n9737), .A(n9672), .B(n9671), .ZN(
        P1_U3219) );
  AOI21_X1 U10557 ( .B1(n9674), .B2(n9673), .A(n9788), .ZN(n9675) );
  NAND2_X1 U10558 ( .A1(n9675), .A2(n5404), .ZN(n9681) );
  NOR2_X1 U10559 ( .A1(n9783), .A2(n9676), .ZN(n9679) );
  OAI22_X1 U10560 ( .A1(n9779), .A2(n9677), .B1(n9781), .B2(n10092), .ZN(n9678) );
  AOI211_X1 U10561 ( .C1(P1_REG3_REG_21__SCAN_IN), .C2(P1_U3086), .A(n9679), 
        .B(n9678), .ZN(n9680) );
  OAI211_X1 U10562 ( .C1(n10319), .C2(n9737), .A(n9681), .B(n9680), .ZN(
        P1_U3223) );
  OAI21_X1 U10563 ( .B1(n9684), .B2(n9682), .A(n9683), .ZN(n9689) );
  AOI22_X1 U10564 ( .A1(n10028), .A2(n9768), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9687) );
  INV_X1 U10565 ( .A(n9685), .ZN(n10023) );
  AOI22_X1 U10566 ( .A1(n10023), .A2(n9769), .B1(n10056), .B2(n9767), .ZN(
        n9686) );
  OAI211_X1 U10567 ( .C1(n10025), .C2(n9737), .A(n9687), .B(n9686), .ZN(n9688)
         );
  AOI21_X1 U10568 ( .B1(n9689), .B2(n9764), .A(n9688), .ZN(n9690) );
  INV_X1 U10569 ( .A(n9690), .ZN(P1_U3225) );
  OAI21_X1 U10570 ( .B1(n9693), .B2(n5069), .A(n9691), .ZN(n9694) );
  NAND2_X1 U10571 ( .A1(n9694), .A2(n9764), .ZN(n9699) );
  OAI22_X1 U10572 ( .A1(n9783), .A2(n9695), .B1(n9781), .B2(n10161), .ZN(n9696) );
  AOI211_X1 U10573 ( .C1(n9768), .C2(n10266), .A(n9697), .B(n9696), .ZN(n9698)
         );
  OAI211_X1 U10574 ( .C1(n10336), .C2(n9737), .A(n9699), .B(n9698), .ZN(
        P1_U3226) );
  INV_X1 U10575 ( .A(n9700), .ZN(n9705) );
  AOI21_X1 U10576 ( .B1(n9704), .B2(n9702), .A(n9701), .ZN(n9703) );
  AOI21_X1 U10577 ( .B1(n9705), .B2(n9704), .A(n9703), .ZN(n9710) );
  OAI21_X1 U10578 ( .B1(n9779), .B2(n10279), .A(n9706), .ZN(n9708) );
  OAI22_X1 U10579 ( .A1(n9783), .A2(n10278), .B1(n9781), .B2(n10150), .ZN(
        n9707) );
  AOI211_X1 U10580 ( .C1(n10282), .C2(n4944), .A(n9708), .B(n9707), .ZN(n9709)
         );
  OAI21_X1 U10581 ( .B1(n9710), .B2(n9788), .A(n9709), .ZN(P1_U3228) );
  NAND2_X1 U10582 ( .A1(n9713), .A2(n9712), .ZN(n9714) );
  XNOR2_X1 U10583 ( .A(n9715), .B(n9714), .ZN(n9720) );
  OAI22_X1 U10584 ( .A1(n10224), .A2(n9779), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9716), .ZN(n9718) );
  OAI22_X1 U10585 ( .A1(n10071), .A2(n9783), .B1(n9781), .B2(n10035), .ZN(
        n9717) );
  AOI211_X1 U10586 ( .C1(n10227), .C2(n4944), .A(n9718), .B(n9717), .ZN(n9719)
         );
  OAI21_X1 U10587 ( .B1(n9720), .B2(n9788), .A(n9719), .ZN(P1_U3229) );
  OAI211_X1 U10588 ( .C1(n9723), .C2(n9722), .A(n9721), .B(n9764), .ZN(n9731)
         );
  INV_X1 U10589 ( .A(n9724), .ZN(n9725) );
  AOI22_X1 U10590 ( .A1(n9767), .A2(n9805), .B1(n9769), .B2(n9725), .ZN(n9730)
         );
  AND2_X1 U10591 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9854) );
  NOR2_X1 U10592 ( .A1(n9779), .A2(n9726), .ZN(n9727) );
  AOI211_X1 U10593 ( .C1(n9728), .C2(n4944), .A(n9854), .B(n9727), .ZN(n9729)
         );
  NAND3_X1 U10594 ( .A1(n9731), .A2(n9730), .A3(n9729), .ZN(P1_U3230) );
  OAI21_X1 U10595 ( .B1(n9734), .B2(n9733), .A(n9732), .ZN(n9739) );
  AOI22_X1 U10596 ( .A1(n9768), .A2(n10249), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9736) );
  AOI22_X1 U10597 ( .A1(n9767), .A2(n10269), .B1(n9769), .B2(n10103), .ZN(
        n9735) );
  OAI211_X1 U10598 ( .C1(n10323), .C2(n9737), .A(n9736), .B(n9735), .ZN(n9738)
         );
  AOI21_X1 U10599 ( .B1(n9739), .B2(n9764), .A(n9738), .ZN(n9740) );
  INV_X1 U10600 ( .A(n9740), .ZN(P1_U3233) );
  INV_X1 U10601 ( .A(n9741), .ZN(n9742) );
  NOR2_X1 U10602 ( .A1(n9743), .A2(n9742), .ZN(n9745) );
  XNOR2_X1 U10603 ( .A(n9745), .B(n9744), .ZN(n9750) );
  OAI22_X1 U10604 ( .A1(n9783), .A2(n10106), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9746), .ZN(n9748) );
  OAI22_X1 U10605 ( .A1(n10071), .A2(n9779), .B1(n9781), .B2(n10067), .ZN(
        n9747) );
  AOI211_X1 U10606 ( .C1(n10077), .C2(n4944), .A(n9748), .B(n9747), .ZN(n9749)
         );
  OAI21_X1 U10607 ( .B1(n9750), .B2(n9788), .A(n9749), .ZN(P1_U3235) );
  INV_X1 U10608 ( .A(n9751), .ZN(n9752) );
  NOR2_X1 U10609 ( .A1(n9753), .A2(n9752), .ZN(n9755) );
  XNOR2_X1 U10610 ( .A(n9755), .B(n9754), .ZN(n9761) );
  NAND2_X1 U10611 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9918) );
  OAI21_X1 U10612 ( .B1(n9779), .B2(n9756), .A(n9918), .ZN(n9758) );
  OAI22_X1 U10613 ( .A1(n9783), .A2(n10137), .B1(n9781), .B2(n10133), .ZN(
        n9757) );
  AOI211_X1 U10614 ( .C1(n10143), .C2(n4944), .A(n9758), .B(n9757), .ZN(n9760)
         );
  OAI21_X1 U10615 ( .B1(n9761), .B2(n9788), .A(n9760), .ZN(P1_U3238) );
  AND2_X1 U10616 ( .A1(n9683), .A2(n9762), .ZN(n9766) );
  OAI211_X1 U10617 ( .C1(n9766), .C2(n9765), .A(n9764), .B(n9763), .ZN(n9773)
         );
  AOI22_X1 U10618 ( .A1(n10005), .A2(n9767), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9772) );
  AOI22_X1 U10619 ( .A1(n10010), .A2(n9769), .B1(n9768), .B2(n10004), .ZN(
        n9771) );
  NAND2_X1 U10620 ( .A1(n10214), .A2(n4944), .ZN(n9770) );
  NAND4_X1 U10621 ( .A1(n9773), .A2(n9772), .A3(n9771), .A4(n9770), .ZN(
        P1_U3240) );
  XNOR2_X1 U10622 ( .A(n9775), .B(n9774), .ZN(n9776) );
  XNOR2_X1 U10623 ( .A(n9777), .B(n9776), .ZN(n9789) );
  OAI21_X1 U10624 ( .B1(n9779), .B2(n10278), .A(n9778), .ZN(n9785) );
  OAI22_X1 U10625 ( .A1(n9783), .A2(n9782), .B1(n9781), .B2(n9780), .ZN(n9784)
         );
  AOI211_X1 U10626 ( .C1(n9786), .C2(n4944), .A(n9785), .B(n9784), .ZN(n9787)
         );
  OAI21_X1 U10627 ( .B1(n9789), .B2(n9788), .A(n9787), .ZN(P1_U3241) );
  MUX2_X1 U10628 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9790), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10629 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9791), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10630 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9792), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10631 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n10004), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10632 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n10028), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10633 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n10005), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10634 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n10056), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10635 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n10086), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10636 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10258), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10637 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10269), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10638 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10257), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10639 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n10266), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10640 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9793), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10641 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n10165), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10642 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9794), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10643 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9795), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10644 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9796), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10645 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9797), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10646 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9798), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10647 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9799), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10648 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9800), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10649 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9801), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10650 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9802), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10651 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9803), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10652 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9804), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10653 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9805), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10654 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9806), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10655 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9807), .S(P1_U3973), .Z(
        P1_U3555) );
  AND2_X1 U10656 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9809) );
  OAI211_X1 U10657 ( .C1(n9810), .C2(n9809), .A(n9944), .B(n9808), .ZN(n9818)
         );
  OAI211_X1 U10658 ( .C1(n9813), .C2(n9812), .A(n9905), .B(n9811), .ZN(n9817)
         );
  AOI22_X1 U10659 ( .A1(n9950), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9816) );
  NAND2_X1 U10660 ( .A1(n9930), .A2(n9814), .ZN(n9815) );
  NAND4_X1 U10661 ( .A1(n9818), .A2(n9817), .A3(n9816), .A4(n9815), .ZN(
        P1_U3244) );
  NAND2_X1 U10662 ( .A1(n9819), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9820) );
  XNOR2_X1 U10663 ( .A(n9820), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9823) );
  NAND2_X1 U10664 ( .A1(n9821), .A2(n9824), .ZN(n9822) );
  OAI211_X1 U10665 ( .C1(n9824), .C2(n9823), .A(n9822), .B(P1_U3973), .ZN(
        n9863) );
  INV_X1 U10666 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9826) );
  OAI22_X1 U10667 ( .A1(n9920), .A2(n9826), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9825), .ZN(n9827) );
  AOI21_X1 U10668 ( .B1(n9828), .B2(n9930), .A(n9827), .ZN(n9837) );
  OAI211_X1 U10669 ( .C1(n9831), .C2(n9830), .A(n9905), .B(n9829), .ZN(n9836)
         );
  OAI211_X1 U10670 ( .C1(n9834), .C2(n9833), .A(n9944), .B(n9832), .ZN(n9835)
         );
  NAND4_X1 U10671 ( .A1(n9863), .A2(n9837), .A3(n9836), .A4(n9835), .ZN(
        P1_U3245) );
  INV_X1 U10672 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9840) );
  INV_X1 U10673 ( .A(n9838), .ZN(n9839) );
  OAI21_X1 U10674 ( .B1(n9920), .B2(n9840), .A(n9839), .ZN(n9841) );
  AOI21_X1 U10675 ( .B1(n9842), .B2(n9930), .A(n9841), .ZN(n9851) );
  OAI211_X1 U10676 ( .C1(n9845), .C2(n9844), .A(n9905), .B(n9843), .ZN(n9850)
         );
  OAI211_X1 U10677 ( .C1(n9848), .C2(n9847), .A(n9944), .B(n9846), .ZN(n9849)
         );
  NAND3_X1 U10678 ( .A1(n9851), .A2(n9850), .A3(n9849), .ZN(P1_U3246) );
  NOR2_X1 U10679 ( .A1(n9947), .A2(n9852), .ZN(n9853) );
  AOI211_X1 U10680 ( .C1(n9950), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n9854), .B(
        n9853), .ZN(n9864) );
  OAI211_X1 U10681 ( .C1(n9857), .C2(n9856), .A(n9944), .B(n9855), .ZN(n9862)
         );
  OAI211_X1 U10682 ( .C1(n9860), .C2(n9859), .A(n9905), .B(n9858), .ZN(n9861)
         );
  NAND4_X1 U10683 ( .A1(n9864), .A2(n9863), .A3(n9862), .A4(n9861), .ZN(
        P1_U3247) );
  AOI211_X1 U10684 ( .C1(n9867), .C2(n9866), .A(n9865), .B(n9895), .ZN(n9868)
         );
  INV_X1 U10685 ( .A(n9868), .ZN(n9878) );
  INV_X1 U10686 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9870) );
  OAI21_X1 U10687 ( .B1(n9920), .B2(n9870), .A(n9869), .ZN(n9871) );
  AOI21_X1 U10688 ( .B1(n9872), .B2(n9930), .A(n9871), .ZN(n9877) );
  OAI211_X1 U10689 ( .C1(n9875), .C2(n9874), .A(n9905), .B(n9873), .ZN(n9876)
         );
  NAND3_X1 U10690 ( .A1(n9878), .A2(n9877), .A3(n9876), .ZN(P1_U3248) );
  AOI211_X1 U10691 ( .C1(n9881), .C2(n9880), .A(n9879), .B(n9895), .ZN(n9882)
         );
  INV_X1 U10692 ( .A(n9882), .ZN(n9893) );
  INV_X1 U10693 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9885) );
  INV_X1 U10694 ( .A(n9883), .ZN(n9884) );
  OAI21_X1 U10695 ( .B1(n9920), .B2(n9885), .A(n9884), .ZN(n9886) );
  AOI21_X1 U10696 ( .B1(n9887), .B2(n9930), .A(n9886), .ZN(n9892) );
  OAI211_X1 U10697 ( .C1(n9890), .C2(n9889), .A(n9905), .B(n9888), .ZN(n9891)
         );
  NAND3_X1 U10698 ( .A1(n9893), .A2(n9892), .A3(n9891), .ZN(P1_U3249) );
  AOI211_X1 U10699 ( .C1(n9897), .C2(n9896), .A(n9895), .B(n9894), .ZN(n9898)
         );
  INV_X1 U10700 ( .A(n9898), .ZN(n9910) );
  INV_X1 U10701 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9901) );
  INV_X1 U10702 ( .A(n9899), .ZN(n9900) );
  OAI21_X1 U10703 ( .B1(n9920), .B2(n9901), .A(n9900), .ZN(n9902) );
  AOI21_X1 U10704 ( .B1(n9903), .B2(n9930), .A(n9902), .ZN(n9909) );
  OAI211_X1 U10705 ( .C1(n9907), .C2(n9906), .A(n9905), .B(n9904), .ZN(n9908)
         );
  NAND3_X1 U10706 ( .A1(n9910), .A2(n9909), .A3(n9908), .ZN(P1_U3251) );
  INV_X1 U10707 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9912) );
  AOI22_X1 U10708 ( .A1(n9914), .A2(n9913), .B1(n9912), .B2(n9911), .ZN(n9917)
         );
  NOR2_X1 U10709 ( .A1(n9915), .A2(n10275), .ZN(n9939) );
  AOI21_X1 U10710 ( .B1(n10275), .B2(n9915), .A(n9939), .ZN(n9916) );
  NAND2_X1 U10711 ( .A1(n9917), .A2(n9916), .ZN(n9941) );
  OAI211_X1 U10712 ( .C1(n9917), .C2(n9916), .A(n9941), .B(n9944), .ZN(n9932)
         );
  INV_X1 U10713 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9919) );
  OAI21_X1 U10714 ( .B1(n9920), .B2(n9919), .A(n9918), .ZN(n9928) );
  NAND2_X1 U10715 ( .A1(n9929), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9934) );
  OAI21_X1 U10716 ( .B1(n9929), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9934), .ZN(
        n9926) );
  INV_X1 U10717 ( .A(n9921), .ZN(n9923) );
  OAI22_X1 U10718 ( .A1(n9924), .A2(n9923), .B1(P1_REG2_REG_17__SCAN_IN), .B2(
        n9922), .ZN(n9925) );
  NOR2_X1 U10719 ( .A1(n9925), .A2(n9926), .ZN(n9936) );
  AOI211_X1 U10720 ( .C1(n9926), .C2(n9925), .A(n9936), .B(n9953), .ZN(n9927)
         );
  AOI211_X1 U10721 ( .C1(n9930), .C2(n9929), .A(n9928), .B(n9927), .ZN(n9931)
         );
  NAND2_X1 U10722 ( .A1(n9932), .A2(n9931), .ZN(P1_U3261) );
  INV_X1 U10723 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9933) );
  MUX2_X1 U10724 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9933), .S(n6137), .Z(n9938) );
  INV_X1 U10725 ( .A(n9934), .ZN(n9935) );
  NOR2_X1 U10726 ( .A1(n9936), .A2(n9935), .ZN(n9937) );
  XOR2_X1 U10727 ( .A(n9938), .B(n9937), .Z(n9954) );
  INV_X1 U10728 ( .A(n9939), .ZN(n9940) );
  NAND2_X1 U10729 ( .A1(n9941), .A2(n9940), .ZN(n9943) );
  XNOR2_X1 U10730 ( .A(n6137), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9942) );
  XNOR2_X1 U10731 ( .A(n9943), .B(n9942), .ZN(n9945) );
  NAND2_X1 U10732 ( .A1(n9945), .A2(n9944), .ZN(n9952) );
  NOR2_X1 U10733 ( .A1(n9947), .A2(n9946), .ZN(n9948) );
  AOI211_X1 U10734 ( .C1(P1_ADDR_REG_19__SCAN_IN), .C2(n9950), .A(n9949), .B(
        n9948), .ZN(n9951) );
  OAI211_X1 U10735 ( .C1(n9954), .C2(n9953), .A(n9952), .B(n9951), .ZN(
        P1_U3262) );
  XOR2_X1 U10736 ( .A(n9955), .B(n10302), .Z(n9956) );
  NAND2_X1 U10737 ( .A1(n10202), .A2(n10814), .ZN(n9959) );
  NOR2_X1 U10738 ( .A1(n10820), .A2(n9957), .ZN(n9961) );
  AOI21_X1 U10739 ( .B1(n10820), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9961), .ZN(
        n9958) );
  OAI211_X1 U10740 ( .C1(n10302), .C2(n10178), .A(n9959), .B(n9958), .ZN(
        P1_U3263) );
  NOR2_X1 U10741 ( .A1(n10732), .A2(n9960), .ZN(n9962) );
  AOI211_X1 U10742 ( .C1(n9963), .C2(n10809), .A(n9962), .B(n9961), .ZN(n9964)
         );
  OAI21_X1 U10743 ( .B1(n9965), .B2(n10184), .A(n9964), .ZN(P1_U3264) );
  NAND2_X1 U10744 ( .A1(n9966), .A2(n10189), .ZN(n9973) );
  OAI22_X1 U10745 ( .A1(n10732), .A2(n9968), .B1(n9967), .B2(n10729), .ZN(
        n9971) );
  NOR2_X1 U10746 ( .A1(n9969), .A2(n10184), .ZN(n9970) );
  AOI211_X1 U10747 ( .C1(n10809), .C2(n6734), .A(n9971), .B(n9970), .ZN(n9972)
         );
  OAI211_X1 U10748 ( .C1(n9974), .C2(n10820), .A(n9973), .B(n9972), .ZN(
        P1_U3356) );
  NAND2_X1 U10749 ( .A1(n9975), .A2(n10189), .ZN(n9985) );
  INV_X1 U10750 ( .A(n9976), .ZN(n9977) );
  AOI22_X1 U10751 ( .A1(n10820), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9977), 
        .B2(n10807), .ZN(n9978) );
  OAI21_X1 U10752 ( .B1(n9979), .B2(n10185), .A(n9978), .ZN(n9982) );
  NOR2_X1 U10753 ( .A1(n9980), .A2(n10184), .ZN(n9981) );
  AOI211_X1 U10754 ( .C1(n10809), .C2(n9983), .A(n9982), .B(n9981), .ZN(n9984)
         );
  OAI211_X1 U10755 ( .C1(n9986), .C2(n10820), .A(n9985), .B(n9984), .ZN(
        P1_U3265) );
  INV_X1 U10756 ( .A(n9987), .ZN(n9988) );
  AOI211_X1 U10757 ( .C1(n9990), .C2(n10009), .A(n10174), .B(n5302), .ZN(
        n10208) );
  NAND2_X1 U10758 ( .A1(n9990), .A2(n10809), .ZN(n9994) );
  INV_X1 U10759 ( .A(n9991), .ZN(n9992) );
  AOI22_X1 U10760 ( .A1(n10820), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n10807), 
        .B2(n9992), .ZN(n9993) );
  OAI211_X1 U10761 ( .C1(n10205), .C2(n10185), .A(n9994), .B(n9993), .ZN(
        n10000) );
  NAND2_X1 U10762 ( .A1(n10002), .A2(n9995), .ZN(n9997) );
  XNOR2_X1 U10763 ( .A(n9997), .B(n9996), .ZN(n9998) );
  NOR2_X1 U10764 ( .A1(n10210), .A2(n10820), .ZN(n9999) );
  OAI21_X1 U10765 ( .B1(n10211), .B2(n10098), .A(n10001), .ZN(P1_U3266) );
  OAI21_X1 U10766 ( .B1(n10007), .B2(n10003), .A(n10002), .ZN(n10006) );
  AOI222_X1 U10767 ( .A1(n10162), .A2(n10006), .B1(n10005), .B2(n10267), .C1(
        n10004), .C2(n10268), .ZN(n10217) );
  NAND2_X1 U10768 ( .A1(n10008), .A2(n10007), .ZN(n10212) );
  NAND3_X1 U10769 ( .A1(n10213), .A2(n10212), .A3(n10189), .ZN(n10016) );
  OAI211_X1 U10770 ( .C1(n10012), .C2(n10022), .A(n10782), .B(n10009), .ZN(
        n10216) );
  INV_X1 U10771 ( .A(n10216), .ZN(n10014) );
  AOI22_X1 U10772 ( .A1(n10010), .A2(n10807), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10820), .ZN(n10011) );
  OAI21_X1 U10773 ( .B1(n10012), .B2(n10178), .A(n10011), .ZN(n10013) );
  AOI21_X1 U10774 ( .B1(n10014), .B2(n10814), .A(n10013), .ZN(n10015) );
  OAI211_X1 U10775 ( .C1(n10820), .C2(n10217), .A(n10016), .B(n10015), .ZN(
        P1_U3267) );
  OR2_X1 U10776 ( .A1(n10017), .A2(n10018), .ZN(n10020) );
  NAND2_X1 U10777 ( .A1(n10020), .A2(n10019), .ZN(n10021) );
  XOR2_X1 U10778 ( .A(n10026), .B(n10021), .Z(n10223) );
  AOI211_X1 U10779 ( .C1(n10220), .C2(n10033), .A(n10174), .B(n10022), .ZN(
        n10219) );
  AOI22_X1 U10780 ( .A1(n10023), .A2(n10807), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10820), .ZN(n10024) );
  OAI21_X1 U10781 ( .B1(n10025), .B2(n10178), .A(n10024), .ZN(n10031) );
  XOR2_X1 U10782 ( .A(n10027), .B(n10026), .Z(n10029) );
  AOI222_X1 U10783 ( .A1(n10162), .A2(n10029), .B1(n10028), .B2(n10268), .C1(
        n10056), .C2(n10267), .ZN(n10222) );
  NOR2_X1 U10784 ( .A1(n10222), .A2(n10820), .ZN(n10030) );
  AOI211_X1 U10785 ( .C1(n10219), .C2(n10814), .A(n10031), .B(n10030), .ZN(
        n10032) );
  OAI21_X1 U10786 ( .B1(n10223), .B2(n10098), .A(n10032), .ZN(P1_U3268) );
  XNOR2_X1 U10787 ( .A(n10017), .B(n10040), .ZN(n10230) );
  INV_X1 U10788 ( .A(n10033), .ZN(n10034) );
  AOI211_X1 U10789 ( .C1(n10227), .C2(n10046), .A(n10174), .B(n10034), .ZN(
        n10225) );
  NAND2_X1 U10790 ( .A1(n10227), .A2(n10809), .ZN(n10038) );
  INV_X1 U10791 ( .A(n10035), .ZN(n10036) );
  AOI22_X1 U10792 ( .A1(P1_REG2_REG_24__SCAN_IN), .A2(n10820), .B1(n10036), 
        .B2(n10807), .ZN(n10037) );
  OAI211_X1 U10793 ( .C1(n10224), .C2(n10185), .A(n10038), .B(n10037), .ZN(
        n10043) );
  XNOR2_X1 U10794 ( .A(n10039), .B(n10040), .ZN(n10041) );
  AOI22_X1 U10795 ( .A1(n10041), .A2(n10162), .B1(n10267), .B2(n10236), .ZN(
        n10229) );
  NOR2_X1 U10796 ( .A1(n10229), .A2(n10820), .ZN(n10042) );
  AOI211_X1 U10797 ( .C1(n10225), .C2(n10814), .A(n10043), .B(n10042), .ZN(
        n10044) );
  OAI21_X1 U10798 ( .B1(n10230), .B2(n10098), .A(n10044), .ZN(P1_U3269) );
  XNOR2_X1 U10799 ( .A(n10045), .B(n10054), .ZN(n10235) );
  INV_X1 U10800 ( .A(n10046), .ZN(n10047) );
  AOI211_X1 U10801 ( .C1(n10232), .C2(n5289), .A(n10174), .B(n10047), .ZN(
        n10231) );
  AOI22_X1 U10802 ( .A1(n10820), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n10048), 
        .B2(n10807), .ZN(n10049) );
  OAI21_X1 U10803 ( .B1(n10050), .B2(n10178), .A(n10049), .ZN(n10059) );
  INV_X1 U10804 ( .A(n10061), .ZN(n10052) );
  NOR2_X1 U10805 ( .A1(n10052), .A2(n10051), .ZN(n10055) );
  OAI21_X1 U10806 ( .B1(n10055), .B2(n10054), .A(n10053), .ZN(n10057) );
  AOI222_X1 U10807 ( .A1(n10162), .A2(n10057), .B1(n10056), .B2(n10268), .C1(
        n10086), .C2(n10267), .ZN(n10234) );
  NOR2_X1 U10808 ( .A1(n10234), .A2(n10820), .ZN(n10058) );
  AOI211_X1 U10809 ( .C1(n10231), .C2(n10814), .A(n10059), .B(n10058), .ZN(
        n10060) );
  OAI21_X1 U10810 ( .B1(n10235), .B2(n10098), .A(n10060), .ZN(P1_U3270) );
  OAI211_X1 U10811 ( .C1(n10063), .C2(n10062), .A(n10061), .B(n10162), .ZN(
        n10239) );
  OAI21_X1 U10812 ( .B1(n10066), .B2(n10065), .A(n10064), .ZN(n10241) );
  NAND2_X1 U10813 ( .A1(n10241), .A2(n10189), .ZN(n10079) );
  INV_X1 U10814 ( .A(n10067), .ZN(n10068) );
  AOI22_X1 U10815 ( .A1(n10820), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n10068), 
        .B2(n10807), .ZN(n10070) );
  NAND2_X1 U10816 ( .A1(n10195), .A2(n10249), .ZN(n10069) );
  OAI211_X1 U10817 ( .C1(n10071), .C2(n10185), .A(n10070), .B(n10069), .ZN(
        n10076) );
  NAND2_X1 U10818 ( .A1(n10077), .A2(n10089), .ZN(n10072) );
  NAND2_X1 U10819 ( .A1(n10072), .A2(n10782), .ZN(n10073) );
  OR2_X1 U10820 ( .A1(n10074), .A2(n10073), .ZN(n10237) );
  NOR2_X1 U10821 ( .A1(n10237), .A2(n10184), .ZN(n10075) );
  AOI211_X1 U10822 ( .C1(n10809), .C2(n10077), .A(n10076), .B(n10075), .ZN(
        n10078) );
  OAI211_X1 U10823 ( .C1(n10820), .C2(n10239), .A(n10079), .B(n10078), .ZN(
        P1_U3271) );
  OAI21_X1 U10824 ( .B1(n10081), .B2(n10084), .A(n10080), .ZN(n10246) );
  INV_X1 U10825 ( .A(n10246), .ZN(n10099) );
  NAND2_X1 U10826 ( .A1(n10083), .A2(n10082), .ZN(n10085) );
  XNOR2_X1 U10827 ( .A(n10085), .B(n10084), .ZN(n10088) );
  AOI22_X1 U10828 ( .A1(n10086), .A2(n10268), .B1(n10267), .B2(n10258), .ZN(
        n10087) );
  OAI21_X1 U10829 ( .B1(n10088), .B2(n10791), .A(n10087), .ZN(n10244) );
  INV_X1 U10830 ( .A(n10089), .ZN(n10090) );
  AOI211_X1 U10831 ( .C1(n10091), .C2(n10107), .A(n10174), .B(n10090), .ZN(
        n10245) );
  NAND2_X1 U10832 ( .A1(n10245), .A2(n10814), .ZN(n10095) );
  INV_X1 U10833 ( .A(n10092), .ZN(n10093) );
  AOI22_X1 U10834 ( .A1(n10820), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n10093), 
        .B2(n10807), .ZN(n10094) );
  OAI211_X1 U10835 ( .C1(n10319), .C2(n10178), .A(n10095), .B(n10094), .ZN(
        n10096) );
  AOI21_X1 U10836 ( .B1(n10732), .B2(n10244), .A(n10096), .ZN(n10097) );
  OAI21_X1 U10837 ( .B1(n10099), .B2(n10098), .A(n10097), .ZN(P1_U3272) );
  XNOR2_X1 U10838 ( .A(n10100), .B(n10101), .ZN(n10252) );
  XNOR2_X1 U10839 ( .A(n10102), .B(n10101), .ZN(n10254) );
  NAND2_X1 U10840 ( .A1(n10254), .A2(n10189), .ZN(n10112) );
  AOI22_X1 U10841 ( .A1(n10820), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n10103), 
        .B2(n10807), .ZN(n10105) );
  NAND2_X1 U10842 ( .A1(n10195), .A2(n10269), .ZN(n10104) );
  OAI211_X1 U10843 ( .C1(n10106), .C2(n10185), .A(n10105), .B(n10104), .ZN(
        n10109) );
  OAI211_X1 U10844 ( .C1(n10323), .C2(n10120), .A(n10782), .B(n10107), .ZN(
        n10250) );
  NOR2_X1 U10845 ( .A1(n10250), .A2(n10184), .ZN(n10108) );
  AOI211_X1 U10846 ( .C1(n10809), .C2(n10110), .A(n10109), .B(n10108), .ZN(
        n10111) );
  OAI211_X1 U10847 ( .C1(n10252), .C2(n10160), .A(n10112), .B(n10111), .ZN(
        P1_U3273) );
  XNOR2_X1 U10848 ( .A(n10114), .B(n10113), .ZN(n10261) );
  XNOR2_X1 U10849 ( .A(n10116), .B(n10115), .ZN(n10263) );
  NAND2_X1 U10850 ( .A1(n10263), .A2(n10189), .ZN(n10127) );
  OAI22_X1 U10851 ( .A1(n10732), .A2(n9933), .B1(n10117), .B2(n10729), .ZN(
        n10118) );
  AOI21_X1 U10852 ( .B1(n10153), .B2(n10258), .A(n10118), .ZN(n10119) );
  OAI21_X1 U10853 ( .B1(n10279), .B2(n10156), .A(n10119), .ZN(n10124) );
  INV_X1 U10854 ( .A(n10140), .ZN(n10122) );
  INV_X1 U10855 ( .A(n10120), .ZN(n10121) );
  OAI211_X1 U10856 ( .C1(n10327), .C2(n10122), .A(n10121), .B(n10782), .ZN(
        n10259) );
  NOR2_X1 U10857 ( .A1(n10259), .A2(n10184), .ZN(n10123) );
  AOI211_X1 U10858 ( .C1(n10809), .C2(n10125), .A(n10124), .B(n10123), .ZN(
        n10126) );
  OAI211_X1 U10859 ( .C1(n10160), .C2(n10261), .A(n10127), .B(n10126), .ZN(
        P1_U3274) );
  NAND2_X1 U10860 ( .A1(n10129), .A2(n10128), .ZN(n10130) );
  XOR2_X1 U10861 ( .A(n10131), .B(n10130), .Z(n10272) );
  XNOR2_X1 U10862 ( .A(n10132), .B(n10131), .ZN(n10274) );
  NAND2_X1 U10863 ( .A1(n10274), .A2(n10189), .ZN(n10145) );
  OAI22_X1 U10864 ( .A1(n10732), .A2(n10134), .B1(n10133), .B2(n10729), .ZN(
        n10135) );
  AOI21_X1 U10865 ( .B1(n10153), .B2(n10269), .A(n10135), .ZN(n10136) );
  OAI21_X1 U10866 ( .B1(n10137), .B2(n10156), .A(n10136), .ZN(n10142) );
  AOI21_X1 U10867 ( .B1(n10143), .B2(n10138), .A(n10174), .ZN(n10139) );
  NAND2_X1 U10868 ( .A1(n10140), .A2(n10139), .ZN(n10270) );
  NOR2_X1 U10869 ( .A1(n10270), .A2(n10184), .ZN(n10141) );
  AOI211_X1 U10870 ( .C1(n10809), .C2(n10143), .A(n10142), .B(n10141), .ZN(
        n10144) );
  OAI211_X1 U10871 ( .C1(n10160), .C2(n10272), .A(n10145), .B(n10144), .ZN(
        P1_U3275) );
  XNOR2_X1 U10872 ( .A(n10146), .B(n10147), .ZN(n10286) );
  AOI21_X1 U10873 ( .B1(n10148), .B2(n10147), .A(n5009), .ZN(n10277) );
  NAND2_X1 U10874 ( .A1(n10277), .A2(n10189), .ZN(n10159) );
  AOI211_X1 U10875 ( .C1(n10282), .C2(n10172), .A(n10174), .B(n10149), .ZN(
        n10280) );
  NAND2_X1 U10876 ( .A1(n10282), .A2(n10809), .ZN(n10155) );
  INV_X1 U10877 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10151) );
  OAI22_X1 U10878 ( .A1(n10732), .A2(n10151), .B1(n10150), .B2(n10729), .ZN(
        n10152) );
  AOI21_X1 U10879 ( .B1(n10153), .B2(n10257), .A(n10152), .ZN(n10154) );
  OAI211_X1 U10880 ( .C1(n10278), .C2(n10156), .A(n10155), .B(n10154), .ZN(
        n10157) );
  AOI21_X1 U10881 ( .B1(n10280), .B2(n10814), .A(n10157), .ZN(n10158) );
  OAI211_X1 U10882 ( .C1(n10286), .C2(n10160), .A(n10159), .B(n10158), .ZN(
        P1_U3276) );
  INV_X1 U10883 ( .A(n10161), .ZN(n10168) );
  OAI211_X1 U10884 ( .C1(n10164), .C2(n10169), .A(n10163), .B(n10162), .ZN(
        n10167) );
  AOI22_X1 U10885 ( .A1(n10267), .A2(n10165), .B1(n10268), .B2(n10266), .ZN(
        n10166) );
  NAND2_X1 U10886 ( .A1(n10167), .A2(n10166), .ZN(n10287) );
  AOI21_X1 U10887 ( .B1(n10168), .B2(n10807), .A(n10287), .ZN(n10182) );
  XNOR2_X1 U10888 ( .A(n10170), .B(n10169), .ZN(n10289) );
  NAND2_X1 U10889 ( .A1(n10289), .A2(n10189), .ZN(n10181) );
  INV_X1 U10890 ( .A(n10171), .ZN(n10175) );
  INV_X1 U10891 ( .A(n10172), .ZN(n10173) );
  AOI211_X1 U10892 ( .C1(n10176), .C2(n10175), .A(n10174), .B(n10173), .ZN(
        n10288) );
  OAI22_X1 U10893 ( .A1(n10336), .A2(n10178), .B1(n10732), .B2(n10177), .ZN(
        n10179) );
  AOI21_X1 U10894 ( .B1(n10288), .B2(n10814), .A(n10179), .ZN(n10180) );
  OAI211_X1 U10895 ( .C1(n10820), .C2(n10182), .A(n10181), .B(n10180), .ZN(
        P1_U3277) );
  OAI22_X1 U10896 ( .A1(n10186), .A2(n10185), .B1(n10184), .B2(n10183), .ZN(
        n10187) );
  AOI21_X1 U10897 ( .B1(n10189), .B2(n10188), .A(n10187), .ZN(n10200) );
  INV_X1 U10898 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10191) );
  OAI22_X1 U10899 ( .A1(n10732), .A2(n10191), .B1(n10190), .B2(n10729), .ZN(
        n10192) );
  AOI21_X1 U10900 ( .B1(n10809), .B2(n10193), .A(n10192), .ZN(n10199) );
  NAND2_X1 U10901 ( .A1(n10195), .A2(n5056), .ZN(n10198) );
  NAND2_X1 U10902 ( .A1(n10732), .A2(n10196), .ZN(n10197) );
  NAND4_X1 U10903 ( .A1(n10200), .A2(n10199), .A3(n10198), .A4(n10197), .ZN(
        P1_U3292) );
  INV_X1 U10904 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10203) );
  NOR2_X1 U10905 ( .A1(n10202), .A2(n10201), .ZN(n10299) );
  MUX2_X1 U10906 ( .A(n10203), .B(n10299), .S(n10831), .Z(n10204) );
  OAI21_X1 U10907 ( .B1(n10302), .B2(n10298), .A(n10204), .ZN(P1_U3553) );
  OAI22_X1 U10908 ( .A1(n10206), .A2(n10824), .B1(n10205), .B2(n10794), .ZN(
        n10207) );
  NOR2_X1 U10909 ( .A1(n10208), .A2(n10207), .ZN(n10209) );
  OAI211_X1 U10910 ( .C1(n10211), .C2(n10735), .A(n10210), .B(n10209), .ZN(
        n10307) );
  MUX2_X1 U10911 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10307), .S(n10831), .Z(
        P1_U3549) );
  NAND3_X1 U10912 ( .A1(n10213), .A2(n10212), .A3(n10828), .ZN(n10218) );
  NAND2_X1 U10913 ( .A1(n10214), .A2(n10283), .ZN(n10215) );
  MUX2_X1 U10914 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10308), .S(n10831), .Z(
        P1_U3548) );
  AOI21_X1 U10915 ( .B1(n10283), .B2(n10220), .A(n10219), .ZN(n10221) );
  OAI211_X1 U10916 ( .C1(n10223), .C2(n10735), .A(n10222), .B(n10221), .ZN(
        n10309) );
  MUX2_X1 U10917 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10309), .S(n10831), .Z(
        P1_U3547) );
  NOR2_X1 U10918 ( .A1(n10224), .A2(n10794), .ZN(n10226) );
  AOI211_X1 U10919 ( .C1(n10283), .C2(n10227), .A(n10226), .B(n10225), .ZN(
        n10228) );
  OAI211_X1 U10920 ( .C1(n10230), .C2(n10735), .A(n10229), .B(n10228), .ZN(
        n10310) );
  MUX2_X1 U10921 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10310), .S(n10831), .Z(
        P1_U3546) );
  AOI21_X1 U10922 ( .B1(n10283), .B2(n10232), .A(n10231), .ZN(n10233) );
  OAI211_X1 U10923 ( .C1(n10235), .C2(n10735), .A(n10234), .B(n10233), .ZN(
        n10311) );
  MUX2_X1 U10924 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10311), .S(n10831), .Z(
        P1_U3545) );
  AOI22_X1 U10925 ( .A1(n10236), .A2(n10268), .B1(n10267), .B2(n10249), .ZN(
        n10238) );
  NAND3_X1 U10926 ( .A1(n10239), .A2(n10238), .A3(n10237), .ZN(n10240) );
  AOI21_X1 U10927 ( .B1(n10241), .B2(n5053), .A(n10240), .ZN(n10312) );
  MUX2_X1 U10928 ( .A(n10242), .B(n10312), .S(n10831), .Z(n10243) );
  OAI21_X1 U10929 ( .B1(n10315), .B2(n10298), .A(n10243), .ZN(P1_U3544) );
  AOI211_X1 U10930 ( .C1(n10246), .C2(n10828), .A(n10245), .B(n10244), .ZN(
        n10316) );
  MUX2_X1 U10931 ( .A(n10247), .B(n10316), .S(n10831), .Z(n10248) );
  OAI21_X1 U10932 ( .B1(n10319), .B2(n10298), .A(n10248), .ZN(P1_U3543) );
  AOI22_X1 U10933 ( .A1(n10249), .A2(n10268), .B1(n10267), .B2(n10269), .ZN(
        n10251) );
  OAI211_X1 U10934 ( .C1(n10252), .C2(n10791), .A(n10251), .B(n10250), .ZN(
        n10253) );
  AOI21_X1 U10935 ( .B1(n10254), .B2(n5053), .A(n10253), .ZN(n10320) );
  MUX2_X1 U10936 ( .A(n10255), .B(n10320), .S(n10831), .Z(n10256) );
  OAI21_X1 U10937 ( .B1(n10323), .B2(n10298), .A(n10256), .ZN(P1_U3542) );
  AOI22_X1 U10938 ( .A1(n10258), .A2(n10268), .B1(n10267), .B2(n10257), .ZN(
        n10260) );
  OAI211_X1 U10939 ( .C1(n10261), .C2(n10791), .A(n10260), .B(n10259), .ZN(
        n10262) );
  AOI21_X1 U10940 ( .B1(n10263), .B2(n5053), .A(n10262), .ZN(n10324) );
  MUX2_X1 U10941 ( .A(n10264), .B(n10324), .S(n10831), .Z(n10265) );
  OAI21_X1 U10942 ( .B1(n10327), .B2(n10298), .A(n10265), .ZN(P1_U3541) );
  AOI22_X1 U10943 ( .A1(n10269), .A2(n10268), .B1(n10267), .B2(n10266), .ZN(
        n10271) );
  OAI211_X1 U10944 ( .C1(n10272), .C2(n10791), .A(n10271), .B(n10270), .ZN(
        n10273) );
  AOI21_X1 U10945 ( .B1(n10274), .B2(n5053), .A(n10273), .ZN(n10328) );
  MUX2_X1 U10946 ( .A(n10275), .B(n10328), .S(n10831), .Z(n10276) );
  OAI21_X1 U10947 ( .B1(n10331), .B2(n10298), .A(n10276), .ZN(P1_U3540) );
  NAND2_X1 U10948 ( .A1(n10277), .A2(n10828), .ZN(n10285) );
  OAI22_X1 U10949 ( .A1(n10279), .A2(n10794), .B1(n10278), .B2(n10796), .ZN(
        n10281) );
  AOI211_X1 U10950 ( .C1(n10283), .C2(n10282), .A(n10281), .B(n10280), .ZN(
        n10284) );
  OAI211_X1 U10951 ( .C1(n10791), .C2(n10286), .A(n10285), .B(n10284), .ZN(
        n10332) );
  MUX2_X1 U10952 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10332), .S(n10831), .Z(
        P1_U3539) );
  AOI211_X1 U10953 ( .C1(n10289), .C2(n10828), .A(n10288), .B(n10287), .ZN(
        n10333) );
  MUX2_X1 U10954 ( .A(n10290), .B(n10333), .S(n10831), .Z(n10291) );
  OAI21_X1 U10955 ( .B1(n10336), .B2(n10298), .A(n10291), .ZN(P1_U3538) );
  INV_X1 U10956 ( .A(n10292), .ZN(n10295) );
  AOI211_X1 U10957 ( .C1(n10295), .C2(n10828), .A(n10294), .B(n10293), .ZN(
        n10337) );
  MUX2_X1 U10958 ( .A(n10296), .B(n10337), .S(n10831), .Z(n10297) );
  OAI21_X1 U10959 ( .B1(n10341), .B2(n10298), .A(n10297), .ZN(P1_U3537) );
  MUX2_X1 U10960 ( .A(n10300), .B(n10299), .S(n10834), .Z(n10301) );
  OAI21_X1 U10961 ( .B1(n10302), .B2(n10340), .A(n10301), .ZN(P1_U3521) );
  MUX2_X1 U10962 ( .A(n10303), .B(P1_REG0_REG_30__SCAN_IN), .S(n6207), .Z(
        n10304) );
  INV_X1 U10963 ( .A(n10304), .ZN(n10305) );
  OAI21_X1 U10964 ( .B1(n10306), .B2(n10340), .A(n10305), .ZN(P1_U3520) );
  MUX2_X1 U10965 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10307), .S(n10834), .Z(
        P1_U3517) );
  MUX2_X1 U10966 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10308), .S(n10834), .Z(
        P1_U3516) );
  MUX2_X1 U10967 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10309), .S(n10834), .Z(
        P1_U3515) );
  MUX2_X1 U10968 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10310), .S(n10834), .Z(
        P1_U3514) );
  MUX2_X1 U10969 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10311), .S(n10834), .Z(
        P1_U3513) );
  INV_X1 U10970 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10313) );
  MUX2_X1 U10971 ( .A(n10313), .B(n10312), .S(n10834), .Z(n10314) );
  OAI21_X1 U10972 ( .B1(n10315), .B2(n10340), .A(n10314), .ZN(P1_U3512) );
  INV_X1 U10973 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10317) );
  MUX2_X1 U10974 ( .A(n10317), .B(n10316), .S(n10834), .Z(n10318) );
  OAI21_X1 U10975 ( .B1(n10319), .B2(n10340), .A(n10318), .ZN(P1_U3511) );
  INV_X1 U10976 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10321) );
  MUX2_X1 U10977 ( .A(n10321), .B(n10320), .S(n10834), .Z(n10322) );
  OAI21_X1 U10978 ( .B1(n10323), .B2(n10340), .A(n10322), .ZN(P1_U3510) );
  INV_X1 U10979 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10325) );
  MUX2_X1 U10980 ( .A(n10325), .B(n10324), .S(n10834), .Z(n10326) );
  OAI21_X1 U10981 ( .B1(n10327), .B2(n10340), .A(n10326), .ZN(P1_U3509) );
  INV_X1 U10982 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10329) );
  MUX2_X1 U10983 ( .A(n10329), .B(n10328), .S(n10834), .Z(n10330) );
  OAI21_X1 U10984 ( .B1(n10331), .B2(n10340), .A(n10330), .ZN(P1_U3507) );
  MUX2_X1 U10985 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10332), .S(n10834), .Z(
        P1_U3504) );
  MUX2_X1 U10986 ( .A(n10334), .B(n10333), .S(n10834), .Z(n10335) );
  OAI21_X1 U10987 ( .B1(n10336), .B2(n10340), .A(n10335), .ZN(P1_U3501) );
  INV_X1 U10988 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10338) );
  MUX2_X1 U10989 ( .A(n10338), .B(n10337), .S(n10834), .Z(n10339) );
  OAI21_X1 U10990 ( .B1(n10341), .B2(n10340), .A(n10339), .ZN(P1_U3498) );
  NAND3_X1 U10991 ( .A1(n10342), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n10348) );
  NAND2_X1 U10992 ( .A1(n10344), .A2(n10343), .ZN(n10347) );
  NAND2_X1 U10993 ( .A1(n10345), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n10346) );
  OAI211_X1 U10994 ( .C1(n10349), .C2(n10348), .A(n10347), .B(n10346), .ZN(
        P1_U3324) );
  OAI222_X1 U10995 ( .A1(n10354), .A2(n10353), .B1(n10352), .B2(P1_U3086), 
        .C1(n10351), .C2(n10350), .ZN(P1_U3326) );
  MUX2_X1 U10996 ( .A(n10355), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U10997 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10356), .ZN(P1_U3323) );
  AND2_X1 U10998 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10356), .ZN(P1_U3322) );
  AND2_X1 U10999 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10356), .ZN(P1_U3321) );
  AND2_X1 U11000 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10356), .ZN(P1_U3320) );
  AND2_X1 U11001 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10356), .ZN(P1_U3319) );
  AND2_X1 U11002 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10356), .ZN(P1_U3318) );
  AND2_X1 U11003 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10356), .ZN(P1_U3317) );
  AND2_X1 U11004 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10356), .ZN(P1_U3316) );
  AND2_X1 U11005 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10356), .ZN(P1_U3315) );
  AND2_X1 U11006 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10356), .ZN(P1_U3314) );
  AND2_X1 U11007 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10356), .ZN(P1_U3313) );
  AND2_X1 U11008 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10356), .ZN(P1_U3312) );
  AND2_X1 U11009 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10356), .ZN(P1_U3311) );
  AND2_X1 U11010 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10356), .ZN(P1_U3310) );
  AND2_X1 U11011 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10356), .ZN(P1_U3309) );
  AND2_X1 U11012 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10356), .ZN(P1_U3308) );
  AND2_X1 U11013 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10356), .ZN(P1_U3307) );
  AND2_X1 U11014 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10356), .ZN(P1_U3306) );
  AND2_X1 U11015 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10356), .ZN(P1_U3305) );
  AND2_X1 U11016 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10356), .ZN(P1_U3304) );
  AND2_X1 U11017 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10356), .ZN(P1_U3303) );
  AND2_X1 U11018 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10356), .ZN(P1_U3302) );
  AND2_X1 U11019 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10356), .ZN(P1_U3301) );
  AND2_X1 U11020 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10356), .ZN(P1_U3300) );
  AND2_X1 U11021 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10356), .ZN(P1_U3299) );
  AND2_X1 U11022 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10356), .ZN(P1_U3298) );
  AND2_X1 U11023 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10356), .ZN(P1_U3297) );
  AND2_X1 U11024 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10356), .ZN(P1_U3296) );
  AND2_X1 U11025 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10356), .ZN(P1_U3295) );
  AND2_X1 U11026 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10356), .ZN(P1_U3294) );
  INV_X1 U11027 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10564) );
  AOI22_X1 U11028 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_122), .B1(
        n10564), .B2(keyinput_125), .ZN(n10357) );
  OAI221_X1 U11029 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_122), .C1(
        n10564), .C2(keyinput_125), .A(n10357), .ZN(n10360) );
  AOI22_X1 U11030 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_123), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_124), .ZN(n10358) );
  OAI221_X1 U11031 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_123), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_124), .A(n10358), .ZN(n10359)
         );
  AOI211_X1 U11032 ( .C1(keyinput_126), .C2(P2_REG3_REG_26__SCAN_IN), .A(
        n10360), .B(n10359), .ZN(n10361) );
  OAI21_X1 U11033 ( .B1(keyinput_126), .B2(P2_REG3_REG_26__SCAN_IN), .A(n10361), .ZN(n10453) );
  AOI22_X1 U11034 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_112), .B1(
        n10460), .B2(keyinput_115), .ZN(n10362) );
  OAI221_X1 U11035 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_112), .C1(
        n10460), .C2(keyinput_115), .A(n10362), .ZN(n10365) );
  AOI22_X1 U11036 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_113), .B1(n10457), .B2(keyinput_114), .ZN(n10363) );
  OAI221_X1 U11037 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_113), .C1(
        n10457), .C2(keyinput_114), .A(n10363), .ZN(n10364) );
  AOI211_X1 U11038 ( .C1(keyinput_116), .C2(P2_REG3_REG_4__SCAN_IN), .A(n10365), .B(n10364), .ZN(n10366) );
  OAI21_X1 U11039 ( .B1(keyinput_116), .B2(P2_REG3_REG_4__SCAN_IN), .A(n10366), 
        .ZN(n10444) );
  INV_X1 U11040 ( .A(keyinput_111), .ZN(n10441) );
  INV_X1 U11041 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10465) );
  OAI22_X1 U11042 ( .A1(n10465), .A2(keyinput_103), .B1(
        P2_REG3_REG_23__SCAN_IN), .B2(keyinput_102), .ZN(n10367) );
  AOI221_X1 U11043 ( .B1(n10465), .B2(keyinput_103), .C1(keyinput_102), .C2(
        P2_REG3_REG_23__SCAN_IN), .A(n10367), .ZN(n10370) );
  OAI22_X1 U11044 ( .A1(n6587), .A2(keyinput_106), .B1(keyinput_104), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n10368) );
  AOI221_X1 U11045 ( .B1(n6587), .B2(keyinput_106), .C1(P2_REG3_REG_3__SCAN_IN), .C2(keyinput_104), .A(n10368), .ZN(n10369) );
  OAI211_X1 U11046 ( .C1(P2_REG3_REG_19__SCAN_IN), .C2(keyinput_105), .A(
        n10370), .B(n10369), .ZN(n10371) );
  AOI21_X1 U11047 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_105), .A(n10371), .ZN(n10439) );
  INV_X1 U11048 ( .A(keyinput_101), .ZN(n10432) );
  INV_X1 U11049 ( .A(keyinput_100), .ZN(n10430) );
  INV_X1 U11050 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10539) );
  INV_X1 U11051 ( .A(SI_10_), .ZN(n10475) );
  OAI22_X1 U11052 ( .A1(n10475), .A2(keyinput_86), .B1(SI_9_), .B2(keyinput_87), .ZN(n10372) );
  AOI221_X1 U11053 ( .B1(n10475), .B2(keyinput_86), .C1(keyinput_87), .C2(
        SI_9_), .A(n10372), .ZN(n10376) );
  OAI22_X1 U11054 ( .A1(n10374), .A2(keyinput_88), .B1(keyinput_85), .B2(
        SI_11_), .ZN(n10373) );
  AOI221_X1 U11055 ( .B1(n10374), .B2(keyinput_88), .C1(SI_11_), .C2(
        keyinput_85), .A(n10373), .ZN(n10375) );
  OAI211_X1 U11056 ( .C1(SI_7_), .C2(keyinput_89), .A(n10376), .B(n10375), 
        .ZN(n10377) );
  AOI21_X1 U11057 ( .B1(SI_7_), .B2(keyinput_89), .A(n10377), .ZN(n10408) );
  INV_X1 U11058 ( .A(keyinput_73), .ZN(n10391) );
  OAI22_X1 U11059 ( .A1(n10379), .A2(keyinput_72), .B1(keyinput_71), .B2(
        SI_25_), .ZN(n10378) );
  AOI221_X1 U11060 ( .B1(n10379), .B2(keyinput_72), .C1(SI_25_), .C2(
        keyinput_71), .A(n10378), .ZN(n10388) );
  INV_X1 U11061 ( .A(keyinput_66), .ZN(n10382) );
  OAI22_X1 U11062 ( .A1(SI_31_), .A2(keyinput_65), .B1(P2_WR_REG_SCAN_IN), 
        .B2(keyinput_64), .ZN(n10380) );
  AOI221_X1 U11063 ( .B1(SI_31_), .B2(keyinput_65), .C1(keyinput_64), .C2(
        P2_WR_REG_SCAN_IN), .A(n10380), .ZN(n10381) );
  AOI221_X1 U11064 ( .B1(SI_30_), .B2(n10382), .C1(n10484), .C2(keyinput_66), 
        .A(n10381), .ZN(n10385) );
  AOI22_X1 U11065 ( .A1(n10491), .A2(keyinput_68), .B1(keyinput_67), .B2(
        n10487), .ZN(n10383) );
  OAI221_X1 U11066 ( .B1(n10491), .B2(keyinput_68), .C1(n10487), .C2(
        keyinput_67), .A(n10383), .ZN(n10384) );
  AOI211_X1 U11067 ( .C1(SI_27_), .C2(keyinput_69), .A(n10385), .B(n10384), 
        .ZN(n10386) );
  OAI21_X1 U11068 ( .B1(SI_27_), .B2(keyinput_69), .A(n10386), .ZN(n10387) );
  OAI211_X1 U11069 ( .C1(SI_26_), .C2(keyinput_70), .A(n10388), .B(n10387), 
        .ZN(n10389) );
  AOI21_X1 U11070 ( .B1(SI_26_), .B2(keyinput_70), .A(n10389), .ZN(n10390) );
  AOI221_X1 U11071 ( .B1(SI_23_), .B2(n10391), .C1(n10498), .C2(keyinput_73), 
        .A(n10390), .ZN(n10406) );
  XNOR2_X1 U11072 ( .A(SI_22_), .B(keyinput_74), .ZN(n10405) );
  OAI22_X1 U11073 ( .A1(n10506), .A2(keyinput_77), .B1(n10393), .B2(
        keyinput_84), .ZN(n10392) );
  AOI221_X1 U11074 ( .B1(n10506), .B2(keyinput_77), .C1(keyinput_84), .C2(
        n10393), .A(n10392), .ZN(n10404) );
  AOI22_X1 U11075 ( .A1(SI_13_), .A2(keyinput_83), .B1(SI_20_), .B2(
        keyinput_76), .ZN(n10394) );
  OAI221_X1 U11076 ( .B1(SI_13_), .B2(keyinput_83), .C1(SI_20_), .C2(
        keyinput_76), .A(n10394), .ZN(n10402) );
  INV_X1 U11077 ( .A(SI_18_), .ZN(n10509) );
  AOI22_X1 U11078 ( .A1(SI_16_), .A2(keyinput_80), .B1(n10509), .B2(
        keyinput_78), .ZN(n10395) );
  OAI221_X1 U11079 ( .B1(SI_16_), .B2(keyinput_80), .C1(n10509), .C2(
        keyinput_78), .A(n10395), .ZN(n10401) );
  AOI22_X1 U11080 ( .A1(n10500), .A2(keyinput_79), .B1(n10397), .B2(
        keyinput_75), .ZN(n10396) );
  OAI221_X1 U11081 ( .B1(n10500), .B2(keyinput_79), .C1(n10397), .C2(
        keyinput_75), .A(n10396), .ZN(n10400) );
  AOI22_X1 U11082 ( .A1(SI_15_), .A2(keyinput_81), .B1(n10504), .B2(
        keyinput_82), .ZN(n10398) );
  OAI221_X1 U11083 ( .B1(SI_15_), .B2(keyinput_81), .C1(n10504), .C2(
        keyinput_82), .A(n10398), .ZN(n10399) );
  NOR4_X1 U11084 ( .A1(n10402), .A2(n10401), .A3(n10400), .A4(n10399), .ZN(
        n10403) );
  OAI211_X1 U11085 ( .C1(n10406), .C2(n10405), .A(n10404), .B(n10403), .ZN(
        n10407) );
  AOI22_X1 U11086 ( .A1(n10408), .A2(n10407), .B1(keyinput_90), .B2(SI_6_), 
        .ZN(n10409) );
  OAI21_X1 U11087 ( .B1(keyinput_90), .B2(SI_6_), .A(n10409), .ZN(n10417) );
  INV_X1 U11088 ( .A(keyinput_91), .ZN(n10410) );
  MUX2_X1 U11089 ( .A(n10410), .B(keyinput_91), .S(SI_5_), .Z(n10416) );
  XNOR2_X1 U11090 ( .A(n10411), .B(keyinput_93), .ZN(n10414) );
  XNOR2_X1 U11091 ( .A(SI_4_), .B(keyinput_92), .ZN(n10413) );
  XNOR2_X1 U11092 ( .A(SI_2_), .B(keyinput_94), .ZN(n10412) );
  NAND3_X1 U11093 ( .A1(n10414), .A2(n10413), .A3(n10412), .ZN(n10415) );
  AOI21_X1 U11094 ( .B1(n10417), .B2(n10416), .A(n10415), .ZN(n10420) );
  INV_X1 U11095 ( .A(keyinput_95), .ZN(n10418) );
  MUX2_X1 U11096 ( .A(keyinput_95), .B(n10418), .S(SI_1_), .Z(n10419) );
  NOR2_X1 U11097 ( .A1(n10420), .A2(n10419), .ZN(n10425) );
  AOI22_X1 U11098 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_98), .B1(n10422), 
        .B2(keyinput_97), .ZN(n10421) );
  OAI221_X1 U11099 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_98), .C1(n10422), 
        .C2(keyinput_97), .A(n10421), .ZN(n10424) );
  XOR2_X1 U11100 ( .A(SI_0_), .B(keyinput_96), .Z(n10423) );
  NOR3_X1 U11101 ( .A1(n10425), .A2(n10424), .A3(n10423), .ZN(n10428) );
  INV_X1 U11102 ( .A(keyinput_99), .ZN(n10426) );
  OAI22_X1 U11103 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(n10426), .B1(keyinput_99), 
        .B2(n6347), .ZN(n10427) );
  OR2_X1 U11104 ( .A1(n10428), .A2(n10427), .ZN(n10429) );
  OAI221_X1 U11105 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(n10430), .C1(n10539), 
        .C2(keyinput_100), .A(n10429), .ZN(n10431) );
  OAI221_X1 U11106 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_101), .C1(
        n10542), .C2(n10432), .A(n10431), .ZN(n10438) );
  INV_X1 U11107 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10434) );
  AOI22_X1 U11108 ( .A1(n10434), .A2(keyinput_107), .B1(n10545), .B2(
        keyinput_110), .ZN(n10433) );
  OAI221_X1 U11109 ( .B1(n10434), .B2(keyinput_107), .C1(n10545), .C2(
        keyinput_110), .A(n10433), .ZN(n10437) );
  AOI22_X1 U11110 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_108), .B1(
        P2_REG3_REG_21__SCAN_IN), .B2(keyinput_109), .ZN(n10435) );
  OAI221_X1 U11111 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_108), .C1(
        P2_REG3_REG_21__SCAN_IN), .C2(keyinput_109), .A(n10435), .ZN(n10436)
         );
  AOI211_X1 U11112 ( .C1(n10439), .C2(n10438), .A(n10437), .B(n10436), .ZN(
        n10440) );
  AOI221_X1 U11113 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n10441), .C1(n6568), 
        .C2(keyinput_111), .A(n10440), .ZN(n10443) );
  NAND2_X1 U11114 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_117), .ZN(n10442) );
  OAI221_X1 U11115 ( .B1(n10444), .B2(n10443), .C1(P2_REG3_REG_9__SCAN_IN), 
        .C2(keyinput_117), .A(n10442), .ZN(n10447) );
  INV_X1 U11116 ( .A(keyinput_118), .ZN(n10445) );
  MUX2_X1 U11117 ( .A(n10445), .B(keyinput_118), .S(P2_REG3_REG_0__SCAN_IN), 
        .Z(n10446) );
  NAND2_X1 U11118 ( .A1(n10447), .A2(n10446), .ZN(n10450) );
  OAI22_X1 U11119 ( .A1(n9093), .A2(keyinput_119), .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_121), .ZN(n10448) );
  AOI221_X1 U11120 ( .B1(n9093), .B2(keyinput_119), .C1(keyinput_121), .C2(
        P2_REG3_REG_22__SCAN_IN), .A(n10448), .ZN(n10449) );
  OAI211_X1 U11121 ( .C1(P2_REG3_REG_13__SCAN_IN), .C2(keyinput_120), .A(
        n10450), .B(n10449), .ZN(n10451) );
  AOI21_X1 U11122 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_120), .A(n10451), .ZN(n10452) );
  OAI22_X1 U11123 ( .A1(n10453), .A2(n10452), .B1(keyinput_127), .B2(
        P2_REG3_REG_15__SCAN_IN), .ZN(n10454) );
  AOI21_X1 U11124 ( .B1(keyinput_127), .B2(P2_REG3_REG_15__SCAN_IN), .A(n10454), .ZN(n10573) );
  AOI22_X1 U11125 ( .A1(n10457), .A2(keyinput_50), .B1(keyinput_52), .B2(
        n10456), .ZN(n10455) );
  OAI221_X1 U11126 ( .B1(n10457), .B2(keyinput_50), .C1(n10456), .C2(
        keyinput_52), .A(n10455), .ZN(n10462) );
  AOI22_X1 U11127 ( .A1(n10460), .A2(keyinput_51), .B1(keyinput_49), .B2(
        n10459), .ZN(n10458) );
  OAI221_X1 U11128 ( .B1(n10460), .B2(keyinput_51), .C1(n10459), .C2(
        keyinput_49), .A(n10458), .ZN(n10461) );
  AOI211_X1 U11129 ( .C1(keyinput_48), .C2(P2_REG3_REG_16__SCAN_IN), .A(n10462), .B(n10461), .ZN(n10463) );
  OAI21_X1 U11130 ( .B1(keyinput_48), .B2(P2_REG3_REG_16__SCAN_IN), .A(n10463), 
        .ZN(n10555) );
  INV_X1 U11131 ( .A(keyinput_47), .ZN(n10552) );
  AOI22_X1 U11132 ( .A1(n10466), .A2(keyinput_40), .B1(n10465), .B2(
        keyinput_39), .ZN(n10464) );
  OAI221_X1 U11133 ( .B1(n10466), .B2(keyinput_40), .C1(n10465), .C2(
        keyinput_39), .A(n10464), .ZN(n10471) );
  OAI22_X1 U11134 ( .A1(n10468), .A2(keyinput_41), .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_38), .ZN(n10467) );
  AOI221_X1 U11135 ( .B1(n10468), .B2(keyinput_41), .C1(keyinput_38), .C2(
        P2_REG3_REG_23__SCAN_IN), .A(n10467), .ZN(n10469) );
  OAI21_X1 U11136 ( .B1(keyinput_42), .B2(P2_REG3_REG_28__SCAN_IN), .A(n10469), 
        .ZN(n10470) );
  AOI211_X1 U11137 ( .C1(keyinput_42), .C2(P2_REG3_REG_28__SCAN_IN), .A(n10471), .B(n10470), .ZN(n10550) );
  INV_X1 U11138 ( .A(keyinput_37), .ZN(n10541) );
  INV_X1 U11139 ( .A(keyinput_36), .ZN(n10538) );
  INV_X1 U11140 ( .A(keyinput_35), .ZN(n10536) );
  AOI22_X1 U11141 ( .A1(SI_0_), .A2(keyinput_32), .B1(P2_RD_REG_SCAN_IN), .B2(
        keyinput_33), .ZN(n10472) );
  OAI221_X1 U11142 ( .B1(SI_0_), .B2(keyinput_32), .C1(P2_RD_REG_SCAN_IN), 
        .C2(keyinput_33), .A(n10472), .ZN(n10533) );
  OAI22_X1 U11143 ( .A1(SI_8_), .A2(keyinput_24), .B1(keyinput_25), .B2(SI_7_), 
        .ZN(n10473) );
  AOI221_X1 U11144 ( .B1(SI_8_), .B2(keyinput_24), .C1(SI_7_), .C2(keyinput_25), .A(n10473), .ZN(n10477) );
  OAI22_X1 U11145 ( .A1(n10475), .A2(keyinput_22), .B1(SI_9_), .B2(keyinput_23), .ZN(n10474) );
  AOI221_X1 U11146 ( .B1(n10475), .B2(keyinput_22), .C1(keyinput_23), .C2(
        SI_9_), .A(n10474), .ZN(n10476) );
  OAI211_X1 U11147 ( .C1(SI_11_), .C2(keyinput_21), .A(n10477), .B(n10476), 
        .ZN(n10478) );
  AOI21_X1 U11148 ( .B1(SI_11_), .B2(keyinput_21), .A(n10478), .ZN(n10519) );
  INV_X1 U11149 ( .A(keyinput_9), .ZN(n10497) );
  OAI22_X1 U11150 ( .A1(n10480), .A2(keyinput_7), .B1(SI_24_), .B2(keyinput_8), 
        .ZN(n10479) );
  AOI221_X1 U11151 ( .B1(n10480), .B2(keyinput_7), .C1(keyinput_8), .C2(SI_24_), .A(n10479), .ZN(n10493) );
  INV_X1 U11152 ( .A(keyinput_2), .ZN(n10483) );
  OAI22_X1 U11153 ( .A1(SI_31_), .A2(keyinput_1), .B1(P2_WR_REG_SCAN_IN), .B2(
        keyinput_0), .ZN(n10481) );
  AOI221_X1 U11154 ( .B1(SI_31_), .B2(keyinput_1), .C1(keyinput_0), .C2(
        P2_WR_REG_SCAN_IN), .A(n10481), .ZN(n10482) );
  AOI221_X1 U11155 ( .B1(SI_30_), .B2(keyinput_2), .C1(n10484), .C2(n10483), 
        .A(n10482), .ZN(n10489) );
  AOI22_X1 U11156 ( .A1(n10487), .A2(keyinput_3), .B1(n10486), .B2(keyinput_5), 
        .ZN(n10485) );
  OAI221_X1 U11157 ( .B1(n10487), .B2(keyinput_3), .C1(n10486), .C2(keyinput_5), .A(n10485), .ZN(n10488) );
  AOI211_X1 U11158 ( .C1(n10491), .C2(keyinput_4), .A(n10489), .B(n10488), 
        .ZN(n10490) );
  OAI21_X1 U11159 ( .B1(n10491), .B2(keyinput_4), .A(n10490), .ZN(n10492) );
  OAI211_X1 U11160 ( .C1(n10495), .C2(keyinput_6), .A(n10493), .B(n10492), 
        .ZN(n10494) );
  AOI21_X1 U11161 ( .B1(n10495), .B2(keyinput_6), .A(n10494), .ZN(n10496) );
  AOI221_X1 U11162 ( .B1(SI_23_), .B2(keyinput_9), .C1(n10498), .C2(n10497), 
        .A(n10496), .ZN(n10517) );
  XOR2_X1 U11163 ( .A(SI_22_), .B(keyinput_10), .Z(n10516) );
  OAI22_X1 U11164 ( .A1(n10501), .A2(keyinput_12), .B1(n10500), .B2(
        keyinput_15), .ZN(n10499) );
  AOI221_X1 U11165 ( .B1(n10501), .B2(keyinput_12), .C1(keyinput_15), .C2(
        n10500), .A(n10499), .ZN(n10515) );
  AOI22_X1 U11166 ( .A1(SI_15_), .A2(keyinput_17), .B1(SI_16_), .B2(
        keyinput_16), .ZN(n10502) );
  OAI221_X1 U11167 ( .B1(SI_15_), .B2(keyinput_17), .C1(SI_16_), .C2(
        keyinput_16), .A(n10502), .ZN(n10513) );
  AOI22_X1 U11168 ( .A1(SI_21_), .A2(keyinput_11), .B1(n10504), .B2(
        keyinput_18), .ZN(n10503) );
  OAI221_X1 U11169 ( .B1(SI_21_), .B2(keyinput_11), .C1(n10504), .C2(
        keyinput_18), .A(n10503), .ZN(n10512) );
  INV_X1 U11170 ( .A(SI_13_), .ZN(n10507) );
  AOI22_X1 U11171 ( .A1(n10507), .A2(keyinput_19), .B1(n10506), .B2(
        keyinput_13), .ZN(n10505) );
  OAI221_X1 U11172 ( .B1(n10507), .B2(keyinput_19), .C1(n10506), .C2(
        keyinput_13), .A(n10505), .ZN(n10511) );
  AOI22_X1 U11173 ( .A1(SI_12_), .A2(keyinput_20), .B1(n10509), .B2(
        keyinput_14), .ZN(n10508) );
  OAI221_X1 U11174 ( .B1(SI_12_), .B2(keyinput_20), .C1(n10509), .C2(
        keyinput_14), .A(n10508), .ZN(n10510) );
  NOR4_X1 U11175 ( .A1(n10513), .A2(n10512), .A3(n10511), .A4(n10510), .ZN(
        n10514) );
  OAI211_X1 U11176 ( .C1(n10517), .C2(n10516), .A(n10515), .B(n10514), .ZN(
        n10518) );
  AOI22_X1 U11177 ( .A1(n10519), .A2(n10518), .B1(keyinput_26), .B2(SI_6_), 
        .ZN(n10520) );
  OAI21_X1 U11178 ( .B1(keyinput_26), .B2(SI_6_), .A(n10520), .ZN(n10528) );
  INV_X1 U11179 ( .A(keyinput_27), .ZN(n10521) );
  MUX2_X1 U11180 ( .A(n10521), .B(keyinput_27), .S(SI_5_), .Z(n10527) );
  XNOR2_X1 U11181 ( .A(n10522), .B(keyinput_30), .ZN(n10525) );
  XNOR2_X1 U11182 ( .A(SI_3_), .B(keyinput_29), .ZN(n10524) );
  XNOR2_X1 U11183 ( .A(SI_4_), .B(keyinput_28), .ZN(n10523) );
  NAND3_X1 U11184 ( .A1(n10525), .A2(n10524), .A3(n10523), .ZN(n10526) );
  AOI21_X1 U11185 ( .B1(n10528), .B2(n10527), .A(n10526), .ZN(n10531) );
  INV_X1 U11186 ( .A(keyinput_31), .ZN(n10529) );
  MUX2_X1 U11187 ( .A(keyinput_31), .B(n10529), .S(SI_1_), .Z(n10530) );
  NOR2_X1 U11188 ( .A1(n10531), .A2(n10530), .ZN(n10532) );
  AOI211_X1 U11189 ( .C1(P2_STATE_REG_SCAN_IN), .C2(keyinput_34), .A(n10533), 
        .B(n10532), .ZN(n10534) );
  OAI21_X1 U11190 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_34), .A(n10534), 
        .ZN(n10535) );
  OAI221_X1 U11191 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_35), .C1(n6347), 
        .C2(n10536), .A(n10535), .ZN(n10537) );
  OAI221_X1 U11192 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_36), .C1(
        n10539), .C2(n10538), .A(n10537), .ZN(n10540) );
  OAI221_X1 U11193 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_37), .C1(
        n10542), .C2(n10541), .A(n10540), .ZN(n10549) );
  AOI22_X1 U11194 ( .A1(n10545), .A2(keyinput_46), .B1(n10544), .B2(
        keyinput_45), .ZN(n10543) );
  OAI221_X1 U11195 ( .B1(n10545), .B2(keyinput_46), .C1(n10544), .C2(
        keyinput_45), .A(n10543), .ZN(n10548) );
  AOI22_X1 U11196 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_43), .B1(n10674), 
        .B2(keyinput_44), .ZN(n10546) );
  OAI221_X1 U11197 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_43), .C1(n10674), .C2(keyinput_44), .A(n10546), .ZN(n10547) );
  AOI211_X1 U11198 ( .C1(n10550), .C2(n10549), .A(n10548), .B(n10547), .ZN(
        n10551) );
  AOI221_X1 U11199 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n10552), .C1(n6568), 
        .C2(keyinput_47), .A(n10551), .ZN(n10554) );
  NAND2_X1 U11200 ( .A1(n6378), .A2(keyinput_53), .ZN(n10553) );
  OAI221_X1 U11201 ( .B1(n10555), .B2(n10554), .C1(n6378), .C2(keyinput_53), 
        .A(n10553), .ZN(n10558) );
  INV_X1 U11202 ( .A(keyinput_54), .ZN(n10556) );
  MUX2_X1 U11203 ( .A(n10556), .B(keyinput_54), .S(P2_REG3_REG_0__SCAN_IN), 
        .Z(n10557) );
  NAND2_X1 U11204 ( .A1(n10558), .A2(n10557), .ZN(n10561) );
  OAI22_X1 U11205 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_55), .B1(
        keyinput_56), .B2(P2_REG3_REG_13__SCAN_IN), .ZN(n10559) );
  AOI221_X1 U11206 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_55), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_56), .A(n10559), .ZN(n10560) );
  OAI211_X1 U11207 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(keyinput_57), .A(n10561), .B(n10560), .ZN(n10562) );
  AOI21_X1 U11208 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_57), .A(n10562), 
        .ZN(n10571) );
  AOI22_X1 U11209 ( .A1(n10693), .A2(keyinput_58), .B1(keyinput_61), .B2(
        n10564), .ZN(n10563) );
  OAI221_X1 U11210 ( .B1(n10693), .B2(keyinput_58), .C1(n10564), .C2(
        keyinput_61), .A(n10563), .ZN(n10568) );
  INV_X1 U11211 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U11212 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_59), .B1(n10566), 
        .B2(keyinput_62), .ZN(n10565) );
  OAI221_X1 U11213 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_59), .C1(n10566), .C2(keyinput_62), .A(n10565), .ZN(n10567) );
  AOI211_X1 U11214 ( .C1(keyinput_60), .C2(P2_REG3_REG_18__SCAN_IN), .A(n10568), .B(n10567), .ZN(n10569) );
  OAI21_X1 U11215 ( .B1(keyinput_60), .B2(P2_REG3_REG_18__SCAN_IN), .A(n10569), 
        .ZN(n10570) );
  OAI22_X1 U11216 ( .A1(n10571), .A2(n10570), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(keyinput_63), .ZN(n10572) );
  AOI211_X1 U11217 ( .C1(P2_REG3_REG_15__SCAN_IN), .C2(keyinput_63), .A(n10573), .B(n10572), .ZN(n10578) );
  MUX2_X1 U11218 ( .A(n10576), .B(n10575), .S(n10574), .Z(n10577) );
  XNOR2_X1 U11219 ( .A(n10578), .B(n10577), .ZN(P2_U3506) );
  XOR2_X1 U11220 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  INV_X1 U11221 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10582) );
  NAND3_X1 U11222 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10581) );
  AND2_X1 U11223 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n10579) );
  NOR2_X1 U11224 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10579), .ZN(n10580) );
  INV_X1 U11225 ( .A(n10580), .ZN(n10584) );
  NAND2_X1 U11226 ( .A1(n10582), .A2(n10581), .ZN(n10583) );
  OAI222_X1 U11227 ( .A1(n10582), .A2(n10581), .B1(n10582), .B2(n10584), .C1(
        n10580), .C2(n10583), .ZN(ADD_1068_U5) );
  NAND2_X1 U11228 ( .A1(n10584), .A2(n10583), .ZN(n10587) );
  NAND2_X1 U11229 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10585) );
  OAI21_X1 U11230 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10585), .ZN(n10586) );
  NOR2_X1 U11231 ( .A1(n10587), .A2(n10586), .ZN(n10588) );
  AOI21_X1 U11232 ( .B1(n10587), .B2(n10586), .A(n10588), .ZN(ADD_1068_U54) );
  AOI21_X1 U11233 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10588), .ZN(n10591) );
  NAND2_X1 U11234 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n10589) );
  OAI21_X1 U11235 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10589), .ZN(n10590) );
  NOR2_X1 U11236 ( .A1(n10591), .A2(n10590), .ZN(n10592) );
  AOI21_X1 U11237 ( .B1(n10591), .B2(n10590), .A(n10592), .ZN(ADD_1068_U53) );
  AOI21_X1 U11238 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10592), .ZN(n10595) );
  NOR2_X1 U11239 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10593) );
  AOI21_X1 U11240 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10593), .ZN(n10594) );
  NAND2_X1 U11241 ( .A1(n10595), .A2(n10594), .ZN(n10597) );
  OAI21_X1 U11242 ( .B1(n10595), .B2(n10594), .A(n10597), .ZN(ADD_1068_U52) );
  NOR2_X1 U11243 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10596) );
  AOI21_X1 U11244 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10596), .ZN(n10599) );
  OAI21_X1 U11245 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10597), .ZN(n10598) );
  NAND2_X1 U11246 ( .A1(n10599), .A2(n10598), .ZN(n10601) );
  OAI21_X1 U11247 ( .B1(n10599), .B2(n10598), .A(n10601), .ZN(ADD_1068_U51) );
  NOR2_X1 U11248 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10600) );
  AOI21_X1 U11249 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10600), .ZN(n10603) );
  OAI21_X1 U11250 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10601), .ZN(n10602) );
  NAND2_X1 U11251 ( .A1(n10603), .A2(n10602), .ZN(n10605) );
  OAI21_X1 U11252 ( .B1(n10603), .B2(n10602), .A(n10605), .ZN(ADD_1068_U50) );
  NOR2_X1 U11253 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10604) );
  AOI21_X1 U11254 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n10604), .ZN(n10607) );
  OAI21_X1 U11255 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10605), .ZN(n10606) );
  NAND2_X1 U11256 ( .A1(n10607), .A2(n10606), .ZN(n10609) );
  OAI21_X1 U11257 ( .B1(n10607), .B2(n10606), .A(n10609), .ZN(ADD_1068_U49) );
  NOR2_X1 U11258 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10608) );
  AOI21_X1 U11259 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n10608), .ZN(n10611) );
  OAI21_X1 U11260 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10609), .ZN(n10610) );
  NAND2_X1 U11261 ( .A1(n10611), .A2(n10610), .ZN(n10613) );
  OAI21_X1 U11262 ( .B1(n10611), .B2(n10610), .A(n10613), .ZN(ADD_1068_U48) );
  NOR2_X1 U11263 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10612) );
  AOI21_X1 U11264 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n10612), .ZN(n10615) );
  OAI21_X1 U11265 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10613), .ZN(n10614) );
  NAND2_X1 U11266 ( .A1(n10615), .A2(n10614), .ZN(n10617) );
  OAI21_X1 U11267 ( .B1(n10615), .B2(n10614), .A(n10617), .ZN(ADD_1068_U47) );
  NOR2_X1 U11268 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10616) );
  AOI21_X1 U11269 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10616), .ZN(n10619) );
  OAI21_X1 U11270 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10617), .ZN(n10618) );
  NAND2_X1 U11271 ( .A1(n10619), .A2(n10618), .ZN(n10621) );
  OAI21_X1 U11272 ( .B1(n10619), .B2(n10618), .A(n10621), .ZN(ADD_1068_U63) );
  NOR2_X1 U11273 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10620) );
  AOI21_X1 U11274 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10620), .ZN(n10623) );
  OAI21_X1 U11275 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10621), .ZN(n10622) );
  NAND2_X1 U11276 ( .A1(n10623), .A2(n10622), .ZN(n10625) );
  OAI21_X1 U11277 ( .B1(n10623), .B2(n10622), .A(n10625), .ZN(ADD_1068_U62) );
  NOR2_X1 U11278 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10624) );
  AOI21_X1 U11279 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10624), .ZN(n10627) );
  OAI21_X1 U11280 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10625), .ZN(n10626) );
  NAND2_X1 U11281 ( .A1(n10627), .A2(n10626), .ZN(n10629) );
  OAI21_X1 U11282 ( .B1(n10627), .B2(n10626), .A(n10629), .ZN(ADD_1068_U61) );
  NOR2_X1 U11283 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10628) );
  AOI21_X1 U11284 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10628), .ZN(n10631) );
  OAI21_X1 U11285 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10629), .ZN(n10630) );
  NAND2_X1 U11286 ( .A1(n10631), .A2(n10630), .ZN(n10633) );
  OAI21_X1 U11287 ( .B1(n10631), .B2(n10630), .A(n10633), .ZN(ADD_1068_U60) );
  NOR2_X1 U11288 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10632) );
  AOI21_X1 U11289 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10632), .ZN(n10635) );
  OAI21_X1 U11290 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10633), .ZN(n10634) );
  NAND2_X1 U11291 ( .A1(n10635), .A2(n10634), .ZN(n10637) );
  OAI21_X1 U11292 ( .B1(n10635), .B2(n10634), .A(n10637), .ZN(ADD_1068_U59) );
  NOR2_X1 U11293 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10636) );
  AOI21_X1 U11294 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10636), .ZN(n10639) );
  OAI21_X1 U11295 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10637), .ZN(n10638) );
  NAND2_X1 U11296 ( .A1(n10639), .A2(n10638), .ZN(n10641) );
  OAI21_X1 U11297 ( .B1(n10639), .B2(n10638), .A(n10641), .ZN(ADD_1068_U58) );
  NOR2_X1 U11298 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10640) );
  AOI21_X1 U11299 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10640), .ZN(n10643) );
  OAI21_X1 U11300 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10641), .ZN(n10642) );
  NAND2_X1 U11301 ( .A1(n10643), .A2(n10642), .ZN(n10645) );
  OAI21_X1 U11302 ( .B1(n10643), .B2(n10642), .A(n10645), .ZN(ADD_1068_U57) );
  NOR2_X1 U11303 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10644) );
  AOI21_X1 U11304 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10644), .ZN(n10647) );
  OAI21_X1 U11305 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10645), .ZN(n10646) );
  NAND2_X1 U11306 ( .A1(n10647), .A2(n10646), .ZN(n10649) );
  OAI21_X1 U11307 ( .B1(n10647), .B2(n10646), .A(n10649), .ZN(ADD_1068_U56) );
  NOR2_X1 U11308 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n10648) );
  AOI21_X1 U11309 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n10648), .ZN(n10651) );
  OAI21_X1 U11310 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10649), .ZN(n10650) );
  NAND2_X1 U11311 ( .A1(n10651), .A2(n10650), .ZN(n10652) );
  OAI21_X1 U11312 ( .B1(n10651), .B2(n10650), .A(n10652), .ZN(ADD_1068_U55) );
  OAI21_X1 U11313 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10652), .ZN(n10654) );
  XOR2_X1 U11314 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .Z(n10653) );
  XNOR2_X1 U11315 ( .A(n10654), .B(n10653), .ZN(ADD_1068_U4) );
  NAND2_X1 U11316 ( .A1(n10676), .A2(n10655), .ZN(n10667) );
  NAND2_X1 U11317 ( .A1(n10698), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n10666) );
  INV_X1 U11318 ( .A(n10656), .ZN(n10657) );
  OAI211_X1 U11319 ( .C1(n10659), .C2(n10658), .A(n10657), .B(n10690), .ZN(
        n10665) );
  AND2_X1 U11320 ( .A1(n10660), .A2(n6250), .ZN(n10662) );
  INV_X1 U11321 ( .A(n10713), .ZN(n10661) );
  OAI21_X1 U11322 ( .B1(n10663), .B2(n10662), .A(n10661), .ZN(n10664) );
  AND4_X1 U11323 ( .A1(n10667), .A2(n10666), .A3(n10665), .A4(n10664), .ZN(
        n10673) );
  INV_X1 U11324 ( .A(n10668), .ZN(n10669) );
  AOI21_X1 U11325 ( .B1(n6246), .B2(n10670), .A(n10669), .ZN(n10671) );
  OR2_X1 U11326 ( .A1(n10682), .A2(n10671), .ZN(n10672) );
  OAI211_X1 U11327 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10674), .A(n10673), .B(
        n10672), .ZN(P2_U3183) );
  AOI22_X1 U11328 ( .A1(n10698), .A2(P2_ADDR_REG_11__SCAN_IN), .B1(n10676), 
        .B2(n10675), .ZN(n10692) );
  OAI21_X1 U11329 ( .B1(n10679), .B2(n10678), .A(n10677), .ZN(n10689) );
  AOI21_X1 U11330 ( .B1(n6401), .B2(n10681), .A(n10680), .ZN(n10683) );
  NOR2_X1 U11331 ( .A1(n10683), .A2(n10682), .ZN(n10688) );
  AOI21_X1 U11332 ( .B1(n6404), .B2(n10685), .A(n10684), .ZN(n10686) );
  NOR2_X1 U11333 ( .A1(n10686), .A2(n10713), .ZN(n10687) );
  AOI211_X1 U11334 ( .C1(n10690), .C2(n10689), .A(n10688), .B(n10687), .ZN(
        n10691) );
  OAI211_X1 U11335 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10693), .A(n10692), .B(
        n10691), .ZN(P2_U3193) );
  INV_X1 U11336 ( .A(n10694), .ZN(n10704) );
  INV_X1 U11337 ( .A(n10705), .ZN(n10696) );
  AOI211_X1 U11338 ( .C1(n10704), .C2(n10703), .A(n10696), .B(n10695), .ZN(
        n10697) );
  AOI21_X1 U11339 ( .B1(n10698), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n10697), 
        .ZN(n10719) );
  NOR2_X1 U11340 ( .A1(n10700), .A2(n10699), .ZN(n10702) );
  XOR2_X1 U11341 ( .A(n10702), .B(n10701), .Z(n10709) );
  NAND3_X1 U11342 ( .A1(n10704), .A2(P2_U3893), .A3(n10703), .ZN(n10707) );
  AOI21_X1 U11343 ( .B1(n10707), .B2(n10706), .A(n10705), .ZN(n10708) );
  AOI21_X1 U11344 ( .B1(n10710), .B2(n10709), .A(n10708), .ZN(n10718) );
  AND2_X1 U11345 ( .A1(n10712), .A2(n10711), .ZN(n10714) );
  XNOR2_X1 U11346 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  NOR2_X1 U11347 ( .A1(n10734), .A2(n10720), .ZN(n10731) );
  NOR2_X1 U11348 ( .A1(n10721), .A2(n10794), .ZN(n10737) );
  INV_X1 U11349 ( .A(n10737), .ZN(n10727) );
  AND2_X1 U11350 ( .A1(n10723), .A2(n10722), .ZN(n10736) );
  INV_X1 U11351 ( .A(n10724), .ZN(n10725) );
  NAND2_X1 U11352 ( .A1(n10736), .A2(n10725), .ZN(n10726) );
  OAI211_X1 U11353 ( .C1(n10729), .C2(n10728), .A(n10727), .B(n10726), .ZN(
        n10730) );
  NOR2_X1 U11354 ( .A1(n10731), .A2(n10730), .ZN(n10733) );
  AOI22_X1 U11355 ( .A1(n10820), .A2(n5734), .B1(n10733), .B2(n10732), .ZN(
        P1_U3293) );
  AOI21_X1 U11356 ( .B1(n10735), .B2(n10791), .A(n10734), .ZN(n10738) );
  NOR3_X1 U11357 ( .A1(n10738), .A2(n10737), .A3(n10736), .ZN(n10740) );
  AOI22_X1 U11358 ( .A1(n10831), .A2(n10740), .B1(n10739), .B2(n10830), .ZN(
        P1_U3522) );
  AOI22_X1 U11359 ( .A1(n10834), .A2(n10740), .B1(n5736), .B2(n6207), .ZN(
        P1_U3453) );
  AOI22_X1 U11360 ( .A1(n10852), .A2(n10741), .B1(n6244), .B2(n10850), .ZN(
        P2_U3393) );
  OAI21_X1 U11361 ( .B1(n10743), .B2(n10824), .A(n10742), .ZN(n10745) );
  AOI211_X1 U11362 ( .C1(n5053), .C2(n10746), .A(n10745), .B(n10744), .ZN(
        n10747) );
  AOI22_X1 U11363 ( .A1(n10831), .A2(n10747), .B1(n6952), .B2(n10830), .ZN(
        P1_U3524) );
  AOI22_X1 U11364 ( .A1(n10834), .A2(n10747), .B1(n5749), .B2(n6207), .ZN(
        P1_U3459) );
  AOI22_X1 U11365 ( .A1(n10852), .A2(n10748), .B1(n6276), .B2(n10850), .ZN(
        P2_U3396) );
  INV_X1 U11366 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U11367 ( .A1(n10852), .A2(n10750), .B1(n10749), .B2(n10850), .ZN(
        P2_U3399) );
  INV_X1 U11368 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10751) );
  AOI22_X1 U11369 ( .A1(n10852), .A2(n10752), .B1(n10751), .B2(n10850), .ZN(
        P2_U3402) );
  INV_X1 U11370 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10753) );
  AOI22_X1 U11371 ( .A1(n10852), .A2(n10754), .B1(n10753), .B2(n10850), .ZN(
        P2_U3405) );
  OAI21_X1 U11372 ( .B1(n10756), .B2(n10824), .A(n10755), .ZN(n10758) );
  AOI211_X1 U11373 ( .C1(n5053), .C2(n10759), .A(n10758), .B(n10757), .ZN(
        n10760) );
  AOI22_X1 U11374 ( .A1(n10831), .A2(n10760), .B1(n5797), .B2(n10830), .ZN(
        P1_U3527) );
  AOI22_X1 U11375 ( .A1(n10834), .A2(n10760), .B1(n5802), .B2(n6207), .ZN(
        P1_U3468) );
  INV_X1 U11376 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10761) );
  AOI22_X1 U11377 ( .A1(n10852), .A2(n10762), .B1(n10761), .B2(n10850), .ZN(
        P2_U3408) );
  INV_X1 U11378 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10763) );
  AOI22_X1 U11379 ( .A1(n10852), .A2(n10764), .B1(n10763), .B2(n10850), .ZN(
        P2_U3414) );
  INV_X1 U11380 ( .A(n10844), .ZN(n10767) );
  OAI21_X1 U11381 ( .B1(n10767), .B2(n10766), .A(n10765), .ZN(n10772) );
  AOI222_X1 U11382 ( .A1(n10846), .A2(n10772), .B1(n10771), .B2(n10770), .C1(
        n10769), .C2(n10768), .ZN(n10773) );
  OAI21_X1 U11383 ( .B1(n10846), .B2(n6376), .A(n10773), .ZN(P2_U3224) );
  INV_X1 U11384 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U11385 ( .A1(n10852), .A2(n10775), .B1(n10774), .B2(n10850), .ZN(
        P2_U3420) );
  INV_X1 U11386 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10776) );
  AOI22_X1 U11387 ( .A1(n10852), .A2(n10777), .B1(n10776), .B2(n10850), .ZN(
        P2_U3423) );
  INV_X1 U11388 ( .A(n10778), .ZN(n10803) );
  XNOR2_X1 U11389 ( .A(n10780), .B(n10779), .ZN(n10816) );
  INV_X1 U11390 ( .A(n10781), .ZN(n10783) );
  OAI211_X1 U11391 ( .C1(n10785), .C2(n10784), .A(n10783), .B(n10782), .ZN(
        n10812) );
  OAI21_X1 U11392 ( .B1(n10785), .B2(n10824), .A(n10812), .ZN(n10802) );
  INV_X1 U11393 ( .A(n10786), .ZN(n10800) );
  INV_X1 U11394 ( .A(n10787), .ZN(n10793) );
  AOI21_X1 U11395 ( .B1(n10790), .B2(n10789), .A(n10788), .ZN(n10792) );
  NOR3_X1 U11396 ( .A1(n10793), .A2(n10792), .A3(n10791), .ZN(n10799) );
  OAI22_X1 U11397 ( .A1(n10797), .A2(n10796), .B1(n10795), .B2(n10794), .ZN(
        n10798) );
  AOI211_X1 U11398 ( .C1(n10816), .C2(n10800), .A(n10799), .B(n10798), .ZN(
        n10819) );
  INV_X1 U11399 ( .A(n10819), .ZN(n10801) );
  AOI211_X1 U11400 ( .C1(n10803), .C2(n10816), .A(n10802), .B(n10801), .ZN(
        n10805) );
  AOI22_X1 U11401 ( .A1(n10831), .A2(n10805), .B1(n7305), .B2(n10830), .ZN(
        P1_U3533) );
  INV_X1 U11402 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10804) );
  AOI22_X1 U11403 ( .A1(n10834), .A2(n10805), .B1(n10804), .B2(n6207), .ZN(
        P1_U3486) );
  INV_X1 U11404 ( .A(n10806), .ZN(n10808) );
  AOI222_X1 U11405 ( .A1(n10810), .A2(n10809), .B1(n10808), .B2(n10807), .C1(
        P1_REG2_REG_11__SCAN_IN), .C2(n10820), .ZN(n10818) );
  NOR2_X1 U11406 ( .A1(n10820), .A2(n10811), .ZN(n10815) );
  INV_X1 U11407 ( .A(n10812), .ZN(n10813) );
  AOI22_X1 U11408 ( .A1(n10816), .A2(n10815), .B1(n10814), .B2(n10813), .ZN(
        n10817) );
  OAI211_X1 U11409 ( .C1(n10820), .C2(n10819), .A(n10818), .B(n10817), .ZN(
        P1_U3282) );
  INV_X1 U11410 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U11411 ( .A1(n10852), .A2(n10822), .B1(n10821), .B2(n10850), .ZN(
        P2_U3426) );
  OAI21_X1 U11412 ( .B1(n10825), .B2(n10824), .A(n10823), .ZN(n10826) );
  AOI211_X1 U11413 ( .C1(n10829), .C2(n5053), .A(n10827), .B(n10826), .ZN(
        n10833) );
  AOI22_X1 U11414 ( .A1(n10831), .A2(n10833), .B1(n5699), .B2(n10830), .ZN(
        P1_U3534) );
  INV_X1 U11415 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10832) );
  AOI22_X1 U11416 ( .A1(n10834), .A2(n10833), .B1(n10832), .B2(n6207), .ZN(
        P1_U3489) );
  INV_X1 U11417 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10835) );
  AOI22_X1 U11418 ( .A1(n10852), .A2(n10836), .B1(n10835), .B2(n10850), .ZN(
        P2_U3429) );
  INV_X1 U11419 ( .A(n10837), .ZN(n10845) );
  OAI22_X1 U11420 ( .A1(n10841), .A2(n10840), .B1(n10839), .B2(n10838), .ZN(
        n10843) );
  AOI211_X1 U11421 ( .C1(n10845), .C2(n10844), .A(n10843), .B(n10842), .ZN(
        n10847) );
  AOI22_X1 U11422 ( .A1(n4949), .A2(n9171), .B1(n10847), .B2(n10846), .ZN(
        P2_U3219) );
  INV_X1 U11423 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10848) );
  AOI22_X1 U11424 ( .A1(n10852), .A2(n10849), .B1(n10848), .B2(n10850), .ZN(
        P2_U3432) );
  AOI22_X1 U11425 ( .A1(n10852), .A2(n10851), .B1(n6462), .B2(n10850), .ZN(
        P2_U3435) );
  XNOR2_X1 U11426 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  CLKBUF_X2 U5024 ( .A(n8600), .Z(n8635) );
  CLKBUF_X1 U5030 ( .A(n7292), .Z(n8630) );
  CLKBUF_X2 U5059 ( .A(n5731), .Z(n6815) );
  CLKBUF_X1 U5068 ( .A(n5767), .Z(n8287) );
  CLKBUF_X1 U5295 ( .A(n6272), .Z(n6766) );
  CLKBUF_X2 U5551 ( .A(n7231), .Z(n4948) );
endmodule

