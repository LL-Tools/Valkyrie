

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
         n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
         n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
         n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038,
         n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054,
         n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
         n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
         n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078,
         n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
         n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
         n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16132;

  AOI211_X1 U7301 ( .C1(n15530), .C2(n15230), .A(n15229), .B(n15228), .ZN(
        n15231) );
  INV_X2 U7302 ( .A(n14285), .ZN(n6557) );
  INV_X4 U7303 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U7304 ( .A1(n14967), .A2(n12434), .ZN(n15007) );
  NAND2_X1 U7305 ( .A1(n7886), .A2(n9069), .ZN(n9451) );
  XNOR2_X1 U7306 ( .A(n8249), .B(n8023), .ZN(n12272) );
  INV_X1 U7307 ( .A(n12862), .ZN(n12799) );
  INV_X1 U7308 ( .A(n11934), .ZN(n10584) );
  NAND2_X1 U7310 ( .A1(n16132), .A2(n6656), .ZN(n13121) );
  INV_X2 U7312 ( .A(n12328), .ZN(n12294) );
  BUF_X1 U7313 ( .A(n11126), .Z(n14792) );
  NAND2_X1 U7314 ( .A1(n9131), .A2(n12242), .ZN(n9436) );
  NAND2_X2 U7315 ( .A1(n8437), .A2(n14587), .ZN(n8945) );
  INV_X1 U7316 ( .A(n8436), .ZN(n14587) );
  INV_X1 U7317 ( .A(n12157), .ZN(n11447) );
  NAND2_X2 U7318 ( .A1(n8381), .A2(n8416), .ZN(n11491) );
  AND2_X1 U7319 ( .A1(n15372), .A2(n10259), .ZN(n11031) );
  INV_X1 U7320 ( .A(n8921), .ZN(n6561) );
  INV_X1 U7322 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7627) );
  NOR2_X1 U7323 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n9103) );
  NOR2_X1 U7324 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n9102) );
  NAND2_X1 U7325 ( .A1(n13229), .A2(n13228), .ZN(n13254) );
  CLKBUF_X3 U7326 ( .A(n8776), .Z(n8997) );
  INV_X1 U7327 ( .A(n11860), .ZN(n12534) );
  INV_X1 U7328 ( .A(n10910), .ZN(n14636) );
  OR2_X1 U7330 ( .A1(n11199), .A2(n11198), .ZN(n11449) );
  CLKBUF_X3 U7331 ( .A(n12947), .Z(n7247) );
  AOI21_X1 U7332 ( .B1(n7580), .B2(n6631), .A(n7579), .ZN(n7578) );
  INV_X2 U7333 ( .A(n9855), .ZN(n9961) );
  INV_X1 U7334 ( .A(n9734), .ZN(n6971) );
  XNOR2_X1 U7335 ( .A(n9078), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n9494) );
  XNOR2_X1 U7336 ( .A(n9451), .B(P1_DATAO_REG_20__SCAN_IN), .ZN(n9450) );
  INV_X1 U7337 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n9199) );
  NAND2_X1 U7338 ( .A1(n11920), .A2(n11919), .ZN(n7744) );
  INV_X1 U7339 ( .A(n8945), .ZN(n8756) );
  INV_X1 U7340 ( .A(n10851), .ZN(n11625) );
  INV_X1 U7341 ( .A(n14789), .ZN(n11153) );
  INV_X1 U7342 ( .A(n11451), .ZN(n12413) );
  NAND2_X1 U7343 ( .A1(n15076), .A2(n15059), .ZN(n15054) );
  INV_X1 U7344 ( .A(n14623), .ZN(n15548) );
  XNOR2_X1 U7345 ( .A(n8064), .B(SI_9_), .ZN(n8174) );
  INV_X2 U7346 ( .A(n8050), .ZN(n10052) );
  NAND2_X1 U7347 ( .A1(n6972), .A2(n6971), .ZN(n9739) );
  NOR2_X1 U7348 ( .A1(n13766), .A2(n12664), .ZN(n13844) );
  OR2_X1 U7349 ( .A1(n8380), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n8416) );
  INV_X1 U7350 ( .A(n14962), .ZN(n15230) );
  NAND2_X1 U7351 ( .A1(n14629), .A2(n12521), .ZN(n14704) );
  NAND2_X2 U7352 ( .A1(n15372), .A2(n15374), .ZN(n10700) );
  NAND2_X1 U7353 ( .A1(n15006), .A2(n14966), .ZN(n15249) );
  CLKBUF_X3 U7354 ( .A(n9748), .Z(n13724) );
  NAND2_X1 U7355 ( .A1(n8681), .A2(n8680), .ZN(n13932) );
  INV_X1 U7356 ( .A(n10260), .ZN(n15372) );
  XNOR2_X1 U7357 ( .A(n7348), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8687) );
  BUF_X1 U7358 ( .A(n8687), .Z(n6562) );
  AND2_X1 U7359 ( .A1(n10376), .A2(n11132), .ZN(n12551) );
  AOI21_X2 U7360 ( .B1(n11572), .B2(n11573), .A(n11574), .ZN(n13123) );
  NAND3_X2 U7361 ( .A1(n10705), .A2(n10704), .A3(n8020), .ZN(n14789) );
  AOI21_X2 U7362 ( .B1(n12416), .B2(n12888), .A(n6668), .ZN(n15194) );
  NAND2_X2 U7363 ( .A1(n12178), .A2(n12177), .ZN(n12416) );
  BUF_X4 U7364 ( .A(n12551), .Z(n6553) );
  AND4_X2 U7365 ( .A1(n8083), .A2(n8082), .A3(n8080), .A4(n8081), .ZN(n7277)
         );
  NAND2_X2 U7366 ( .A1(n11642), .A2(n11641), .ZN(n11920) );
  INV_X2 U7367 ( .A(n7528), .ZN(n8779) );
  OAI21_X2 U7368 ( .B1(n9423), .B2(n7883), .A(n6738), .ZN(n9466) );
  NAND2_X2 U7369 ( .A1(n9068), .A2(n9067), .ZN(n9423) );
  OAI222_X1 U7370 ( .A1(n14590), .A2(n12239), .B1(P2_U3088), .B2(n8399), .C1(
        n14594), .C2(n15378), .ZN(P2_U3300) );
  OAI21_X2 U7372 ( .B1(n6936), .B2(n10356), .A(n12688), .ZN(n11175) );
  NAND2_X2 U7373 ( .A1(n10265), .A2(n10264), .ZN(n10356) );
  AND2_X1 U7374 ( .A1(n10672), .A2(n10384), .ZN(n10673) );
  AND3_X2 U7375 ( .A1(n7174), .A2(n8093), .A3(n7774), .ZN(n8393) );
  NAND2_X2 U7376 ( .A1(n13408), .A2(n13407), .ZN(n13410) );
  BUF_X4 U7377 ( .A(n12133), .Z(n6554) );
  INV_X1 U7378 ( .A(n10379), .ZN(n12133) );
  NAND2_X1 U7379 ( .A1(n10463), .A2(n15473), .ZN(n6555) );
  NAND4_X4 U7380 ( .A1(n8451), .A2(n8450), .A3(n8449), .A4(n8448), .ZN(n8788)
         );
  OAI222_X1 U7381 ( .A1(n14594), .A2(n15373), .B1(P2_U3088), .B2(n8395), .C1(
        n12595), .C2(n14590), .ZN(P2_U3297) );
  NAND2_X2 U7383 ( .A1(n8775), .A2(n8774), .ZN(n8921) );
  NAND2_X2 U7384 ( .A1(n8398), .A2(n8399), .ZN(n8111) );
  OR2_X2 U7385 ( .A1(n9654), .A2(n9652), .ZN(n7441) );
  BUF_X4 U7386 ( .A(n10587), .Z(n12947) );
  NAND2_X2 U7387 ( .A1(n9483), .A2(n9077), .ZN(n9078) );
  NAND2_X2 U7388 ( .A1(n14580), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8392) );
  XNOR2_X1 U7389 ( .A(n12053), .B(n7247), .ZN(n11746) );
  XNOR2_X2 U7390 ( .A(n13035), .B(n13036), .ZN(n13037) );
  NAND2_X1 U7391 ( .A1(n10011), .A2(n10010), .ZN(n10022) );
  NOR2_X1 U7392 ( .A1(n14973), .A2(n14972), .ZN(n14971) );
  NAND2_X1 U7393 ( .A1(n9695), .A2(n9694), .ZN(n12996) );
  AOI21_X1 U7394 ( .B1(n12654), .B2(n6585), .A(n6692), .ZN(n7364) );
  NAND2_X1 U7395 ( .A1(n7686), .A2(n7689), .ZN(n7685) );
  AND2_X1 U7396 ( .A1(n13287), .A2(n6613), .ZN(n7686) );
  OAI21_X1 U7397 ( .B1(n13441), .B2(n7925), .A(n9664), .ZN(n7924) );
  NAND2_X1 U7398 ( .A1(n9459), .A2(n9458), .ZN(n13434) );
  AOI21_X1 U7399 ( .B1(n13165), .B2(n13163), .A(n13164), .ZN(n13182) );
  NAND2_X1 U7400 ( .A1(n11004), .A2(n11003), .ZN(n11271) );
  NAND2_X1 U7401 ( .A1(n7286), .A2(n7130), .ZN(n11434) );
  NAND2_X1 U7402 ( .A1(n8237), .A2(n8236), .ZN(n14469) );
  INV_X2 U7403 ( .A(n10587), .ZN(n12995) );
  INV_X1 U7404 ( .A(n12708), .ZN(n11186) );
  XNOR2_X1 U7405 ( .A(n14788), .B(n12699), .ZN(n12872) );
  AND2_X1 U7406 ( .A1(n9610), .A2(n9611), .ZN(n11464) );
  INV_X1 U7407 ( .A(n9824), .ZN(n13703) );
  INV_X1 U7408 ( .A(n12552), .ZN(n10699) );
  INV_X1 U7409 ( .A(n12552), .ZN(n12463) );
  INV_X4 U7410 ( .A(n10379), .ZN(n12552) );
  INV_X4 U7411 ( .A(n6553), .ZN(n14638) );
  INV_X1 U7412 ( .A(n14338), .ZN(n10010) );
  NAND4_X1 U7413 ( .A1(n8464), .A2(n8463), .A3(n8462), .A4(n8461), .ZN(n13955)
         );
  INV_X4 U7414 ( .A(n9436), .ZN(n9554) );
  AND2_X1 U7415 ( .A1(n8687), .A2(n11283), .ZN(n10009) );
  NAND2_X1 U7416 ( .A1(n8388), .A2(n7347), .ZN(n11283) );
  XNOR2_X1 U7418 ( .A(n6897), .B(n9130), .ZN(n12242) );
  INV_X2 U7419 ( .A(n8050), .ZN(n8097) );
  NAND3_X1 U7420 ( .A1(n6971), .A2(n9738), .A3(n9737), .ZN(n9815) );
  INV_X2 U7421 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9811) );
  OR2_X1 U7422 ( .A1(n14413), .A2(n12591), .ZN(n7101) );
  NAND2_X1 U7423 ( .A1(n7142), .A2(n12579), .ZN(n14648) );
  NAND2_X1 U7424 ( .A1(n14956), .A2(n14955), .ZN(n14954) );
  OAI21_X1 U7425 ( .B1(n9524), .B2(n7913), .A(n7911), .ZN(n9871) );
  NOR2_X1 U7426 ( .A1(n7398), .A2(n7720), .ZN(n9720) );
  NOR2_X1 U7427 ( .A1(n13351), .A2(n13355), .ZN(n13350) );
  AND2_X1 U7428 ( .A1(n13334), .A2(n13333), .ZN(n7253) );
  NAND2_X1 U7429 ( .A1(n7364), .A2(n7363), .ZN(n13767) );
  NAND2_X1 U7430 ( .A1(n13002), .A2(n13352), .ZN(n9694) );
  NAND2_X1 U7431 ( .A1(n7549), .A2(n7551), .ZN(n14127) );
  NAND2_X1 U7432 ( .A1(n12944), .A2(n13047), .ZN(n13005) );
  AOI21_X1 U7433 ( .B1(n8917), .B2(n7843), .A(n7840), .ZN(n8926) );
  NAND2_X1 U7434 ( .A1(n9541), .A2(n9540), .ZN(n13002) );
  NAND2_X1 U7435 ( .A1(n9528), .A2(n9527), .ZN(n13566) );
  NAND2_X1 U7436 ( .A1(n6974), .A2(n13332), .ZN(n7254) );
  NAND2_X1 U7437 ( .A1(n7962), .A2(n7959), .ZN(n15068) );
  AND2_X1 U7438 ( .A1(n7921), .A2(n6949), .ZN(n6950) );
  INV_X1 U7439 ( .A(n7010), .ZN(n12984) );
  OAI21_X1 U7440 ( .B1(n9526), .B2(n6610), .A(n9084), .ZN(n9539) );
  NAND2_X1 U7441 ( .A1(n15108), .A2(n15109), .ZN(n15107) );
  NAND2_X1 U7442 ( .A1(n9673), .A2(n9672), .ZN(n13390) );
  AOI21_X1 U7443 ( .B1(n7238), .B2(n7236), .A(n7806), .ZN(n7235) );
  INV_X1 U7444 ( .A(n7924), .ZN(n7923) );
  CLKBUF_X1 U7445 ( .A(n13020), .Z(n6774) );
  AOI21_X1 U7446 ( .B1(n13020), .B2(n6570), .A(n7011), .ZN(n7010) );
  NAND2_X1 U7447 ( .A1(n12929), .A2(n12928), .ZN(n13020) );
  NOR2_X1 U7448 ( .A1(n14999), .A2(n7239), .ZN(n7238) );
  NAND2_X1 U7449 ( .A1(n7920), .A2(n7918), .ZN(n13470) );
  NAND2_X1 U7450 ( .A1(n14156), .A2(n6659), .ZN(n8729) );
  NAND2_X1 U7451 ( .A1(n7887), .A2(n7125), .ZN(n7124) );
  NAND2_X1 U7452 ( .A1(n9496), .A2(n9495), .ZN(n13396) );
  AOI21_X1 U7453 ( .B1(n13194), .B2(n7671), .A(n13204), .ZN(n13220) );
  INV_X1 U7454 ( .A(n14111), .ZN(n13797) );
  AOI21_X1 U7455 ( .B1(n15029), .B2(n7815), .A(n6672), .ZN(n7814) );
  AND2_X1 U7456 ( .A1(n8353), .A2(n8352), .ZN(n14111) );
  OR2_X1 U7457 ( .A1(n9078), .A2(n11790), .ZN(n9079) );
  AOI21_X1 U7458 ( .B1(n7928), .B2(n7931), .A(n13499), .ZN(n7927) );
  AOI21_X1 U7459 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n13183), .A(n13182), .ZN(
        n13185) );
  OAI21_X1 U7460 ( .B1(n14333), .B2(n8711), .A(n8713), .ZN(n14315) );
  NOR2_X1 U7461 ( .A1(n12631), .A2(n7387), .ZN(n7386) );
  NAND2_X1 U7462 ( .A1(n6769), .A2(n6768), .ZN(n8840) );
  NAND2_X1 U7463 ( .A1(n7663), .A2(n7665), .ZN(n13170) );
  NAND2_X1 U7464 ( .A1(n8310), .A2(n8309), .ZN(n14182) );
  OR2_X1 U7465 ( .A1(n9450), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9453) );
  NAND2_X1 U7466 ( .A1(n13255), .A2(n7560), .ZN(n13259) );
  INV_X1 U7467 ( .A(n14537), .ZN(n14167) );
  OR2_X1 U7468 ( .A1(n13597), .A2(n13490), .ZN(n13454) );
  XNOR2_X1 U7469 ( .A(n8308), .B(n8307), .ZN(n12340) );
  NOR2_X1 U7470 ( .A1(n13530), .A2(n7739), .ZN(n7738) );
  OR2_X1 U7471 ( .A1(n15175), .A2(n15314), .ZN(n15176) );
  NAND2_X1 U7472 ( .A1(n9416), .A2(n9415), .ZN(n13597) );
  NOR2_X1 U7473 ( .A1(n12886), .A2(n7221), .ZN(n7223) );
  NAND2_X1 U7474 ( .A1(n8217), .A2(n8216), .ZN(n14306) );
  NAND2_X1 U7475 ( .A1(n12252), .A2(n12251), .ZN(n15308) );
  NAND2_X1 U7476 ( .A1(n12284), .A2(n12283), .ZN(n15294) );
  NOR2_X1 U7477 ( .A1(n12365), .A2(n12353), .ZN(n7283) );
  OR2_X1 U7478 ( .A1(n14325), .A2(n13944), .ZN(n7786) );
  AND2_X1 U7479 ( .A1(n11549), .A2(n11548), .ZN(n7963) );
  NOR2_X1 U7480 ( .A1(n11571), .A2(n6775), .ZN(n11806) );
  OR2_X1 U7481 ( .A1(n8815), .A2(n8814), .ZN(n8820) );
  NAND2_X1 U7482 ( .A1(n12263), .A2(n12262), .ZN(n15302) );
  NAND2_X1 U7483 ( .A1(n7464), .A2(n7462), .ZN(n8326) );
  AND2_X1 U7484 ( .A1(n11570), .A2(n11807), .ZN(n6775) );
  NAND2_X1 U7485 ( .A1(n12329), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n12343) );
  NAND2_X1 U7486 ( .A1(n9342), .A2(n9341), .ZN(n13555) );
  NAND2_X1 U7487 ( .A1(n8201), .A2(n8200), .ZN(n14357) );
  NAND2_X1 U7488 ( .A1(n8105), .A2(n8104), .ZN(n14481) );
  NAND2_X1 U7489 ( .A1(n9371), .A2(n9370), .ZN(n13685) );
  AOI21_X1 U7490 ( .B1(n8238), .B2(n8024), .A(n7451), .ZN(n7448) );
  NAND2_X1 U7491 ( .A1(n11496), .A2(n11495), .ZN(n15336) );
  NAND2_X1 U7492 ( .A1(n8183), .A2(n8182), .ZN(n14575) );
  NAND2_X1 U7493 ( .A1(n11517), .A2(n11516), .ZN(n15499) );
  XNOR2_X1 U7494 ( .A(n9350), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9349) );
  XNOR2_X1 U7495 ( .A(n10608), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n15385) );
  NAND2_X1 U7496 ( .A1(n7097), .A2(n8486), .ZN(n11651) );
  NAND2_X1 U7497 ( .A1(n7457), .A2(n7456), .ZN(n8225) );
  OR2_X1 U7498 ( .A1(n11080), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n6994) );
  NAND2_X1 U7499 ( .A1(n6783), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n12304) );
  NAND2_X1 U7500 ( .A1(n8173), .A2(n8172), .ZN(n14519) );
  NAND2_X1 U7501 ( .A1(n7873), .A2(n9053), .ZN(n9350) );
  OR2_X1 U7502 ( .A1(n8190), .A2(n8189), .ZN(n7802) );
  NAND2_X1 U7503 ( .A1(n11513), .A2(n11512), .ZN(n12724) );
  OAI21_X1 U7504 ( .B1(n8190), .B2(n7461), .A(n7458), .ZN(n8219) );
  NAND2_X1 U7505 ( .A1(n10409), .A2(n10410), .ZN(n10408) );
  NAND2_X1 U7506 ( .A1(n10400), .A2(n10017), .ZN(n10409) );
  NAND2_X1 U7507 ( .A1(n8165), .A2(n8164), .ZN(n11683) );
  AOI21_X1 U7508 ( .B1(n10674), .B2(n11860), .A(n10673), .ZN(n10688) );
  NAND2_X1 U7509 ( .A1(n10773), .A2(n10774), .ZN(n10772) );
  NAND2_X1 U7510 ( .A1(n10401), .A2(n10402), .ZN(n10400) );
  AND2_X1 U7511 ( .A1(n10378), .A2(n10377), .ZN(n10384) );
  AND2_X1 U7512 ( .A1(n10013), .A2(n10012), .ZN(n10402) );
  AND2_X1 U7513 ( .A1(n9262), .A2(n9261), .ZN(n11720) );
  NAND4_X1 U7514 ( .A1(n11036), .A2(n11035), .A3(n11034), .A4(n11033), .ZN(
        n14786) );
  NAND2_X1 U7515 ( .A1(n9173), .A2(n7429), .ZN(n7706) );
  AND2_X1 U7516 ( .A1(n6696), .A2(n6927), .ZN(n6564) );
  OR2_X1 U7517 ( .A1(n13116), .A2(n11427), .ZN(n9610) );
  NAND2_X1 U7518 ( .A1(n8056), .A2(n8055), .ZN(n8161) );
  NAND2_X1 U7519 ( .A1(n10516), .A2(n9766), .ZN(n11055) );
  AND2_X2 U7520 ( .A1(n10667), .A2(n7601), .ZN(n11133) );
  INV_X2 U7521 ( .A(n8776), .ZN(n8960) );
  OAI211_X1 U7522 ( .C1(n10897), .C2(n10890), .A(n10889), .B(n10888), .ZN(
        n14623) );
  INV_X1 U7523 ( .A(n11269), .ZN(n15769) );
  NAND4_X1 U7524 ( .A1(n10363), .A2(n10362), .A3(n10361), .A4(n10360), .ZN(
        n11126) );
  AND3_X1 U7525 ( .A1(n9167), .A2(n9166), .A3(n9165), .ZN(n11046) );
  INV_X2 U7526 ( .A(n8921), .ZN(n8776) );
  AND3_X1 U7527 ( .A1(n9225), .A2(n9224), .A3(n9223), .ZN(n11269) );
  NAND2_X1 U7528 ( .A1(n8688), .A2(n10011), .ZN(n15715) );
  INV_X2 U7529 ( .A(n9256), .ZN(n9550) );
  INV_X1 U7530 ( .A(n9202), .ZN(n9429) );
  NAND2_X1 U7531 ( .A1(n9150), .A2(n6647), .ZN(n13120) );
  BUF_X2 U7532 ( .A(n11031), .Z(n11451) );
  CLKBUF_X1 U7533 ( .A(n12157), .Z(n12158) );
  CLKBUF_X1 U7534 ( .A(n10185), .Z(n12588) );
  NAND4_X2 U7535 ( .A1(n8459), .A2(n8458), .A3(n8457), .A4(n8456), .ZN(n13956)
         );
  AOI21_X1 U7536 ( .B1(n7803), .B2(n7800), .A(n7799), .ZN(n7798) );
  NAND2_X1 U7537 ( .A1(n9260), .A2(n9276), .ZN(n11568) );
  NAND2_X1 U7538 ( .A1(n6560), .A2(n10052), .ZN(n9256) );
  OR2_X1 U7539 ( .A1(n8550), .A2(n8549), .ZN(n8558) );
  NAND2_X1 U7540 ( .A1(n9741), .A2(n9739), .ZN(n12057) );
  NAND2_X1 U7541 ( .A1(n9747), .A2(n9748), .ZN(n8022) );
  NAND2_X2 U7542 ( .A1(n10463), .A2(n15473), .ZN(n12328) );
  AND2_X1 U7543 ( .A1(n10260), .A2(n10259), .ZN(n12157) );
  INV_X1 U7544 ( .A(n10011), .ZN(n8775) );
  NAND2_X1 U7545 ( .A1(n6779), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n11521) );
  XNOR2_X1 U7546 ( .A(n8108), .B(n8107), .ZN(n10663) );
  INV_X2 U7547 ( .A(n8468), .ZN(n8757) );
  OAI21_X1 U7548 ( .B1(n9951), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9946) );
  NAND2_X1 U7549 ( .A1(n10225), .A2(n10226), .ZN(n15473) );
  NAND2_X1 U7550 ( .A1(n7218), .A2(n6934), .ZN(n10260) );
  NAND2_X1 U7551 ( .A1(n8272), .A2(n8384), .ZN(n10011) );
  INV_X1 U7552 ( .A(n11519), .ZN(n6779) );
  NAND2_X1 U7553 ( .A1(n9184), .A2(n9183), .ZN(n9186) );
  NAND2_X1 U7554 ( .A1(n9945), .A2(n9944), .ZN(n9951) );
  MUX2_X1 U7555 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10224), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n10225) );
  NAND2_X1 U7556 ( .A1(n9744), .A2(n9743), .ZN(n11892) );
  NAND2_X1 U7557 ( .A1(n6780), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11519) );
  AOI21_X1 U7558 ( .B1(n8271), .B2(n8270), .A(n8269), .ZN(n8272) );
  AOI21_X1 U7559 ( .B1(n10257), .B2(n6591), .A(n6935), .ZN(n6934) );
  INV_X1 U7560 ( .A(n11449), .ZN(n6780) );
  NAND2_X1 U7561 ( .A1(n8233), .A2(n8232), .ZN(n8271) );
  NAND2_X1 U7562 ( .A1(n7964), .A2(n7965), .ZN(n10257) );
  NAND2_X1 U7563 ( .A1(n8387), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7348) );
  NAND2_X1 U7564 ( .A1(n9201), .A2(n9232), .ZN(n10991) );
  AND2_X1 U7565 ( .A1(n8198), .A2(n7747), .ZN(n8233) );
  INV_X1 U7566 ( .A(n10642), .ZN(n7964) );
  INV_X1 U7567 ( .A(n9815), .ZN(n6558) );
  NAND2_X1 U7568 ( .A1(n8390), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8096) );
  AOI21_X1 U7569 ( .B1(n7105), .B2(n7108), .A(n6679), .ZN(n7104) );
  AND2_X1 U7570 ( .A1(n8195), .A2(n8101), .ZN(n8198) );
  NOR2_X1 U7571 ( .A1(n8098), .A2(n8100), .ZN(n8195) );
  NAND3_X2 U7572 ( .A1(n9196), .A2(n7661), .A3(n6621), .ZN(n10106) );
  NOR2_X1 U7573 ( .A1(n8092), .A2(n8091), .ZN(n8093) );
  AND2_X1 U7574 ( .A1(n9037), .A2(n9036), .ZN(n9203) );
  AND2_X1 U7575 ( .A1(n9039), .A2(n9038), .ZN(n9218) );
  AND2_X1 U7576 ( .A1(n9568), .A2(n9100), .ZN(n7260) );
  AND3_X1 U7577 ( .A1(n7092), .A2(n7091), .A3(n7090), .ZN(n8099) );
  CLKBUF_X1 U7578 ( .A(n9729), .Z(n16100) );
  AND3_X1 U7579 ( .A1(n9102), .A2(n9103), .A3(n9101), .ZN(n9325) );
  AND2_X1 U7580 ( .A1(n8084), .A2(n8085), .ZN(n7521) );
  AND3_X1 U7581 ( .A1(n9097), .A2(n9096), .A3(n9384), .ZN(n9569) );
  AND2_X1 U7582 ( .A1(n7089), .A2(n7088), .ZN(n7522) );
  NAND2_X1 U7583 ( .A1(n9028), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9161) );
  AND3_X1 U7584 ( .A1(n9099), .A2(n7630), .A3(n9098), .ZN(n9568) );
  NOR2_X1 U7585 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n9942) );
  INV_X1 U7586 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n10205) );
  INV_X1 U7587 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8383) );
  NOR2_X1 U7588 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n7089) );
  NOR2_X1 U7589 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7088) );
  NOR2_X1 U7590 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n10217) );
  INV_X1 U7591 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n15963) );
  NOR2_X1 U7592 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n8081) );
  INV_X1 U7593 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8401) );
  INV_X1 U7594 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n10096) );
  NOR2_X2 U7595 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n9101) );
  INV_X4 U7596 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7597 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8417) );
  INV_X1 U7598 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7662) );
  INV_X1 U7599 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n15826) );
  INV_X1 U7600 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8084) );
  NOR2_X1 U7601 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n8082) );
  NOR2_X1 U7602 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n8080) );
  INV_X4 U7603 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7604 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n9934) );
  NOR2_X1 U7605 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n9935) );
  NOR2_X1 U7606 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7090) );
  INV_X1 U7607 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9729) );
  NOR2_X1 U7608 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7092) );
  NOR2_X1 U7609 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7091) );
  INV_X1 U7610 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7792) );
  INV_X1 U7611 ( .A(n13122), .ZN(n10516) );
  INV_X2 U7612 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6932) );
  OAI21_X2 U7613 ( .B1(n7333), .B2(n6940), .A(n6938), .ZN(n15127) );
  INV_X1 U7614 ( .A(n12872), .ZN(n11344) );
  NAND2_X1 U7615 ( .A1(n11133), .A2(n11126), .ZN(n12687) );
  AND2_X2 U7617 ( .A1(n12696), .A2(n12697), .ZN(n12874) );
  NAND2_X1 U7618 ( .A1(n11153), .A2(n14623), .ZN(n12696) );
  AOI21_X2 U7619 ( .B1(n13744), .B2(n13743), .A(n13742), .ZN(n13902) );
  OAI21_X2 U7620 ( .B1(n9245), .B2(n9244), .A(n9042), .ZN(n9253) );
  NAND2_X2 U7621 ( .A1(n15491), .A2(n15494), .ZN(n12092) );
  NAND2_X2 U7622 ( .A1(n7211), .A2(n11514), .ZN(n15491) );
  NOR2_X1 U7623 ( .A1(n10642), .A2(n7329), .ZN(n10223) );
  NAND2_X1 U7624 ( .A1(n9747), .A2(n9748), .ZN(n6559) );
  NAND2_X1 U7625 ( .A1(n9747), .A2(n9748), .ZN(n6560) );
  INV_X2 U7626 ( .A(n13445), .ZN(n13441) );
  XNOR2_X2 U7627 ( .A(n10222), .B(n10253), .ZN(n10463) );
  NOR2_X2 U7628 ( .A1(n15243), .A2(n12435), .ZN(n14973) );
  NOR2_X2 U7629 ( .A1(n14974), .A2(n15230), .ZN(n14957) );
  OAI21_X2 U7630 ( .B1(n9186), .B2(n7880), .A(n7877), .ZN(n9219) );
  NAND2_X4 U7631 ( .A1(n13714), .A2(n12242), .ZN(n9211) );
  NAND2_X1 U7632 ( .A1(n15068), .A2(n12311), .ZN(n15049) );
  NOR2_X1 U7633 ( .A1(n9636), .A2(n9635), .ZN(n9640) );
  AOI21_X1 U7634 ( .B1(n7445), .B2(n7444), .A(n7442), .ZN(n9636) );
  AOI21_X1 U7635 ( .B1(n6563), .B2(n15105), .A(n12790), .ZN(n7594) );
  AND3_X1 U7636 ( .A1(n9682), .A2(n9704), .A3(n9681), .ZN(n9693) );
  INV_X1 U7637 ( .A(n9659), .ZN(n7925) );
  INV_X1 U7638 ( .A(n12242), .ZN(n9132) );
  NAND2_X1 U7639 ( .A1(n7265), .A2(n7264), .ZN(n7270) );
  NOR2_X1 U7640 ( .A1(n13220), .A2(n13219), .ZN(n13221) );
  OR2_X1 U7641 ( .A1(n13580), .A2(n13069), .ZN(n9674) );
  AND2_X1 U7642 ( .A1(n6729), .A2(n8720), .ZN(n7021) );
  INV_X1 U7643 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U7644 ( .A1(n6624), .A2(n7807), .ZN(n7806) );
  INV_X1 U7645 ( .A(n7815), .ZN(n7236) );
  INV_X1 U7646 ( .A(n12435), .ZN(n7807) );
  OAI21_X1 U7647 ( .B1(n8341), .B2(n12055), .A(n8340), .ZN(n8343) );
  OAI21_X1 U7648 ( .B1(n8335), .B2(n8334), .A(n8336), .ZN(n8341) );
  XNOR2_X1 U7649 ( .A(n8219), .B(SI_14_), .ZN(n8208) );
  INV_X1 U7650 ( .A(n9177), .ZN(n9547) );
  NAND2_X1 U7651 ( .A1(n9970), .A2(n10739), .ZN(n7581) );
  NOR2_X1 U7652 ( .A1(n13352), .A2(n13533), .ZN(n9865) );
  NAND2_X1 U7653 ( .A1(n13416), .A2(n9667), .ZN(n9479) );
  NAND2_X1 U7654 ( .A1(n9848), .A2(n9884), .ZN(n10534) );
  AND2_X1 U7655 ( .A1(n10501), .A2(n10081), .ZN(n10535) );
  AND2_X1 U7656 ( .A1(n10500), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10081) );
  NAND2_X1 U7657 ( .A1(n11491), .A2(n10009), .ZN(n8773) );
  NAND2_X1 U7658 ( .A1(n8395), .A2(n8436), .ZN(n8455) );
  AOI21_X1 U7659 ( .B1(n7554), .B2(n7552), .A(n6669), .ZN(n7551) );
  INV_X1 U7660 ( .A(n15662), .ZN(n14375) );
  NAND2_X1 U7661 ( .A1(n12328), .A2(n10885), .ZN(n10897) );
  INV_X1 U7662 ( .A(n15482), .ZN(n6869) );
  NOR2_X1 U7663 ( .A1(n12438), .A2(n12440), .ZN(n14933) );
  NOR2_X1 U7664 ( .A1(n12781), .A2(n12300), .ZN(n7959) );
  OR2_X1 U7665 ( .A1(n15294), .A2(n15131), .ZN(n12779) );
  INV_X1 U7666 ( .A(n14933), .ZN(n14935) );
  NAND2_X1 U7667 ( .A1(n6944), .A2(n6945), .ZN(n14930) );
  INV_X1 U7668 ( .A(n6946), .ZN(n6944) );
  NAND3_X1 U7669 ( .A1(n6948), .A2(n12385), .A3(n6943), .ZN(n6945) );
  OAI211_X1 U7670 ( .C1(n7706), .C2(n9855), .A(n9585), .B(n7427), .ZN(n9592)
         );
  NAND2_X1 U7671 ( .A1(n7428), .A2(n9855), .ZN(n7427) );
  INV_X1 U7672 ( .A(n9708), .ZN(n7428) );
  NAND2_X1 U7673 ( .A1(n7405), .A2(n9855), .ZN(n7404) );
  OAI21_X1 U7674 ( .B1(n7437), .B2(n7441), .A(n7440), .ZN(n7436) );
  NAND2_X1 U7675 ( .A1(n9657), .A2(n9656), .ZN(n7440) );
  NOR2_X1 U7676 ( .A1(n6667), .A2(n7598), .ZN(n7597) );
  NAND2_X1 U7677 ( .A1(n8910), .A2(n7865), .ZN(n7864) );
  AND2_X1 U7678 ( .A1(n8918), .A2(n7854), .ZN(n7853) );
  INV_X1 U7679 ( .A(n8920), .ZN(n7854) );
  INV_X1 U7680 ( .A(n12791), .ZN(n7591) );
  AOI21_X1 U7681 ( .B1(n7594), .B2(n7595), .A(n12792), .ZN(n7593) );
  NAND2_X1 U7682 ( .A1(n7592), .A2(n7595), .ZN(n7323) );
  INV_X1 U7683 ( .A(n13363), .ZN(n9704) );
  MUX2_X1 U7684 ( .A(n9686), .B(n9685), .S(n9961), .Z(n9687) );
  NAND2_X1 U7685 ( .A1(n7455), .A2(n7454), .ZN(n12838) );
  NAND2_X1 U7686 ( .A1(n12814), .A2(n12799), .ZN(n7454) );
  NAND2_X1 U7687 ( .A1(n14923), .A2(n12862), .ZN(n7455) );
  INV_X1 U7688 ( .A(n8300), .ZN(n7468) );
  NAND2_X1 U7689 ( .A1(n8211), .A2(SI_15_), .ZN(n8222) );
  NAND2_X1 U7690 ( .A1(n9697), .A2(n9855), .ZN(n7266) );
  INV_X1 U7691 ( .A(n9696), .ZN(n7268) );
  AOI21_X1 U7692 ( .B1(n7738), .B2(n7736), .A(n7735), .ZN(n7734) );
  INV_X1 U7693 ( .A(n7741), .ZN(n7736) );
  INV_X1 U7694 ( .A(n13516), .ZN(n7735) );
  AND2_X1 U7695 ( .A1(n6566), .A2(n6858), .ZN(n6856) );
  AND2_X1 U7696 ( .A1(n7057), .A2(n8707), .ZN(n7769) );
  NOR2_X1 U7697 ( .A1(n7770), .A2(n7058), .ZN(n7057) );
  INV_X1 U7698 ( .A(n8705), .ZN(n7058) );
  INV_X1 U7699 ( .A(n8703), .ZN(n7770) );
  NOR2_X1 U7700 ( .A1(n14306), .A2(n14481), .ZN(n7514) );
  AND2_X1 U7701 ( .A1(n7949), .A2(n6709), .ZN(n7947) );
  NAND2_X1 U7702 ( .A1(n12248), .A2(n7950), .ZN(n7949) );
  NAND2_X1 U7703 ( .A1(n15314), .A2(n14758), .ZN(n12757) );
  OAI21_X1 U7704 ( .B1(n8024), .B2(n7451), .A(n8023), .ZN(n7450) );
  AND2_X1 U7705 ( .A1(n7804), .A2(n8029), .ZN(n7803) );
  NAND2_X1 U7706 ( .A1(n8072), .A2(n10183), .ZN(n8074) );
  INV_X1 U7707 ( .A(n8062), .ZN(n7319) );
  INV_X1 U7708 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10126) );
  NAND2_X1 U7709 ( .A1(n7192), .A2(n7189), .ZN(n10133) );
  AND2_X1 U7710 ( .A1(n7190), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n7189) );
  NOR2_X1 U7711 ( .A1(n13029), .A2(n7633), .ZN(n7632) );
  INV_X1 U7712 ( .A(n12932), .ZN(n7633) );
  AND2_X1 U7713 ( .A1(n10984), .A2(n9957), .ZN(n10733) );
  NAND2_X1 U7714 ( .A1(n13183), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7668) );
  INV_X1 U7715 ( .A(n9804), .ZN(n7724) );
  NAND2_X1 U7716 ( .A1(n9127), .A2(n9126), .ZN(n9893) );
  NAND3_X1 U7717 ( .A1(n6893), .A2(n6891), .A3(n6649), .ZN(n13351) );
  NAND2_X1 U7718 ( .A1(n6892), .A2(n6634), .ZN(n6891) );
  OR2_X1 U7719 ( .A1(n13434), .A2(n13446), .ZN(n9663) );
  OR2_X1 U7720 ( .A1(n13118), .A2(n15769), .ZN(n9603) );
  NAND2_X1 U7721 ( .A1(n9796), .A2(n6650), .ZN(n7752) );
  NAND2_X1 U7722 ( .A1(n7869), .A2(n7867), .ZN(n9684) );
  NOR2_X1 U7723 ( .A1(n13353), .A2(n7868), .ZN(n7867) );
  INV_X1 U7724 ( .A(n9518), .ZN(n7868) );
  NOR2_X1 U7725 ( .A1(n13431), .A2(n7754), .ZN(n7753) );
  INV_X1 U7726 ( .A(n9795), .ZN(n7754) );
  NAND2_X1 U7727 ( .A1(n7930), .A2(n9379), .ZN(n7929) );
  OAI22_X1 U7728 ( .A1(n7734), .A2(n6888), .B1(n7737), .B2(n6882), .ZN(n6887)
         );
  NAND2_X1 U7729 ( .A1(n13515), .A2(n12103), .ZN(n6882) );
  INV_X1 U7730 ( .A(n7738), .ZN(n7737) );
  OR2_X1 U7731 ( .A1(n13689), .A2(n13548), .ZN(n9632) );
  INV_X1 U7732 ( .A(n11110), .ZN(n9764) );
  AND2_X1 U7733 ( .A1(n11892), .A2(n9817), .ZN(n9818) );
  INV_X1 U7734 ( .A(n7120), .ZN(n7119) );
  OAI21_X1 U7735 ( .B1(n7122), .B2(n7121), .A(n7894), .ZN(n7120) );
  INV_X1 U7736 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9128) );
  INV_X1 U7737 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n9106) );
  AND2_X1 U7738 ( .A1(n9727), .A2(n9726), .ZN(n9732) );
  INV_X1 U7739 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n9726) );
  AND2_X2 U7740 ( .A1(n9980), .A2(n7662), .ZN(n9326) );
  NAND2_X1 U7741 ( .A1(n6678), .A2(n6594), .ZN(n7370) );
  NAND2_X1 U7742 ( .A1(n14111), .A2(n7520), .ZN(n7519) );
  OR2_X1 U7743 ( .A1(n13797), .A2(n9917), .ZN(n9907) );
  OR2_X1 U7744 ( .A1(n14194), .A2(n13801), .ZN(n14157) );
  NAND2_X1 U7745 ( .A1(n8724), .A2(n7758), .ZN(n7757) );
  INV_X1 U7746 ( .A(n8723), .ZN(n7758) );
  AND2_X1 U7747 ( .A1(n8717), .A2(n6701), .ZN(n7337) );
  NAND2_X1 U7748 ( .A1(n11729), .A2(n11730), .ZN(n8708) );
  NAND2_X1 U7749 ( .A1(n7977), .A2(n7980), .ZN(n7975) );
  INV_X1 U7750 ( .A(n14696), .ZN(n7980) );
  AOI21_X1 U7751 ( .B1(n14696), .B2(n7979), .A(n7978), .ZN(n7977) );
  AND2_X1 U7752 ( .A1(n12544), .A2(n12543), .ZN(n12546) );
  INV_X1 U7753 ( .A(n7995), .ZN(n7994) );
  OAI21_X1 U7754 ( .B1(n7998), .B2(n7996), .A(n12508), .ZN(n7995) );
  OAI21_X1 U7755 ( .B1(n10656), .B2(n10657), .A(n6748), .ZN(n7081) );
  INV_X1 U7756 ( .A(n7238), .ZN(n7237) );
  INV_X1 U7757 ( .A(n12433), .ZN(n7816) );
  NAND2_X1 U7758 ( .A1(n14619), .A2(n7477), .ZN(n7476) );
  NOR2_X1 U7759 ( .A1(n15253), .A2(n15267), .ZN(n7477) );
  NOR2_X1 U7760 ( .A1(n7482), .A2(n15287), .ZN(n7481) );
  INV_X1 U7761 ( .A(n7483), .ZN(n7482) );
  AOI21_X1 U7762 ( .B1(n6567), .B2(n7809), .A(n6670), .ZN(n7808) );
  INV_X1 U7763 ( .A(n7812), .ZN(n7809) );
  INV_X1 U7764 ( .A(n7231), .ZN(n7230) );
  OAI21_X1 U7765 ( .B1(n7794), .B2(n7232), .A(n15149), .ZN(n7231) );
  NAND2_X1 U7766 ( .A1(n12063), .A2(n11547), .ZN(n6941) );
  NAND2_X1 U7767 ( .A1(n12687), .A2(n6937), .ZN(n6936) );
  INV_X1 U7768 ( .A(n6849), .ZN(n6848) );
  OR2_X1 U7769 ( .A1(n10135), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n10137) );
  OR2_X1 U7770 ( .A1(n12958), .A2(n13375), .ZN(n12959) );
  OR2_X1 U7771 ( .A1(n13084), .A2(n7036), .ZN(n7034) );
  NAND2_X1 U7772 ( .A1(n6570), .A2(n7015), .ZN(n7012) );
  NAND2_X1 U7773 ( .A1(n11586), .A2(n11585), .ZN(n11593) );
  OR2_X1 U7774 ( .A1(n9852), .A2(n9851), .ZN(n10532) );
  NAND2_X1 U7775 ( .A1(n6684), .A2(n9721), .ZN(n6957) );
  AND2_X1 U7776 ( .A1(n9515), .A2(n9514), .ZN(n13085) );
  INV_X1 U7777 ( .A(n9175), .ZN(n9553) );
  OAI21_X1 U7778 ( .B1(n6685), .B2(n6575), .A(n7570), .ZN(n7569) );
  NAND2_X1 U7779 ( .A1(n13134), .A2(n13153), .ZN(n13147) );
  NAND2_X1 U7780 ( .A1(n7667), .A2(n13128), .ZN(n7666) );
  NAND2_X1 U7781 ( .A1(n13221), .A2(n7675), .ZN(n7673) );
  NAND2_X1 U7782 ( .A1(n13256), .A2(n7675), .ZN(n7672) );
  NAND2_X1 U7783 ( .A1(n13271), .A2(n7559), .ZN(n13275) );
  OR2_X1 U7784 ( .A1(n13272), .A2(n13273), .ZN(n7559) );
  NAND2_X1 U7785 ( .A1(n13275), .A2(n13274), .ZN(n13299) );
  XNOR2_X1 U7786 ( .A(n13327), .B(n13302), .ZN(n13304) );
  NAND2_X1 U7787 ( .A1(n13410), .A2(n9674), .ZN(n13385) );
  OR2_X1 U7788 ( .A1(n9417), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9432) );
  INV_X1 U7789 ( .A(n9780), .ZN(n11843) );
  OR2_X1 U7790 ( .A1(n13117), .A2(n11411), .ZN(n9609) );
  INV_X1 U7791 ( .A(n10631), .ZN(n13324) );
  OR2_X1 U7792 ( .A1(n8022), .A2(n11102), .ZN(n9165) );
  NAND2_X1 U7793 ( .A1(n7923), .A2(n9706), .ZN(n6951) );
  AND2_X1 U7794 ( .A1(n6952), .A2(n9706), .ZN(n13442) );
  NAND2_X1 U7795 ( .A1(n13470), .A2(n9649), .ZN(n6952) );
  NAND2_X1 U7796 ( .A1(n9961), .A2(n9749), .ZN(n13533) );
  INV_X1 U7797 ( .A(n13533), .ZN(n13549) );
  AOI21_X1 U7798 ( .B1(n6625), .B2(n7902), .A(n7901), .ZN(n7900) );
  INV_X1 U7799 ( .A(n9288), .ZN(n7902) );
  INV_X1 U7800 ( .A(n9621), .ZN(n7901) );
  XNOR2_X1 U7801 ( .A(n9129), .B(P3_IR_REG_30__SCAN_IN), .ZN(n9131) );
  AOI21_X1 U7802 ( .B1(n9290), .B2(n7107), .A(n7106), .ZN(n7105) );
  INV_X1 U7803 ( .A(n9048), .ZN(n7106) );
  INV_X1 U7804 ( .A(n9046), .ZN(n7107) );
  INV_X1 U7805 ( .A(n9290), .ZN(n7108) );
  NAND2_X1 U7806 ( .A1(n7275), .A2(n9277), .ZN(n9308) );
  NAND2_X1 U7807 ( .A1(n9272), .A2(n9271), .ZN(n9274) );
  INV_X1 U7808 ( .A(n9203), .ZN(n7880) );
  AOI21_X1 U7809 ( .B1(n9203), .B2(n7879), .A(n7878), .ZN(n7877) );
  INV_X1 U7810 ( .A(n9035), .ZN(n7879) );
  NAND2_X1 U7811 ( .A1(n10056), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9035) );
  AND2_X1 U7812 ( .A1(n12638), .A2(n12637), .ZN(n13834) );
  NOR2_X1 U7813 ( .A1(n15697), .A2(n11616), .ZN(n10040) );
  AND4_X1 U7814 ( .A1(n8546), .A2(n8545), .A3(n8544), .A4(n8543), .ZN(n13812)
         );
  OR2_X1 U7815 ( .A1(n8739), .A2(n8438), .ZN(n8441) );
  INV_X1 U7816 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8101) );
  NOR2_X1 U7817 ( .A1(n8765), .A2(n6652), .ZN(n7160) );
  AOI21_X1 U7818 ( .B1(n7555), .B2(n8655), .A(n6676), .ZN(n7554) );
  NAND2_X1 U7819 ( .A1(n14189), .A2(n8646), .ZN(n14174) );
  NAND2_X1 U7820 ( .A1(n14548), .A2(n12655), .ZN(n7535) );
  OAI21_X1 U7821 ( .B1(n14261), .B2(n7112), .A(n7109), .ZN(n7534) );
  INV_X1 U7822 ( .A(n9013), .ZN(n7112) );
  AND2_X1 U7823 ( .A1(n6715), .A2(n7110), .ZN(n7109) );
  AND2_X1 U7824 ( .A1(n8723), .A2(n8722), .ZN(n14222) );
  NAND2_X1 U7825 ( .A1(n7543), .A2(n7547), .ZN(n7540) );
  INV_X1 U7826 ( .A(n10428), .ZN(n8274) );
  INV_X1 U7827 ( .A(n8376), .ZN(n8235) );
  OR2_X1 U7828 ( .A1(n15701), .A2(n10028), .ZN(n11616) );
  NAND2_X1 U7829 ( .A1(n8339), .A2(n8338), .ZN(n14130) );
  BUF_X1 U7830 ( .A(n8111), .Z(n10428) );
  OAI21_X1 U7831 ( .B1(n11491), .B2(n10009), .A(n8773), .ZN(n8688) );
  XOR2_X1 U7832 ( .A(n11788), .B(n15938), .Z(n8413) );
  OR2_X1 U7833 ( .A1(n8393), .A2(n6809), .ZN(n8394) );
  OR2_X1 U7834 ( .A1(n8405), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n8408) );
  NAND2_X1 U7835 ( .A1(n12225), .A2(n12224), .ZN(n12228) );
  INV_X1 U7836 ( .A(n11866), .ZN(n11868) );
  NAND2_X1 U7837 ( .A1(n7285), .A2(n8001), .ZN(n12225) );
  AOI21_X1 U7838 ( .B1(n8003), .B2(n8005), .A(n8002), .ZN(n8001) );
  NAND2_X1 U7839 ( .A1(n11866), .A2(n8003), .ZN(n7285) );
  INV_X1 U7840 ( .A(n12142), .ZN(n8002) );
  INV_X1 U7841 ( .A(n7283), .ZN(n12375) );
  NAND2_X1 U7842 ( .A1(n7283), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n12400) );
  NOR2_X1 U7843 ( .A1(n12853), .A2(n12852), .ZN(n7322) );
  NAND2_X1 U7844 ( .A1(n11031), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10703) );
  INV_X1 U7845 ( .A(n7498), .ZN(n6874) );
  NAND2_X1 U7846 ( .A1(n10898), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7302) );
  INV_X1 U7847 ( .A(n10824), .ZN(n7077) );
  NAND2_X1 U7848 ( .A1(n6878), .A2(n6875), .ZN(n14867) );
  NOR2_X1 U7849 ( .A1(n7504), .A2(n6876), .ZN(n6875) );
  INV_X1 U7850 ( .A(n14855), .ZN(n6876) );
  INV_X1 U7851 ( .A(n6860), .ZN(n6859) );
  NAND2_X1 U7852 ( .A1(n6863), .A2(n6870), .ZN(n6862) );
  OAI21_X1 U7853 ( .B1(n7492), .B2(n6866), .A(n6861), .ZN(n6860) );
  NOR2_X1 U7854 ( .A1(n14954), .A2(n12437), .ZN(n7214) );
  XNOR2_X1 U7855 ( .A(n15236), .B(n14990), .ZN(n14969) );
  NAND2_X1 U7856 ( .A1(n7954), .A2(n6660), .ZN(n7953) );
  OR2_X1 U7857 ( .A1(n15044), .A2(n15051), .ZN(n12339) );
  NOR2_X1 U7858 ( .A1(n15100), .A2(n7961), .ZN(n7960) );
  INV_X1 U7859 ( .A(n12779), .ZN(n7961) );
  NAND2_X1 U7860 ( .A1(n15127), .A2(n12767), .ZN(n15108) );
  NOR2_X1 U7861 ( .A1(n7487), .A2(n15331), .ZN(n7486) );
  AND2_X1 U7862 ( .A1(n12075), .A2(n12011), .ZN(n12885) );
  NAND2_X1 U7863 ( .A1(n12155), .A2(n12154), .ZN(n15319) );
  AND2_X1 U7864 ( .A1(n10220), .A2(n7966), .ZN(n7965) );
  AND2_X1 U7865 ( .A1(n7967), .A2(n10253), .ZN(n7966) );
  XNOR2_X1 U7866 ( .A(n8375), .B(n8374), .ZN(n14579) );
  NAND2_X1 U7867 ( .A1(n8372), .A2(n8371), .ZN(n8375) );
  XNOR2_X1 U7868 ( .A(n8349), .B(n8344), .ZN(n12394) );
  OAI211_X1 U7869 ( .C1(n8208), .C2(n6834), .A(n6831), .B(n6830), .ZN(n12250)
         );
  NAND2_X1 U7870 ( .A1(n8208), .A2(n6837), .ZN(n6830) );
  AOI21_X1 U7871 ( .B1(n15383), .B2(n15384), .A(n10160), .ZN(n10162) );
  AND2_X1 U7872 ( .A1(n10159), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n10160) );
  NAND2_X1 U7873 ( .A1(n12043), .A2(n12042), .ZN(n12196) );
  OR2_X1 U7874 ( .A1(n12041), .A2(n12040), .ZN(n12043) );
  AND2_X1 U7875 ( .A1(n15392), .A2(n15391), .ZN(n15401) );
  AND2_X1 U7876 ( .A1(n7640), .A2(n15451), .ZN(n7202) );
  INV_X1 U7877 ( .A(n13106), .ZN(n13433) );
  INV_X1 U7878 ( .A(n13375), .ZN(n13353) );
  AND2_X1 U7879 ( .A1(n9536), .A2(n9535), .ZN(n13089) );
  NAND2_X1 U7880 ( .A1(n10511), .A2(n13479), .ZN(n13102) );
  INV_X1 U7881 ( .A(n13089), .ZN(n9803) );
  NOR2_X1 U7882 ( .A1(n8012), .A2(n11741), .ZN(n7827) );
  NOR2_X1 U7883 ( .A1(n8389), .A2(n14338), .ZN(n14088) );
  OAI21_X1 U7884 ( .B1(n7343), .B2(n14375), .A(n14137), .ZN(n14415) );
  XNOR2_X1 U7885 ( .A(n14135), .B(n7344), .ZN(n7343) );
  INV_X1 U7886 ( .A(n14136), .ZN(n7344) );
  OAI21_X1 U7887 ( .B1(n14143), .B2(n8730), .A(n6623), .ZN(n14135) );
  OAI21_X1 U7888 ( .B1(n14162), .B2(n14375), .A(n14161), .ZN(n14425) );
  NAND2_X1 U7889 ( .A1(n7500), .A2(n7499), .ZN(n7498) );
  NAND2_X1 U7890 ( .A1(n6568), .A2(n10235), .ZN(n10267) );
  NOR2_X1 U7891 ( .A1(n14905), .A2(n6905), .ZN(n6903) );
  NAND2_X1 U7892 ( .A1(n14930), .A2(n6590), .ZN(n7941) );
  AOI21_X1 U7893 ( .B1(n7942), .B2(n7939), .A(n15213), .ZN(n7334) );
  INV_X1 U7894 ( .A(n12692), .ZN(n7607) );
  INV_X1 U7895 ( .A(n8800), .ZN(n7821) );
  OR2_X1 U7896 ( .A1(n7615), .A2(n12710), .ZN(n7614) );
  INV_X1 U7897 ( .A(n12709), .ZN(n7615) );
  OR2_X1 U7898 ( .A1(n7618), .A2(n12722), .ZN(n7617) );
  INV_X1 U7899 ( .A(n12721), .ZN(n7618) );
  NAND2_X1 U7900 ( .A1(n6773), .A2(n6772), .ZN(n6771) );
  INV_X1 U7901 ( .A(n8818), .ZN(n6772) );
  NAND2_X1 U7902 ( .A1(n7610), .A2(n7609), .ZN(n12740) );
  NAND2_X1 U7903 ( .A1(n12733), .A2(n12735), .ZN(n7609) );
  NAND2_X1 U7904 ( .A1(n7424), .A2(n9596), .ZN(n7421) );
  NAND2_X1 U7905 ( .A1(n9588), .A2(n9855), .ZN(n7425) );
  NOR2_X1 U7906 ( .A1(n11240), .A2(n11361), .ZN(n7418) );
  NAND2_X1 U7907 ( .A1(n8835), .A2(n8834), .ZN(n6768) );
  NOR2_X1 U7908 ( .A1(n8834), .A2(n8835), .ZN(n7839) );
  INV_X1 U7909 ( .A(n8844), .ZN(n7836) );
  INV_X1 U7910 ( .A(n7438), .ZN(n7437) );
  AOI21_X1 U7911 ( .B1(n7314), .B2(n12799), .A(n7313), .ZN(n7312) );
  NAND2_X1 U7912 ( .A1(n12785), .A2(n12780), .ZN(n7314) );
  NOR2_X1 U7913 ( .A1(n12779), .A2(n12799), .ZN(n7313) );
  AOI21_X1 U7914 ( .B1(n7403), .B2(n9645), .A(n9644), .ZN(n9646) );
  OAI21_X1 U7915 ( .B1(n9642), .B2(n13515), .A(n7404), .ZN(n7403) );
  AND2_X1 U7916 ( .A1(n7594), .A2(n12792), .ZN(n7592) );
  NAND2_X1 U7917 ( .A1(n7863), .A2(n8909), .ZN(n7862) );
  NAND2_X1 U7918 ( .A1(n8907), .A2(n7859), .ZN(n7861) );
  AOI21_X1 U7919 ( .B1(n7850), .B2(n7848), .A(n7847), .ZN(n7846) );
  INV_X1 U7920 ( .A(n8924), .ZN(n7847) );
  INV_X1 U7921 ( .A(n7852), .ZN(n7848) );
  AND2_X1 U7922 ( .A1(n7852), .A2(n8923), .ZN(n7851) );
  NOR2_X1 U7923 ( .A1(n11731), .A2(n7153), .ZN(n7152) );
  NAND2_X1 U7924 ( .A1(n14391), .A2(n14363), .ZN(n7153) );
  NOR2_X1 U7925 ( .A1(n11955), .A2(n7171), .ZN(n9012) );
  NOR2_X1 U7926 ( .A1(n9011), .A2(n7173), .ZN(n7172) );
  NAND2_X1 U7927 ( .A1(n8691), .A2(n9010), .ZN(n7173) );
  NAND2_X1 U7928 ( .A1(n7846), .A2(n7849), .ZN(n7842) );
  INV_X1 U7929 ( .A(n7850), .ZN(n7849) );
  NAND2_X1 U7930 ( .A1(n7851), .A2(n7853), .ZN(n7841) );
  INV_X1 U7931 ( .A(n7846), .ZN(n7845) );
  INV_X1 U7932 ( .A(n7851), .ZN(n7844) );
  NAND2_X1 U7933 ( .A1(n15037), .A2(n15075), .ZN(n7282) );
  NAND2_X1 U7934 ( .A1(n12840), .A2(n12838), .ZN(n7453) );
  INV_X1 U7935 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9932) );
  NOR2_X1 U7936 ( .A1(n9716), .A2(n13390), .ZN(n7401) );
  INV_X1 U7937 ( .A(n7909), .ZN(n7908) );
  OAI21_X1 U7938 ( .B1(n11399), .B2(n7910), .A(n11464), .ZN(n7909) );
  INV_X1 U7939 ( .A(n9609), .ZN(n7910) );
  INV_X1 U7940 ( .A(n12421), .ZN(n7810) );
  NOR2_X1 U7941 ( .A1(n15294), .A2(n15298), .ZN(n7483) );
  AOI21_X1 U7942 ( .B1(n7466), .B2(n7468), .A(n7463), .ZN(n7462) );
  INV_X1 U7943 ( .A(n8320), .ZN(n7463) );
  NAND2_X1 U7944 ( .A1(n7449), .A2(n6928), .ZN(n6927) );
  INV_X1 U7945 ( .A(n8224), .ZN(n6928) );
  NAND2_X1 U7946 ( .A1(n8075), .A2(n10281), .ZN(n8078) );
  OAI21_X1 U7947 ( .B1(n10885), .B2(n10119), .A(n6846), .ZN(n6845) );
  NAND2_X1 U7948 ( .A1(n10885), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n6846) );
  NAND2_X1 U7949 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(n7191), .ZN(n7190) );
  INV_X1 U7950 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7191) );
  NAND2_X1 U7951 ( .A1(n7193), .A2(n6674), .ZN(n7192) );
  INV_X1 U7952 ( .A(n12993), .ZN(n7031) );
  INV_X1 U7953 ( .A(n9693), .ZN(n7412) );
  AOI21_X1 U7954 ( .B1(n7410), .B2(n9855), .A(n6598), .ZN(n7409) );
  NAND2_X1 U7955 ( .A1(n7890), .A2(n7888), .ZN(n7891) );
  NOR2_X1 U7956 ( .A1(n13336), .A2(n7889), .ZN(n7888) );
  OR2_X1 U7957 ( .A1(n13622), .A2(n12004), .ZN(n9718) );
  NAND2_X1 U7958 ( .A1(n6988), .A2(n6987), .ZN(n7265) );
  INV_X1 U7959 ( .A(n10746), .ZN(n6988) );
  OAI211_X1 U7960 ( .C1(n10986), .C2(n10985), .A(n7669), .B(n6683), .ZN(n7670)
         );
  NAND2_X1 U7961 ( .A1(n11568), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7297) );
  AND2_X1 U7962 ( .A1(n13198), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7678) );
  AOI21_X1 U7963 ( .B1(n13197), .B2(n13198), .A(n7680), .ZN(n6992) );
  INV_X1 U7964 ( .A(n13227), .ZN(n7680) );
  OR2_X1 U7965 ( .A1(n13269), .A2(n13279), .ZN(n7701) );
  AND2_X1 U7966 ( .A1(n9121), .A2(n7397), .ZN(n7396) );
  INV_X1 U7967 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n7397) );
  INV_X1 U7968 ( .A(n9432), .ZN(n9122) );
  AND2_X1 U7969 ( .A1(n9119), .A2(n9118), .ZN(n9394) );
  INV_X1 U7970 ( .A(n9395), .ZN(n9119) );
  INV_X1 U7971 ( .A(n9343), .ZN(n9117) );
  NOR2_X1 U7972 ( .A1(n9299), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7391) );
  INV_X1 U7973 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n7394) );
  OR2_X1 U7974 ( .A1(n9773), .A2(n6633), .ZN(n6858) );
  INV_X1 U7975 ( .A(n11382), .ZN(n10521) );
  NAND2_X1 U7976 ( .A1(n11046), .A2(n13121), .ZN(n9708) );
  OR2_X1 U7977 ( .A1(n9894), .A2(n12999), .ZN(n9703) );
  INV_X1 U7978 ( .A(n6964), .ZN(n6963) );
  OAI21_X1 U7979 ( .B1(n6622), .B2(n9676), .A(n13370), .ZN(n6964) );
  OR2_X1 U7980 ( .A1(n13649), .A2(n13433), .ZN(n9666) );
  NAND2_X1 U7981 ( .A1(n6884), .A2(n6883), .ZN(n7715) );
  AND2_X1 U7982 ( .A1(n6885), .A2(n7717), .ZN(n6884) );
  AND2_X1 U7983 ( .A1(n6691), .A2(n9789), .ZN(n7717) );
  INV_X1 U7984 ( .A(n7734), .ZN(n6889) );
  INV_X1 U7985 ( .A(n9787), .ZN(n7739) );
  NAND2_X1 U7986 ( .A1(n9786), .A2(n7741), .ZN(n7740) );
  AOI21_X1 U7987 ( .B1(n6566), .B2(n9775), .A(n7746), .ZN(n7745) );
  INV_X1 U7988 ( .A(n9779), .ZN(n7746) );
  OR2_X1 U7989 ( .A1(n12003), .A2(n13112), .ZN(n9624) );
  AND2_X1 U7990 ( .A1(n11372), .A2(n9777), .ZN(n11773) );
  NAND3_X1 U7991 ( .A1(n9094), .A2(n9199), .A3(n9093), .ZN(n9323) );
  INV_X1 U7992 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9099) );
  INV_X1 U7993 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9098) );
  NOR2_X1 U7994 ( .A1(n9070), .A2(n7885), .ZN(n7884) );
  INV_X1 U7995 ( .A(n9069), .ZN(n7885) );
  NAND2_X1 U7996 ( .A1(n7884), .A2(n7882), .ZN(n7881) );
  INV_X1 U7997 ( .A(n9422), .ZN(n7882) );
  NOR2_X1 U7998 ( .A1(n9570), .A2(n9735), .ZN(n9574) );
  AND2_X1 U7999 ( .A1(n9574), .A2(n9573), .ZN(n9727) );
  INV_X1 U8000 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9573) );
  INV_X1 U8001 ( .A(n7875), .ZN(n7874) );
  OAI21_X1 U8002 ( .B1(n9051), .B2(n7876), .A(n9055), .ZN(n7875) );
  INV_X1 U8003 ( .A(n9053), .ZN(n7876) );
  AND3_X1 U8004 ( .A1(n9324), .A2(n7625), .A3(n7624), .ZN(n9424) );
  AND2_X1 U8005 ( .A1(n9980), .A2(n9103), .ZN(n7624) );
  AND4_X1 U8006 ( .A1(n7626), .A2(n9102), .A3(n9101), .A4(n7662), .ZN(n7625)
         );
  AND2_X1 U8007 ( .A1(n7630), .A2(n7627), .ZN(n7626) );
  INV_X1 U8008 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9052) );
  NOR2_X1 U8009 ( .A1(n9259), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7275) );
  NAND2_X1 U8010 ( .A1(n10119), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9044) );
  INV_X1 U8011 ( .A(n7116), .ZN(n7115) );
  OAI21_X1 U8012 ( .B1(n9218), .B2(n7117), .A(n9040), .ZN(n7116) );
  INV_X1 U8013 ( .A(n9039), .ZN(n7117) );
  NOR2_X1 U8014 ( .A1(n9232), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n7309) );
  NAND2_X1 U8015 ( .A1(n10067), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9037) );
  INV_X1 U8016 ( .A(n11226), .ZN(n7354) );
  AND2_X1 U8017 ( .A1(n11922), .A2(n11921), .ZN(n7743) );
  NOR2_X1 U8018 ( .A1(n12600), .A2(n7362), .ZN(n7361) );
  INV_X1 U8019 ( .A(n12028), .ZN(n7362) );
  NOR2_X1 U8020 ( .A1(n8664), .A2(n8662), .ZN(n8673) );
  NAND2_X1 U8021 ( .A1(n7147), .A2(n14222), .ZN(n9017) );
  AND2_X1 U8022 ( .A1(n14240), .A2(n6583), .ZN(n7147) );
  INV_X1 U8023 ( .A(n14272), .ZN(n7148) );
  INV_X1 U8024 ( .A(n7778), .ZN(n7777) );
  OAI22_X1 U8025 ( .A1(n6573), .A2(n7785), .B1(n9019), .B2(n7782), .ZN(n7778)
         );
  NOR2_X1 U8026 ( .A1(n14167), .A2(n14194), .ZN(n7507) );
  NAND2_X1 U8027 ( .A1(n7021), .A2(n8721), .ZN(n7019) );
  AND2_X1 U8028 ( .A1(n7514), .A2(n7513), .ZN(n7512) );
  INV_X1 U8029 ( .A(n14469), .ZN(n7513) );
  INV_X1 U8030 ( .A(n7042), .ZN(n7037) );
  NAND2_X1 U8031 ( .A1(n7042), .A2(n7040), .ZN(n7039) );
  INV_X1 U8032 ( .A(n7786), .ZN(n7040) );
  OR2_X1 U8033 ( .A1(n14469), .A2(n13942), .ZN(n8590) );
  NAND2_X1 U8034 ( .A1(n7539), .A2(n7538), .ZN(n7537) );
  NOR2_X1 U8035 ( .A1(n7542), .A2(n8565), .ZN(n7538) );
  NOR2_X1 U8036 ( .A1(n8021), .A2(n14357), .ZN(n14337) );
  INV_X1 U8037 ( .A(n8547), .ZN(n7544) );
  NOR2_X1 U8038 ( .A1(n8512), .A2(n11681), .ZN(n7180) );
  INV_X1 U8039 ( .A(n7769), .ZN(n7768) );
  AND2_X1 U8040 ( .A1(n7056), .A2(n7054), .ZN(n7766) );
  NAND2_X1 U8041 ( .A1(n7509), .A2(n14513), .ZN(n7508) );
  INV_X1 U8042 ( .A(n7510), .ZN(n7509) );
  NOR2_X1 U8043 ( .A1(n8704), .A2(n7773), .ZN(n7772) );
  INV_X1 U8044 ( .A(n8701), .ZN(n7773) );
  NOR2_X1 U8045 ( .A1(n11934), .A2(n10558), .ZN(n6819) );
  NAND2_X1 U8046 ( .A1(n14223), .A2(n8723), .ZN(n14204) );
  INV_X1 U8047 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8086) );
  INV_X1 U8048 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8085) );
  NOR2_X2 U8049 ( .A1(n12343), .A2(n14614), .ZN(n6778) );
  AND2_X1 U8050 ( .A1(n14656), .A2(n6642), .ZN(n7990) );
  AOI21_X1 U8051 ( .B1(n7990), .B2(n7988), .A(n14725), .ZN(n7987) );
  INV_X1 U8052 ( .A(n14703), .ZN(n7988) );
  INV_X1 U8053 ( .A(n7990), .ZN(n7989) );
  INV_X1 U8054 ( .A(n12139), .ZN(n8006) );
  AND2_X1 U8055 ( .A1(n12551), .A2(n15538), .ZN(n10910) );
  AND2_X1 U8056 ( .A1(n6916), .A2(n12803), .ZN(n6915) );
  OR2_X1 U8057 ( .A1(n15253), .A2(n14989), .ZN(n14967) );
  NOR2_X1 U8058 ( .A1(n7958), .A2(n7957), .ZN(n7956) );
  INV_X1 U8059 ( .A(n12324), .ZN(n7958) );
  AND2_X1 U8060 ( .A1(n12270), .A2(n12760), .ZN(n7331) );
  NAND2_X1 U8061 ( .A1(n12248), .A2(n12886), .ZN(n7951) );
  AND2_X1 U8062 ( .A1(n15164), .A2(n12417), .ZN(n7794) );
  NAND2_X1 U8063 ( .A1(n7278), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11528) );
  INV_X1 U8064 ( .A(n11521), .ZN(n7278) );
  NOR2_X1 U8065 ( .A1(n15499), .A2(n12724), .ZN(n7489) );
  AND2_X1 U8066 ( .A1(n10354), .A2(n11280), .ZN(n12683) );
  NAND2_X1 U8067 ( .A1(n11027), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n11199) );
  INV_X1 U8068 ( .A(n11029), .ZN(n11027) );
  INV_X1 U8069 ( .A(n14787), .ZN(n11195) );
  NOR2_X1 U8070 ( .A1(n10356), .A2(n11317), .ZN(n12679) );
  INV_X1 U8071 ( .A(n7480), .ZN(n7478) );
  INV_X1 U8072 ( .A(n7814), .ZN(n7239) );
  NAND2_X1 U8073 ( .A1(n15142), .A2(n7483), .ZN(n15113) );
  INV_X1 U8074 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n10208) );
  NAND2_X1 U8075 ( .A1(n8363), .A2(n8362), .ZN(n8366) );
  OAI22_X1 U8076 ( .A1(n8356), .A2(n8355), .B1(SI_28_), .B2(n8354), .ZN(n8360)
         );
  XNOR2_X1 U8077 ( .A(n8279), .B(SI_18_), .ZN(n8256) );
  INV_X1 U8078 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10196) );
  OR2_X1 U8079 ( .A1(n10118), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n10198) );
  INV_X1 U8080 ( .A(n8071), .ZN(n7800) );
  INV_X1 U8081 ( .A(n8074), .ZN(n7799) );
  INV_X1 U8082 ( .A(n7803), .ZN(n7801) );
  AOI21_X1 U8083 ( .B1(n8063), .B2(n7319), .A(n6680), .ZN(n7316) );
  INV_X1 U8084 ( .A(n7315), .ZN(n7318) );
  OAI21_X1 U8085 ( .B1(n8061), .B2(n7319), .A(n8063), .ZN(n7315) );
  NAND2_X1 U8086 ( .A1(n6845), .A2(SI_8_), .ZN(n8062) );
  XNOR2_X1 U8087 ( .A(n6845), .B(SI_8_), .ZN(n8166) );
  INV_X1 U8088 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n10070) );
  OR2_X1 U8089 ( .A1(n10130), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n7649) );
  NAND2_X1 U8090 ( .A1(n10130), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n10131) );
  NAND2_X1 U8091 ( .A1(n10623), .A2(n10622), .ZN(n10941) );
  OR2_X1 U8092 ( .A1(n15410), .A2(n15409), .ZN(n15412) );
  INV_X1 U8093 ( .A(n13013), .ZN(n7032) );
  INV_X1 U8094 ( .A(n11596), .ZN(n7622) );
  NAND2_X1 U8095 ( .A1(n6774), .A2(n13019), .ZN(n12933) );
  NAND2_X1 U8096 ( .A1(n12933), .A2(n7632), .ZN(n13026) );
  INV_X1 U8097 ( .A(n7632), .ZN(n7015) );
  NAND2_X1 U8098 ( .A1(n7632), .A2(n7014), .ZN(n7013) );
  INV_X1 U8099 ( .A(n13019), .ZN(n7014) );
  NAND2_X1 U8100 ( .A1(n12957), .A2(n13085), .ZN(n7036) );
  OR2_X1 U8101 ( .A1(n9893), .A2(n9177), .ZN(n9560) );
  NAND2_X1 U8102 ( .A1(n7270), .A2(n10063), .ZN(n10984) );
  NAND2_X1 U8103 ( .A1(n10733), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10986) );
  NAND2_X1 U8104 ( .A1(n7576), .A2(n7581), .ZN(n7575) );
  INV_X1 U8105 ( .A(n10730), .ZN(n7576) );
  NAND2_X1 U8106 ( .A1(n9987), .A2(n10115), .ZN(n9990) );
  NAND2_X1 U8107 ( .A1(n7694), .A2(n9990), .ZN(n10783) );
  INV_X1 U8108 ( .A(n7695), .ZN(n7694) );
  AOI21_X1 U8109 ( .B1(n7567), .B2(n9977), .A(n7566), .ZN(n7565) );
  INV_X1 U8110 ( .A(n10968), .ZN(n7566) );
  NAND2_X1 U8111 ( .A1(n10950), .A2(n10963), .ZN(n6995) );
  NOR2_X1 U8112 ( .A1(n10950), .A2(n10963), .ZN(n11080) );
  AOI21_X1 U8113 ( .B1(n7565), .B2(n7568), .A(n7563), .ZN(n7562) );
  INV_X1 U8114 ( .A(n11069), .ZN(n7563) );
  INV_X1 U8115 ( .A(n7565), .ZN(n7564) );
  OR2_X1 U8116 ( .A1(n11561), .A2(n11569), .ZN(n6991) );
  NAND2_X1 U8117 ( .A1(n7562), .A2(n7564), .ZN(n6976) );
  AND2_X1 U8118 ( .A1(n13147), .A2(n6753), .ZN(n7664) );
  NOR2_X1 U8119 ( .A1(n13185), .A2(n13184), .ZN(n13193) );
  NOR2_X1 U8120 ( .A1(n7587), .A2(n13212), .ZN(n7583) );
  OR2_X1 U8121 ( .A1(n13174), .A2(n7584), .ZN(n13206) );
  NAND2_X1 U8122 ( .A1(n13176), .A2(n7585), .ZN(n7584) );
  INV_X1 U8123 ( .A(n7588), .ZN(n7585) );
  NAND2_X1 U8124 ( .A1(n13299), .A2(n6973), .ZN(n13327) );
  OR2_X1 U8125 ( .A1(n13300), .A2(n13301), .ZN(n6973) );
  OAI21_X1 U8126 ( .B1(n7723), .B2(n7720), .A(n8027), .ZN(n7719) );
  AND2_X1 U8127 ( .A1(n13351), .A2(n13355), .ZN(n7259) );
  NAND2_X1 U8128 ( .A1(n9124), .A2(n9123), .ZN(n9509) );
  INV_X1 U8129 ( .A(n9497), .ZN(n9124) );
  NAND2_X1 U8130 ( .A1(n9122), .A2(n9121), .ZN(n9442) );
  NAND2_X1 U8131 ( .A1(n9117), .A2(n7392), .ZN(n9395) );
  AND2_X1 U8132 ( .A1(n6606), .A2(n15910), .ZN(n7392) );
  NAND2_X1 U8133 ( .A1(n9117), .A2(n9116), .ZN(n9361) );
  NAND2_X1 U8134 ( .A1(n8009), .A2(n11373), .ZN(n11372) );
  NAND2_X1 U8135 ( .A1(n6857), .A2(n6858), .ZN(n8009) );
  AND4_X1 U8136 ( .A1(n9287), .A2(n9286), .A3(n9285), .A4(n9284), .ZN(n11845)
         );
  NAND2_X1 U8137 ( .A1(n6959), .A2(n9603), .ZN(n11400) );
  AND2_X1 U8138 ( .A1(n9763), .A2(n9827), .ZN(n13394) );
  NAND2_X1 U8139 ( .A1(n7912), .A2(n9695), .ZN(n7911) );
  NAND2_X1 U8140 ( .A1(n9695), .A2(n13355), .ZN(n7913) );
  NAND2_X1 U8141 ( .A1(n9696), .A2(n7914), .ZN(n7912) );
  NOR2_X1 U8142 ( .A1(n7709), .A2(n13407), .ZN(n6895) );
  INV_X1 U8143 ( .A(n7751), .ZN(n7750) );
  AOI21_X1 U8144 ( .B1(n7710), .B2(n7708), .A(n6695), .ZN(n7707) );
  INV_X1 U8145 ( .A(n9800), .ZN(n7708) );
  NAND2_X1 U8146 ( .A1(n9683), .A2(n9684), .ZN(n13363) );
  NOR2_X2 U8147 ( .A1(n13370), .A2(n7711), .ZN(n7710) );
  INV_X1 U8148 ( .A(n9801), .ZN(n7711) );
  NAND2_X1 U8149 ( .A1(n7712), .A2(n9801), .ZN(n13371) );
  NAND2_X1 U8150 ( .A1(n13410), .A2(n6622), .ZN(n13383) );
  NAND2_X1 U8151 ( .A1(n13443), .A2(n7753), .ZN(n13428) );
  AND2_X1 U8152 ( .A1(n9666), .A2(n9667), .ZN(n13417) );
  INV_X1 U8153 ( .A(n13108), .ZN(n13476) );
  NAND2_X1 U8154 ( .A1(n13442), .A2(n13441), .ZN(n13440) );
  AND2_X1 U8155 ( .A1(n9449), .A2(n9448), .ZN(n13460) );
  NOR2_X1 U8156 ( .A1(n13473), .A2(n7919), .ZN(n7918) );
  INV_X1 U8157 ( .A(n9652), .ZN(n7919) );
  AOI21_X1 U8158 ( .B1(n13477), .B2(n9547), .A(n9421), .ZN(n13490) );
  AOI21_X1 U8159 ( .B1(n7927), .B2(n6661), .A(n6968), .ZN(n6967) );
  NAND2_X1 U8160 ( .A1(n12104), .A2(n6965), .ZN(n6966) );
  INV_X1 U8161 ( .A(n9645), .ZN(n6968) );
  AND2_X1 U8162 ( .A1(n9410), .A2(n9409), .ZN(n13504) );
  NAND2_X1 U8163 ( .A1(n9639), .A2(n9638), .ZN(n7937) );
  INV_X1 U8164 ( .A(n7929), .ZN(n7928) );
  NAND2_X1 U8165 ( .A1(n6970), .A2(n9629), .ZN(n13545) );
  AND2_X1 U8166 ( .A1(n9961), .A2(n9765), .ZN(n13547) );
  NAND2_X1 U8167 ( .A1(n9289), .A2(n9288), .ZN(n7904) );
  NAND2_X1 U8168 ( .A1(n9821), .A2(n9822), .ZN(n10082) );
  INV_X1 U8169 ( .A(n12057), .ZN(n9821) );
  AOI21_X1 U8170 ( .B1(n6610), .B2(n7894), .A(n6758), .ZN(n7892) );
  OAI21_X1 U8171 ( .B1(n7124), .B2(n7121), .A(n7119), .ZN(n7893) );
  INV_X1 U8172 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n9130) );
  XNOR2_X1 U8173 ( .A(n9104), .B(n9128), .ZN(n9747) );
  NAND2_X1 U8174 ( .A1(n7756), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9104) );
  INV_X1 U8175 ( .A(n9739), .ZN(n9105) );
  XNOR2_X1 U8176 ( .A(n9107), .B(n9106), .ZN(n9748) );
  NAND2_X1 U8177 ( .A1(n9739), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9107) );
  NAND2_X1 U8178 ( .A1(n7118), .A2(n9083), .ZN(n9526) );
  NAND2_X1 U8179 ( .A1(n7124), .A2(n7122), .ZN(n7118) );
  NAND2_X1 U8180 ( .A1(n6558), .A2(n7245), .ZN(n9743) );
  INV_X1 U8181 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7245) );
  INV_X1 U8182 ( .A(n9727), .ZN(n9582) );
  NOR2_X1 U8183 ( .A1(n9426), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n7639) );
  AND2_X1 U8184 ( .A1(n9048), .A2(n9047), .ZN(n9290) );
  AND2_X1 U8185 ( .A1(n9046), .A2(n9045), .ZN(n9271) );
  OR2_X1 U8186 ( .A1(n9257), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n9259) );
  NAND2_X1 U8187 ( .A1(n10069), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9039) );
  NAND2_X1 U8188 ( .A1(n9219), .A2(n9218), .ZN(n9221) );
  NAND2_X1 U8189 ( .A1(n9200), .A2(n9199), .ZN(n9232) );
  INV_X1 U8190 ( .A(n9198), .ZN(n9200) );
  AND2_X1 U8191 ( .A1(n9035), .A2(n9034), .ZN(n9183) );
  XNOR2_X1 U8192 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7093) );
  INV_X1 U8193 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n9953) );
  AND2_X1 U8194 ( .A1(n12623), .A2(n12616), .ZN(n7729) );
  OR2_X1 U8195 ( .A1(n8601), .A2(n13894), .ZN(n8610) );
  AOI21_X1 U8196 ( .B1(n7358), .B2(n7360), .A(n7356), .ZN(n7355) );
  INV_X1 U8197 ( .A(n13881), .ZN(n7356) );
  INV_X1 U8198 ( .A(n7353), .ZN(n7352) );
  OAI21_X1 U8199 ( .B1(n10854), .B2(n7354), .A(n11225), .ZN(n7353) );
  INV_X1 U8200 ( .A(n12631), .ZN(n7385) );
  NAND2_X1 U8201 ( .A1(n7371), .A2(n7370), .ZN(n13729) );
  NAND2_X1 U8202 ( .A1(n8519), .A2(n8518), .ZN(n8530) );
  NAND2_X1 U8203 ( .A1(n8608), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8619) );
  INV_X1 U8204 ( .A(n8610), .ZN(n8608) );
  INV_X1 U8205 ( .A(n13834), .ZN(n7387) );
  AND2_X1 U8206 ( .A1(n11262), .A2(n11255), .ZN(n7733) );
  NAND2_X1 U8207 ( .A1(n8673), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8734) );
  AND2_X2 U8208 ( .A1(n13755), .A2(n12624), .ZN(n13823) );
  AND2_X1 U8209 ( .A1(n8782), .A2(n6562), .ZN(n10427) );
  AOI21_X1 U8210 ( .B1(n14014), .B2(n6806), .A(n6628), .ZN(n6805) );
  INV_X1 U8211 ( .A(n10421), .ZN(n6806) );
  INV_X1 U8212 ( .A(n14014), .ZN(n6807) );
  NAND2_X1 U8213 ( .A1(n6801), .A2(n6800), .ZN(n10716) );
  INV_X1 U8214 ( .A(n10719), .ZN(n6800) );
  INV_X1 U8215 ( .A(n10718), .ZN(n6801) );
  NAND2_X1 U8216 ( .A1(n6799), .A2(n6798), .ZN(n10865) );
  INV_X1 U8217 ( .A(n10868), .ZN(n6798) );
  INV_X1 U8218 ( .A(n10867), .ZN(n6799) );
  NOR2_X1 U8219 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n7749) );
  OR2_X1 U8220 ( .A1(n11881), .A2(n6788), .ZN(n6787) );
  INV_X1 U8221 ( .A(n11823), .ZN(n6788) );
  NAND2_X1 U8222 ( .A1(n11882), .A2(n11881), .ZN(n11880) );
  AND2_X1 U8223 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n8270) );
  AND2_X1 U8224 ( .A1(n8744), .A2(n8743), .ZN(n9917) );
  INV_X1 U8225 ( .A(n7558), .ZN(n7556) );
  NAND2_X1 U8226 ( .A1(n14541), .A2(n13731), .ZN(n7558) );
  OR2_X1 U8227 ( .A1(n14174), .A2(n8655), .ZN(n7557) );
  NAND2_X1 U8228 ( .A1(n7531), .A2(n6592), .ZN(n14189) );
  OR2_X1 U8229 ( .A1(n6572), .A2(n8721), .ZN(n7020) );
  INV_X1 U8230 ( .A(n9016), .ZN(n14213) );
  OR2_X1 U8231 ( .A1(n14230), .A2(n14214), .ZN(n14216) );
  OR2_X1 U8232 ( .A1(n14456), .A2(n13939), .ZN(n9014) );
  NAND2_X1 U8233 ( .A1(n7175), .A2(n8606), .ZN(n14261) );
  AND2_X1 U8234 ( .A1(n7337), .A2(n7043), .ZN(n7042) );
  NAND2_X1 U8235 ( .A1(n7786), .A2(n8714), .ZN(n7043) );
  NAND2_X1 U8236 ( .A1(n14315), .A2(n7786), .ZN(n7038) );
  AOI21_X1 U8237 ( .B1(n7337), .B2(n8715), .A(n6640), .ZN(n7336) );
  NAND2_X1 U8238 ( .A1(n7041), .A2(n7786), .ZN(n14299) );
  OR2_X1 U8239 ( .A1(n14315), .A2(n8714), .ZN(n7041) );
  CLKBUF_X1 U8240 ( .A(n14281), .Z(n14303) );
  NAND2_X1 U8241 ( .A1(n7005), .A2(n7003), .ZN(n14333) );
  INV_X1 U8242 ( .A(n7004), .ZN(n7003) );
  NAND2_X1 U8243 ( .A1(n8708), .A2(n7760), .ZN(n7005) );
  OAI21_X1 U8244 ( .B1(n7761), .B2(n8709), .A(n6689), .ZN(n7004) );
  INV_X1 U8245 ( .A(n8538), .ZN(n7548) );
  OR2_X1 U8246 ( .A1(n8541), .A2(n8540), .ZN(n8550) );
  NAND2_X1 U8247 ( .A1(n11973), .A2(n8692), .ZN(n11707) );
  OR2_X1 U8248 ( .A1(n8781), .A2(n7528), .ZN(n8453) );
  OR2_X1 U8249 ( .A1(n15716), .A2(n6562), .ZN(n10035) );
  NAND2_X1 U8250 ( .A1(n8788), .A2(n10558), .ZN(n11969) );
  AND2_X1 U8251 ( .A1(n6814), .A2(n6705), .ZN(n14100) );
  NAND2_X1 U8252 ( .A1(n9903), .A2(n9922), .ZN(n6814) );
  NAND2_X1 U8253 ( .A1(n8288), .A2(n8287), .ZN(n14451) );
  OAI211_X1 U8254 ( .C1(n10428), .C2(n13977), .A(n8139), .B(n8138), .ZN(n10851) );
  OR3_X1 U8255 ( .A1(n12119), .A2(n11788), .A3(n11895), .ZN(n9929) );
  XNOR2_X1 U8256 ( .A(n8418), .B(n8417), .ZN(n10426) );
  AND2_X1 U8257 ( .A1(n14695), .A2(n12549), .ZN(n14608) );
  NAND2_X1 U8258 ( .A1(n14704), .A2(n14703), .ZN(n7991) );
  AND2_X1 U8259 ( .A1(n12570), .A2(n12569), .ZN(n14665) );
  AND2_X1 U8260 ( .A1(n7999), .A2(n12489), .ZN(n7998) );
  AND2_X1 U8261 ( .A1(n7997), .A2(n7999), .ZN(n7996) );
  INV_X1 U8262 ( .A(n12505), .ZN(n7997) );
  NAND2_X1 U8263 ( .A1(n12550), .A2(n14608), .ZN(n14610) );
  AND2_X1 U8264 ( .A1(n14664), .A2(n12561), .ZN(n14696) );
  NAND2_X1 U8265 ( .A1(n14734), .A2(n6662), .ZN(n14629) );
  AND2_X1 U8266 ( .A1(n14607), .A2(n12541), .ZN(n14724) );
  OAI22_X1 U8267 ( .A1(n14636), .A2(n11353), .B1(n15537), .B2(n10699), .ZN(
        n10880) );
  INV_X1 U8268 ( .A(n11323), .ZN(n7133) );
  NAND2_X1 U8269 ( .A1(n6841), .A2(n6839), .ZN(n14745) );
  AOI21_X1 U8270 ( .B1(n6617), .B2(n6844), .A(n6840), .ZN(n6839) );
  INV_X1 U8271 ( .A(n12570), .ZN(n6840) );
  AND2_X1 U8272 ( .A1(n12359), .A2(n12358), .ZN(n14748) );
  AND2_X1 U8273 ( .A1(n12349), .A2(n12348), .ZN(n14729) );
  OAI21_X1 U8274 ( .B1(n7080), .B2(n7077), .A(n7079), .ZN(n7076) );
  NOR2_X1 U8275 ( .A1(n11117), .A2(n7083), .ZN(n7079) );
  NAND2_X1 U8276 ( .A1(n7074), .A2(n7073), .ZN(n11113) );
  NAND2_X1 U8277 ( .A1(n11477), .A2(n6879), .ZN(n6878) );
  NAND2_X1 U8278 ( .A1(n14869), .A2(n7502), .ZN(n6867) );
  NOR2_X1 U8279 ( .A1(n14903), .A2(n14911), .ZN(n15805) );
  XNOR2_X1 U8280 ( .A(n12678), .B(n14772), .ZN(n14999) );
  AND2_X1 U8281 ( .A1(n12382), .A2(n12381), .ZN(n14990) );
  OR2_X1 U8282 ( .A1(n14976), .A2(n11447), .ZN(n12382) );
  AND2_X1 U8283 ( .A1(n12323), .A2(n12322), .ZN(n15071) );
  NOR2_X1 U8284 ( .A1(n12422), .A2(n7813), .ZN(n7812) );
  INV_X1 U8285 ( .A(n12419), .ZN(n7813) );
  AND2_X1 U8286 ( .A1(n12292), .A2(n12291), .ZN(n15131) );
  NAND2_X1 U8287 ( .A1(n7229), .A2(n12418), .ZN(n7228) );
  OR2_X1 U8288 ( .A1(n15308), .A2(n14681), .ZN(n12760) );
  NOR2_X1 U8289 ( .A1(n15308), .A2(n15176), .ZN(n15169) );
  INV_X1 U8290 ( .A(n7284), .ZN(n12265) );
  OR2_X1 U8291 ( .A1(n15314), .A2(n14758), .ZN(n15163) );
  NAND2_X1 U8292 ( .A1(n15192), .A2(n7794), .ZN(n15157) );
  OR2_X1 U8293 ( .A1(n6584), .A2(n6565), .ZN(n7220) );
  NAND2_X1 U8294 ( .A1(n7489), .A2(n7488), .ZN(n7487) );
  INV_X1 U8295 ( .A(n7327), .ZN(n7326) );
  NAND2_X1 U8296 ( .A1(n6942), .A2(n6665), .ZN(n7325) );
  OAI21_X1 U8297 ( .B1(n7328), .B2(n12883), .A(n12014), .ZN(n7327) );
  NAND2_X1 U8298 ( .A1(n12061), .A2(n11547), .ZN(n15493) );
  NAND2_X1 U8299 ( .A1(n12871), .A2(n11175), .ZN(n11159) );
  OR2_X1 U8300 ( .A1(n15538), .A2(n15819), .ZN(n11130) );
  NAND2_X1 U8301 ( .A1(n8015), .A2(n15212), .ZN(n15213) );
  OR2_X1 U8302 ( .A1(n15207), .A2(n15538), .ZN(n8015) );
  INV_X1 U8303 ( .A(n14980), .ZN(n15236) );
  INV_X1 U8304 ( .A(n15059), .ZN(n15271) );
  NAND2_X1 U8305 ( .A1(n12010), .A2(n12009), .ZN(n15331) );
  OR2_X1 U8306 ( .A1(n11320), .A2(n12672), .ZN(n15566) );
  OR2_X1 U8307 ( .A1(n10386), .A2(n10385), .ZN(n15599) );
  NAND2_X1 U8308 ( .A1(n15566), .A2(n15565), .ZN(n15561) );
  OR3_X1 U8309 ( .A1(n10187), .A2(n10186), .A3(n12588), .ZN(n10349) );
  XNOR2_X1 U8310 ( .A(n10258), .B(P1_IR_REG_29__SCAN_IN), .ZN(n10259) );
  XNOR2_X1 U8311 ( .A(n8341), .B(n8337), .ZN(n12372) );
  INV_X1 U8312 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9944) );
  INV_X1 U8313 ( .A(n9949), .ZN(n9945) );
  XNOR2_X1 U8314 ( .A(n10203), .B(P1_IR_REG_21__SCAN_IN), .ZN(n10354) );
  NAND2_X1 U8315 ( .A1(n10202), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10203) );
  XNOR2_X1 U8316 ( .A(n8293), .B(n8292), .ZN(n12312) );
  XNOR2_X1 U8317 ( .A(n10331), .B(P1_IR_REG_20__SCAN_IN), .ZN(n12675) );
  XNOR2_X1 U8318 ( .A(n8208), .B(n8079), .ZN(n12244) );
  AND2_X1 U8319 ( .A1(n10551), .A2(n10314), .ZN(n14859) );
  XNOR2_X1 U8320 ( .A(n8190), .B(n8189), .ZN(n12007) );
  XNOR2_X1 U8321 ( .A(n8155), .B(n8156), .ZN(n11189) );
  NAND2_X1 U8322 ( .A1(n10050), .A2(n9931), .ZN(n10093) );
  INV_X1 U8323 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7305) );
  NOR2_X1 U8324 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n10050) );
  NAND2_X1 U8325 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7306) );
  NAND2_X1 U8326 ( .A1(n10137), .A2(n10136), .ZN(n10159) );
  NAND2_X1 U8327 ( .A1(n12047), .A2(n12192), .ZN(n7655) );
  NAND2_X1 U8328 ( .A1(n7274), .A2(n7621), .ZN(n11607) );
  AND2_X1 U8329 ( .A1(n11592), .A2(n7622), .ZN(n7621) );
  NAND2_X1 U8330 ( .A1(n7706), .A2(n12947), .ZN(n7252) );
  OAI21_X1 U8331 ( .B1(n12952), .B2(n12951), .A(n12950), .ZN(n12953) );
  CLKBUF_X1 U8332 ( .A(n11593), .Z(n7274) );
  AOI21_X1 U8333 ( .B1(n13435), .B2(n9547), .A(n9464), .ZN(n13446) );
  AND2_X1 U8334 ( .A1(n9492), .A2(n9491), .ZN(n13069) );
  AND2_X1 U8335 ( .A1(n9237), .A2(n9236), .ZN(n11411) );
  NAND2_X1 U8336 ( .A1(n10536), .A2(n10535), .ZN(n13104) );
  NAND2_X1 U8337 ( .A1(n10512), .A2(n10514), .ZN(n13099) );
  AOI21_X1 U8338 ( .B1(n13343), .B2(n9547), .A(n9546), .ZN(n13352) );
  NAND2_X1 U8339 ( .A1(n9523), .A2(n9522), .ZN(n13375) );
  INV_X1 U8340 ( .A(n13069), .ZN(n13421) );
  NAND2_X1 U8341 ( .A1(n9478), .A2(n9477), .ZN(n13106) );
  INV_X1 U8342 ( .A(n13460), .ZN(n13107) );
  NAND4_X1 U8343 ( .A1(n9231), .A2(n9230), .A3(n9229), .A4(n9228), .ZN(n13117)
         );
  NOR2_X1 U8344 ( .A1(n6982), .A2(n10106), .ZN(n7579) );
  NAND2_X1 U8345 ( .A1(n9196), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9182) );
  NAND2_X1 U8346 ( .A1(n11071), .A2(n11070), .ZN(n11553) );
  NOR2_X1 U8347 ( .A1(n13173), .A2(n13613), .ZN(n13199) );
  NAND2_X1 U8348 ( .A1(n13259), .A2(n13258), .ZN(n13271) );
  INV_X1 U8349 ( .A(n7677), .ZN(n13250) );
  INV_X1 U8350 ( .A(n13002), .ZN(n13345) );
  XNOR2_X1 U8351 ( .A(n9755), .B(n9754), .ZN(n13342) );
  NAND2_X1 U8352 ( .A1(n7287), .A2(n6737), .ZN(n13347) );
  NAND2_X1 U8353 ( .A1(n10535), .A2(n9888), .ZN(n13479) );
  NAND2_X1 U8354 ( .A1(n9298), .A2(n9297), .ZN(n12053) );
  NAND2_X1 U8355 ( .A1(n9280), .A2(n9279), .ZN(n11985) );
  NAND2_X1 U8356 ( .A1(n15804), .A2(n13598), .ZN(n13610) );
  AOI21_X1 U8357 ( .B1(n13342), .B2(n15755), .A(n13347), .ZN(n9861) );
  OR2_X1 U8358 ( .A1(n15788), .A2(n15770), .ZN(n13688) );
  NAND2_X1 U8359 ( .A1(n8188), .A2(n8187), .ZN(n14367) );
  NAND2_X1 U8360 ( .A1(n8207), .A2(n8206), .ZN(n14339) );
  INV_X1 U8361 ( .A(n14545), .ZN(n14194) );
  NAND2_X1 U8362 ( .A1(n10037), .A2(n14398), .ZN(n13923) );
  XNOR2_X1 U8363 ( .A(n7163), .B(n14086), .ZN(n9022) );
  NAND2_X1 U8364 ( .A1(n9021), .A2(n7164), .ZN(n7163) );
  AND2_X1 U8365 ( .A1(n9020), .A2(n6586), .ZN(n7164) );
  NAND2_X1 U8366 ( .A1(n8670), .A2(n8669), .ZN(n13933) );
  INV_X1 U8367 ( .A(n13893), .ZN(n13939) );
  INV_X1 U8368 ( .A(n12639), .ZN(n13940) );
  OR3_X1 U8369 ( .A1(n8600), .A2(n8599), .A3(n8598), .ZN(n13941) );
  OR2_X1 U8370 ( .A1(n10424), .A2(n10425), .ZN(n10477) );
  OR2_X1 U8371 ( .A1(n10481), .A2(n10482), .ZN(n10842) );
  AND2_X1 U8372 ( .A1(n8199), .A2(n8203), .ZN(n10495) );
  NAND2_X1 U8373 ( .A1(n6794), .A2(n6793), .ZN(n6792) );
  NAND2_X1 U8374 ( .A1(n14084), .A2(n15644), .ZN(n6793) );
  NAND2_X1 U8375 ( .A1(n14085), .A2(n15653), .ZN(n6794) );
  OAI21_X1 U8376 ( .B1(n14085), .B2(n15623), .A(n6797), .ZN(n6796) );
  NOR2_X1 U8377 ( .A1(n6589), .A2(n15651), .ZN(n6797) );
  OR2_X1 U8378 ( .A1(n15658), .A2(n8037), .ZN(n6790) );
  NAND2_X1 U8379 ( .A1(n7160), .A2(n9900), .ZN(n7158) );
  NAND2_X1 U8380 ( .A1(n7296), .A2(n13750), .ZN(n14124) );
  OR2_X1 U8381 ( .A1(n8748), .A2(n14375), .ZN(n7296) );
  INV_X1 U8382 ( .A(n7781), .ZN(n8752) );
  AND2_X1 U8383 ( .A1(n8323), .A2(n8322), .ZN(n14537) );
  NAND2_X1 U8384 ( .A1(n8378), .A2(n8377), .ZN(n8995) );
  NOR2_X1 U8385 ( .A1(n14108), .A2(n8770), .ZN(n12589) );
  INV_X1 U8386 ( .A(n14113), .ZN(n8768) );
  NAND2_X1 U8387 ( .A1(n8346), .A2(n8345), .ZN(n13752) );
  NOR2_X1 U8388 ( .A1(n14124), .A2(n7102), .ZN(n14413) );
  NAND2_X1 U8389 ( .A1(n7295), .A2(n7294), .ZN(n7102) );
  INV_X1 U8390 ( .A(n14119), .ZN(n7294) );
  NAND2_X1 U8391 ( .A1(n14118), .A2(n15740), .ZN(n7295) );
  INV_X1 U8392 ( .A(n14130), .ZN(n14530) );
  NAND2_X1 U8393 ( .A1(n7342), .A2(n7341), .ZN(n7340) );
  INV_X1 U8394 ( .A(n14416), .ZN(n7341) );
  OR2_X1 U8395 ( .A1(n14425), .A2(n7049), .ZN(n7048) );
  AOI21_X1 U8396 ( .B1(n14427), .B2(n15740), .A(n14426), .ZN(n7050) );
  NAND2_X1 U8397 ( .A1(n8421), .A2(n8420), .ZN(n15701) );
  OR2_X1 U8398 ( .A1(n8385), .A2(n8386), .ZN(n8388) );
  NAND2_X1 U8399 ( .A1(n11434), .A2(n11433), .ZN(n7970) );
  INV_X1 U8400 ( .A(n15179), .ZN(n14681) );
  AND2_X1 U8401 ( .A1(n12342), .A2(n12341), .ZN(n14619) );
  NAND2_X1 U8402 ( .A1(n12296), .A2(n12295), .ZN(n15287) );
  AOI21_X1 U8403 ( .B1(n7971), .B2(n7973), .A(n6648), .ZN(n7969) );
  NAND2_X1 U8404 ( .A1(n11434), .A2(n7971), .ZN(n7968) );
  AND2_X1 U8405 ( .A1(n12310), .A2(n12309), .ZN(n15090) );
  INV_X1 U8406 ( .A(n14773), .ZN(n14989) );
  AND3_X1 U8407 ( .A1(n12280), .A2(n12279), .A3(n12278), .ZN(n14680) );
  NAND2_X1 U8408 ( .A1(n12392), .A2(n12391), .ZN(n14770) );
  INV_X1 U8409 ( .A(n14748), .ZN(n14772) );
  INV_X1 U8410 ( .A(n14729), .ZN(n14774) );
  NAND2_X1 U8411 ( .A1(n12337), .A2(n12336), .ZN(n15051) );
  OR2_X1 U8412 ( .A1(n15040), .A2(n11447), .ZN(n12337) );
  INV_X1 U8413 ( .A(n15071), .ZN(n14775) );
  INV_X1 U8414 ( .A(n15090), .ZN(n15050) );
  INV_X1 U8415 ( .A(n14680), .ZN(n15151) );
  OAI21_X1 U8416 ( .B1(P1_REG1_REG_1__SCAN_IN), .B2(n10666), .A(n7307), .ZN(
        n14802) );
  NAND2_X1 U8417 ( .A1(n10666), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7307) );
  AND2_X1 U8418 ( .A1(n6759), .A2(n10267), .ZN(n10294) );
  AND2_X1 U8419 ( .A1(n7065), .A2(n7062), .ZN(n14848) );
  NOR2_X1 U8420 ( .A1(n10291), .A2(n7063), .ZN(n7062) );
  NOR2_X1 U8421 ( .A1(n10321), .A2(n7064), .ZN(n7063) );
  NAND2_X1 U8422 ( .A1(n11119), .A2(n11120), .ZN(n11477) );
  XNOR2_X1 U8423 ( .A(n10552), .B(P1_IR_REG_14__SCAN_IN), .ZN(n14868) );
  NAND2_X1 U8424 ( .A1(n6869), .A2(n6751), .ZN(n6864) );
  AND2_X1 U8425 ( .A1(n6867), .A2(n6866), .ZN(n6865) );
  INV_X1 U8426 ( .A(n7491), .ZN(n14901) );
  NAND2_X1 U8427 ( .A1(n7087), .A2(n12672), .ZN(n7497) );
  NAND2_X1 U8428 ( .A1(n12445), .A2(n7213), .ZN(n15214) );
  INV_X1 U8429 ( .A(n12442), .ZN(n12443) );
  XNOR2_X1 U8430 ( .A(n14930), .B(n14935), .ZN(n15218) );
  NAND2_X1 U8431 ( .A1(n15214), .A2(n15561), .ZN(n7789) );
  NAND2_X1 U8432 ( .A1(n15606), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7945) );
  AND2_X1 U8433 ( .A1(n7941), .A2(n6588), .ZN(n7939) );
  NAND2_X1 U8434 ( .A1(n7946), .A2(n7943), .ZN(n7942) );
  NOR2_X1 U8435 ( .A1(n12441), .A2(n6619), .ZN(n7943) );
  INV_X1 U8436 ( .A(n10257), .ZN(n10255) );
  INV_X1 U8437 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n10254) );
  NAND2_X1 U8438 ( .A1(n10163), .A2(n10164), .ZN(n10165) );
  NAND2_X1 U8439 ( .A1(n10165), .A2(n13984), .ZN(n7651) );
  NAND2_X1 U8440 ( .A1(n10161), .A2(n10162), .ZN(n10603) );
  AND2_X1 U8441 ( .A1(n11302), .A2(n7658), .ZN(n7659) );
  INV_X1 U8442 ( .A(n11308), .ZN(n7658) );
  NAND2_X1 U8443 ( .A1(n11309), .A2(n11308), .ZN(n11670) );
  NAND2_X1 U8444 ( .A1(n15403), .A2(n15402), .ZN(n15408) );
  NAND2_X1 U8445 ( .A1(n15399), .A2(n15398), .ZN(n15407) );
  NAND2_X1 U8446 ( .A1(n15401), .A2(n15400), .ZN(n15403) );
  NAND2_X1 U8447 ( .A1(n15433), .A2(n15432), .ZN(n15435) );
  NAND2_X1 U8448 ( .A1(n15430), .A2(n15429), .ZN(n15434) );
  NAND3_X1 U8449 ( .A1(n15454), .A2(n7199), .A3(n7197), .ZN(n15452) );
  INV_X1 U8450 ( .A(n15451), .ZN(n7201) );
  NOR2_X1 U8451 ( .A1(n15452), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n15456) );
  OR2_X1 U8452 ( .A1(n6561), .A2(n15660), .ZN(n8783) );
  NAND2_X1 U8453 ( .A1(n7820), .A2(n7817), .ZN(n8806) );
  INV_X1 U8454 ( .A(n8824), .ZN(n7855) );
  NOR2_X1 U8455 ( .A1(n8824), .A2(n7857), .ZN(n7856) );
  AOI21_X1 U8456 ( .B1(n9602), .B2(n7423), .A(n6597), .ZN(n7422) );
  INV_X1 U8457 ( .A(n12742), .ZN(n7612) );
  INV_X1 U8458 ( .A(n8845), .ZN(n7834) );
  NAND2_X1 U8459 ( .A1(n12755), .A2(n12756), .ZN(n7599) );
  INV_X1 U8460 ( .A(n12763), .ZN(n7600) );
  NAND2_X1 U8461 ( .A1(n7446), .A2(n6646), .ZN(n7445) );
  NAND2_X1 U8462 ( .A1(n7443), .A2(n9630), .ZN(n7442) );
  INV_X1 U8463 ( .A(n9631), .ZN(n7444) );
  NAND2_X1 U8464 ( .A1(n6699), .A2(n7831), .ZN(n7830) );
  NAND2_X1 U8465 ( .A1(n7838), .A2(n8845), .ZN(n7831) );
  NAND2_X1 U8466 ( .A1(n8874), .A2(n7832), .ZN(n7829) );
  NAND2_X1 U8467 ( .A1(n7833), .A2(n7837), .ZN(n7832) );
  INV_X1 U8468 ( .A(n8875), .ZN(n7837) );
  OR2_X1 U8469 ( .A1(n7835), .A2(n6728), .ZN(n7833) );
  INV_X1 U8470 ( .A(n12762), .ZN(n7598) );
  NAND2_X1 U8471 ( .A1(n9665), .A2(n13417), .ZN(n7439) );
  INV_X1 U8472 ( .A(n7434), .ZN(n7433) );
  INV_X1 U8473 ( .A(n7436), .ZN(n7435) );
  AND2_X1 U8474 ( .A1(n7864), .A2(n8908), .ZN(n7859) );
  INV_X1 U8475 ( .A(n8910), .ZN(n7863) );
  NAND2_X1 U8476 ( .A1(n8920), .A2(n8919), .ZN(n7852) );
  OAI21_X1 U8477 ( .B1(n7592), .B2(n7590), .A(n12778), .ZN(n7324) );
  AND2_X1 U8478 ( .A1(n7594), .A2(n12791), .ZN(n7590) );
  AOI21_X1 U8479 ( .B1(n7853), .B2(n7852), .A(n8923), .ZN(n7850) );
  AOI21_X1 U8480 ( .B1(n7798), .B2(n7801), .A(n7797), .ZN(n7796) );
  NAND2_X1 U8481 ( .A1(n12800), .A2(n12801), .ZN(n6922) );
  NAND2_X1 U8482 ( .A1(n12816), .A2(n12674), .ZN(n12808) );
  INV_X1 U8483 ( .A(n12151), .ZN(n7950) );
  INV_X1 U8484 ( .A(n7467), .ZN(n7466) );
  OAI21_X1 U8485 ( .B1(n6577), .B2(n7468), .A(n8313), .ZN(n7467) );
  NAND2_X1 U8486 ( .A1(n7449), .A2(n7451), .ZN(n7447) );
  AOI21_X1 U8487 ( .B1(n7796), .B2(n7460), .A(n7459), .ZN(n7458) );
  INV_X1 U8488 ( .A(n8078), .ZN(n7459) );
  INV_X1 U8489 ( .A(n7798), .ZN(n7460) );
  INV_X1 U8490 ( .A(n7796), .ZN(n7461) );
  INV_X1 U8491 ( .A(n8134), .ZN(n7469) );
  NOR2_X1 U8492 ( .A1(n12996), .A2(n9691), .ZN(n7413) );
  INV_X1 U8493 ( .A(n9108), .ZN(n7889) );
  NAND2_X1 U8494 ( .A1(n6887), .A2(n6889), .ZN(n6885) );
  NOR2_X1 U8495 ( .A1(n7150), .A2(n14326), .ZN(n7149) );
  AND2_X1 U8496 ( .A1(n14332), .A2(n7152), .ZN(n7151) );
  NAND2_X1 U8497 ( .A1(n7845), .A2(n7844), .ZN(n7843) );
  NAND2_X1 U8498 ( .A1(n7842), .A2(n7841), .ZN(n7840) );
  NOR2_X1 U8499 ( .A1(n6573), .A2(n7780), .ZN(n7779) );
  INV_X1 U8500 ( .A(n8728), .ZN(n7780) );
  AND2_X1 U8501 ( .A1(n8582), .A2(n8581), .ZN(n8594) );
  INV_X1 U8502 ( .A(n7772), .ZN(n7767) );
  INV_X1 U8503 ( .A(n14373), .ZN(n7055) );
  NOR2_X1 U8504 ( .A1(n15007), .A2(n7282), .ZN(n7281) );
  NAND2_X1 U8505 ( .A1(n6917), .A2(n12802), .ZN(n6916) );
  INV_X1 U8506 ( .A(n6922), .ZN(n6917) );
  AND2_X1 U8507 ( .A1(n6922), .A2(n6919), .ZN(n6914) );
  NOR2_X1 U8508 ( .A1(n7602), .A2(n6919), .ZN(n6918) );
  NOR2_X1 U8509 ( .A1(n12847), .A2(n12822), .ZN(n12831) );
  AND2_X1 U8510 ( .A1(n12757), .A2(n12246), .ZN(n12248) );
  NOR2_X1 U8511 ( .A1(n15220), .A2(n15230), .ZN(n7480) );
  NAND2_X1 U8512 ( .A1(n8329), .A2(n11891), .ZN(n8336) );
  INV_X1 U8513 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n10204) );
  AOI21_X1 U8514 ( .B1(n8284), .B2(n8283), .A(n8282), .ZN(n8285) );
  NOR2_X1 U8515 ( .A1(n8280), .A2(SI_18_), .ZN(n8284) );
  AND2_X1 U8516 ( .A1(n15826), .A2(n7146), .ZN(n8007) );
  NAND2_X1 U8517 ( .A1(n6924), .A2(n6564), .ZN(n8279) );
  NAND2_X1 U8518 ( .A1(n15823), .A2(n9933), .ZN(n6930) );
  INV_X1 U8519 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9933) );
  NAND2_X1 U8520 ( .A1(n8240), .A2(n10395), .ZN(n8250) );
  NAND2_X1 U8521 ( .A1(n8226), .A2(n10307), .ZN(n8239) );
  OAI21_X1 U8522 ( .B1(n10052), .B2(n10084), .A(n7320), .ZN(n8054) );
  OAI21_X1 U8523 ( .B1(n12325), .B2(n10076), .A(n6777), .ZN(n8142) );
  NAND2_X1 U8524 ( .A1(n12325), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6777) );
  OAI21_X1 U8525 ( .B1(n8050), .B2(n10890), .A(n7346), .ZN(n8124) );
  NAND2_X1 U8526 ( .A1(n8050), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7346) );
  INV_X1 U8527 ( .A(P2_RD_REG_SCAN_IN), .ZN(n8034) );
  INV_X1 U8528 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8036) );
  INV_X1 U8529 ( .A(n13073), .ZN(n7634) );
  NAND2_X1 U8530 ( .A1(n7402), .A2(n7399), .ZN(n7398) );
  INV_X1 U8531 ( .A(n9870), .ZN(n7402) );
  NOR2_X1 U8532 ( .A1(n12996), .A2(n7400), .ZN(n7399) );
  OR2_X1 U8533 ( .A1(n11091), .A2(n9955), .ZN(n6987) );
  NOR2_X1 U8534 ( .A1(n6575), .A2(n7572), .ZN(n7571) );
  INV_X1 U8535 ( .A(n7581), .ZN(n7572) );
  INV_X1 U8536 ( .A(n10975), .ZN(n7573) );
  INV_X1 U8537 ( .A(n13286), .ZN(n7690) );
  OR2_X1 U8538 ( .A1(n13345), .A2(n13352), .ZN(n8027) );
  NOR2_X1 U8539 ( .A1(n13566), .A2(n9803), .ZN(n9804) );
  OR2_X1 U8540 ( .A1(n13396), .A2(n13406), .ZN(n9673) );
  INV_X1 U8541 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n7393) );
  INV_X1 U8542 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9116) );
  OR2_X1 U8543 ( .A1(n11241), .A2(n10810), .ZN(n9594) );
  NAND2_X1 U8544 ( .A1(n13355), .A2(n9686), .ZN(n7914) );
  NAND2_X1 U8545 ( .A1(n13403), .A2(n13404), .ZN(n13388) );
  AOI21_X1 U8546 ( .B1(n7923), .B2(n7925), .A(n7922), .ZN(n7921) );
  INV_X1 U8547 ( .A(n9663), .ZN(n7922) );
  INV_X1 U8548 ( .A(n9629), .ZN(n6969) );
  OR2_X1 U8549 ( .A1(n11363), .A2(n6727), .ZN(n6857) );
  INV_X1 U8550 ( .A(n6856), .ZN(n6854) );
  AOI21_X1 U8551 ( .B1(n7908), .B2(n7910), .A(n7906), .ZN(n7905) );
  INV_X1 U8552 ( .A(n9610), .ZN(n7906) );
  INV_X1 U8553 ( .A(n9083), .ZN(n7121) );
  AND2_X1 U8554 ( .A1(n9084), .A2(n6755), .ZN(n7894) );
  NOR2_X1 U8555 ( .A1(n9082), .A2(n7123), .ZN(n7122) );
  INV_X1 U8556 ( .A(n9081), .ZN(n7123) );
  NAND2_X1 U8557 ( .A1(n10100), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9042) );
  INV_X1 U8558 ( .A(n9037), .ZN(n7878) );
  NOR2_X1 U8559 ( .A1(n8558), .A2(n10873), .ZN(n8567) );
  AND2_X1 U8560 ( .A1(n8567), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8582) );
  BUF_X1 U8561 ( .A(n11633), .Z(n12649) );
  NAND2_X1 U8562 ( .A1(n6786), .A2(n6785), .ZN(n14068) );
  AOI21_X1 U8563 ( .B1(n6609), .B2(n6788), .A(n6752), .ZN(n6785) );
  NAND2_X1 U8564 ( .A1(n14142), .A2(n14136), .ZN(n7784) );
  AOI21_X1 U8565 ( .B1(n14136), .B2(n7783), .A(n6698), .ZN(n7782) );
  INV_X1 U8566 ( .A(n6623), .ZN(n7783) );
  INV_X1 U8567 ( .A(n14174), .ZN(n7155) );
  INV_X1 U8568 ( .A(n8672), .ZN(n7553) );
  NOR2_X1 U8569 ( .A1(n8672), .A2(n7555), .ZN(n7552) );
  NAND2_X1 U8570 ( .A1(n9013), .A2(n7111), .ZN(n7110) );
  INV_X1 U8571 ( .A(n8607), .ZN(n7111) );
  OAI21_X1 U8572 ( .B1(n11726), .B2(n7762), .A(n8710), .ZN(n7761) );
  INV_X1 U8573 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U8574 ( .A1(n6824), .A2(n6820), .ZN(n8021) );
  INV_X1 U8575 ( .A(n7508), .ZN(n6824) );
  AND2_X1 U8576 ( .A1(n14570), .A2(n6821), .ZN(n6820) );
  NOR2_X1 U8577 ( .A1(n11958), .A2(n6822), .ZN(n6821) );
  OR2_X1 U8578 ( .A1(n14575), .A2(n11645), .ZN(n8707) );
  NAND2_X1 U8579 ( .A1(n7170), .A2(n6639), .ZN(n8511) );
  NAND2_X1 U8580 ( .A1(n11696), .A2(n7511), .ZN(n7510) );
  NAND2_X1 U8581 ( .A1(n7169), .A2(n8173), .ZN(n8705) );
  AND2_X1 U8582 ( .A1(n13950), .A2(n8172), .ZN(n7169) );
  NAND2_X1 U8583 ( .A1(n14519), .A2(n11388), .ZN(n14371) );
  NAND2_X1 U8584 ( .A1(n14318), .A2(n7514), .ZN(n14304) );
  OR2_X1 U8585 ( .A1(n15659), .A2(n11283), .ZN(n10034) );
  NAND2_X1 U8586 ( .A1(n7775), .A2(n7349), .ZN(n8384) );
  INV_X1 U8587 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8265) );
  INV_X1 U8588 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8102) );
  AND2_X1 U8589 ( .A1(n12564), .A2(n12563), .ZN(n12566) );
  AND2_X1 U8590 ( .A1(n12126), .A2(n12125), .ZN(n12183) );
  NOR2_X1 U8591 ( .A1(n12276), .A2(n12275), .ZN(n6783) );
  OR2_X1 U8592 ( .A1(n10271), .A2(n10272), .ZN(n7069) );
  INV_X1 U8593 ( .A(n14885), .ZN(n6861) );
  INV_X1 U8594 ( .A(n6867), .ZN(n6863) );
  NAND2_X1 U8595 ( .A1(n14902), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7490) );
  NOR2_X1 U8596 ( .A1(n15807), .A2(n6905), .ZN(n6898) );
  NAND2_X1 U8597 ( .A1(n7480), .A2(n15210), .ZN(n7479) );
  AND2_X1 U8598 ( .A1(n15220), .A2(n14769), .ZN(n12440) );
  NOR2_X1 U8599 ( .A1(n15220), .A2(n14769), .ZN(n12438) );
  NAND2_X1 U8600 ( .A1(n15029), .A2(n7955), .ZN(n7954) );
  INV_X1 U8601 ( .A(n12339), .ZN(n7955) );
  INV_X1 U8602 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n12275) );
  NAND2_X1 U8603 ( .A1(n7284), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n12276) );
  INV_X1 U8604 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n15981) );
  INV_X1 U8605 ( .A(n15181), .ZN(n12754) );
  NAND2_X1 U8606 ( .A1(n12060), .A2(n11547), .ZN(n6942) );
  INV_X1 U8607 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n11198) );
  NAND2_X1 U8608 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n10921) );
  INV_X1 U8609 ( .A(n11126), .ZN(n7298) );
  INV_X1 U8610 ( .A(n7215), .ZN(n6935) );
  OAI21_X1 U8611 ( .B1(n7217), .B2(P1_IR_REG_30__SCAN_IN), .A(n7216), .ZN(
        n7215) );
  NAND2_X1 U8612 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n7216) );
  NOR2_X1 U8613 ( .A1(n10254), .A2(n10221), .ZN(n7217) );
  INV_X1 U8614 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7967) );
  OAI21_X1 U8615 ( .B1(n8349), .B2(n8348), .A(n8351), .ZN(n8356) );
  NAND2_X1 U8616 ( .A1(n8328), .A2(n8327), .ZN(n8335) );
  NAND2_X1 U8617 ( .A1(n8325), .A2(n8324), .ZN(n8328) );
  NAND2_X1 U8618 ( .A1(n6926), .A2(n6925), .ZN(n8286) );
  AOI21_X1 U8619 ( .B1(n6564), .B2(n7450), .A(n8278), .ZN(n6925) );
  NOR2_X1 U8620 ( .A1(n10206), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n10212) );
  NAND2_X1 U8621 ( .A1(n8286), .A2(n8285), .ZN(n8301) );
  NAND2_X1 U8622 ( .A1(n8008), .A2(n8007), .ZN(n10330) );
  INV_X1 U8623 ( .A(n8239), .ZN(n7451) );
  OR2_X1 U8624 ( .A1(n8213), .A2(n8220), .ZN(n6838) );
  AND2_X1 U8625 ( .A1(n8213), .A2(n8220), .ZN(n6837) );
  NAND2_X1 U8626 ( .A1(n8068), .A2(n10166), .ZN(n8071) );
  NAND2_X1 U8627 ( .A1(n6929), .A2(SI_12_), .ZN(n8073) );
  INV_X1 U8628 ( .A(n8072), .ZN(n6929) );
  OR2_X1 U8629 ( .A1(n10073), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n10543) );
  NAND2_X1 U8630 ( .A1(n8124), .A2(SI_3_), .ZN(n8134) );
  NAND2_X1 U8631 ( .A1(n8050), .A2(n10053), .ZN(n7280) );
  NAND2_X1 U8632 ( .A1(n11090), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n7195) );
  NAND2_X1 U8633 ( .A1(n14794), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10125) );
  INV_X1 U8634 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10127) );
  AND2_X1 U8635 ( .A1(n7192), .A2(n7190), .ZN(n10132) );
  OR2_X1 U8636 ( .A1(n10134), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n7646) );
  OAI21_X1 U8637 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n10614), .A(n10613), .ZN(
        n10621) );
  NAND2_X1 U8638 ( .A1(n10943), .A2(n10942), .ZN(n11304) );
  AND2_X1 U8639 ( .A1(n15425), .A2(n15424), .ZN(n15439) );
  OR2_X1 U8640 ( .A1(n15423), .A2(n15422), .ZN(n15425) );
  NAND2_X1 U8641 ( .A1(n7643), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n7640) );
  NOR2_X1 U8642 ( .A1(n7030), .A2(n6681), .ZN(n7028) );
  NOR2_X1 U8643 ( .A1(n6618), .A2(n7031), .ZN(n7030) );
  NAND2_X1 U8644 ( .A1(n11046), .A2(n7244), .ZN(n10519) );
  INV_X1 U8645 ( .A(n13121), .ZN(n7244) );
  AND2_X1 U8646 ( .A1(n12948), .A2(n12949), .ZN(n7246) );
  OR2_X1 U8647 ( .A1(n13038), .A2(n13406), .ZN(n12948) );
  AND2_X1 U8648 ( .A1(n6712), .A2(n11945), .ZN(n7052) );
  NAND2_X1 U8649 ( .A1(n6635), .A2(n9111), .ZN(n9238) );
  AND4_X1 U8650 ( .A1(n9338), .A2(n9337), .A3(n9336), .A4(n9335), .ZN(n13059)
         );
  OR2_X1 U8651 ( .A1(n9211), .A2(n9168), .ZN(n9170) );
  NOR2_X1 U8652 ( .A1(n11092), .A2(n15789), .ZN(n11091) );
  XNOR2_X1 U8653 ( .A(n10106), .B(P3_REG1_REG_2__SCAN_IN), .ZN(n10746) );
  INV_X1 U8654 ( .A(n7265), .ZN(n10744) );
  INV_X1 U8655 ( .A(n6987), .ZN(n10745) );
  OR2_X1 U8656 ( .A1(n13724), .A2(n10770), .ZN(n6984) );
  NAND2_X1 U8657 ( .A1(n13724), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n6983) );
  NAND2_X1 U8658 ( .A1(n7682), .A2(n10978), .ZN(n10732) );
  NAND2_X1 U8659 ( .A1(n7682), .A2(n6611), .ZN(n10980) );
  NAND2_X1 U8660 ( .A1(n9958), .A2(n10779), .ZN(n6998) );
  AOI21_X1 U8661 ( .B1(n10778), .B2(n6999), .A(n9959), .ZN(n10948) );
  NAND2_X1 U8662 ( .A1(n7670), .A2(n10115), .ZN(n6999) );
  NAND2_X1 U8663 ( .A1(n7693), .A2(n11072), .ZN(n10956) );
  NAND2_X1 U8664 ( .A1(n7693), .A2(n6750), .ZN(n11074) );
  AOI21_X1 U8665 ( .B1(n10772), .B2(n10776), .A(n9977), .ZN(n10970) );
  AND2_X1 U8666 ( .A1(n6990), .A2(n6989), .ZN(n13132) );
  AND2_X1 U8667 ( .A1(n9103), .A2(n9102), .ZN(n7631) );
  NAND2_X1 U8668 ( .A1(n7272), .A2(n13196), .ZN(n13173) );
  NOR2_X1 U8669 ( .A1(n7589), .A2(n13171), .ZN(n7588) );
  NAND2_X1 U8670 ( .A1(n13224), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7705) );
  NAND2_X1 U8671 ( .A1(n6992), .A2(n6993), .ZN(n13223) );
  OR2_X1 U8672 ( .A1(n13221), .A2(n13256), .ZN(n7677) );
  NAND2_X1 U8673 ( .A1(n7687), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n13288) );
  NAND2_X1 U8674 ( .A1(n7699), .A2(n7702), .ZN(n7698) );
  NAND3_X1 U8675 ( .A1(n7701), .A2(n13292), .A3(n6612), .ZN(n7700) );
  INV_X1 U8676 ( .A(n12996), .ZN(n9754) );
  NAND2_X1 U8677 ( .A1(n7310), .A2(n7722), .ZN(n9862) );
  NOR2_X1 U8678 ( .A1(n13350), .A2(n9804), .ZN(n9806) );
  OR2_X1 U8679 ( .A1(n9529), .A2(n9125), .ZN(n9542) );
  NAND2_X1 U8680 ( .A1(n13356), .A2(n13355), .ZN(n13354) );
  OR2_X1 U8681 ( .A1(n9509), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9529) );
  OR2_X1 U8682 ( .A1(n9486), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9497) );
  INV_X1 U8683 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n7395) );
  OR2_X1 U8684 ( .A1(n9472), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9486) );
  NAND2_X1 U8685 ( .A1(n9122), .A2(n7396), .ZN(n9460) );
  NAND2_X1 U8686 ( .A1(n9394), .A2(n9120), .ZN(n9417) );
  NAND2_X1 U8687 ( .A1(n9117), .A2(n6606), .ZN(n9372) );
  NAND2_X1 U8688 ( .A1(n7389), .A2(n9115), .ZN(n9343) );
  INV_X1 U8689 ( .A(n9332), .ZN(n7389) );
  NAND2_X1 U8690 ( .A1(n7391), .A2(n7390), .ZN(n9332) );
  INV_X1 U8691 ( .A(n7391), .ZN(n9314) );
  NAND2_X1 U8692 ( .A1(n9114), .A2(n9113), .ZN(n9299) );
  INV_X1 U8693 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9113) );
  INV_X1 U8694 ( .A(n9281), .ZN(n9114) );
  INV_X1 U8695 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n9112) );
  OR2_X1 U8696 ( .A1(n9263), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9281) );
  NAND2_X1 U8697 ( .A1(n9111), .A2(n9110), .ZN(n9226) );
  NAND2_X1 U8698 ( .A1(n10811), .A2(n9109), .ZN(n9212) );
  INV_X1 U8699 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n9109) );
  NAND2_X1 U8700 ( .A1(n11047), .A2(n10519), .ZN(n10761) );
  INV_X1 U8701 ( .A(n9585), .ZN(n10760) );
  NAND2_X1 U8702 ( .A1(n10761), .A2(n10760), .ZN(n10804) );
  NAND2_X1 U8703 ( .A1(n11056), .A2(n11048), .ZN(n11047) );
  NAND2_X1 U8704 ( .A1(n7706), .A2(n9708), .ZN(n11056) );
  OR2_X1 U8705 ( .A1(n10082), .A2(n9842), .ZN(n9884) );
  AND2_X1 U8706 ( .A1(n9847), .A2(n9852), .ZN(n9886) );
  NOR2_X1 U8707 ( .A1(n13336), .A2(n13335), .ZN(n13619) );
  NAND2_X1 U8708 ( .A1(n9552), .A2(n9551), .ZN(n9894) );
  AOI21_X1 U8709 ( .B1(n6963), .B2(n9676), .A(n6962), .ZN(n6961) );
  INV_X1 U8710 ( .A(n9680), .ZN(n6962) );
  NAND2_X1 U8711 ( .A1(n13388), .A2(n9800), .ZN(n7712) );
  NOR2_X1 U8712 ( .A1(n7716), .A2(n7714), .ZN(n7713) );
  INV_X1 U8713 ( .A(n13458), .ZN(n7714) );
  AND2_X1 U8714 ( .A1(n7715), .A2(n9793), .ZN(n13459) );
  INV_X1 U8715 ( .A(n15770), .ZN(n13598) );
  OR2_X1 U8716 ( .A1(n12105), .A2(n6889), .ZN(n6886) );
  INV_X1 U8717 ( .A(n9632), .ZN(n13511) );
  AND3_X1 U8718 ( .A1(n9376), .A2(n9375), .A3(n9374), .ZN(n13536) );
  NAND2_X1 U8719 ( .A1(n7740), .A2(n9787), .ZN(n13531) );
  NAND2_X1 U8720 ( .A1(n7934), .A2(n9637), .ZN(n13526) );
  NAND2_X1 U8721 ( .A1(n7936), .A2(n7935), .ZN(n7934) );
  INV_X1 U8722 ( .A(n13545), .ZN(n7936) );
  NAND2_X1 U8723 ( .A1(n12105), .A2(n12103), .ZN(n9786) );
  NAND2_X1 U8724 ( .A1(n7895), .A2(n7896), .ZN(n12104) );
  AOI21_X1 U8725 ( .B1(n6571), .B2(n7903), .A(n7897), .ZN(n7896) );
  INV_X1 U8726 ( .A(n9624), .ZN(n7897) );
  NAND2_X1 U8727 ( .A1(n11372), .A2(n6566), .ZN(n11772) );
  NOR2_X1 U8728 ( .A1(n7126), .A2(n9080), .ZN(n7125) );
  INV_X1 U8729 ( .A(n9079), .ZN(n7126) );
  CLKBUF_X1 U8730 ( .A(n9736), .Z(n9737) );
  XNOR2_X1 U8731 ( .A(n9730), .B(n16100), .ZN(n10500) );
  INV_X1 U8732 ( .A(n7884), .ZN(n7883) );
  AND2_X1 U8733 ( .A1(n9075), .A2(n9074), .ZN(n9465) );
  INV_X1 U8734 ( .A(n9571), .ZN(n7637) );
  AOI21_X1 U8735 ( .B1(n7874), .B2(n7876), .A(n7871), .ZN(n7870) );
  INV_X1 U8736 ( .A(n9058), .ZN(n7871) );
  NAND2_X1 U8737 ( .A1(n9322), .A2(n9051), .ZN(n7873) );
  INV_X1 U8738 ( .A(n7275), .ZN(n9276) );
  AND2_X1 U8739 ( .A1(n9044), .A2(n9043), .ZN(n9252) );
  AOI21_X1 U8740 ( .B1(n7115), .B2(n7117), .A(n6687), .ZN(n7114) );
  NAND2_X1 U8741 ( .A1(n7309), .A2(n9247), .ZN(n9257) );
  INV_X1 U8742 ( .A(n7309), .ZN(n9246) );
  INV_X1 U8743 ( .A(n13950), .ZN(n11388) );
  NAND2_X1 U8744 ( .A1(n7367), .A2(n13733), .ZN(n7366) );
  NAND2_X1 U8745 ( .A1(n7368), .A2(n7373), .ZN(n7365) );
  INV_X1 U8746 ( .A(n7370), .ZN(n7367) );
  OR2_X1 U8747 ( .A1(n7379), .A2(n13890), .ZN(n7376) );
  NOR2_X1 U8748 ( .A1(n7727), .A2(n7726), .ZN(n7725) );
  INV_X1 U8749 ( .A(n13851), .ZN(n7727) );
  INV_X1 U8750 ( .A(n12648), .ZN(n7726) );
  NAND2_X1 U8751 ( .A1(n10408), .A2(n7755), .ZN(n10853) );
  INV_X1 U8752 ( .A(n10032), .ZN(n10030) );
  NAND2_X1 U8753 ( .A1(n7744), .A2(n7743), .ZN(n12029) );
  OR2_X1 U8754 ( .A1(n8619), .A2(n13854), .ZN(n8630) );
  NAND2_X1 U8755 ( .A1(n8628), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8639) );
  INV_X1 U8756 ( .A(n8630), .ZN(n8628) );
  AOI21_X1 U8757 ( .B1(n7359), .B2(n7361), .A(n6686), .ZN(n7358) );
  INV_X1 U8758 ( .A(n7743), .ZN(n7359) );
  INV_X1 U8759 ( .A(n7361), .ZN(n7360) );
  AOI21_X1 U8760 ( .B1(n7386), .B2(n7384), .A(n7383), .ZN(n7382) );
  INV_X1 U8761 ( .A(n12638), .ZN(n7383) );
  INV_X1 U8762 ( .A(n12632), .ZN(n7384) );
  CLKBUF_X3 U8763 ( .A(n10022), .Z(n12612) );
  NOR2_X1 U8764 ( .A1(n9019), .A2(n7167), .ZN(n7166) );
  AND2_X1 U8765 ( .A1(n8998), .A2(n8958), .ZN(n9021) );
  AND2_X1 U8766 ( .A1(n8617), .A2(n8616), .ZN(n13893) );
  AND3_X1 U8767 ( .A1(n8605), .A2(n8604), .A3(n8603), .ZN(n12639) );
  OR2_X1 U8768 ( .A1(n10872), .A2(n10871), .ZN(n10869) );
  OR2_X1 U8769 ( .A1(n14061), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n14077) );
  NOR2_X1 U8770 ( .A1(n8767), .A2(n7519), .ZN(n14093) );
  NOR2_X1 U8771 ( .A1(n7517), .A2(n14097), .ZN(n7516) );
  NAND2_X1 U8772 ( .A1(n7518), .A2(n14414), .ZN(n7517) );
  INV_X1 U8773 ( .A(n7519), .ZN(n7518) );
  AOI21_X1 U8774 ( .B1(n7162), .B2(n9900), .A(n9899), .ZN(n7157) );
  AND2_X1 U8775 ( .A1(n13797), .A2(n13930), .ZN(n9899) );
  AND2_X1 U8776 ( .A1(n8736), .A2(n8735), .ZN(n14101) );
  NAND2_X1 U8777 ( .A1(n10427), .A2(n8745), .ZN(n13915) );
  AND2_X1 U8778 ( .A1(n9911), .A2(n15662), .ZN(n9912) );
  OR2_X1 U8779 ( .A1(n8767), .A2(n13797), .ZN(n9903) );
  NOR3_X1 U8780 ( .A1(n14216), .A2(n6828), .A3(n6569), .ZN(n14128) );
  NAND2_X1 U8781 ( .A1(n14530), .A2(n14534), .ZN(n6828) );
  NOR3_X1 U8782 ( .A1(n14216), .A2(n6569), .A3(n14146), .ZN(n14149) );
  NAND2_X1 U8783 ( .A1(n8637), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8647) );
  INV_X1 U8784 ( .A(n8639), .ZN(n8637) );
  XNOR2_X1 U8785 ( .A(n14182), .B(n13731), .ZN(n14175) );
  OR2_X1 U8786 ( .A1(n14176), .A2(n14175), .ZN(n14178) );
  NAND2_X1 U8787 ( .A1(n7534), .A2(n7532), .ZN(n7531) );
  NOR2_X1 U8788 ( .A1(n14213), .A2(n7533), .ZN(n7532) );
  INV_X1 U8789 ( .A(n8627), .ZN(n7533) );
  NOR2_X1 U8790 ( .A1(n7018), .A2(n6572), .ZN(n7017) );
  NAND2_X1 U8791 ( .A1(n7019), .A2(n14191), .ZN(n7018) );
  NAND2_X1 U8792 ( .A1(n7759), .A2(n14222), .ZN(n14223) );
  OAI21_X1 U8793 ( .B1(n14241), .B2(n8721), .A(n8720), .ZN(n14225) );
  NOR2_X1 U8794 ( .A1(n14456), .A2(n14451), .ZN(n6827) );
  AOI21_X1 U8795 ( .B1(n7524), .B2(n7526), .A(n6682), .ZN(n7177) );
  AND3_X1 U8796 ( .A1(n14318), .A2(n7512), .A3(n14555), .ZN(n14273) );
  NAND2_X1 U8797 ( .A1(n7044), .A2(n8718), .ZN(n14254) );
  OAI21_X1 U8798 ( .B1(n6578), .B2(n7096), .A(n7095), .ZN(n14327) );
  AND2_X1 U8799 ( .A1(n7537), .A2(n8564), .ZN(n7095) );
  NAND2_X1 U8800 ( .A1(n8539), .A2(n7540), .ZN(n7096) );
  NAND2_X1 U8801 ( .A1(n14318), .A2(n14325), .ZN(n14319) );
  NAND2_X1 U8802 ( .A1(n8708), .A2(n11726), .ZN(n11733) );
  INV_X1 U8803 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U8804 ( .A1(n8528), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8541) );
  AND2_X1 U8805 ( .A1(n7764), .A2(n14363), .ZN(n7763) );
  NAND2_X1 U8806 ( .A1(n7766), .A2(n7768), .ZN(n7764) );
  NAND2_X1 U8807 ( .A1(n6826), .A2(n14504), .ZN(n6825) );
  NOR2_X1 U8808 ( .A1(n11986), .A2(n11683), .ZN(n11987) );
  NOR2_X1 U8809 ( .A1(n11986), .A2(n7510), .ZN(n14396) );
  NAND2_X1 U8810 ( .A1(n8702), .A2(n7772), .ZN(n7771) );
  NAND2_X1 U8811 ( .A1(n8497), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8517) );
  NAND2_X1 U8812 ( .A1(n11655), .A2(n11656), .ZN(n8702) );
  NAND2_X1 U8813 ( .A1(n10790), .A2(n10788), .ZN(n10789) );
  NAND2_X1 U8814 ( .A1(n11715), .A2(n11625), .ZN(n11957) );
  AND3_X1 U8815 ( .A1(n6819), .A2(n15707), .A3(n15717), .ZN(n11715) );
  INV_X1 U8816 ( .A(n10577), .ZN(n11706) );
  NAND2_X1 U8817 ( .A1(n8779), .A2(n15660), .ZN(n11970) );
  NAND2_X1 U8818 ( .A1(n6819), .A2(n15707), .ZN(n11716) );
  XNOR2_X1 U8819 ( .A(n13956), .B(n10584), .ZN(n10577) );
  NAND2_X1 U8820 ( .A1(n10575), .A2(n10577), .ZN(n10576) );
  AND2_X1 U8821 ( .A1(n8951), .A2(n8782), .ZN(n9924) );
  INV_X1 U8822 ( .A(n14338), .ZN(n14470) );
  INV_X1 U8823 ( .A(n15740), .ZN(n14484) );
  AND3_X1 U8824 ( .A1(n10005), .A2(P2_STATE_REG_SCAN_IN), .A3(n10007), .ZN(
        n11617) );
  AND3_X1 U8825 ( .A1(n7277), .A2(n8099), .A3(n8095), .ZN(n7174) );
  NAND2_X1 U8826 ( .A1(n8384), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8385) );
  AND2_X1 U8827 ( .A1(n7749), .A2(n7748), .ZN(n7747) );
  INV_X1 U8828 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7748) );
  OR2_X1 U8829 ( .A1(n8168), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8170) );
  OR2_X1 U8830 ( .A1(n8170), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8177) );
  INV_X1 U8831 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8129) );
  NAND2_X1 U8832 ( .A1(n8115), .A2(n6808), .ZN(n10433) );
  AOI22_X1 U8833 ( .A1(n6690), .A2(P2_IR_REG_0__SCAN_IN), .B1(n6810), .B2(
        n6809), .ZN(n6808) );
  INV_X1 U8834 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6810) );
  NAND2_X1 U8835 ( .A1(n8050), .A2(SI_0_), .ZN(n9159) );
  NAND2_X1 U8836 ( .A1(n14744), .A2(n12578), .ZN(n7142) );
  INV_X1 U8837 ( .A(n7972), .ZN(n7971) );
  OAI21_X1 U8838 ( .B1(n11433), .B2(n7973), .A(n11853), .ZN(n7972) );
  INV_X1 U8839 ( .A(n11438), .ZN(n7973) );
  INV_X1 U8840 ( .A(n12315), .ZN(n12316) );
  NAND2_X1 U8841 ( .A1(n7977), .A2(n6843), .ZN(n6842) );
  AND2_X1 U8842 ( .A1(n7975), .A2(n14665), .ZN(n7974) );
  INV_X1 U8843 ( .A(n14608), .ZN(n6843) );
  INV_X1 U8844 ( .A(n7977), .ZN(n6844) );
  AOI22_X1 U8845 ( .A1(n10380), .A2(P1_IR_REG_0__SCAN_IN), .B1(n6937), .B2(
        n12552), .ZN(n10377) );
  INV_X1 U8846 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14705) );
  AND2_X1 U8847 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n12077) );
  INV_X1 U8848 ( .A(n12330), .ZN(n12329) );
  NAND2_X1 U8849 ( .A1(n7986), .A2(n7984), .ZN(n14606) );
  AOI21_X1 U8850 ( .B1(n7987), .B2(n7989), .A(n7985), .ZN(n7984) );
  INV_X1 U8851 ( .A(n14724), .ZN(n7985) );
  NAND2_X1 U8852 ( .A1(n10910), .A2(n14792), .ZN(n7129) );
  NAND2_X1 U8853 ( .A1(n14792), .A2(n6554), .ZN(n10670) );
  INV_X1 U8854 ( .A(n6783), .ZN(n12286) );
  NAND2_X1 U8855 ( .A1(n14598), .A2(n7994), .ZN(n7137) );
  AOI21_X1 U8856 ( .B1(n7994), .B2(n7996), .A(n6671), .ZN(n7992) );
  INV_X1 U8857 ( .A(n14770), .ZN(n14939) );
  NAND2_X1 U8858 ( .A1(n14598), .A2(n12489), .ZN(n14673) );
  INV_X1 U8859 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14794) );
  OR2_X1 U8860 ( .A1(n10247), .A2(n10246), .ZN(n10273) );
  NAND2_X1 U8861 ( .A1(n7066), .A2(n7069), .ZN(n10323) );
  NAND2_X1 U8862 ( .A1(n7061), .A2(n10321), .ZN(n10320) );
  NAND2_X1 U8863 ( .A1(n7066), .A2(n7067), .ZN(n7061) );
  AND2_X1 U8864 ( .A1(n11440), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7301) );
  NOR2_X1 U8865 ( .A1(n7068), .A2(n10322), .ZN(n7067) );
  INV_X1 U8866 ( .A(n7069), .ZN(n7068) );
  OR2_X1 U8867 ( .A1(n7070), .A2(n10247), .ZN(n7066) );
  NAND2_X1 U8868 ( .A1(n7072), .A2(n7071), .ZN(n7070) );
  INV_X1 U8869 ( .A(n10246), .ZN(n7071) );
  INV_X1 U8870 ( .A(n10271), .ZN(n7072) );
  INV_X1 U8871 ( .A(n10292), .ZN(n7064) );
  OR2_X1 U8872 ( .A1(n14842), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7501) );
  NAND2_X1 U8873 ( .A1(n11118), .A2(n7262), .ZN(n11119) );
  OR2_X1 U8874 ( .A1(n12008), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7262) );
  OR2_X1 U8875 ( .A1(n14868), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7503) );
  NAND2_X1 U8876 ( .A1(n15479), .A2(n6657), .ZN(n14890) );
  INV_X1 U8877 ( .A(n14877), .ZN(n7084) );
  NAND2_X1 U8878 ( .A1(n6869), .A2(n12258), .ZN(n6868) );
  INV_X1 U8879 ( .A(n14871), .ZN(n6866) );
  INV_X1 U8880 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n6905) );
  XNOR2_X1 U8881 ( .A(n7085), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n15816) );
  OAI21_X1 U8882 ( .B1(n15810), .B2(n7086), .A(n15811), .ZN(n7085) );
  INV_X1 U8883 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n7086) );
  OAI211_X1 U8884 ( .C1(n6903), .C2(n6902), .A(n6901), .B(n6900), .ZN(n15818)
         );
  NAND2_X1 U8885 ( .A1(n6899), .A2(n6898), .ZN(n6900) );
  OR2_X1 U8886 ( .A1(n15805), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6902) );
  NAND2_X1 U8887 ( .A1(n15805), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6901) );
  NAND2_X1 U8888 ( .A1(n12857), .A2(n12856), .ZN(n14916) );
  NAND2_X1 U8889 ( .A1(n12813), .A2(n12812), .ZN(n14923) );
  OR2_X1 U8890 ( .A1(n14974), .A2(n7479), .ZN(n14922) );
  NOR3_X1 U8891 ( .A1(n14974), .A2(n14923), .A3(n7479), .ZN(n14924) );
  NAND2_X1 U8892 ( .A1(n12409), .A2(n12408), .ZN(n12819) );
  NOR2_X1 U8893 ( .A1(n12400), .A2(n12399), .ZN(n12456) );
  NAND2_X1 U8894 ( .A1(n14972), .A2(n6624), .ZN(n7805) );
  NAND2_X1 U8895 ( .A1(n7235), .A2(n7237), .ZN(n7233) );
  AND2_X1 U8896 ( .A1(n12678), .A2(n14772), .ZN(n12435) );
  NOR2_X1 U8897 ( .A1(n7476), .A2(n12678), .ZN(n7475) );
  OR2_X2 U8898 ( .A1(n14994), .A2(n15236), .ZN(n14974) );
  AND2_X1 U8899 ( .A1(n12375), .A2(n12354), .ZN(n14995) );
  INV_X1 U8900 ( .A(n15007), .ZN(n14966) );
  NOR3_X1 U8901 ( .A1(n15054), .A2(n15259), .A3(n15267), .ZN(n15025) );
  NOR2_X1 U8902 ( .A1(n15054), .A2(n7476), .ZN(n15010) );
  AND2_X1 U8903 ( .A1(n15142), .A2(n6704), .ZN(n15076) );
  NAND2_X1 U8904 ( .A1(n15142), .A2(n7481), .ZN(n15088) );
  AND2_X1 U8905 ( .A1(n7962), .A2(n12785), .ZN(n15069) );
  AOI21_X1 U8906 ( .B1(n6581), .B2(n7232), .A(n7227), .ZN(n7226) );
  INV_X1 U8907 ( .A(n7808), .ZN(n7227) );
  INV_X1 U8908 ( .A(n7331), .ZN(n6940) );
  INV_X1 U8909 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n12253) );
  NAND2_X1 U8910 ( .A1(n7333), .A2(n6579), .ZN(n15166) );
  AND2_X1 U8911 ( .A1(n12169), .A2(n15325), .ZN(n12170) );
  NAND2_X1 U8912 ( .A1(n12152), .A2(n12151), .ZN(n12249) );
  OR2_X1 U8913 ( .A1(n15331), .A2(n12214), .ZN(n12075) );
  INV_X1 U8914 ( .A(n12882), .ZN(n11549) );
  NAND2_X1 U8915 ( .A1(n12066), .A2(n7489), .ZN(n15501) );
  OR2_X1 U8916 ( .A1(n12060), .A2(n12063), .ZN(n12061) );
  AND2_X1 U8917 ( .A1(n12066), .A2(n15592), .ZN(n15502) );
  INV_X1 U8918 ( .A(n12878), .ZN(n15508) );
  OR2_X1 U8919 ( .A1(n11337), .A2(n12708), .ZN(n11210) );
  NAND2_X1 U8920 ( .A1(n7471), .A2(n7470), .ZN(n11337) );
  INV_X1 U8921 ( .A(n11351), .ZN(n7471) );
  NOR2_X1 U8922 ( .A1(n11172), .A2(n12691), .ZN(n11349) );
  INV_X1 U8923 ( .A(n15180), .ZN(n15128) );
  AND2_X1 U8924 ( .A1(n10358), .A2(n10357), .ZN(n12684) );
  AND2_X1 U8925 ( .A1(n15382), .A2(n12328), .ZN(n15267) );
  AND2_X1 U8926 ( .A1(n15048), .A2(n12324), .ZN(n15036) );
  NAND2_X1 U8927 ( .A1(n15142), .A2(n15137), .ZN(n15112) );
  XNOR2_X1 U8928 ( .A(n9939), .B(P1_IR_REG_23__SCAN_IN), .ZN(n10333) );
  OAI21_X1 U8929 ( .B1(n10202), .B2(n9938), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9939) );
  XNOR2_X1 U8930 ( .A(n8366), .B(n8367), .ZN(n12811) );
  XNOR2_X1 U8931 ( .A(n8360), .B(n8359), .ZN(n14586) );
  INV_X1 U8932 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n10253) );
  XNOR2_X1 U8933 ( .A(n8356), .B(n8355), .ZN(n12461) );
  XNOR2_X1 U8934 ( .A(n8321), .B(n8324), .ZN(n12360) );
  NAND2_X1 U8935 ( .A1(n7465), .A2(n8300), .ZN(n8314) );
  NAND2_X1 U8936 ( .A1(n8286), .A2(n6577), .ZN(n7465) );
  OR2_X1 U8937 ( .A1(n10198), .A2(n10197), .ZN(n10572) );
  NAND2_X1 U8938 ( .A1(n7798), .A2(n7795), .ZN(n8202) );
  OR2_X1 U8939 ( .A1(n8190), .A2(n7801), .ZN(n7795) );
  OAI21_X1 U8940 ( .B1(n10572), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10311) );
  NAND2_X1 U8941 ( .A1(n7316), .A2(n6850), .ZN(n8185) );
  NAND2_X1 U8942 ( .A1(n7318), .A2(n8167), .ZN(n6850) );
  NAND2_X1 U8943 ( .A1(n8167), .A2(n8061), .ZN(n7317) );
  AND2_X1 U8944 ( .A1(n9931), .A2(n15823), .ZN(n6908) );
  OAI21_X1 U8945 ( .B1(n9159), .B2(n9028), .A(n10048), .ZN(n8106) );
  NAND2_X1 U8946 ( .A1(n7649), .A2(n10131), .ZN(n7648) );
  NAND2_X1 U8947 ( .A1(n7651), .A2(n10603), .ZN(n10608) );
  NOR2_X1 U8948 ( .A1(n15386), .A2(n7185), .ZN(n7184) );
  INV_X1 U8949 ( .A(n15385), .ZN(n7182) );
  AND2_X1 U8950 ( .A1(n10610), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7181) );
  NAND2_X1 U8951 ( .A1(n10619), .A2(n10618), .ZN(n10938) );
  NAND2_X1 U8952 ( .A1(n15387), .A2(n15388), .ZN(n10619) );
  NAND2_X1 U8953 ( .A1(n10935), .A2(n14026), .ZN(n7205) );
  NAND2_X1 U8954 ( .A1(n7029), .A2(n6618), .ZN(n12994) );
  NAND2_X1 U8955 ( .A1(n9485), .A2(n9484), .ZN(n13580) );
  NAND2_X1 U8956 ( .A1(n7012), .A2(n12938), .ZN(n7011) );
  OAI21_X1 U8957 ( .B1(n7035), .B2(n7028), .A(n7024), .ZN(n7023) );
  NAND2_X1 U8958 ( .A1(n7025), .A2(n7028), .ZN(n7024) );
  OR2_X1 U8959 ( .A1(n6636), .A2(n7035), .ZN(n7025) );
  NAND2_X1 U8960 ( .A1(n7028), .A2(n12997), .ZN(n7027) );
  AND2_X1 U8961 ( .A1(n6636), .A2(n7035), .ZN(n7026) );
  NAND2_X1 U8962 ( .A1(n10529), .A2(n10527), .ZN(n10590) );
  NAND2_X1 U8963 ( .A1(n11946), .A2(n11945), .ZN(n7053) );
  NAND2_X1 U8964 ( .A1(n11271), .A2(n11270), .ZN(n11272) );
  NAND2_X1 U8965 ( .A1(n12933), .A2(n12932), .ZN(n13028) );
  AND4_X1 U8966 ( .A1(n9348), .A2(n9347), .A3(n9346), .A4(n9345), .ZN(n13534)
         );
  NOR2_X1 U8967 ( .A1(n11606), .A2(n7620), .ZN(n7619) );
  AND2_X1 U8968 ( .A1(n11592), .A2(n6710), .ZN(n7261) );
  INV_X1 U8969 ( .A(n11747), .ZN(n7620) );
  CLKBUF_X1 U8970 ( .A(n10595), .Z(n10632) );
  NAND2_X1 U8971 ( .A1(n13026), .A2(n12935), .ZN(n13074) );
  OAI21_X1 U8972 ( .B1(n6774), .B2(n7015), .A(n6570), .ZN(n13075) );
  NAND2_X1 U8973 ( .A1(n10509), .A2(n10508), .ZN(n13095) );
  INV_X1 U8974 ( .A(n7036), .ZN(n7033) );
  AND2_X1 U8975 ( .A1(n9560), .A2(n9559), .ZN(n12999) );
  NAND2_X1 U8976 ( .A1(n9503), .A2(n9502), .ZN(n13374) );
  NAND2_X1 U8977 ( .A1(n9439), .A2(n9438), .ZN(n13108) );
  INV_X1 U8978 ( .A(n13534), .ZN(n12106) );
  INV_X1 U8979 ( .A(n13059), .ZN(n13550) );
  NOR2_X1 U8980 ( .A1(n10501), .A2(n13702), .ZN(n13115) );
  OAI211_X1 U8981 ( .C1(n9175), .C2(n10371), .A(n7915), .B(n7916), .ZN(n13122)
         );
  OR2_X1 U8982 ( .A1(n9436), .A2(n10713), .ZN(n7915) );
  INV_X1 U8983 ( .A(n7917), .ZN(n7916) );
  OAI22_X1 U8984 ( .A1(n9211), .A2(n9157), .B1(n9177), .B2(n11062), .ZN(n7917)
         );
  INV_X1 U8985 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n11090) );
  AOI21_X1 U8986 ( .B1(n10986), .B2(n10984), .A(n10985), .ZN(n10988) );
  NAND2_X1 U8987 ( .A1(n7574), .A2(n7575), .ZN(n10976) );
  NAND2_X1 U8988 ( .A1(n7696), .A2(n9990), .ZN(n10781) );
  NAND2_X1 U8989 ( .A1(n10772), .A2(n7567), .ZN(n7561) );
  NOR2_X1 U8990 ( .A1(n11080), .A2(n15802), .ZN(n6996) );
  OR2_X1 U8991 ( .A1(n11080), .A2(n6997), .ZN(n10951) );
  INV_X1 U8992 ( .A(n6995), .ZN(n6997) );
  OAI211_X1 U8993 ( .C1(n6995), .C2(n11080), .A(n6994), .B(n11079), .ZN(n11558) );
  NAND2_X1 U8994 ( .A1(n11553), .A2(n6980), .ZN(n11801) );
  NAND2_X1 U8995 ( .A1(n11562), .A2(n6991), .ZN(n11811) );
  NAND2_X1 U8996 ( .A1(n6979), .A2(n6978), .ZN(n11805) );
  NAND2_X1 U8997 ( .A1(n6981), .A2(n11802), .ZN(n6978) );
  NAND2_X1 U8998 ( .A1(n13147), .A2(n7666), .ZN(n13135) );
  OAI21_X1 U8999 ( .B1(n13199), .B2(n13197), .A(n13198), .ZN(n13222) );
  INV_X1 U9000 ( .A(n13193), .ZN(n7671) );
  NAND2_X1 U9001 ( .A1(n13206), .A2(n7586), .ZN(n13211) );
  NAND2_X1 U9002 ( .A1(n7704), .A2(n13242), .ZN(n13243) );
  INV_X1 U9003 ( .A(n7705), .ZN(n7704) );
  AND2_X1 U9004 ( .A1(n13242), .A2(n13224), .ZN(n13225) );
  NOR2_X1 U9005 ( .A1(n7676), .A2(n7675), .ZN(n13251) );
  NAND2_X1 U9006 ( .A1(n13254), .A2(n13235), .ZN(n7560) );
  AND3_X1 U9007 ( .A1(n13288), .A2(n13287), .A3(n13286), .ZN(n13289) );
  AND2_X1 U9008 ( .A1(n9996), .A2(n9993), .ZN(n13318) );
  NAND2_X1 U9009 ( .A1(n7700), .A2(n7698), .ZN(n13311) );
  XNOR2_X1 U9010 ( .A(n6975), .B(n13331), .ZN(n6974) );
  NAND2_X1 U9011 ( .A1(n13325), .A2(n7582), .ZN(n6975) );
  AND2_X1 U9012 ( .A1(n9996), .A2(n13724), .ZN(n13313) );
  NOR2_X1 U9013 ( .A1(n9866), .A2(n9865), .ZN(n9867) );
  NOR2_X1 U9014 ( .A1(n12004), .A2(n13335), .ZN(n9866) );
  INV_X1 U9015 ( .A(n7257), .ZN(n7256) );
  OAI21_X1 U9016 ( .B1(n13350), .B2(n7259), .A(n13552), .ZN(n7258) );
  OAI22_X1 U9017 ( .A1(n13352), .A2(n13535), .B1(n13533), .B2(n13353), .ZN(
        n7257) );
  NAND2_X1 U9018 ( .A1(n13440), .A2(n9659), .ZN(n13427) );
  NAND2_X1 U9019 ( .A1(n13443), .A2(n9795), .ZN(n13430) );
  INV_X1 U9020 ( .A(n13553), .ZN(n13540) );
  AND2_X1 U9021 ( .A1(n11429), .A2(n13598), .ZN(n13558) );
  NAND2_X1 U9022 ( .A1(n11400), .A2(n11399), .ZN(n7907) );
  NOR2_X1 U9023 ( .A1(n13540), .A2(n10759), .ZN(n13400) );
  INV_X1 U9024 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10811) );
  INV_X1 U9025 ( .A(n13479), .ZN(n13557) );
  INV_X1 U9026 ( .A(n13558), .ZN(n13456) );
  NAND2_X1 U9027 ( .A1(n9140), .A2(n9139), .ZN(n13622) );
  NAND2_X1 U9028 ( .A1(n13403), .A2(n6895), .ZN(n6894) );
  NAND2_X1 U9029 ( .A1(n13383), .A2(n9672), .ZN(n13369) );
  NAND2_X1 U9030 ( .A1(n9471), .A2(n9470), .ZN(n13649) );
  NAND2_X1 U9031 ( .A1(n13428), .A2(n9796), .ZN(n13419) );
  NAND2_X1 U9032 ( .A1(n9403), .A2(n9402), .ZN(n13672) );
  NAND2_X1 U9033 ( .A1(n9393), .A2(n9392), .ZN(n13679) );
  NAND2_X1 U9034 ( .A1(n7926), .A2(n7928), .ZN(n13500) );
  NAND2_X1 U9035 ( .A1(n13545), .A2(n7932), .ZN(n7926) );
  NAND2_X1 U9036 ( .A1(n9331), .A2(n9330), .ZN(n12113) );
  NAND2_X1 U9037 ( .A1(n7898), .A2(n7900), .ZN(n11783) );
  NAND2_X1 U9038 ( .A1(n7899), .A2(n6625), .ZN(n7898) );
  INV_X1 U9039 ( .A(n11720), .ZN(n11767) );
  INV_X1 U9040 ( .A(n13688), .ZN(n13695) );
  INV_X1 U9041 ( .A(n9766), .ZN(n10715) );
  AND2_X1 U9042 ( .A1(n9826), .A2(n9825), .ZN(n13701) );
  OR2_X1 U9043 ( .A1(n10082), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9826) );
  INV_X1 U9044 ( .A(n10081), .ZN(n13702) );
  OAI21_X1 U9045 ( .B1(n6896), .B2(n9734), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n6897) );
  INV_X1 U9046 ( .A(SI_24_), .ZN(n11701) );
  NAND2_X1 U9047 ( .A1(n7251), .A2(n7249), .ZN(n11703) );
  NOR2_X1 U9048 ( .A1(n6558), .A2(n7250), .ZN(n7249) );
  OR2_X1 U9049 ( .A1(n9733), .A2(n9812), .ZN(n7251) );
  NOR2_X1 U9050 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), .ZN(
        n7250) );
  INV_X1 U9051 ( .A(SI_23_), .ZN(n11314) );
  XNOR2_X1 U9052 ( .A(n9583), .B(P3_IR_REG_22__SCAN_IN), .ZN(n11110) );
  NAND2_X1 U9053 ( .A1(n9575), .A2(n9582), .ZN(n11382) );
  INV_X1 U9054 ( .A(SI_20_), .ZN(n11250) );
  OAI21_X1 U9055 ( .B1(n7639), .B2(n7638), .A(n7635), .ZN(n11251) );
  NAND2_X1 U9056 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_20__SCAN_IN), 
        .ZN(n7638) );
  NOR2_X1 U9057 ( .A1(n7637), .A2(n7636), .ZN(n7635) );
  NOR2_X1 U9058 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7636) );
  INV_X1 U9059 ( .A(SI_19_), .ZN(n10630) );
  NAND2_X1 U9060 ( .A1(n9427), .A2(n9567), .ZN(n10631) );
  INV_X1 U9061 ( .A(n7639), .ZN(n9567) );
  INV_X1 U9062 ( .A(SI_18_), .ZN(n10549) );
  INV_X1 U9063 ( .A(SI_17_), .ZN(n10395) );
  INV_X1 U9064 ( .A(SI_13_), .ZN(n10281) );
  INV_X1 U9065 ( .A(SI_12_), .ZN(n10183) );
  INV_X1 U9066 ( .A(SI_11_), .ZN(n10166) );
  OAI21_X1 U9067 ( .B1(n9274), .B2(n7108), .A(n7105), .ZN(n9307) );
  NAND2_X1 U9068 ( .A1(n9291), .A2(n9290), .ZN(n9293) );
  XNOR2_X1 U9069 ( .A(n9295), .B(n9294), .ZN(n13124) );
  NAND2_X1 U9070 ( .A1(n9221), .A2(n9039), .ZN(n9235) );
  NAND2_X1 U9071 ( .A1(n9204), .A2(n9203), .ZN(n9206) );
  NAND2_X1 U9072 ( .A1(n9186), .A2(n9035), .ZN(n9204) );
  INV_X1 U9073 ( .A(n7093), .ZN(n9162) );
  NAND2_X1 U9074 ( .A1(n9953), .A2(n9811), .ZN(n6986) );
  AND2_X1 U9075 ( .A1(n10426), .A2(n9930), .ZN(n10430) );
  NAND2_X1 U9076 ( .A1(n7350), .A2(n7730), .ZN(n11642) );
  INV_X1 U9077 ( .A(n7731), .ZN(n7730) );
  OAI21_X1 U9078 ( .B1(n7733), .B2(n7732), .A(n11385), .ZN(n7731) );
  NAND2_X1 U9079 ( .A1(n11384), .A2(n11383), .ZN(n11386) );
  NAND2_X1 U9080 ( .A1(n12617), .A2(n12616), .ZN(n13757) );
  NAND2_X1 U9081 ( .A1(n12029), .A2(n12028), .ZN(n12601) );
  NAND2_X1 U9082 ( .A1(n10408), .A2(n10021), .ZN(n10033) );
  NAND2_X1 U9083 ( .A1(n12654), .A2(n13850), .ZN(n13800) );
  NAND2_X1 U9084 ( .A1(n7351), .A2(n7352), .ZN(n11256) );
  NAND2_X1 U9085 ( .A1(n7388), .A2(n7386), .ZN(n13833) );
  AND2_X1 U9086 ( .A1(n7388), .A2(n7385), .ZN(n13835) );
  NAND2_X1 U9087 ( .A1(n13823), .A2(n12632), .ZN(n7388) );
  NAND2_X1 U9088 ( .A1(n10855), .A2(n10854), .ZN(n11228) );
  NAND2_X1 U9089 ( .A1(n7744), .A2(n11921), .ZN(n11924) );
  AND2_X1 U9090 ( .A1(n13775), .A2(n12648), .ZN(n13852) );
  OAI21_X1 U9091 ( .B1(n7744), .B2(n7360), .A(n7358), .ZN(n13882) );
  NAND2_X1 U9092 ( .A1(n12007), .A2(n8264), .ZN(n7345) );
  NAND2_X1 U9093 ( .A1(n7380), .A2(n7382), .ZN(n13891) );
  NAND2_X1 U9094 ( .A1(n7381), .A2(n7386), .ZN(n7380) );
  INV_X1 U9095 ( .A(n13823), .ZN(n7381) );
  NAND2_X1 U9096 ( .A1(n8255), .A2(n8254), .ZN(n14460) );
  NAND2_X1 U9097 ( .A1(n11256), .A2(n7733), .ZN(n11384) );
  AND2_X1 U9098 ( .A1(n10397), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13859) );
  INV_X1 U9099 ( .A(n13855), .ZN(n13919) );
  INV_X1 U9100 ( .A(n13859), .ZN(n13921) );
  NAND2_X1 U9101 ( .A1(n10040), .A2(n10029), .ZN(n13925) );
  NAND2_X1 U9102 ( .A1(n8686), .A2(n8685), .ZN(n13931) );
  NAND4_X1 U9103 ( .A1(n8474), .A2(n8473), .A3(n8472), .A4(n8471), .ZN(n13954)
         );
  OR2_X1 U9104 ( .A1(n8944), .A2(n10417), .ZN(n8462) );
  OR2_X1 U9105 ( .A1(n8468), .A2(n8439), .ZN(n8440) );
  OR2_X1 U9106 ( .A1(n8945), .A2(n11977), .ZN(n8442) );
  OR2_X1 U9107 ( .A1(n8945), .A2(n8447), .ZN(n8448) );
  NAND2_X1 U9108 ( .A1(n14001), .A2(n10421), .ZN(n14013) );
  NAND2_X1 U9109 ( .A1(n14013), .A2(n14014), .ZN(n14012) );
  AOI21_X1 U9110 ( .B1(n6805), .B2(n6807), .A(n6804), .ZN(n6803) );
  INV_X1 U9111 ( .A(n14031), .ZN(n6804) );
  OAI21_X1 U9112 ( .B1(n14001), .B2(n6807), .A(n6805), .ZN(n14032) );
  NAND2_X1 U9113 ( .A1(n10477), .A2(n10476), .ZN(n10718) );
  NAND2_X1 U9114 ( .A1(n10716), .A2(n10478), .ZN(n14044) );
  NAND2_X1 U9115 ( .A1(n10842), .A2(n10841), .ZN(n10867) );
  NAND2_X1 U9116 ( .A1(n10865), .A2(n10844), .ZN(n10847) );
  NAND2_X1 U9117 ( .A1(n8198), .A2(n7749), .ZN(n8229) );
  NAND2_X1 U9118 ( .A1(n11880), .A2(n11823), .ZN(n11825) );
  NAND2_X1 U9119 ( .A1(n6784), .A2(n6609), .ZN(n14066) );
  OR2_X1 U9120 ( .A1(n11882), .A2(n6788), .ZN(n6784) );
  OR2_X1 U9121 ( .A1(n14071), .A2(n14070), .ZN(n14080) );
  AND2_X1 U9122 ( .A1(n10454), .A2(n8399), .ZN(n15644) );
  INV_X1 U9123 ( .A(n7160), .ZN(n7159) );
  XNOR2_X1 U9124 ( .A(n7127), .B(n8765), .ZN(n14118) );
  OAI21_X1 U9125 ( .B1(n14127), .B2(n6652), .A(n6580), .ZN(n7127) );
  NAND2_X1 U9126 ( .A1(n7550), .A2(n7554), .ZN(n14141) );
  NAND2_X1 U9127 ( .A1(n14174), .A2(n7555), .ZN(n7550) );
  AND2_X1 U9128 ( .A1(n6765), .A2(n14165), .ZN(n14427) );
  NAND2_X1 U9129 ( .A1(n7557), .A2(n7555), .ZN(n14165) );
  NAND2_X1 U9130 ( .A1(n7557), .A2(n7558), .ZN(n14164) );
  NAND2_X1 U9131 ( .A1(n7534), .A2(n8627), .ZN(n14212) );
  NAND2_X1 U9132 ( .A1(n14239), .A2(n9013), .ZN(n8618) );
  INV_X1 U9133 ( .A(n14460), .ZN(n14260) );
  NAND2_X1 U9134 ( .A1(n7335), .A2(n7336), .ZN(n14268) );
  NAND2_X1 U9135 ( .A1(n7038), .A2(n7042), .ZN(n7335) );
  NAND2_X1 U9136 ( .A1(n14303), .A2(n8589), .ZN(n7523) );
  OAI21_X1 U9137 ( .B1(n14299), .B2(n8715), .A(n8717), .ZN(n14286) );
  OAI21_X1 U9138 ( .B1(n8539), .B2(n7539), .A(n7541), .ZN(n14331) );
  NAND2_X1 U9139 ( .A1(n7545), .A2(n8547), .ZN(n14346) );
  NAND2_X1 U9140 ( .A1(n8539), .A2(n7546), .ZN(n7545) );
  NAND2_X1 U9141 ( .A1(n8539), .A2(n8538), .ZN(n11727) );
  INV_X1 U9142 ( .A(n14401), .ZN(n14370) );
  INV_X1 U9143 ( .A(n14399), .ZN(n14368) );
  INV_X1 U9144 ( .A(n10035), .ZN(n10036) );
  INV_X1 U9145 ( .A(n14398), .ZN(n15666) );
  OR2_X1 U9146 ( .A1(n8376), .A2(n10053), .ZN(n8119) );
  OR2_X1 U9147 ( .A1(n10428), .A2(n13964), .ZN(n8120) );
  NAND2_X1 U9148 ( .A1(n6817), .A2(n6816), .ZN(n6815) );
  INV_X1 U9149 ( .A(n14105), .ZN(n6816) );
  AND2_X1 U9150 ( .A1(n8303), .A2(n8302), .ZN(n14545) );
  AND2_X1 U9151 ( .A1(n8295), .A2(n8294), .ZN(n14548) );
  INV_X1 U9152 ( .A(n14339), .ZN(n14564) );
  NOR2_X1 U9153 ( .A1(n15670), .A2(n15699), .ZN(n15694) );
  INV_X1 U9155 ( .A(n15702), .ZN(n15699) );
  AND2_X1 U9156 ( .A1(n10426), .A2(n9024), .ZN(n15702) );
  AND2_X1 U9157 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9929), .ZN(n9024) );
  INV_X1 U9158 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n14581) );
  INV_X1 U9159 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n16023) );
  NAND2_X1 U9160 ( .A1(n8412), .A2(n8411), .ZN(n12119) );
  INV_X1 U9161 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11898) );
  NAND2_X1 U9162 ( .A1(n8406), .A2(n8408), .ZN(n11895) );
  INV_X1 U9163 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11284) );
  INV_X1 U9164 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n15896) );
  INV_X1 U9165 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n15888) );
  INV_X1 U9166 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10641) );
  INV_X1 U9167 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10554) );
  INV_X1 U9168 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10309) );
  INV_X1 U9169 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10286) );
  INV_X1 U9170 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n16097) );
  INV_X1 U9171 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10168) );
  INV_X1 U9172 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10121) );
  INV_X1 U9173 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10124) );
  INV_X1 U9174 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10069) );
  INV_X1 U9175 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10067) );
  INV_X1 U9176 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10056) );
  AND2_X1 U9177 ( .A1(n12407), .A2(n12406), .ZN(n14959) );
  OR2_X1 U9178 ( .A1(n14944), .A2(n11447), .ZN(n12407) );
  NOR2_X1 U9179 ( .A1(n7143), .A2(n7140), .ZN(n7139) );
  INV_X1 U9180 ( .A(n7144), .ZN(n7140) );
  NAND2_X1 U9181 ( .A1(n7144), .A2(n7145), .ZN(n7141) );
  CLKBUF_X1 U9182 ( .A(n11017), .Z(n14620) );
  NAND2_X1 U9183 ( .A1(n14734), .A2(n12516), .ZN(n14631) );
  AND2_X1 U9184 ( .A1(n7991), .A2(n6642), .ZN(n14657) );
  NAND2_X1 U9185 ( .A1(n7983), .A2(n12230), .ZN(n12474) );
  INV_X1 U9186 ( .A(n12228), .ZN(n7983) );
  INV_X1 U9187 ( .A(n7996), .ZN(n6851) );
  NAND2_X1 U9188 ( .A1(n14598), .A2(n7998), .ZN(n7993) );
  NAND2_X1 U9189 ( .A1(n14610), .A2(n14695), .ZN(n7976) );
  NAND2_X1 U9190 ( .A1(n12301), .A2(n12393), .ZN(n7311) );
  OR2_X1 U9191 ( .A1(n14737), .A2(n15128), .ZN(n14715) );
  NAND2_X1 U9192 ( .A1(n7128), .A2(n7981), .ZN(n14712) );
  AND2_X1 U9193 ( .A1(n14713), .A2(n7982), .ZN(n7981) );
  NAND2_X1 U9194 ( .A1(n12228), .A2(n12473), .ZN(n7128) );
  NAND2_X1 U9195 ( .A1(n12229), .A2(n12473), .ZN(n7982) );
  NAND2_X1 U9196 ( .A1(n12474), .A2(n12473), .ZN(n14714) );
  NAND2_X1 U9197 ( .A1(n8000), .A2(n8003), .ZN(n12141) );
  NAND2_X1 U9198 ( .A1(n11868), .A2(n8004), .ZN(n8000) );
  NAND2_X1 U9199 ( .A1(n7131), .A2(n7132), .ZN(n7130) );
  NAND2_X1 U9200 ( .A1(n11325), .A2(n11324), .ZN(n7286) );
  AOI21_X1 U9201 ( .B1(n6627), .B2(n7134), .A(n7133), .ZN(n7132) );
  NAND2_X1 U9202 ( .A1(n11192), .A2(n11191), .ZN(n12712) );
  AND2_X1 U9203 ( .A1(n10918), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14690) );
  AND2_X1 U9204 ( .A1(n11042), .A2(n15530), .ZN(n14740) );
  INV_X1 U9205 ( .A(n14690), .ZN(n14759) );
  AND2_X1 U9206 ( .A1(n10389), .A2(n10388), .ZN(n14753) );
  NOR2_X1 U9207 ( .A1(n10915), .A2(P1_U3086), .ZN(n12913) );
  INV_X1 U9208 ( .A(n12864), .ZN(n12865) );
  INV_X1 U9209 ( .A(n14959), .ZN(n14769) );
  OR2_X1 U9210 ( .A1(n15012), .A2(n11447), .ZN(n12371) );
  OR2_X1 U9211 ( .A1(n12260), .A2(n12259), .ZN(n15179) );
  NAND4_X1 U9212 ( .A1(n10926), .A2(n10925), .A3(n10924), .A4(n10923), .ZN(
        n14787) );
  OR2_X1 U9213 ( .A1(n10700), .A2(n10701), .ZN(n10704) );
  NAND3_X2 U9214 ( .A1(n10680), .A2(n10679), .A3(n10678), .ZN(n14790) );
  CLKBUF_X2 U9215 ( .A(P1_U4016), .Z(n14791) );
  NAND2_X1 U9216 ( .A1(n14802), .A2(n14801), .ZN(n14800) );
  XNOR2_X1 U9217 ( .A(n10054), .B(P1_IR_REG_3__SCAN_IN), .ZN(n14828) );
  NAND2_X1 U9218 ( .A1(n6731), .A2(n6874), .ZN(n6873) );
  AND2_X1 U9219 ( .A1(n10231), .A2(n10228), .ZN(n15475) );
  AOI21_X1 U9220 ( .B1(n14846), .B2(n10657), .A(n10656), .ZN(n10826) );
  AND2_X1 U9221 ( .A1(n6906), .A2(n6607), .ZN(n10819) );
  INV_X1 U9222 ( .A(n7078), .ZN(n11482) );
  OAI21_X1 U9223 ( .B1(n14846), .B2(n6664), .A(n7075), .ZN(n7078) );
  NAND2_X1 U9224 ( .A1(n11113), .A2(n7082), .ZN(n11116) );
  OR2_X1 U9225 ( .A1(n12071), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6881) );
  AND2_X1 U9226 ( .A1(n6878), .A2(n6877), .ZN(n14854) );
  XNOR2_X1 U9227 ( .A(n14869), .B(n7502), .ZN(n15482) );
  NAND2_X1 U9228 ( .A1(n15479), .A2(n14876), .ZN(n14878) );
  NAND2_X1 U9229 ( .A1(n6868), .A2(n6867), .ZN(n14870) );
  NAND2_X1 U9230 ( .A1(n7494), .A2(n15819), .ZN(n7493) );
  OAI22_X1 U9231 ( .A1(n15818), .A2(n15817), .B1(n15816), .B2(n15815), .ZN(
        n7494) );
  INV_X1 U9232 ( .A(n7496), .ZN(n7495) );
  OAI21_X1 U9233 ( .B1(n15821), .B2(n16058), .A(n15820), .ZN(n7496) );
  INV_X1 U9234 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n16119) );
  INV_X1 U9235 ( .A(n14916), .ZN(n15201) );
  INV_X1 U9236 ( .A(n14923), .ZN(n15206) );
  NAND2_X1 U9237 ( .A1(n12441), .A2(n6619), .ZN(n7944) );
  INV_X1 U9238 ( .A(n12819), .ZN(n15210) );
  AND2_X1 U9239 ( .A1(n12396), .A2(n12395), .ZN(n14962) );
  AOI21_X1 U9240 ( .B1(n6948), .B2(n12385), .A(n12386), .ZN(n14953) );
  AND2_X1 U9241 ( .A1(n12374), .A2(n12373), .ZN(n14980) );
  NAND2_X1 U9242 ( .A1(n7240), .A2(n7814), .ZN(n15000) );
  NAND2_X1 U9243 ( .A1(n15261), .A2(n12433), .ZN(n15005) );
  NAND2_X1 U9244 ( .A1(n15035), .A2(n12339), .ZN(n15020) );
  OR2_X1 U9245 ( .A1(n15030), .A2(n15029), .ZN(n15261) );
  INV_X1 U9246 ( .A(n15267), .ZN(n15044) );
  AND2_X1 U9247 ( .A1(n12314), .A2(n12313), .ZN(n15059) );
  AND2_X1 U9248 ( .A1(n15053), .A2(n15052), .ZN(n15274) );
  OR2_X1 U9249 ( .A1(n15060), .A2(n15075), .ZN(n15277) );
  INV_X1 U9250 ( .A(n15287), .ZN(n15095) );
  NAND2_X1 U9251 ( .A1(n15107), .A2(n12779), .ZN(n15087) );
  NAND2_X1 U9252 ( .A1(n7811), .A2(n12421), .ZN(n15106) );
  NAND2_X1 U9253 ( .A1(n12420), .A2(n7812), .ZN(n7811) );
  NAND2_X1 U9254 ( .A1(n11105), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10332) );
  NAND2_X1 U9255 ( .A1(n12420), .A2(n12419), .ZN(n15123) );
  NAND2_X1 U9256 ( .A1(n12250), .A2(n12393), .ZN(n12252) );
  NAND2_X1 U9257 ( .A1(n15192), .A2(n12417), .ZN(n15159) );
  NAND2_X1 U9258 ( .A1(n12244), .A2(n12393), .ZN(n7788) );
  INV_X1 U9259 ( .A(n15319), .ZN(n14723) );
  OAI21_X1 U9260 ( .B1(n12092), .B2(n7222), .A(n7224), .ZN(n12176) );
  INV_X1 U9261 ( .A(n7220), .ZN(n7224) );
  NAND2_X1 U9262 ( .A1(n12066), .A2(n7485), .ZN(n12022) );
  INV_X1 U9263 ( .A(n7487), .ZN(n7485) );
  OR2_X1 U9264 ( .A1(n15525), .A2(n11141), .ZN(n15147) );
  NAND2_X1 U9265 ( .A1(n6740), .A2(n11548), .ZN(n11550) );
  NAND2_X1 U9266 ( .A1(n11442), .A2(n11441), .ZN(n15516) );
  INV_X1 U9267 ( .A(n15189), .ZN(n15513) );
  INV_X1 U9268 ( .A(n15082), .ZN(n15521) );
  INV_X1 U9269 ( .A(n15147), .ZN(n15515) );
  OR2_X1 U9270 ( .A1(n11131), .A2(n11130), .ZN(n15189) );
  INV_X1 U9271 ( .A(n15195), .ZN(n15101) );
  AND2_X1 U9272 ( .A1(n15224), .A2(n15223), .ZN(n15225) );
  AND2_X1 U9273 ( .A1(n15222), .A2(n15221), .ZN(n15223) );
  OR2_X1 U9274 ( .A1(n10333), .A2(P1_U3086), .ZN(n10191) );
  CLKBUF_X1 U9275 ( .A(n15473), .Z(n6762) );
  INV_X1 U9276 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11894) );
  NAND2_X1 U9277 ( .A1(n9951), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U9278 ( .A1(n9951), .A2(n9952), .ZN(n11786) );
  INV_X1 U9279 ( .A(n10354), .ZN(n12917) );
  INV_X1 U9280 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11281) );
  INV_X1 U9281 ( .A(n12675), .ZN(n11280) );
  INV_X1 U9282 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n16042) );
  INV_X1 U9283 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10545) );
  INV_X1 U9284 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10201) );
  INV_X1 U9285 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10179) );
  INV_X1 U9286 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10174) );
  INV_X1 U9287 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10100) );
  INV_X1 U9288 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10087) );
  INV_X1 U9289 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16025) );
  XNOR2_X1 U9290 ( .A(n10089), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10898) );
  NAND2_X1 U9291 ( .A1(n10088), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10089) );
  NAND2_X1 U9292 ( .A1(n7506), .A2(n7505), .ZN(n10094) );
  NAND2_X1 U9293 ( .A1(n9931), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7505) );
  NAND2_X1 U9294 ( .A1(n7059), .A2(n10092), .ZN(n10666) );
  INV_X1 U9295 ( .A(n10050), .ZN(n10092) );
  NAND2_X1 U9296 ( .A1(n7305), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7304) );
  OR2_X1 U9297 ( .A1(n10152), .A2(n10151), .ZN(n15468) );
  XNOR2_X1 U9298 ( .A(n10159), .B(n10138), .ZN(n15384) );
  XNOR2_X1 U9299 ( .A(n10938), .B(n10936), .ZN(n10935) );
  NAND2_X1 U9300 ( .A1(n7205), .A2(n7203), .ZN(n11301) );
  AND2_X1 U9301 ( .A1(n10939), .A2(n7204), .ZN(n7203) );
  INV_X1 U9302 ( .A(n10945), .ZN(n7204) );
  INV_X1 U9303 ( .A(n11679), .ZN(n7208) );
  NAND2_X1 U9304 ( .A1(n7209), .A2(n11679), .ZN(n12038) );
  NAND2_X1 U9305 ( .A1(n11671), .A2(n11670), .ZN(n7209) );
  AND2_X1 U9306 ( .A1(n7655), .A2(n7653), .ZN(n7652) );
  INV_X1 U9307 ( .A(n12202), .ZN(n7653) );
  INV_X1 U9308 ( .A(n15415), .ZN(n7656) );
  CLKBUF_X2 U9309 ( .A(n13115), .Z(P3_U3897) );
  NAND2_X1 U9310 ( .A1(n11607), .A2(n11606), .ZN(n11748) );
  NAND2_X1 U9311 ( .A1(n7274), .A2(n11592), .ZN(n11595) );
  NAND2_X1 U9312 ( .A1(n7578), .A2(n7577), .ZN(n10729) );
  NOR2_X1 U9313 ( .A1(n7289), .A2(n6653), .ZN(n7288) );
  NOR2_X1 U9314 ( .A1(n15804), .A2(n9846), .ZN(n7289) );
  NOR2_X1 U9315 ( .A1(n7292), .A2(n6654), .ZN(n7291) );
  NOR2_X1 U9316 ( .A1(n15786), .A2(n16000), .ZN(n7292) );
  AOI21_X1 U9317 ( .B1(n9023), .B2(n9010), .A(n9027), .ZN(n7826) );
  AND2_X1 U9318 ( .A1(n6790), .A2(n14087), .ZN(n6789) );
  NAND2_X1 U9319 ( .A1(n6796), .A2(n8775), .ZN(n6795) );
  NAND2_X1 U9320 ( .A1(n6792), .A2(n14086), .ZN(n6791) );
  MUX2_X1 U9321 ( .A(n15880), .B(n14406), .S(n15750), .Z(n14407) );
  NAND2_X1 U9322 ( .A1(n6813), .A2(n6811), .ZN(P2_U3528) );
  NOR2_X1 U9323 ( .A1(n6812), .A2(n6651), .ZN(n6811) );
  OR2_X1 U9324 ( .A1(n9927), .A2(n12591), .ZN(n6813) );
  NOR2_X1 U9325 ( .A1(n15750), .A2(n9928), .ZN(n6812) );
  NAND2_X1 U9326 ( .A1(n7101), .A2(n7099), .ZN(P2_U3526) );
  INV_X1 U9327 ( .A(n7100), .ZN(n7099) );
  OAI22_X1 U9328 ( .A1(n14414), .A2(n14514), .B1(n15750), .B2(n16101), .ZN(
        n7100) );
  MUX2_X1 U9329 ( .A(n14428), .B(n14535), .S(n15750), .Z(n14429) );
  INV_X1 U9330 ( .A(n7048), .ZN(n14535) );
  AND2_X1 U9331 ( .A1(n8031), .A2(n8013), .ZN(n8772) );
  NAND2_X1 U9332 ( .A1(n7339), .A2(n7338), .ZN(n14529) );
  NAND2_X1 U9333 ( .A1(n15741), .A2(n14528), .ZN(n7338) );
  NAND2_X1 U9334 ( .A1(n14527), .A2(n15743), .ZN(n7339) );
  NAND2_X1 U9335 ( .A1(n7047), .A2(n7045), .ZN(P2_U3491) );
  AOI21_X1 U9336 ( .B1(n14167), .B2(n8433), .A(n7046), .ZN(n7045) );
  NAND2_X1 U9337 ( .A1(n7048), .A2(n15743), .ZN(n7047) );
  NOR2_X1 U9338 ( .A1(n15743), .A2(n14536), .ZN(n7046) );
  NAND2_X1 U9339 ( .A1(n10267), .A2(n7498), .ZN(n10268) );
  OAI21_X1 U9340 ( .B1(n6865), .B2(n7492), .A(n6864), .ZN(n14886) );
  AND2_X1 U9341 ( .A1(n6904), .A2(n6903), .ZN(n15806) );
  NAND2_X1 U9342 ( .A1(n15620), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n7241) );
  NAND2_X1 U9343 ( .A1(n7789), .A2(n7334), .ZN(n7243) );
  OAI211_X1 U9344 ( .C1(n7789), .C2(n15606), .A(n6781), .B(n7940), .ZN(
        P1_U3525) );
  INV_X1 U9345 ( .A(n6782), .ZN(n6781) );
  OAI21_X1 U9346 ( .B1(n7790), .B2(n15606), .A(n7945), .ZN(n6782) );
  NAND2_X1 U9347 ( .A1(n10255), .A2(n10254), .ZN(n15365) );
  NAND2_X1 U9348 ( .A1(n7650), .A2(n10603), .ZN(n10604) );
  INV_X1 U9349 ( .A(n7651), .ZN(n7650) );
  NAND2_X1 U9350 ( .A1(n12045), .A2(n12046), .ZN(n12193) );
  OR2_X1 U9351 ( .A1(n12045), .A2(n12046), .ZN(n12194) );
  NAND2_X1 U9352 ( .A1(n7642), .A2(n15441), .ZN(n15443) );
  NAND2_X1 U9353 ( .A1(n15435), .A2(n15434), .ZN(n7642) );
  NOR2_X1 U9354 ( .A1(n15456), .A2(n15455), .ZN(n15464) );
  AND3_X1 U9355 ( .A1(n7312), .A2(n15075), .A3(n6576), .ZN(n6563) );
  NAND2_X1 U9356 ( .A1(n7522), .A2(n7521), .ZN(n8098) );
  XNOR2_X1 U9357 ( .A(n13752), .B(n8764), .ZN(n9019) );
  INV_X1 U9358 ( .A(n9019), .ZN(n8765) );
  NOR2_X1 U9359 ( .A1(n15331), .A2(n14781), .ZN(n6565) );
  NAND2_X1 U9360 ( .A1(n8008), .A2(n6596), .ZN(n10202) );
  NAND2_X1 U9361 ( .A1(n6740), .A2(n7963), .ZN(n12015) );
  AND2_X1 U9362 ( .A1(n9778), .A2(n9777), .ZN(n6566) );
  NOR2_X1 U9363 ( .A1(n12423), .A2(n7810), .ZN(n6567) );
  AND2_X1 U9364 ( .A1(n7303), .A2(n7302), .ZN(n6568) );
  NAND2_X1 U9365 ( .A1(n14541), .A2(n7507), .ZN(n6569) );
  XNOR2_X1 U9366 ( .A(n15259), .B(n14774), .ZN(n15029) );
  AND2_X1 U9367 ( .A1(n6694), .A2(n7013), .ZN(n6570) );
  AND2_X1 U9368 ( .A1(n7900), .A2(n11779), .ZN(n6571) );
  NAND2_X1 U9369 ( .A1(n6677), .A2(n7757), .ZN(n6572) );
  OR2_X1 U9370 ( .A1(n9019), .A2(n7784), .ZN(n6573) );
  AND2_X1 U9371 ( .A1(n7267), .A2(n7266), .ZN(n6574) );
  INV_X1 U9372 ( .A(n14619), .ZN(n15259) );
  NOR2_X1 U9373 ( .A1(n9971), .A2(n10991), .ZN(n6575) );
  NAND2_X1 U9374 ( .A1(n15095), .A2(n14776), .ZN(n6576) );
  AND2_X1 U9375 ( .A1(n8285), .A2(n6666), .ZN(n6577) );
  OR2_X1 U9376 ( .A1(n13593), .A2(n13108), .ZN(n9706) );
  INV_X1 U9377 ( .A(n8709), .ZN(n7762) );
  OR2_X1 U9378 ( .A1(n7542), .A2(n8565), .ZN(n6578) );
  NAND2_X1 U9379 ( .A1(n7771), .A2(n8703), .ZN(n11687) );
  BUF_X1 U9380 ( .A(n8779), .Z(n15707) );
  XNOR2_X1 U9381 ( .A(n9922), .B(n9006), .ZN(n9910) );
  INV_X1 U9382 ( .A(n9910), .ZN(n7165) );
  AND2_X1 U9383 ( .A1(n7952), .A2(n7332), .ZN(n6579) );
  NAND2_X1 U9384 ( .A1(n14130), .A2(n13932), .ZN(n6580) );
  AND2_X1 U9385 ( .A1(n7230), .A2(n6567), .ZN(n6581) );
  INV_X1 U9386 ( .A(n7450), .ZN(n7449) );
  AND2_X1 U9387 ( .A1(n14555), .A2(n14260), .ZN(n6582) );
  AND4_X1 U9388 ( .A1(n7154), .A2(n14264), .A3(n7149), .A4(n7148), .ZN(n6583)
         );
  INV_X1 U9389 ( .A(n12802), .ZN(n6919) );
  AND2_X1 U9390 ( .A1(n12095), .A2(n6714), .ZN(n6584) );
  NAND2_X1 U9391 ( .A1(n15166), .A2(n7331), .ZN(n15150) );
  AND2_X1 U9392 ( .A1(n7372), .A2(n13733), .ZN(n6585) );
  NAND2_X1 U9393 ( .A1(n8358), .A2(n8357), .ZN(n9922) );
  INV_X1 U9394 ( .A(n9922), .ZN(n7520) );
  AND4_X1 U9395 ( .A1(n7168), .A2(n7166), .A3(n9018), .A4(n7165), .ZN(n6586)
         );
  AND2_X1 U9396 ( .A1(n8636), .A2(n8635), .ZN(n12655) );
  OR3_X1 U9397 ( .A1(n14216), .A2(n14182), .A3(n14194), .ZN(n6587) );
  AND2_X1 U9398 ( .A1(n7944), .A2(n15552), .ZN(n6588) );
  AND2_X1 U9399 ( .A1(n14083), .A2(n15644), .ZN(n6589) );
  AND2_X1 U9400 ( .A1(n12441), .A2(n14935), .ZN(n6590) );
  NAND2_X1 U9401 ( .A1(n9326), .A2(n9325), .ZN(n9734) );
  AND2_X1 U9402 ( .A1(n10256), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6591) );
  AND2_X1 U9403 ( .A1(n9015), .A2(n7535), .ZN(n6592) );
  AND2_X1 U9404 ( .A1(n7701), .A2(n13292), .ZN(n6593) );
  NAND2_X1 U9405 ( .A1(n13871), .A2(n12656), .ZN(n6594) );
  OR2_X1 U9406 ( .A1(n12755), .A2(n12756), .ZN(n6595) );
  AND2_X1 U9407 ( .A1(n8007), .A2(n10204), .ZN(n6596) );
  NAND2_X1 U9408 ( .A1(n6697), .A2(n8006), .ZN(n8003) );
  INV_X1 U9409 ( .A(n8098), .ZN(n7349) );
  NAND2_X1 U9410 ( .A1(n9145), .A2(n7891), .ZN(n9701) );
  NOR2_X1 U9411 ( .A1(n9604), .A2(n9855), .ZN(n6597) );
  NAND2_X1 U9412 ( .A1(n9718), .A2(n9703), .ZN(n6598) );
  AND2_X1 U9413 ( .A1(n11563), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n6599) );
  AND2_X1 U9414 ( .A1(n8475), .A2(n8466), .ZN(n6600) );
  NAND2_X1 U9415 ( .A1(n12046), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6601) );
  NAND2_X1 U9416 ( .A1(n10965), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n6602) );
  NAND2_X1 U9417 ( .A1(n12641), .A2(n12640), .ZN(n6603) );
  AND2_X1 U9418 ( .A1(n13147), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n6604) );
  NAND2_X1 U9419 ( .A1(n15185), .A2(n6595), .ZN(n6605) );
  OR2_X1 U9420 ( .A1(n7508), .A2(n6825), .ZN(n11735) );
  AND2_X1 U9421 ( .A1(n7540), .A2(n8556), .ZN(n7541) );
  AND2_X1 U9422 ( .A1(n9116), .A2(n7393), .ZN(n6606) );
  INV_X1 U9423 ( .A(n14695), .ZN(n7979) );
  NAND2_X1 U9424 ( .A1(n11868), .A2(n11867), .ZN(n12124) );
  NAND2_X1 U9425 ( .A1(n15287), .A2(n15070), .ZN(n12785) );
  INV_X1 U9426 ( .A(n7963), .ZN(n7328) );
  NAND2_X1 U9427 ( .A1(n11494), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6607) );
  INV_X1 U9428 ( .A(n12883), .ZN(n15494) );
  AND2_X1 U9429 ( .A1(n11562), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n6608) );
  AND2_X1 U9430 ( .A1(n6787), .A2(n11824), .ZN(n6609) );
  AND2_X1 U9431 ( .A1(n15380), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6610) );
  INV_X1 U9432 ( .A(n11324), .ZN(n7134) );
  AND2_X1 U9433 ( .A1(n10978), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n6611) );
  AND2_X1 U9434 ( .A1(n7702), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n6612) );
  AND2_X1 U9435 ( .A1(n7690), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n6613) );
  XNOR2_X1 U9436 ( .A(n10332), .B(P1_IR_REG_19__SCAN_IN), .ZN(n12672) );
  NAND2_X2 U9437 ( .A1(n11619), .A2(n14398), .ZN(n14285) );
  INV_X1 U9438 ( .A(n12103), .ZN(n6890) );
  NAND2_X1 U9439 ( .A1(n9360), .A2(n9359), .ZN(n13689) );
  NAND2_X1 U9440 ( .A1(n8109), .A2(n8084), .ZN(n8117) );
  NOR2_X1 U9441 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n8109) );
  AND2_X1 U9442 ( .A1(n12124), .A2(n12123), .ZN(n6614) );
  NAND2_X1 U9443 ( .A1(n15107), .A2(n7960), .ZN(n7962) );
  XNOR2_X1 U9444 ( .A(n9182), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10739) );
  INV_X1 U9445 ( .A(n15441), .ZN(n7643) );
  AND2_X1 U9446 ( .A1(n7976), .A2(n14696), .ZN(n6615) );
  NAND2_X1 U9447 ( .A1(n7740), .A2(n7738), .ZN(n13514) );
  AND2_X1 U9448 ( .A1(n7258), .A2(n7256), .ZN(n6616) );
  AND2_X1 U9449 ( .A1(n7974), .A2(n6842), .ZN(n6617) );
  INV_X1 U9450 ( .A(n12886), .ZN(n12175) );
  XNOR2_X1 U9451 ( .A(n12745), .B(n14780), .ZN(n12886) );
  AND2_X1 U9452 ( .A1(n7034), .A2(n12959), .ZN(n6618) );
  AND2_X1 U9453 ( .A1(n15220), .A2(n14959), .ZN(n6619) );
  AND2_X1 U9454 ( .A1(n13518), .A2(n9789), .ZN(n6620) );
  NAND2_X1 U9455 ( .A1(n9811), .A2(n7662), .ZN(n6621) );
  AND2_X1 U9456 ( .A1(n9663), .A2(n9664), .ZN(n13431) );
  AND2_X1 U9457 ( .A1(n9504), .A2(n9674), .ZN(n6622) );
  OR2_X1 U9458 ( .A1(n14534), .A2(n13933), .ZN(n6623) );
  NAND2_X1 U9459 ( .A1(n15236), .A2(n14771), .ZN(n6624) );
  NAND2_X1 U9460 ( .A1(n7228), .A2(n7230), .ZN(n12420) );
  AND2_X1 U9461 ( .A1(n11843), .A2(n7904), .ZN(n6625) );
  AND2_X1 U9462 ( .A1(n10260), .A2(n15374), .ZN(n10902) );
  NAND2_X1 U9463 ( .A1(n14274), .A2(n13892), .ZN(n6626) );
  AND2_X1 U9464 ( .A1(n11015), .A2(n11014), .ZN(n6627) );
  AND2_X1 U9465 ( .A1(n14020), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6628) );
  AND2_X1 U9466 ( .A1(n10882), .A2(n10881), .ZN(n6629) );
  OR2_X1 U9467 ( .A1(n15054), .A2(n15267), .ZN(n6630) );
  AND2_X1 U9468 ( .A1(n9967), .A2(n9968), .ZN(n6631) );
  NOR2_X1 U9469 ( .A1(n13084), .A2(n7032), .ZN(n6632) );
  AND2_X1 U9470 ( .A1(n11472), .A2(n13116), .ZN(n6633) );
  NAND2_X1 U9471 ( .A1(n14261), .A2(n8607), .ZN(n14239) );
  NAND2_X1 U9472 ( .A1(n7311), .A2(n12302), .ZN(n15278) );
  OAI21_X1 U9473 ( .B1(n13470), .B2(n6951), .A(n6950), .ZN(n13416) );
  NAND2_X1 U9474 ( .A1(n7993), .A2(n6851), .ZN(n14686) );
  NAND2_X1 U9475 ( .A1(n8248), .A2(n8247), .ZN(n14274) );
  OR2_X1 U9476 ( .A1(n13629), .A2(n13375), .ZN(n6634) );
  NAND2_X1 U9477 ( .A1(n8618), .A2(n9014), .ZN(n14221) );
  NAND2_X1 U9478 ( .A1(n15157), .A2(n12418), .ZN(n15141) );
  NAND2_X1 U9479 ( .A1(n8593), .A2(n7523), .ZN(n14271) );
  NAND2_X1 U9480 ( .A1(n10901), .A2(n10900), .ZN(n12699) );
  INV_X1 U9481 ( .A(n12699), .ZN(n7470) );
  INV_X1 U9482 ( .A(n13404), .ZN(n13407) );
  INV_X1 U9483 ( .A(n12880), .ZN(n12063) );
  AND2_X1 U9484 ( .A1(n9110), .A2(n7394), .ZN(n6635) );
  AND2_X1 U9485 ( .A1(n12993), .A2(n6632), .ZN(n6636) );
  AND2_X1 U9486 ( .A1(n6894), .A2(n7707), .ZN(n6637) );
  NAND2_X1 U9487 ( .A1(n8333), .A2(n8332), .ZN(n14146) );
  INV_X1 U9488 ( .A(n14146), .ZN(n14534) );
  AND2_X1 U9489 ( .A1(n9615), .A2(n9616), .ZN(n9775) );
  NAND2_X1 U9490 ( .A1(n8654), .A2(n8653), .ZN(n13935) );
  INV_X1 U9491 ( .A(n13935), .ZN(n13731) );
  AND4_X1 U9492 ( .A1(n11688), .A2(n9012), .A3(n11656), .A4(n11992), .ZN(n6638) );
  AND2_X1 U9493 ( .A1(n11683), .A2(n13951), .ZN(n6639) );
  INV_X1 U9494 ( .A(n8909), .ZN(n7865) );
  NAND2_X1 U9495 ( .A1(n7137), .A2(n7992), .ZN(n14733) );
  AND2_X1 U9496 ( .A1(n14469), .A2(n13918), .ZN(n6640) );
  AND2_X1 U9497 ( .A1(n7666), .A2(n6604), .ZN(n6641) );
  NAND2_X1 U9498 ( .A1(n15150), .A2(n12271), .ZN(n15125) );
  NAND2_X1 U9499 ( .A1(n12528), .A2(n12527), .ZN(n6642) );
  AND2_X1 U9500 ( .A1(n7956), .A2(n15029), .ZN(n6643) );
  AND2_X1 U9501 ( .A1(n15386), .A2(n7185), .ZN(n6644) );
  NAND2_X1 U9502 ( .A1(n13629), .A2(n13353), .ZN(n9683) );
  OR2_X1 U9503 ( .A1(n14451), .A2(n13938), .ZN(n6645) );
  AND3_X1 U9504 ( .A1(n11779), .A2(n9622), .A3(n9623), .ZN(n6646) );
  INV_X1 U9505 ( .A(n7504), .ZN(n6877) );
  AND2_X1 U9506 ( .A1(n14859), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7504) );
  AND3_X1 U9507 ( .A1(n9148), .A2(n9147), .A3(n9149), .ZN(n6647) );
  INV_X1 U9508 ( .A(n13544), .ZN(n7443) );
  AND2_X1 U9509 ( .A1(n8276), .A2(n8275), .ZN(n14251) );
  INV_X1 U9510 ( .A(n14251), .ZN(n14456) );
  NAND2_X1 U9511 ( .A1(n7531), .A2(n7535), .ZN(n14187) );
  INV_X1 U9512 ( .A(n7568), .ZN(n7567) );
  OAI21_X1 U9513 ( .B1(n9977), .B2(n10776), .A(n10962), .ZN(n7568) );
  INV_X1 U9514 ( .A(n13355), .ZN(n7720) );
  AND2_X1 U9515 ( .A1(n11857), .A2(n11856), .ZN(n6648) );
  OR2_X1 U9516 ( .A1(n9802), .A2(n13353), .ZN(n6649) );
  OR2_X1 U9517 ( .A1(n13649), .A2(n13106), .ZN(n6650) );
  INV_X1 U9518 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6809) );
  AND2_X1 U9519 ( .A1(n12398), .A2(n12397), .ZN(n14947) );
  INV_X1 U9520 ( .A(n14947), .ZN(n15220) );
  NOR2_X1 U9521 ( .A1(n7520), .A2(n14514), .ZN(n6651) );
  INV_X1 U9522 ( .A(n15253), .ZN(n15016) );
  NAND2_X1 U9523 ( .A1(n12362), .A2(n12361), .ZN(n15253) );
  AND2_X1 U9524 ( .A1(n14530), .A2(n8746), .ZN(n6652) );
  INV_X1 U9525 ( .A(n11383), .ZN(n7732) );
  NOR2_X1 U9526 ( .A1(n13345), .A2(n13610), .ZN(n6653) );
  NOR2_X1 U9527 ( .A1(n13345), .A2(n13688), .ZN(n6654) );
  AND2_X1 U9528 ( .A1(n15166), .A2(n12760), .ZN(n6655) );
  OR2_X1 U9529 ( .A1(n9436), .A2(n11054), .ZN(n6656) );
  AND2_X1 U9530 ( .A1(n14876), .A2(n7084), .ZN(n6657) );
  NAND2_X1 U9531 ( .A1(n7674), .A2(n7677), .ZN(n7676) );
  OR2_X1 U9532 ( .A1(n9662), .A2(n7437), .ZN(n6658) );
  AND2_X1 U9533 ( .A1(n14158), .A2(n8725), .ZN(n6659) );
  AND2_X1 U9534 ( .A1(n9705), .A2(n13454), .ZN(n9649) );
  OR2_X1 U9535 ( .A1(n14619), .A2(n14774), .ZN(n6660) );
  INV_X1 U9536 ( .A(n12418), .ZN(n7232) );
  OR2_X1 U9537 ( .A1(n7929), .A2(n6969), .ZN(n6661) );
  INV_X1 U9538 ( .A(n10902), .ZN(n12161) );
  INV_X1 U9539 ( .A(n8005), .ZN(n8004) );
  NAND2_X1 U9540 ( .A1(n8006), .A2(n11867), .ZN(n8005) );
  AND2_X1 U9541 ( .A1(n12518), .A2(n12516), .ZN(n6662) );
  NAND3_X1 U9542 ( .A1(n8902), .A2(n8901), .A3(n8900), .ZN(n6663) );
  AND2_X1 U9543 ( .A1(n12339), .A2(n12338), .ZN(n15037) );
  INV_X1 U9544 ( .A(n15037), .ZN(n7957) );
  OR2_X1 U9545 ( .A1(n10656), .A2(n7077), .ZN(n6664) );
  INV_X1 U9546 ( .A(n6625), .ZN(n7903) );
  AND2_X1 U9547 ( .A1(n8365), .A2(n8364), .ZN(n14526) );
  AND2_X1 U9548 ( .A1(n7963), .A2(n6941), .ZN(n6665) );
  AND2_X1 U9549 ( .A1(n8032), .A2(n8025), .ZN(n6666) );
  INV_X1 U9550 ( .A(n9637), .ZN(n7933) );
  NOR2_X1 U9551 ( .A1(n12800), .A2(n12801), .ZN(n7602) );
  AND2_X1 U9552 ( .A1(n7600), .A2(n6605), .ZN(n6667) );
  AND2_X1 U9553 ( .A1(n12352), .A2(n12351), .ZN(n15245) );
  INV_X1 U9554 ( .A(n15245), .ZN(n12678) );
  INV_X1 U9555 ( .A(n7373), .ZN(n7372) );
  NAND2_X1 U9556 ( .A1(n6678), .A2(n13850), .ZN(n7373) );
  NOR2_X1 U9557 ( .A1(n15319), .A2(n15181), .ZN(n6668) );
  NOR2_X1 U9558 ( .A1(n14146), .A2(n13933), .ZN(n6669) );
  NOR2_X1 U9559 ( .A1(n15294), .A2(n14777), .ZN(n6670) );
  NOR2_X1 U9560 ( .A1(n14687), .A2(n14688), .ZN(n6671) );
  NOR2_X1 U9561 ( .A1(n15253), .A2(n14773), .ZN(n6672) );
  INV_X1 U9562 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11518) );
  INV_X1 U9563 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n11448) );
  INV_X1 U9564 ( .A(n6563), .ZN(n7595) );
  INV_X1 U9565 ( .A(n7547), .ZN(n7546) );
  OR2_X1 U9566 ( .A1(n8548), .A2(n7548), .ZN(n7547) );
  INV_X1 U9567 ( .A(n7083), .ZN(n7082) );
  NOR2_X1 U9568 ( .A1(n11114), .A2(n11115), .ZN(n7083) );
  OR2_X1 U9569 ( .A1(n14414), .A2(n8764), .ZN(n6673) );
  INV_X1 U9570 ( .A(n13515), .ZN(n6888) );
  INV_X1 U9571 ( .A(n8213), .ZN(n6835) );
  NAND2_X1 U9572 ( .A1(n7647), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n6674) );
  AND2_X1 U9573 ( .A1(n13431), .A2(n9661), .ZN(n6675) );
  INV_X1 U9574 ( .A(n13530), .ZN(n13527) );
  AND2_X1 U9575 ( .A1(n9632), .A2(n9639), .ZN(n13530) );
  AND2_X1 U9576 ( .A1(n14167), .A2(n13934), .ZN(n6676) );
  OR2_X1 U9577 ( .A1(n14548), .A2(n13937), .ZN(n6677) );
  INV_X1 U9578 ( .A(n14548), .ZN(n14214) );
  INV_X1 U9579 ( .A(n8010), .ZN(n7785) );
  NAND2_X1 U9580 ( .A1(n7194), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n10144) );
  NAND2_X1 U9581 ( .A1(n13454), .A2(n9655), .ZN(n13473) );
  NAND2_X1 U9582 ( .A1(n15163), .A2(n12757), .ZN(n15193) );
  INV_X1 U9583 ( .A(n15193), .ZN(n15185) );
  AND2_X1 U9584 ( .A1(n12663), .A2(n12662), .ZN(n6678) );
  AND2_X1 U9585 ( .A1(n10194), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n6679) );
  AND2_X1 U9586 ( .A1(n8064), .A2(SI_9_), .ZN(n6680) );
  AND2_X1 U9587 ( .A1(n12992), .A2(n13089), .ZN(n6681) );
  AND2_X1 U9588 ( .A1(n14274), .A2(n13941), .ZN(n6682) );
  INV_X1 U9589 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10076) );
  INV_X1 U9590 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10119) );
  INV_X1 U9591 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10084) );
  INV_X1 U9592 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10890) );
  INV_X1 U9593 ( .A(n7162), .ZN(n7161) );
  OAI21_X1 U9594 ( .B1(n8765), .B2(n6580), .A(n6673), .ZN(n7162) );
  NAND2_X1 U9595 ( .A1(n10991), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n6683) );
  AND2_X1 U9596 ( .A1(n9563), .A2(n9562), .ZN(n6684) );
  AND2_X1 U9597 ( .A1(n7575), .A2(n7573), .ZN(n6685) );
  AND2_X1 U9598 ( .A1(n12599), .A2(n12598), .ZN(n6686) );
  AND2_X1 U9599 ( .A1(n10084), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6687) );
  AND2_X1 U9600 ( .A1(n11070), .A2(n11802), .ZN(n6688) );
  NAND2_X1 U9601 ( .A1(n14357), .A2(n13864), .ZN(n6689) );
  INV_X1 U9602 ( .A(n14182), .ZN(n14541) );
  NAND2_X1 U9603 ( .A1(n7991), .A2(n7990), .ZN(n14655) );
  INV_X1 U9604 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10095) );
  AND2_X1 U9605 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6690) );
  INV_X1 U9606 ( .A(n9015), .ZN(n14191) );
  AND2_X1 U9607 ( .A1(n13471), .A2(n13473), .ZN(n6691) );
  NAND2_X1 U9608 ( .A1(n7365), .A2(n7366), .ZN(n6692) );
  AND2_X1 U9609 ( .A1(n7414), .A2(n9754), .ZN(n6693) );
  AND2_X1 U9610 ( .A1(n7634), .A2(n12935), .ZN(n6694) );
  INV_X1 U9611 ( .A(n6981), .ZN(n6980) );
  NOR2_X1 U9612 ( .A1(n11554), .A2(n11568), .ZN(n6981) );
  AND2_X1 U9613 ( .A1(n13636), .A2(n13386), .ZN(n6695) );
  NAND2_X1 U9614 ( .A1(n7345), .A2(n8193), .ZN(n13887) );
  INV_X1 U9615 ( .A(n13887), .ZN(n14570) );
  INV_X1 U9616 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10256) );
  INV_X1 U9617 ( .A(n12386), .ZN(n6947) );
  AND2_X1 U9618 ( .A1(n15236), .A2(n14990), .ZN(n12386) );
  XNOR2_X1 U9619 ( .A(n15278), .B(n15090), .ZN(n12781) );
  INV_X1 U9620 ( .A(n12781), .ZN(n15075) );
  AND2_X1 U9621 ( .A1(n7447), .A2(n8250), .ZN(n6696) );
  NAND2_X1 U9622 ( .A1(n12140), .A2(n12123), .ZN(n6697) );
  AND2_X1 U9623 ( .A1(n14130), .A2(n8746), .ZN(n6698) );
  INV_X1 U9624 ( .A(n7838), .ZN(n7835) );
  NAND2_X1 U9625 ( .A1(n8851), .A2(n8850), .ZN(n7838) );
  XNOR2_X1 U9626 ( .A(n12819), .B(n14768), .ZN(n12895) );
  OR2_X1 U9627 ( .A1(n7835), .A2(n7836), .ZN(n6699) );
  AND2_X1 U9628 ( .A1(n7554), .A2(n7553), .ZN(n6700) );
  OR2_X1 U9629 ( .A1(n14469), .A2(n13918), .ZN(n6701) );
  INV_X1 U9630 ( .A(n9633), .ZN(n7935) );
  NAND2_X1 U9631 ( .A1(n12996), .A2(n7724), .ZN(n7723) );
  INV_X1 U9632 ( .A(n7723), .ZN(n7722) );
  AND2_X1 U9633 ( .A1(n13306), .A2(n13307), .ZN(n6702) );
  NAND2_X1 U9634 ( .A1(n9907), .A2(n9905), .ZN(n9900) );
  INV_X1 U9635 ( .A(n9900), .ZN(n7168) );
  AND2_X1 U9636 ( .A1(n7336), .A2(n6626), .ZN(n6703) );
  AND2_X1 U9637 ( .A1(n7481), .A2(n12782), .ZN(n6704) );
  NOR2_X1 U9638 ( .A1(n14093), .A2(n14338), .ZN(n6705) );
  OR2_X1 U9639 ( .A1(n12830), .A2(n12825), .ZN(n6706) );
  INV_X1 U9640 ( .A(n11361), .ZN(n7423) );
  AND2_X1 U9641 ( .A1(n7712), .A2(n7710), .ZN(n6707) );
  OR2_X1 U9642 ( .A1(n11073), .A2(n7692), .ZN(n6708) );
  NAND2_X1 U9643 ( .A1(n15048), .A2(n7956), .ZN(n15035) );
  BUF_X1 U9644 ( .A(n8465), .Z(n11717) );
  AND2_X1 U9645 ( .A1(n12247), .A2(n15163), .ZN(n6709) );
  AND2_X1 U9646 ( .A1(n7622), .A2(n11747), .ZN(n6710) );
  AND2_X1 U9647 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(n10254), .ZN(n6711) );
  NAND2_X1 U9648 ( .A1(n12919), .A2(n13550), .ZN(n6712) );
  AND2_X1 U9649 ( .A1(n12281), .A2(n12271), .ZN(n6713) );
  NAND2_X1 U9650 ( .A1(n12091), .A2(n12090), .ZN(n6714) );
  AND2_X1 U9651 ( .A1(n9014), .A2(n6645), .ZN(n6715) );
  OR2_X1 U9652 ( .A1(n12735), .A2(n12733), .ZN(n6716) );
  NAND2_X1 U9653 ( .A1(n8218), .A2(n8222), .ZN(n6717) );
  AND2_X1 U9654 ( .A1(n9706), .A2(n9650), .ZN(n6718) );
  OR2_X1 U9655 ( .A1(n12742), .A2(n12744), .ZN(n6719) );
  OR2_X1 U9656 ( .A1(n12723), .A2(n12721), .ZN(n6720) );
  OR2_X1 U9657 ( .A1(n12711), .A2(n12709), .ZN(n6721) );
  AND2_X1 U9658 ( .A1(n10216), .A2(n7146), .ZN(n6722) );
  INV_X1 U9659 ( .A(n6829), .ZN(n14166) );
  NOR2_X1 U9660 ( .A1(n14216), .A2(n6569), .ZN(n6829) );
  NOR2_X1 U9661 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n8090) );
  OR2_X1 U9662 ( .A1(n7612), .A2(n12743), .ZN(n6723) );
  INV_X1 U9663 ( .A(n9793), .ZN(n7716) );
  AND2_X1 U9664 ( .A1(n7352), .A2(n11383), .ZN(n6724) );
  AND2_X1 U9665 ( .A1(n7938), .A2(n9130), .ZN(n6725) );
  INV_X1 U9666 ( .A(n8475), .ZN(n7530) );
  AND2_X1 U9667 ( .A1(n7600), .A2(n7599), .ZN(n6726) );
  INV_X1 U9668 ( .A(n9695), .ZN(n9697) );
  OR2_X1 U9669 ( .A1(n13002), .A2(n13352), .ZN(n9695) );
  OR2_X1 U9670 ( .A1(n9774), .A2(n6633), .ZN(n6727) );
  INV_X1 U9671 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7146) );
  INV_X1 U9672 ( .A(n7369), .ZN(n7368) );
  NAND2_X1 U9673 ( .A1(n7370), .A2(n13726), .ZN(n7369) );
  OR2_X1 U9674 ( .A1(n7836), .A2(n7834), .ZN(n6728) );
  INV_X1 U9675 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8095) );
  INV_X1 U9676 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8386) );
  AND2_X1 U9677 ( .A1(n14222), .A2(n8724), .ZN(n6729) );
  INV_X1 U9678 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n9094) );
  AND2_X1 U9679 ( .A1(n9106), .A2(n9128), .ZN(n7938) );
  INV_X1 U9680 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7630) );
  AND2_X1 U9681 ( .A1(n8386), .A2(n6809), .ZN(n6730) );
  NAND2_X1 U9682 ( .A1(n14362), .A2(n14374), .ZN(n8539) );
  INV_X1 U9683 ( .A(n14298), .ZN(n7154) );
  INV_X1 U9684 ( .A(n15336), .ZN(n7488) );
  AND2_X2 U9685 ( .A1(n9860), .A2(n9859), .ZN(n15788) );
  XNOR2_X1 U9686 ( .A(n9310), .B(n9309), .ZN(n13153) );
  AND2_X1 U9687 ( .A1(n14337), .A2(n14564), .ZN(n14318) );
  NOR2_X1 U9688 ( .A1(n11986), .A2(n7508), .ZN(n14364) );
  NAND2_X1 U9689 ( .A1(n7763), .A2(n7765), .ZN(n11729) );
  NAND2_X1 U9690 ( .A1(n8198), .A2(n8102), .ZN(n8214) );
  NAND2_X1 U9691 ( .A1(n11806), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n11572) );
  NAND2_X1 U9692 ( .A1(n7527), .A2(n8496), .ZN(n11650) );
  NAND2_X1 U9693 ( .A1(n11190), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6731) );
  OR2_X1 U9694 ( .A1(n15203), .A2(n10350), .ZN(n15606) );
  INV_X1 U9695 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9030) );
  INV_X1 U9696 ( .A(n7170), .ZN(n11688) );
  NAND2_X1 U9697 ( .A1(n14371), .A2(n8705), .ZN(n7170) );
  INV_X1 U9698 ( .A(n7207), .ZN(n12045) );
  NAND2_X1 U9699 ( .A1(n6966), .A2(n6967), .ZN(n13484) );
  NAND2_X1 U9700 ( .A1(n11733), .A2(n8709), .ZN(n14347) );
  NAND2_X1 U9701 ( .A1(n7907), .A2(n9609), .ZN(n11417) );
  NAND2_X1 U9702 ( .A1(n7970), .A2(n11438), .ZN(n11854) );
  OR2_X1 U9703 ( .A1(n12999), .A2(n13535), .ZN(n6732) );
  NOR2_X1 U9704 ( .A1(n11958), .A2(n11661), .ZN(n6826) );
  INV_X1 U9705 ( .A(n14664), .ZN(n7978) );
  AND3_X1 U9706 ( .A1(n6582), .A2(n14318), .A3(n7512), .ZN(n14244) );
  NAND2_X1 U9707 ( .A1(n12074), .A2(n12886), .ZN(n12152) );
  AND2_X1 U9708 ( .A1(n6608), .A2(n6991), .ZN(n6733) );
  NAND2_X1 U9709 ( .A1(n12760), .A2(n12761), .ZN(n15164) );
  INV_X1 U9710 ( .A(n15164), .ZN(n7952) );
  NOR2_X1 U9711 ( .A1(n10652), .A2(n6907), .ZN(n6734) );
  INV_X1 U9712 ( .A(n7932), .ZN(n7931) );
  NAND2_X1 U9713 ( .A1(n7920), .A2(n9652), .ZN(n13468) );
  INV_X1 U9714 ( .A(n13752), .ZN(n14414) );
  NOR2_X1 U9715 ( .A1(n8557), .A2(n7544), .ZN(n7543) );
  INV_X1 U9716 ( .A(n7543), .ZN(n7539) );
  NAND2_X1 U9717 ( .A1(n7512), .A2(n14318), .ZN(n7515) );
  INV_X1 U9718 ( .A(n7587), .ZN(n7586) );
  AND2_X1 U9719 ( .A1(n6904), .A2(n6899), .ZN(n6735) );
  AND2_X1 U9720 ( .A1(n6865), .A2(n6868), .ZN(n6736) );
  AND2_X1 U9721 ( .A1(n9807), .A2(n6732), .ZN(n6737) );
  AND2_X1 U9722 ( .A1(n7881), .A2(n9072), .ZN(n6738) );
  AND2_X1 U9723 ( .A1(n6995), .A2(n6996), .ZN(n6739) );
  OR2_X1 U9724 ( .A1(n15493), .A2(n15494), .ZN(n6740) );
  AND3_X1 U9725 ( .A1(n9980), .A2(n9101), .A3(n7662), .ZN(n6741) );
  AND2_X1 U9726 ( .A1(n6607), .A2(n10820), .ZN(n6742) );
  NOR2_X1 U9727 ( .A1(n13174), .A2(n7588), .ZN(n6743) );
  INV_X1 U9728 ( .A(n8556), .ZN(n7542) );
  NOR2_X1 U9729 ( .A1(n12973), .A2(n13106), .ZN(n6744) );
  OR2_X1 U9730 ( .A1(n13140), .A2(n13133), .ZN(n6745) );
  AND2_X1 U9731 ( .A1(n11256), .A2(n11255), .ZN(n6746) );
  AND2_X1 U9732 ( .A1(n7396), .A2(n7395), .ZN(n6747) );
  INV_X1 U9733 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n15910) );
  OR2_X1 U9734 ( .A1(n13685), .A2(n13536), .ZN(n9638) );
  INV_X1 U9735 ( .A(n11683), .ZN(n7511) );
  OR2_X1 U9736 ( .A1(n15203), .A2(n15202), .ZN(n15620) );
  INV_X1 U9737 ( .A(n15484), .ZN(n7502) );
  INV_X1 U9738 ( .A(n11661), .ZN(n6823) );
  AND2_X1 U9739 ( .A1(n14887), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7492) );
  NAND2_X1 U9740 ( .A1(n14835), .A2(n6734), .ZN(n6906) );
  INV_X1 U9741 ( .A(n7081), .ZN(n7080) );
  AND2_X2 U9742 ( .A1(n9886), .A2(n9845), .ZN(n15804) );
  NAND2_X1 U9743 ( .A1(n10789), .A2(n8475), .ZN(n11954) );
  OR2_X1 U9744 ( .A1(n10822), .A2(n10821), .ZN(n6748) );
  NAND2_X1 U9745 ( .A1(n8467), .A2(n8466), .ZN(n10788) );
  AND2_X1 U9746 ( .A1(n9805), .A2(n9849), .ZN(n13502) );
  AND2_X1 U9747 ( .A1(n7561), .A2(n7565), .ZN(n6749) );
  AND2_X1 U9748 ( .A1(n11072), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n6750) );
  AND2_X1 U9749 ( .A1(n6870), .A2(n12258), .ZN(n6751) );
  INV_X1 U9750 ( .A(n7492), .ZN(n6870) );
  INV_X1 U9751 ( .A(n13291), .ZN(n7702) );
  AND2_X1 U9752 ( .A1(n14065), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6752) );
  AND2_X1 U9753 ( .A1(n13148), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n6753) );
  AND2_X1 U9754 ( .A1(n13249), .A2(n7672), .ZN(n6754) );
  NAND2_X1 U9755 ( .A1(n9085), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6755) );
  AND2_X1 U9756 ( .A1(n6998), .A2(n6999), .ZN(n6756) );
  INV_X1 U9757 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n7390) );
  INV_X1 U9758 ( .A(n11020), .ZN(n7500) );
  INV_X1 U9759 ( .A(n8775), .ZN(n14086) );
  INV_X1 U9760 ( .A(n11283), .ZN(n9010) );
  AND2_X1 U9761 ( .A1(n9002), .A2(n8773), .ZN(n6757) );
  AND2_X1 U9762 ( .A1(n12462), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6758) );
  INV_X1 U9763 ( .A(n12672), .ZN(n15819) );
  NOR2_X1 U9764 ( .A1(n10269), .A2(n6874), .ZN(n6759) );
  AND2_X1 U9765 ( .A1(n10165), .A2(n10603), .ZN(n6760) );
  OR2_X1 U9766 ( .A1(n6757), .A2(n11741), .ZN(n6761) );
  INV_X1 U9767 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n7675) );
  INV_X1 U9768 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7499) );
  OR2_X1 U9769 ( .A1(n10955), .A2(n10965), .ZN(n7693) );
  NAND2_X1 U9770 ( .A1(n10955), .A2(n10965), .ZN(n11072) );
  NOR2_X1 U9771 ( .A1(n10965), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7692) );
  NAND2_X1 U9772 ( .A1(n11508), .A2(n11507), .ZN(n15506) );
  NAND2_X1 U9773 ( .A1(n7225), .A2(n7226), .ZN(n15099) );
  NAND2_X1 U9774 ( .A1(n12431), .A2(n12430), .ZN(n15034) );
  NAND2_X1 U9775 ( .A1(n11157), .A2(n11156), .ZN(n11185) );
  NAND2_X1 U9776 ( .A1(n7212), .A2(n11509), .ZN(n12058) );
  NAND2_X1 U9777 ( .A1(n11152), .A2(n11151), .ZN(n11348) );
  BUF_X2 U9778 ( .A(n11032), .Z(n12410) );
  INV_X1 U9779 ( .A(n10700), .ZN(n11032) );
  NAND2_X2 U9780 ( .A1(n15194), .A2(n15193), .ZN(n15192) );
  INV_X1 U9781 ( .A(n12092), .ZN(n7219) );
  NAND2_X1 U9782 ( .A1(n6763), .A2(n14922), .ZN(n15207) );
  OR2_X1 U9783 ( .A1(n14937), .A2(n15210), .ZN(n6763) );
  NAND2_X1 U9784 ( .A1(n11349), .A2(n15548), .ZN(n11351) );
  NAND2_X1 U9785 ( .A1(n8043), .A2(n8042), .ZN(n8113) );
  INV_X1 U9786 ( .A(n7448), .ZN(n8249) );
  INV_X1 U9787 ( .A(n7375), .ZN(n7374) );
  INV_X1 U9788 ( .A(n7382), .ZN(n7379) );
  AND2_X1 U9789 ( .A1(n12891), .A2(n7281), .ZN(n12892) );
  NOR2_X1 U9790 ( .A1(n13767), .A2(n8018), .ZN(n13766) );
  NAND2_X1 U9791 ( .A1(n8048), .A2(n7006), .ZN(n8141) );
  NAND2_X1 U9792 ( .A1(n7802), .A2(n8071), .ZN(n8194) );
  XNOR2_X1 U9793 ( .A(n7279), .B(n15819), .ZN(n12908) );
  NAND3_X1 U9794 ( .A1(n6764), .A2(n7183), .A3(n7186), .ZN(n15387) );
  NAND2_X1 U9795 ( .A1(n7181), .A2(n7182), .ZN(n6764) );
  NAND2_X1 U9796 ( .A1(n7198), .A2(n7201), .ZN(n7197) );
  NAND2_X1 U9797 ( .A1(n7660), .A2(n7659), .ZN(n11669) );
  NAND2_X1 U9798 ( .A1(n10125), .A2(n7195), .ZN(n10145) );
  NAND2_X1 U9799 ( .A1(n12038), .A2(n7206), .ZN(n7207) );
  NAND3_X1 U9800 ( .A1(n7657), .A2(n15428), .A3(n15420), .ZN(n15433) );
  NAND2_X1 U9801 ( .A1(n14164), .A2(n14163), .ZN(n6765) );
  NAND2_X1 U9802 ( .A1(n8113), .A2(n8114), .ZN(n7008) );
  OAI21_X1 U9803 ( .B1(n11651), .B2(n11656), .A(n7180), .ZN(n7179) );
  INV_X1 U9804 ( .A(n7050), .ZN(n7049) );
  OR2_X1 U9805 ( .A1(n10663), .A2(n8121), .ZN(n6818) );
  NAND2_X1 U9806 ( .A1(n6766), .A2(n7829), .ZN(n7828) );
  NAND3_X1 U9807 ( .A1(n8846), .A2(n8874), .A3(n7830), .ZN(n6766) );
  NAND2_X1 U9808 ( .A1(n8792), .A2(n8791), .ZN(n6767) );
  OR3_X2 U9809 ( .A1(n8829), .A2(n8832), .A3(n7839), .ZN(n6769) );
  OR2_X2 U9810 ( .A1(n8808), .A2(n8807), .ZN(n8813) );
  NAND2_X1 U9811 ( .A1(n8820), .A2(n8819), .ZN(n6773) );
  NAND2_X1 U9812 ( .A1(n6770), .A2(n6771), .ZN(n7858) );
  OAI21_X1 U9813 ( .B1(n8929), .B2(n8928), .A(n8927), .ZN(n8943) );
  AOI21_X1 U9814 ( .B1(n8921), .B2(n8781), .A(n8780), .ZN(n8794) );
  AOI21_X1 U9815 ( .B1(n8843), .B2(n8842), .A(n8841), .ZN(n8846) );
  NAND2_X1 U9816 ( .A1(n6767), .A2(n8797), .ZN(n7823) );
  NOR2_X1 U9817 ( .A1(n7828), .A2(n6663), .ZN(n8905) );
  OR2_X1 U9818 ( .A1(n8820), .A2(n8819), .ZN(n6770) );
  NAND2_X1 U9819 ( .A1(n9050), .A2(n9049), .ZN(n9322) );
  NAND2_X1 U9820 ( .A1(n9692), .A2(n9691), .ZN(n7414) );
  NAND2_X1 U9821 ( .A1(n12054), .A2(n9550), .ZN(n7869) );
  INV_X1 U9822 ( .A(n6955), .ZN(n6954) );
  AND2_X1 U9823 ( .A1(n10518), .A2(n10519), .ZN(n10524) );
  NAND2_X1 U9824 ( .A1(n7308), .A2(n7252), .ZN(n10529) );
  NAND2_X1 U9825 ( .A1(n7051), .A2(n12921), .ZN(n13055) );
  OAI21_X1 U9826 ( .B1(n9725), .B2(n11052), .A(n9724), .ZN(n6955) );
  NAND2_X1 U9827 ( .A1(n7124), .A2(n9081), .ZN(n9517) );
  INV_X1 U9828 ( .A(n8019), .ZN(n7797) );
  XNOR2_X1 U9829 ( .A(n8263), .B(n8262), .ZN(n12293) );
  OAI211_X1 U9830 ( .C1(n7593), .C2(n7591), .A(n7324), .B(n7323), .ZN(n12793)
         );
  OAI21_X1 U9831 ( .B1(n12854), .B2(n6706), .A(n7322), .ZN(n7452) );
  NAND3_X1 U9832 ( .A1(n13308), .A2(n13309), .A3(n6702), .ZN(P3_U3200) );
  INV_X1 U9833 ( .A(n13267), .ZN(n7687) );
  AOI21_X1 U9834 ( .B1(n7691), .B2(n6602), .A(n6708), .ZN(n11567) );
  NAND2_X1 U9835 ( .A1(n7683), .A2(n10739), .ZN(n7682) );
  XNOR2_X1 U9836 ( .A(n13185), .B(n13207), .ZN(n13186) );
  NAND2_X1 U9837 ( .A1(n7696), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7695) );
  NAND2_X1 U9838 ( .A1(n7682), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7681) );
  NAND2_X1 U9839 ( .A1(n7271), .A2(n10977), .ZN(n10982) );
  INV_X1 U9840 ( .A(n10955), .ZN(n7691) );
  INV_X1 U9841 ( .A(n9984), .ZN(n7683) );
  AOI21_X1 U9842 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n11568), .A(n11567), .ZN(
        n11570) );
  NOR2_X1 U9843 ( .A1(n13161), .A2(n13126), .ZN(n13127) );
  NAND2_X1 U9844 ( .A1(n7688), .A2(n7690), .ZN(n7684) );
  NAND2_X1 U9845 ( .A1(n7317), .A2(n8062), .ZN(n8175) );
  NOR2_X1 U9846 ( .A1(n6815), .A2(n14100), .ZN(n9927) );
  INV_X1 U9847 ( .A(n7156), .ZN(n9902) );
  NAND2_X1 U9848 ( .A1(n14099), .A2(n15740), .ZN(n6817) );
  NAND2_X1 U9849 ( .A1(n9062), .A2(n9061), .ZN(n9382) );
  NAND2_X1 U9850 ( .A1(n7866), .A2(n9065), .ZN(n9412) );
  NAND2_X1 U9851 ( .A1(n9154), .A2(n9153), .ZN(n9152) );
  INV_X1 U9852 ( .A(n9687), .ZN(n9688) );
  NAND2_X1 U9853 ( .A1(n7413), .A2(n7414), .ZN(n7416) );
  NAND2_X1 U9854 ( .A1(n13355), .A2(n9688), .ZN(n9692) );
  NAND2_X1 U9855 ( .A1(n7412), .A2(n7417), .ZN(n7411) );
  NAND2_X1 U9856 ( .A1(n7947), .A2(n7951), .ZN(n7332) );
  NAND2_X1 U9857 ( .A1(n7094), .A2(n9063), .ZN(n9400) );
  NAND2_X1 U9858 ( .A1(n6776), .A2(n7432), .ZN(n9669) );
  AOI21_X1 U9859 ( .B1(n7433), .B2(n6658), .A(n7439), .ZN(n6776) );
  NAND2_X1 U9860 ( .A1(n6953), .A2(n9731), .ZN(n9752) );
  NAND2_X1 U9861 ( .A1(n7093), .A2(n9029), .ZN(n9163) );
  INV_X1 U9862 ( .A(n6939), .ZN(n6938) );
  NAND2_X1 U9863 ( .A1(n7176), .A2(n7177), .ZN(n14263) );
  NAND2_X1 U9864 ( .A1(n7155), .A2(n6700), .ZN(n7549) );
  NAND2_X1 U9865 ( .A1(n7178), .A2(n8526), .ZN(n14362) );
  NOR2_X1 U9866 ( .A1(n14415), .A2(n7340), .ZN(n14527) );
  NAND2_X1 U9867 ( .A1(n14417), .A2(n15740), .ZN(n7342) );
  INV_X1 U9868 ( .A(n6778), .ZN(n12363) );
  NAND2_X1 U9869 ( .A1(n6778), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n12365) );
  NAND2_X1 U9870 ( .A1(n12315), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n12330) );
  NAND2_X1 U9871 ( .A1(n11882), .A2(n6609), .ZN(n6786) );
  NAND3_X1 U9872 ( .A1(n6795), .A2(n6791), .A3(n6789), .ZN(P2_U3233) );
  NAND2_X1 U9873 ( .A1(n14001), .A2(n6805), .ZN(n6802) );
  NAND2_X1 U9874 ( .A1(n6802), .A2(n6803), .ZN(n14030) );
  MUX2_X1 U9875 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n10415), .S(n10433), .Z(
        n15631) );
  OAI211_X2 U9876 ( .C1(n9030), .C2(n8376), .A(n6818), .B(n8110), .ZN(n7528)
         );
  NAND2_X1 U9877 ( .A1(n14504), .A2(n6823), .ZN(n6822) );
  INV_X1 U9878 ( .A(n6826), .ZN(n11986) );
  NAND4_X1 U9879 ( .A1(n6582), .A2(n14318), .A3(n7512), .A4(n14251), .ZN(
        n14229) );
  NAND4_X1 U9880 ( .A1(n6582), .A2(n14318), .A3(n7512), .A4(n6827), .ZN(n14230) );
  NAND2_X1 U9881 ( .A1(n6833), .A2(n6832), .ZN(n6831) );
  NAND2_X1 U9882 ( .A1(n8210), .A2(n6838), .ZN(n6832) );
  NAND2_X1 U9883 ( .A1(n6836), .A2(n6835), .ZN(n6833) );
  NAND2_X1 U9884 ( .A1(n8210), .A2(n6835), .ZN(n6834) );
  INV_X1 U9885 ( .A(n8210), .ZN(n6836) );
  OAI21_X1 U9886 ( .B1(n12550), .B2(n6844), .A(n6617), .ZN(n14666) );
  NAND2_X1 U9887 ( .A1(n12550), .A2(n6617), .ZN(n6841) );
  OAI21_X1 U9888 ( .B1(n7316), .B2(n8184), .A(n8067), .ZN(n6849) );
  NAND2_X2 U9889 ( .A1(n6847), .A2(n6848), .ZN(n8190) );
  NAND3_X1 U9890 ( .A1(n7318), .A2(n8167), .A3(n8065), .ZN(n6847) );
  NAND3_X1 U9891 ( .A1(n7137), .A2(n12511), .A3(n7992), .ZN(n14734) );
  NAND2_X1 U9892 ( .A1(n6852), .A2(n7745), .ZN(n11844) );
  NAND2_X1 U9893 ( .A1(n6857), .A2(n6856), .ZN(n6852) );
  OAI211_X1 U9894 ( .C1(n6857), .C2(n6855), .A(n9780), .B(n6853), .ZN(n9782)
         );
  NAND2_X1 U9895 ( .A1(n6854), .A2(n7745), .ZN(n6853) );
  INV_X1 U9896 ( .A(n7745), .ZN(n6855) );
  NAND3_X1 U9897 ( .A1(n6864), .A2(n6862), .A3(n6859), .ZN(n7491) );
  NAND3_X1 U9898 ( .A1(n6873), .A2(n6872), .A3(n6871), .ZN(n10319) );
  NAND2_X1 U9899 ( .A1(n10269), .A2(n6731), .ZN(n6871) );
  NAND3_X1 U9900 ( .A1(n6568), .A2(n6731), .A3(n10235), .ZN(n6872) );
  INV_X2 U9901 ( .A(n13121), .ZN(n7429) );
  NAND2_X1 U9902 ( .A1(n11477), .A2(n6881), .ZN(n11478) );
  INV_X1 U9903 ( .A(n6878), .ZN(n14853) );
  NOR2_X1 U9904 ( .A1(n11479), .A2(n6880), .ZN(n6879) );
  INV_X1 U9905 ( .A(n6881), .ZN(n6880) );
  NAND2_X1 U9906 ( .A1(n12105), .A2(n6887), .ZN(n6883) );
  NAND2_X1 U9907 ( .A1(n6886), .A2(n6887), .ZN(n13518) );
  INV_X1 U9908 ( .A(n7707), .ZN(n6892) );
  NAND3_X1 U9909 ( .A1(n13403), .A2(n6634), .A3(n6895), .ZN(n6893) );
  AND3_X2 U9910 ( .A1(n9736), .A2(n9569), .A3(n7260), .ZN(n6972) );
  NAND4_X1 U9911 ( .A1(n9736), .A2(n9569), .A3(n7260), .A4(n7938), .ZN(n6896)
         );
  INV_X1 U9912 ( .A(n14905), .ZN(n6899) );
  INV_X1 U9913 ( .A(n15805), .ZN(n6904) );
  NAND2_X1 U9914 ( .A1(n6906), .A2(n6742), .ZN(n11118) );
  NAND2_X1 U9915 ( .A1(n14835), .A2(n7501), .ZN(n10651) );
  INV_X1 U9916 ( .A(n6906), .ZN(n10818) );
  INV_X1 U9917 ( .A(n7501), .ZN(n6907) );
  NAND2_X1 U9918 ( .A1(n6908), .A2(n10050), .ZN(n10088) );
  NAND2_X1 U9919 ( .A1(n6909), .A2(n12916), .ZN(P1_U3242) );
  NAND2_X1 U9920 ( .A1(n6910), .A2(n12911), .ZN(n6909) );
  OAI211_X1 U9921 ( .C1(n7452), .C2(n12865), .A(n6911), .B(n12910), .ZN(n6910)
         );
  NAND2_X1 U9922 ( .A1(n7452), .A2(n12867), .ZN(n6911) );
  NAND3_X1 U9923 ( .A1(n7603), .A2(n7604), .A3(n6923), .ZN(n6913) );
  NAND2_X1 U9924 ( .A1(n6912), .A2(n6915), .ZN(n6921) );
  NAND3_X1 U9925 ( .A1(n7603), .A2(n6918), .A3(n7604), .ZN(n6912) );
  NAND2_X1 U9926 ( .A1(n6913), .A2(n6914), .ZN(n6920) );
  AND2_X1 U9927 ( .A1(n6921), .A2(n6920), .ZN(n12804) );
  INV_X1 U9928 ( .A(n7602), .ZN(n6923) );
  OR2_X1 U9929 ( .A1(n8225), .A2(n7450), .ZN(n6924) );
  NAND2_X1 U9930 ( .A1(n8225), .A2(n6564), .ZN(n6926) );
  NAND2_X1 U9931 ( .A1(n8225), .A2(n8224), .ZN(n8238) );
  MUX2_X1 U9932 ( .A(n9052), .B(n10286), .S(n8050), .Z(n8072) );
  NOR2_X2 U9933 ( .A1(n6931), .A2(n6930), .ZN(n7330) );
  NAND4_X1 U9934 ( .A1(n6933), .A2(n9932), .A3(n9931), .A4(n6932), .ZN(n6931)
         );
  NOR2_X2 U9935 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6933) );
  NAND2_X2 U9936 ( .A1(n15049), .A2(n15062), .ZN(n15048) );
  INV_X1 U9937 ( .A(n11317), .ZN(n6937) );
  OAI21_X1 U9938 ( .B1(n6579), .B2(n6940), .A(n6713), .ZN(n6939) );
  NAND2_X1 U9939 ( .A1(n15006), .A2(n8016), .ZN(n6948) );
  OAI22_X1 U9940 ( .A1(n14955), .A2(n6947), .B1(n14962), .B2(n14770), .ZN(
        n6946) );
  INV_X1 U9941 ( .A(n14955), .ZN(n6943) );
  NAND2_X1 U9942 ( .A1(n7923), .A2(n6718), .ZN(n6949) );
  NAND3_X1 U9943 ( .A1(n6956), .A2(n7269), .A3(n6954), .ZN(n6953) );
  NAND3_X1 U9944 ( .A1(n6957), .A2(n9580), .A3(n9579), .ZN(n6956) );
  NAND2_X1 U9945 ( .A1(n6958), .A2(n7905), .ZN(n11371) );
  NAND2_X1 U9946 ( .A1(n11400), .A2(n7908), .ZN(n6958) );
  NAND2_X1 U9947 ( .A1(n11360), .A2(n7423), .ZN(n6959) );
  NAND2_X1 U9948 ( .A1(n13410), .A2(n6963), .ZN(n6960) );
  NAND2_X1 U9949 ( .A1(n6960), .A2(n6961), .ZN(n13362) );
  AND2_X1 U9950 ( .A1(n7927), .A2(n6890), .ZN(n6965) );
  NAND2_X1 U9951 ( .A1(n12104), .A2(n6890), .ZN(n6970) );
  NAND3_X1 U9952 ( .A1(n6971), .A2(n6972), .A3(n6725), .ZN(n13707) );
  OAI21_X1 U9953 ( .B1(n10772), .B2(n7564), .A(n7562), .ZN(n11071) );
  NAND3_X1 U9954 ( .A1(n6977), .A2(n6976), .A3(n6688), .ZN(n6979) );
  NAND2_X1 U9955 ( .A1(n10772), .A2(n7562), .ZN(n6977) );
  XNOR2_X1 U9956 ( .A(n6982), .B(n10106), .ZN(n10743) );
  NAND2_X1 U9957 ( .A1(n6984), .A2(n6983), .ZN(n6982) );
  OAI211_X2 U9958 ( .C1(P3_IR_REG_1__SCAN_IN), .C2(P3_IR_REG_0__SCAN_IN), .A(
        n6986), .B(n6985), .ZN(n11102) );
  NAND3_X1 U9959 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n6985) );
  NAND3_X1 U9960 ( .A1(n6991), .A2(n11562), .A3(n6599), .ZN(n6989) );
  NAND2_X1 U9961 ( .A1(n11564), .A2(n11563), .ZN(n6990) );
  NAND3_X1 U9962 ( .A1(n6992), .A2(n6993), .A3(n13256), .ZN(n13224) );
  NAND2_X1 U9963 ( .A1(n7679), .A2(n7678), .ZN(n6993) );
  NAND3_X1 U9964 ( .A1(n6998), .A2(P3_REG1_REG_5__SCAN_IN), .A3(n6999), .ZN(
        n10778) );
  AOI21_X2 U9965 ( .B1(n7261), .B2(n11593), .A(n7619), .ZN(n11942) );
  NAND2_X2 U9966 ( .A1(n11272), .A2(n11273), .ZN(n11586) );
  NAND2_X1 U9967 ( .A1(n7000), .A2(n8038), .ZN(n10048) );
  INV_X1 U9968 ( .A(n8050), .ZN(n7000) );
  NAND2_X4 U9969 ( .A1(n7002), .A2(n7001), .ZN(n8050) );
  NAND2_X1 U9970 ( .A1(n7793), .A2(n7792), .ZN(n7001) );
  NAND2_X1 U9971 ( .A1(n7791), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n7002) );
  INV_X1 U9972 ( .A(n8046), .ZN(n7009) );
  NAND2_X1 U9973 ( .A1(n7007), .A2(n7008), .ZN(n7006) );
  NOR2_X1 U9974 ( .A1(n7009), .A2(n7469), .ZN(n7007) );
  NAND2_X1 U9975 ( .A1(n7008), .A2(n8046), .ZN(n7787) );
  XNOR2_X1 U9976 ( .A(n8044), .B(SI_2_), .ZN(n8114) );
  NAND2_X1 U9977 ( .A1(n7017), .A2(n7016), .ZN(n14190) );
  NAND2_X1 U9978 ( .A1(n14241), .A2(n7021), .ZN(n7016) );
  OAI22_X1 U9979 ( .A1(n7020), .A2(n14241), .B1(n6572), .B2(n7021), .ZN(n14156) );
  NAND2_X1 U9980 ( .A1(n13012), .A2(n7026), .ZN(n7022) );
  OAI211_X1 U9981 ( .C1(n13012), .C2(n7027), .A(n7023), .B(n7022), .ZN(n13004)
         );
  AOI21_X1 U9982 ( .B1(n13012), .B2(n13013), .A(n7033), .ZN(n13083) );
  NAND2_X1 U9983 ( .A1(n13012), .A2(n6632), .ZN(n7029) );
  INV_X1 U9984 ( .A(n12997), .ZN(n7035) );
  OAI211_X1 U9985 ( .C1(n14315), .C2(n7037), .A(n7039), .B(n6703), .ZN(n7044)
         );
  NAND2_X1 U9986 ( .A1(n11946), .A2(n7052), .ZN(n7051) );
  XNOR2_X1 U9987 ( .A(n7053), .B(n11947), .ZN(n11953) );
  AOI21_X1 U9988 ( .B1(n8707), .B2(n8706), .A(n7055), .ZN(n7054) );
  NAND2_X1 U9989 ( .A1(n7769), .A2(n7767), .ZN(n7056) );
  OAI21_X1 U9990 ( .B1(n12975), .B2(n6744), .A(n7246), .ZN(n12955) );
  OAI21_X2 U9991 ( .B1(n13005), .B2(n13006), .A(n12946), .ZN(n12975) );
  MUX2_X1 U9992 ( .A(n11140), .B(P1_REG2_REG_1__SCAN_IN), .S(n10666), .Z(
        n14799) );
  NAND2_X1 U9993 ( .A1(n7060), .A2(n7304), .ZN(n7059) );
  NAND2_X1 U9994 ( .A1(n7306), .A2(P1_IR_REG_1__SCAN_IN), .ZN(n7060) );
  NAND3_X1 U9995 ( .A1(n7066), .A2(n7067), .A3(n10292), .ZN(n7065) );
  AOI21_X1 U9996 ( .B1(n7080), .B2(n10656), .A(n7077), .ZN(n7073) );
  NAND2_X1 U9997 ( .A1(n14846), .A2(n7080), .ZN(n7074) );
  INV_X1 U9998 ( .A(n7076), .ZN(n7075) );
  NAND2_X1 U9999 ( .A1(n15481), .A2(n15480), .ZN(n15479) );
  NAND2_X1 U10000 ( .A1(n14890), .A2(n14889), .ZN(n14892) );
  NAND3_X1 U10001 ( .A1(n7276), .A2(n15814), .A3(n15813), .ZN(n7087) );
  NAND3_X1 U10002 ( .A1(n7775), .A2(n8093), .A3(n7774), .ZN(n8390) );
  AND3_X2 U10003 ( .A1(n7522), .A2(n7521), .A3(n8386), .ZN(n7774) );
  AND2_X2 U10004 ( .A1(n7277), .A2(n8099), .ZN(n7775) );
  NAND2_X1 U10005 ( .A1(n9400), .A2(n9064), .ZN(n7866) );
  NAND2_X1 U10006 ( .A1(n9382), .A2(n9380), .ZN(n7094) );
  NAND3_X1 U10007 ( .A1(n7098), .A2(n8485), .A3(n7529), .ZN(n7097) );
  NAND2_X1 U10008 ( .A1(n8467), .A2(n6600), .ZN(n7098) );
  NAND2_X1 U10009 ( .A1(n9274), .A2(n7105), .ZN(n7103) );
  NAND2_X1 U10010 ( .A1(n7103), .A2(n7104), .ZN(n9050) );
  NAND2_X1 U10011 ( .A1(n9274), .A2(n9046), .ZN(n9291) );
  NAND2_X1 U10012 ( .A1(n9219), .A2(n7115), .ZN(n7113) );
  NAND2_X1 U10013 ( .A1(n7113), .A2(n7114), .ZN(n9245) );
  NAND2_X4 U10014 ( .A1(n8111), .A2(n8097), .ZN(n8376) );
  XNOR2_X2 U10015 ( .A(n8096), .B(n8095), .ZN(n8398) );
  NAND2_X1 U10016 ( .A1(n7887), .A2(n9079), .ZN(n9506) );
  OAI21_X1 U10017 ( .B1(n11133), .B2(n10699), .A(n7129), .ZN(n10685) );
  NAND2_X1 U10018 ( .A1(n7135), .A2(n11017), .ZN(n7131) );
  INV_X1 U10019 ( .A(n11016), .ZN(n7136) );
  AOI21_X2 U10020 ( .B1(n11017), .B2(n11016), .A(n6627), .ZN(n11325) );
  NOR2_X1 U10021 ( .A1(n7136), .A2(n11324), .ZN(n7135) );
  NAND2_X1 U10022 ( .A1(n14744), .A2(n7139), .ZN(n7138) );
  OAI211_X1 U10023 ( .C1(n14744), .C2(n7141), .A(n7138), .B(n14753), .ZN(
        n12585) );
  NOR2_X1 U10024 ( .A1(n12579), .A2(n12577), .ZN(n7143) );
  NAND2_X1 U10025 ( .A1(n12579), .A2(n12577), .ZN(n7144) );
  INV_X1 U10026 ( .A(n12579), .ZN(n7145) );
  NAND2_X1 U10027 ( .A1(n7330), .A2(n10540), .ZN(n10642) );
  NAND3_X1 U10028 ( .A1(n7330), .A2(n10540), .A3(n10216), .ZN(n11103) );
  AND3_X2 U10029 ( .A1(n7330), .A2(n10541), .A3(n6722), .ZN(n9940) );
  NAND4_X1 U10030 ( .A1(n14287), .A2(n7151), .A3(n14348), .A4(n6638), .ZN(
        n7150) );
  OAI21_X1 U10031 ( .B1(n14127), .B2(n7159), .A(n7161), .ZN(n9901) );
  OAI21_X1 U10032 ( .B1(n14127), .B2(n7158), .A(n7157), .ZN(n7156) );
  NAND3_X1 U10033 ( .A1(n14136), .A2(n14142), .A3(n14163), .ZN(n7167) );
  NAND4_X1 U10034 ( .A1(n10792), .A2(n7172), .A3(n15661), .A4(n11706), .ZN(
        n7171) );
  INV_X1 U10035 ( .A(n14263), .ZN(n7175) );
  NAND2_X1 U10036 ( .A1(n14281), .A2(n7524), .ZN(n7176) );
  NAND2_X1 U10037 ( .A1(n8525), .A2(n7179), .ZN(n7178) );
  NAND2_X1 U10038 ( .A1(n7657), .A2(n15420), .ZN(n15430) );
  NAND2_X1 U10039 ( .A1(n15385), .A2(n15386), .ZN(n7188) );
  AOI22_X1 U10040 ( .A1(n15385), .A2(n6644), .B1(n10610), .B2(n7184), .ZN(
        n7183) );
  INV_X1 U10041 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7185) );
  NAND2_X1 U10042 ( .A1(n7188), .A2(n10610), .ZN(n10617) );
  NAND2_X1 U10043 ( .A1(n7187), .A2(n7185), .ZN(n7186) );
  INV_X1 U10044 ( .A(n10610), .ZN(n7187) );
  INV_X1 U10045 ( .A(n10130), .ZN(n7193) );
  NAND3_X1 U10046 ( .A1(n7649), .A2(n7647), .A3(n10131), .ZN(n10140) );
  INV_X1 U10047 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7194) );
  INV_X1 U10048 ( .A(n10144), .ZN(n7196) );
  NAND3_X1 U10049 ( .A1(n7196), .A2(n10125), .A3(n7195), .ZN(n10147) );
  NAND2_X1 U10050 ( .A1(n7641), .A2(n7640), .ZN(n7198) );
  NAND2_X1 U10051 ( .A1(n7200), .A2(n7201), .ZN(n7199) );
  INV_X1 U10052 ( .A(n15444), .ZN(n7200) );
  NAND3_X1 U10053 ( .A1(n15444), .A2(n7641), .A3(n7202), .ZN(n15454) );
  NAND2_X1 U10054 ( .A1(n7205), .A2(n10939), .ZN(n10946) );
  NAND2_X1 U10055 ( .A1(n12037), .A2(n14049), .ZN(n7206) );
  NAND3_X1 U10056 ( .A1(n11670), .A2(n11671), .A3(n7208), .ZN(n12037) );
  NAND2_X1 U10057 ( .A1(n7207), .A2(n6601), .ZN(n7654) );
  NAND2_X1 U10058 ( .A1(n7210), .A2(n11171), .ZN(n11152) );
  XNOR2_X1 U10059 ( .A(n7210), .B(n11171), .ZN(n15542) );
  NAND2_X1 U10060 ( .A1(n11150), .A2(n11149), .ZN(n7210) );
  NAND2_X1 U10061 ( .A1(n12058), .A2(n12063), .ZN(n7211) );
  NAND2_X1 U10062 ( .A1(n15506), .A2(n15508), .ZN(n7212) );
  NOR2_X1 U10063 ( .A1(n7214), .A2(n12443), .ZN(n7213) );
  NAND2_X1 U10064 ( .A1(n10255), .A2(n6711), .ZN(n7218) );
  OAI21_X1 U10065 ( .B1(n7220), .B2(n7219), .A(n7223), .ZN(n12178) );
  INV_X1 U10066 ( .A(n12095), .ZN(n7222) );
  NOR2_X1 U10067 ( .A1(n12095), .A2(n6565), .ZN(n7221) );
  INV_X1 U10068 ( .A(n15192), .ZN(n7229) );
  NAND2_X1 U10069 ( .A1(n6581), .A2(n15192), .ZN(n7225) );
  NAND2_X1 U10070 ( .A1(n15030), .A2(n7235), .ZN(n7234) );
  NAND2_X1 U10071 ( .A1(n15030), .A2(n7815), .ZN(n7240) );
  NAND3_X1 U10072 ( .A1(n7234), .A2(n7805), .A3(n7233), .ZN(n14956) );
  AND2_X2 U10073 ( .A1(n7240), .A2(n7238), .ZN(n15243) );
  NAND2_X1 U10074 ( .A1(n7242), .A2(n7241), .ZN(P1_U3557) );
  NAND2_X1 U10075 ( .A1(n7243), .A2(n15622), .ZN(n7242) );
  NAND2_X1 U10076 ( .A1(n10590), .A2(n10589), .ZN(n10633) );
  OAI22_X2 U10077 ( .A1(n13055), .A2(n12922), .B1(n13534), .B2(n13056), .ZN(
        n12966) );
  NAND2_X1 U10078 ( .A1(n10524), .A2(n12995), .ZN(n7308) );
  NAND3_X1 U10079 ( .A1(n15435), .A2(n15434), .A3(n7643), .ZN(n15444) );
  INV_X1 U10080 ( .A(n11588), .ZN(n11755) );
  NAND2_X1 U10081 ( .A1(n10595), .A2(n10594), .ZN(n10998) );
  NAND2_X1 U10082 ( .A1(n10633), .A2(n10634), .ZN(n10595) );
  OAI21_X2 U10083 ( .B1(n10082), .B2(P3_D_REG_0__SCAN_IN), .A(n9823), .ZN(
        n9824) );
  NAND2_X1 U10084 ( .A1(n7248), .A2(n12432), .ZN(n15030) );
  NAND2_X1 U10085 ( .A1(n15034), .A2(n7957), .ZN(n7248) );
  NAND2_X2 U10086 ( .A1(n7299), .A2(n7298), .ZN(n12688) );
  NAND4_X2 U10087 ( .A1(n10906), .A2(n10905), .A3(n10904), .A4(n10903), .ZN(
        n14788) );
  NAND2_X1 U10088 ( .A1(n12955), .A2(n12954), .ZN(n13012) );
  NAND2_X1 U10089 ( .A1(n13707), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9129) );
  XNOR2_X1 U10091 ( .A(n8326), .B(n11701), .ZN(n8325) );
  NAND2_X1 U10092 ( .A1(n12820), .A2(n7453), .ZN(n12847) );
  NAND2_X2 U10093 ( .A1(n8060), .A2(n8059), .ZN(n8167) );
  NAND2_X1 U10094 ( .A1(n8341), .A2(n12055), .ZN(n8342) );
  NAND3_X1 U10095 ( .A1(n7255), .A2(n7254), .A3(n7253), .ZN(P3_U3201) );
  NAND2_X1 U10096 ( .A1(n13314), .A2(n13313), .ZN(n7255) );
  NAND2_X1 U10097 ( .A1(n11301), .A2(n11300), .ZN(n7660) );
  OAI21_X1 U10098 ( .B1(n8589), .B2(n7526), .A(n14272), .ZN(n7525) );
  NAND2_X1 U10099 ( .A1(n9253), .A2(n9252), .ZN(n9255) );
  NAND2_X1 U10100 ( .A1(n7872), .A2(n7870), .ZN(n9368) );
  NAND2_X1 U10101 ( .A1(n9466), .A2(n9465), .ZN(n9468) );
  NAND2_X1 U10102 ( .A1(n7408), .A2(n9693), .ZN(n7406) );
  NAND2_X1 U10103 ( .A1(n7491), .A2(n7490), .ZN(n14904) );
  NAND2_X1 U10104 ( .A1(n10469), .A2(n10470), .ZN(n7303) );
  NOR2_X1 U10105 ( .A1(n10317), .A2(n7301), .ZN(n10295) );
  NAND2_X1 U10106 ( .A1(n13484), .A2(n13485), .ZN(n7920) );
  NAND2_X1 U10107 ( .A1(n7932), .A2(n9633), .ZN(n7930) );
  NOR2_X1 U10108 ( .A1(n7937), .A2(n7933), .ZN(n7932) );
  NAND2_X1 U10109 ( .A1(n9255), .A2(n9044), .ZN(n9272) );
  NAND3_X1 U10110 ( .A1(n15408), .A2(n15407), .A3(n7656), .ZN(n15419) );
  NAND2_X1 U10111 ( .A1(n7263), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n7644) );
  NAND2_X1 U10112 ( .A1(n7646), .A2(n10605), .ZN(n7263) );
  XNOR2_X2 U10113 ( .A(n11464), .B(n7247), .ZN(n11588) );
  OAI22_X1 U10114 ( .A1(n13037), .A2(n13421), .B1(n13036), .B2(n13035), .ZN(
        n13040) );
  INV_X1 U10115 ( .A(n7719), .ZN(n7718) );
  OR2_X1 U10116 ( .A1(n7415), .A2(n6693), .ZN(n7407) );
  INV_X1 U10117 ( .A(n7270), .ZN(n9956) );
  NAND2_X1 U10118 ( .A1(n10106), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7264) );
  NAND3_X1 U10119 ( .A1(n9695), .A2(n9961), .A3(n7268), .ZN(n7267) );
  NAND2_X1 U10120 ( .A1(n7664), .A2(n7666), .ZN(n7663) );
  NAND2_X1 U10121 ( .A1(n9725), .A2(n9760), .ZN(n7269) );
  NAND2_X1 U10122 ( .A1(n7893), .A2(n7892), .ZN(n9549) );
  NAND2_X1 U10123 ( .A1(n13132), .A2(n6745), .ZN(n13134) );
  OR2_X1 U10124 ( .A1(n10984), .A2(n10985), .ZN(n7669) );
  NAND4_X1 U10125 ( .A1(n10217), .A2(n10216), .A3(n15963), .A4(n7146), .ZN(
        n10219) );
  INV_X1 U10126 ( .A(n11133), .ZN(n7299) );
  NAND2_X1 U10127 ( .A1(n10220), .A2(n7967), .ZN(n7329) );
  NAND2_X1 U10129 ( .A1(n7697), .A2(n10779), .ZN(n7696) );
  NAND2_X1 U10130 ( .A1(n7681), .A2(n10978), .ZN(n7271) );
  INV_X1 U10131 ( .A(n13287), .ZN(n7688) );
  NAND2_X1 U10132 ( .A1(n7629), .A2(n7628), .ZN(n9570) );
  INV_X1 U10133 ( .A(n13173), .ZN(n7679) );
  NAND2_X1 U10134 ( .A1(n7273), .A2(n13184), .ZN(n7272) );
  INV_X1 U10135 ( .A(n13172), .ZN(n7273) );
  NAND2_X1 U10136 ( .A1(n13149), .A2(n13148), .ZN(n7665) );
  NAND2_X1 U10137 ( .A1(n8306), .A2(n8305), .ZN(n8308) );
  INV_X1 U10138 ( .A(n13292), .ZN(n7699) );
  INV_X1 U10139 ( .A(n9326), .ZN(n9196) );
  NAND2_X1 U10140 ( .A1(n9326), .A2(n9094), .ZN(n9198) );
  INV_X1 U10141 ( .A(n14904), .ZN(n14903) );
  NAND2_X1 U10142 ( .A1(n10295), .A2(n10296), .ZN(n10649) );
  NAND2_X1 U10143 ( .A1(n15818), .A2(n15486), .ZN(n7276) );
  NOR2_X1 U10144 ( .A1(n10319), .A2(n10318), .ZN(n10317) );
  NAND2_X1 U10145 ( .A1(n6574), .A2(n7416), .ZN(n7410) );
  NAND2_X1 U10146 ( .A1(n15408), .A2(n15407), .ZN(n15416) );
  NAND2_X1 U10147 ( .A1(n9494), .A2(n11787), .ZN(n7887) );
  NAND2_X1 U10148 ( .A1(n9871), .A2(n9703), .ZN(n9563) );
  INV_X1 U10149 ( .A(n8593), .ZN(n7526) );
  NAND2_X1 U10150 ( .A1(n8189), .A2(n8071), .ZN(n7804) );
  INV_X1 U10151 ( .A(n7525), .ZN(n7524) );
  AOI21_X1 U10152 ( .B1(n7458), .B2(n7461), .A(n6717), .ZN(n7456) );
  NAND2_X1 U10153 ( .A1(n10919), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n11029) );
  NAND2_X1 U10154 ( .A1(n12078), .A2(n12077), .ZN(n12159) );
  NAND4_X1 U10155 ( .A1(n12896), .A2(n12897), .A3(n12894), .A4(n12895), .ZN(
        n7279) );
  OR4_X2 U10156 ( .A1(n12889), .A2(n15105), .A3(n15126), .A4(n15164), .ZN(
        n12890) );
  OAI21_X1 U10157 ( .B1(n8050), .B2(P2_DATAO_REG_2__SCAN_IN), .A(n7280), .ZN(
        n8044) );
  INV_X1 U10158 ( .A(n12909), .ZN(n12910) );
  NOR2_X2 U10159 ( .A1(n12254), .A2(n12253), .ZN(n7284) );
  NOR3_X2 U10160 ( .A1(n12304), .A2(n12303), .A3(n14705), .ZN(n12315) );
  NAND2_X2 U10161 ( .A1(n7968), .A2(n7969), .ZN(n11866) );
  NAND2_X1 U10162 ( .A1(n7703), .A2(n13244), .ZN(n13268) );
  NAND3_X1 U10163 ( .A1(n7663), .A2(n7665), .A3(n7668), .ZN(n13172) );
  NAND3_X1 U10164 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), 
        .A3(n9151), .ZN(n7661) );
  NAND2_X1 U10165 ( .A1(n11558), .A2(n7297), .ZN(n11561) );
  NAND2_X1 U10166 ( .A1(n11155), .A2(n11154), .ZN(n11345) );
  OR2_X1 U10167 ( .A1(n14792), .A2(n10668), .ZN(n11149) );
  NAND2_X1 U10168 ( .A1(n14867), .A2(n7503), .ZN(n14869) );
  OAI211_X1 U10169 ( .C1(n9806), .C2(n12996), .A(n9862), .B(n13552), .ZN(n7287) );
  NAND2_X1 U10170 ( .A1(n7290), .A2(n7288), .ZN(P3_U3487) );
  OR2_X1 U10171 ( .A1(n9861), .A2(n15801), .ZN(n7290) );
  NAND2_X1 U10172 ( .A1(n7293), .A2(n7291), .ZN(P3_U3455) );
  OR2_X1 U10173 ( .A1(n9861), .A2(n15788), .ZN(n7293) );
  INV_X1 U10174 ( .A(n13350), .ZN(n7310) );
  NAND2_X1 U10175 ( .A1(n9423), .A2(n9422), .ZN(n7886) );
  NAND2_X1 U10176 ( .A1(n9152), .A2(n9033), .ZN(n9184) );
  OAI22_X1 U10177 ( .A1(n7753), .A2(n7752), .B1(n9797), .B2(n13433), .ZN(n7751) );
  NAND4_X1 U10178 ( .A1(n7407), .A2(n7406), .A3(n7411), .A4(n7409), .ZN(n9700)
         );
  NAND2_X1 U10179 ( .A1(n9481), .A2(n9480), .ZN(n9483) );
  INV_X1 U10180 ( .A(n7415), .ZN(n7408) );
  OAI21_X1 U10181 ( .B1(n14143), .B2(n7784), .A(n7782), .ZN(n7781) );
  NAND2_X1 U10182 ( .A1(n11669), .A2(n11668), .ZN(n11671) );
  NAND2_X1 U10183 ( .A1(n15419), .A2(n15418), .ZN(n7657) );
  NAND2_X1 U10184 ( .A1(n6593), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n13293) );
  INV_X1 U10185 ( .A(n7472), .ZN(n7601) );
  NOR2_X2 U10186 ( .A1(n10218), .A2(n10219), .ZN(n10220) );
  NAND4_X1 U10187 ( .A1(n9942), .A2(n9941), .A3(n15826), .A4(n10205), .ZN(
        n10218) );
  NOR2_X2 U10188 ( .A1(n7300), .A2(n9936), .ZN(n10540) );
  NAND3_X1 U10189 ( .A1(n9934), .A2(n10195), .A3(n9935), .ZN(n7300) );
  NAND2_X1 U10190 ( .A1(n9105), .A2(n9106), .ZN(n7756) );
  XNOR2_X1 U10191 ( .A(n11589), .B(n13114), .ZN(n11758) );
  AOI21_X1 U10192 ( .B1(P3_REG1_REG_6__SCAN_IN), .B2(n10949), .A(n10948), .ZN(
        n10950) );
  NAND2_X1 U10193 ( .A1(n12966), .A2(n12965), .ZN(n12925) );
  INV_X1 U10194 ( .A(n7710), .ZN(n7709) );
  NAND2_X1 U10195 ( .A1(n9468), .A2(n9075), .ZN(n9481) );
  NAND2_X1 U10196 ( .A1(n9412), .A2(n9066), .ZN(n9068) );
  NAND2_X1 U10197 ( .A1(n10052), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7320) );
  NAND2_X2 U10198 ( .A1(n7321), .A2(P3_U3151), .ZN(n13723) );
  NAND2_X2 U10199 ( .A1(n7321), .A2(P1_U3086), .ZN(n15370) );
  INV_X1 U10200 ( .A(n10052), .ZN(n7321) );
  MUX2_X1 U10201 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n10052), .Z(n8211) );
  MUX2_X1 U10202 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n10052), .Z(n8298) );
  MUX2_X1 U10203 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n10052), .Z(n8260) );
  MUX2_X1 U10204 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n10052), .Z(n8324) );
  MUX2_X1 U10205 ( .A(n16023), .B(n12586), .S(n10052), .Z(n8340) );
  MUX2_X1 U10206 ( .A(n14589), .B(n15376), .S(n10052), .Z(n8361) );
  MUX2_X1 U10207 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n10052), .Z(n8373) );
  NAND2_X1 U10208 ( .A1(n7326), .A2(n7325), .ZN(n12016) );
  AOI21_X2 U10209 ( .B1(n15048), .B2(n6643), .A(n7953), .ZN(n15006) );
  NAND2_X1 U10210 ( .A1(n7948), .A2(n7947), .ZN(n7333) );
  INV_X4 U10211 ( .A(n10897), .ZN(n12855) );
  AOI21_X2 U10212 ( .B1(n8729), .B2(n8728), .A(n8010), .ZN(n14143) );
  INV_X1 U10213 ( .A(n7761), .ZN(n7760) );
  NAND2_X1 U10214 ( .A1(n10853), .A2(n10852), .ZN(n10857) );
  NOR2_X1 U10215 ( .A1(n8382), .A2(n6730), .ZN(n7347) );
  NAND2_X1 U10216 ( .A1(n7351), .A2(n6724), .ZN(n7350) );
  OR2_X2 U10217 ( .A1(n10855), .A2(n7354), .ZN(n7351) );
  NAND2_X1 U10218 ( .A1(n7744), .A2(n7358), .ZN(n7357) );
  NAND2_X1 U10219 ( .A1(n7357), .A2(n7355), .ZN(n12606) );
  NAND2_X1 U10220 ( .A1(n12654), .A2(n7372), .ZN(n7371) );
  OR2_X2 U10221 ( .A1(n12654), .A2(n7369), .ZN(n7363) );
  NAND2_X1 U10222 ( .A1(n13823), .A2(n7378), .ZN(n7377) );
  INV_X1 U10223 ( .A(n7376), .ZN(n7378) );
  NAND2_X1 U10224 ( .A1(n7377), .A2(n7374), .ZN(n13778) );
  OAI21_X1 U10225 ( .B1(n7376), .B2(n7386), .A(n6603), .ZN(n7375) );
  NAND3_X1 U10226 ( .A1(n6635), .A2(n9112), .A3(n9111), .ZN(n9263) );
  NAND2_X1 U10227 ( .A1(n9122), .A2(n6747), .ZN(n9472) );
  NAND3_X1 U10228 ( .A1(n9704), .A2(n7401), .A3(n13370), .ZN(n7400) );
  NAND3_X1 U10229 ( .A1(n9641), .A2(n9638), .A3(n9581), .ZN(n7405) );
  NAND3_X1 U10230 ( .A1(n7416), .A2(n6574), .A3(n9961), .ZN(n7415) );
  AND2_X1 U10231 ( .A1(n6693), .A2(n9855), .ZN(n7417) );
  NAND3_X1 U10232 ( .A1(n7419), .A2(n7421), .A3(n7418), .ZN(n7420) );
  NAND2_X1 U10233 ( .A1(n9597), .A2(n9596), .ZN(n7419) );
  NAND2_X1 U10234 ( .A1(n7420), .A2(n7422), .ZN(n9608) );
  NAND2_X1 U10235 ( .A1(n7426), .A2(n7425), .ZN(n7424) );
  NAND2_X1 U10236 ( .A1(n9587), .A2(n9961), .ZN(n7426) );
  XNOR2_X1 U10237 ( .A(n13120), .B(n10765), .ZN(n9585) );
  NAND2_X1 U10239 ( .A1(n9653), .A2(n7433), .ZN(n7432) );
  OAI21_X1 U10240 ( .B1(n7435), .B2(n9662), .A(n6675), .ZN(n7434) );
  AOI21_X1 U10241 ( .B1(n7441), .B2(n13487), .A(n13473), .ZN(n7438) );
  NAND4_X1 U10242 ( .A1(n9618), .A2(n11843), .A3(n9617), .A4(n11771), .ZN(
        n7446) );
  NAND2_X1 U10243 ( .A1(n8190), .A2(n7458), .ZN(n7457) );
  NAND2_X1 U10244 ( .A1(n8286), .A2(n7466), .ZN(n7464) );
  NOR2_X2 U10245 ( .A1(n11210), .A2(n12712), .ZN(n15519) );
  INV_X1 U10246 ( .A(n10463), .ZN(n10692) );
  INV_X1 U10247 ( .A(n15473), .ZN(n12912) );
  OAI21_X1 U10248 ( .B1(n6555), .B2(n10666), .A(n7473), .ZN(n7472) );
  NAND2_X1 U10249 ( .A1(n6555), .A2(n10665), .ZN(n7473) );
  INV_X1 U10250 ( .A(n15054), .ZN(n7474) );
  NAND2_X1 U10251 ( .A1(n7474), .A2(n7475), .ZN(n14994) );
  NOR2_X1 U10252 ( .A1(n14974), .A2(n7478), .ZN(n14937) );
  NAND2_X1 U10253 ( .A1(n7484), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10224) );
  NAND2_X1 U10254 ( .A1(n7964), .A2(n10220), .ZN(n7484) );
  AND2_X2 U10255 ( .A1(n7486), .A2(n12066), .ZN(n12169) );
  NAND3_X1 U10256 ( .A1(n7497), .A2(n7495), .A3(n7493), .ZN(n16121) );
  OAI21_X1 U10257 ( .B1(n10050), .B2(n10221), .A(P1_IR_REG_2__SCAN_IN), .ZN(
        n7506) );
  MUX2_X1 U10258 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n7000), .Z(n8107) );
  MUX2_X1 U10259 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n10052), .Z(n8317) );
  NOR2_X1 U10260 ( .A1(n14216), .A2(n14194), .ZN(n14197) );
  INV_X1 U10261 ( .A(n7515), .ZN(n14291) );
  NAND2_X1 U10262 ( .A1(n7516), .A2(n14128), .ZN(n14092) );
  NAND2_X1 U10263 ( .A1(n14128), .A2(n14414), .ZN(n8767) );
  INV_X1 U10264 ( .A(n11651), .ZN(n7527) );
  XNOR2_X2 U10265 ( .A(n8781), .B(n7528), .ZN(n8691) );
  OR2_X1 U10266 ( .A1(n10790), .A2(n7530), .ZN(n7529) );
  NAND2_X1 U10267 ( .A1(n7536), .A2(n8088), .ZN(n8094) );
  NAND4_X1 U10268 ( .A1(n7774), .A2(n7775), .A3(n8090), .A4(n8087), .ZN(n7536)
         );
  NAND3_X1 U10269 ( .A1(n7774), .A2(n7775), .A3(n8087), .ZN(n8405) );
  AND2_X2 U10270 ( .A1(n7774), .A2(n7775), .ZN(n8382) );
  NOR2_X1 U10271 ( .A1(n14163), .A2(n7556), .ZN(n7555) );
  NOR2_X4 U10272 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n9980) );
  INV_X1 U10273 ( .A(n10743), .ZN(n7580) );
  NAND3_X1 U10274 ( .A1(n7577), .A2(n7578), .A3(n7581), .ZN(n7574) );
  INV_X1 U10275 ( .A(n7569), .ZN(n10773) );
  NAND3_X1 U10276 ( .A1(n7577), .A2(n7578), .A3(n7571), .ZN(n7570) );
  NAND2_X1 U10277 ( .A1(n11093), .A2(n7580), .ZN(n7577) );
  NOR2_X1 U10278 ( .A1(n11093), .A2(n6631), .ZN(n10742) );
  OR2_X1 U10279 ( .A1(n13327), .A2(n13326), .ZN(n7582) );
  NAND2_X1 U10280 ( .A1(n13206), .A2(n7583), .ZN(n13229) );
  NOR2_X1 U10281 ( .A1(n13208), .A2(n13207), .ZN(n7587) );
  INV_X1 U10282 ( .A(n13175), .ZN(n7589) );
  NAND3_X1 U10283 ( .A1(n12753), .A2(n12752), .A3(n6726), .ZN(n7596) );
  NAND2_X1 U10284 ( .A1(n7596), .A2(n7597), .ZN(n12769) );
  INV_X4 U10285 ( .A(n12681), .ZN(n12862) );
  NAND2_X2 U10286 ( .A1(n12808), .A2(n12677), .ZN(n12681) );
  AND2_X1 U10287 ( .A1(n12687), .A2(n12862), .ZN(n12680) );
  INV_X1 U10288 ( .A(n12796), .ZN(n7603) );
  NAND2_X1 U10289 ( .A1(n12798), .A2(n12797), .ZN(n7604) );
  NAND2_X1 U10290 ( .A1(n12693), .A2(n12692), .ZN(n7608) );
  NAND3_X1 U10291 ( .A1(n7606), .A2(n12698), .A3(n7605), .ZN(n12702) );
  NAND3_X1 U10292 ( .A1(n12874), .A2(n12694), .A3(n7607), .ZN(n7605) );
  NAND4_X1 U10293 ( .A1(n12689), .A2(n7608), .A3(n12690), .A4(n12874), .ZN(
        n7606) );
  NAND3_X1 U10294 ( .A1(n12732), .A2(n12731), .A3(n6716), .ZN(n7610) );
  NAND2_X1 U10295 ( .A1(n7611), .A2(n6723), .ZN(n12748) );
  NAND3_X1 U10296 ( .A1(n12741), .A2(n8026), .A3(n6719), .ZN(n7611) );
  NAND2_X1 U10297 ( .A1(n7613), .A2(n7614), .ZN(n12715) );
  NAND3_X1 U10298 ( .A1(n12707), .A2(n6721), .A3(n12706), .ZN(n7613) );
  NAND2_X1 U10299 ( .A1(n7616), .A2(n7617), .ZN(n12727) );
  NAND3_X1 U10300 ( .A1(n12720), .A2(n6720), .A3(n12719), .ZN(n7616) );
  XNOR2_X2 U10301 ( .A(n12975), .B(n12973), .ZN(n13064) );
  AND2_X1 U10302 ( .A1(n9324), .A2(n7631), .ZN(n7628) );
  AND2_X1 U10303 ( .A1(n7627), .A2(n7662), .ZN(n7623) );
  AND3_X1 U10304 ( .A1(n9101), .A2(n7623), .A3(n9980), .ZN(n7629) );
  NAND3_X1 U10305 ( .A1(n9324), .A2(n6741), .A3(n7631), .ZN(n9328) );
  NAND3_X1 U10306 ( .A1(n15435), .A2(n15434), .A3(P2_ADDR_REG_17__SCAN_IN), 
        .ZN(n7641) );
  NAND3_X1 U10307 ( .A1(n7646), .A2(n7645), .A3(n10605), .ZN(n10606) );
  NAND2_X1 U10308 ( .A1(n10606), .A2(n7644), .ZN(n10164) );
  INV_X1 U10309 ( .A(n10164), .ZN(n10161) );
  INV_X1 U10310 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7645) );
  INV_X1 U10311 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7647) );
  NAND2_X1 U10312 ( .A1(n7648), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n10139) );
  NAND2_X1 U10313 ( .A1(n7654), .A2(n7655), .ZN(n12203) );
  NAND2_X1 U10314 ( .A1(n7654), .A2(n7652), .ZN(n15390) );
  NAND2_X1 U10315 ( .A1(n7660), .A2(n11302), .ZN(n11309) );
  NAND2_X1 U10316 ( .A1(n8149), .A2(n8148), .ZN(n11958) );
  INV_X1 U10317 ( .A(n11103), .ZN(n8008) );
  INV_X1 U10318 ( .A(n10330), .ZN(n9937) );
  NAND2_X1 U10319 ( .A1(n10215), .A2(n10214), .ZN(n12673) );
  OR2_X2 U10320 ( .A1(n12740), .A2(n12739), .ZN(n8026) );
  INV_X1 U10321 ( .A(n15213), .ZN(n7790) );
  OAI21_X1 U10322 ( .B1(n14327), .B2(n8574), .A(n9007), .ZN(n14281) );
  NAND2_X1 U10323 ( .A1(n8452), .A2(n11969), .ZN(n11968) );
  NAND2_X1 U10324 ( .A1(n8094), .A2(n8390), .ZN(n8399) );
  XNOR2_X1 U10325 ( .A(n10106), .B(n10770), .ZN(n10749) );
  INV_X1 U10326 ( .A(n13134), .ZN(n7667) );
  INV_X1 U10327 ( .A(n7670), .ZN(n9958) );
  NAND2_X1 U10328 ( .A1(n13186), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n13194) );
  NAND2_X1 U10329 ( .A1(n13221), .A2(n13256), .ZN(n7674) );
  NAND3_X1 U10330 ( .A1(n7674), .A2(n7673), .A3(n6754), .ZN(n13264) );
  NAND3_X1 U10331 ( .A1(n7685), .A2(n13315), .A3(n7684), .ZN(n13317) );
  NAND2_X1 U10332 ( .A1(n7689), .A2(n13287), .ZN(n13267) );
  NAND2_X1 U10333 ( .A1(n7684), .A2(n7685), .ZN(n13316) );
  OR2_X1 U10334 ( .A1(n13265), .A2(n13279), .ZN(n7689) );
  NAND2_X1 U10335 ( .A1(n7695), .A2(n9990), .ZN(n9988) );
  INV_X1 U10336 ( .A(n9987), .ZN(n7697) );
  NAND3_X1 U10337 ( .A1(n7700), .A2(n7698), .A3(n13310), .ZN(n13312) );
  NAND2_X1 U10338 ( .A1(n7705), .A2(n13242), .ZN(n7703) );
  NAND2_X1 U10339 ( .A1(n10526), .A2(n7706), .ZN(n10758) );
  AOI21_X1 U10340 ( .B1(n9593), .B2(n7706), .A(n9592), .ZN(n9597) );
  NAND2_X1 U10341 ( .A1(n7715), .A2(n7713), .ZN(n13457) );
  NAND2_X1 U10342 ( .A1(n7721), .A2(n7718), .ZN(n9863) );
  NAND2_X1 U10343 ( .A1(n13351), .A2(n7722), .ZN(n7721) );
  NAND2_X2 U10344 ( .A1(n13775), .A2(n7725), .ZN(n12654) );
  NAND2_X2 U10345 ( .A1(n7728), .A2(n12647), .ZN(n13775) );
  INV_X1 U10346 ( .A(n13778), .ZN(n7728) );
  NAND2_X1 U10347 ( .A1(n12617), .A2(n7729), .ZN(n13755) );
  NAND2_X1 U10348 ( .A1(n9786), .A2(n9785), .ZN(n13546) );
  NOR2_X1 U10349 ( .A1(n9788), .A2(n7742), .ZN(n7741) );
  INV_X1 U10350 ( .A(n9785), .ZN(n7742) );
  OAI21_X2 U10351 ( .B1(n13443), .B2(n7752), .A(n7750), .ZN(n13403) );
  AND2_X1 U10352 ( .A1(n10030), .A2(n10021), .ZN(n7755) );
  INV_X1 U10353 ( .A(n14225), .ZN(n7759) );
  NAND2_X1 U10354 ( .A1(n8702), .A2(n7766), .ZN(n7765) );
  NAND2_X1 U10355 ( .A1(n8702), .A2(n8701), .ZN(n11993) );
  NAND2_X1 U10356 ( .A1(n8729), .A2(n7779), .ZN(n7776) );
  NAND2_X1 U10357 ( .A1(n7776), .A2(n7777), .ZN(n9906) );
  NAND2_X1 U10358 ( .A1(n8133), .A2(n7787), .ZN(n8135) );
  XNOR2_X1 U10359 ( .A(n8132), .B(n7787), .ZN(n10886) );
  NAND2_X2 U10360 ( .A1(n7788), .A2(n12245), .ZN(n15314) );
  NAND3_X1 U10361 ( .A1(n8035), .A2(n8036), .A3(n8037), .ZN(n7791) );
  NAND3_X1 U10362 ( .A1(n8034), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7793) );
  NOR2_X2 U10363 ( .A1(n14966), .A2(n7816), .ZN(n7815) );
  AOI21_X1 U10364 ( .B1(n8806), .B2(n8805), .A(n8804), .ZN(n8808) );
  NAND2_X1 U10365 ( .A1(n7819), .A2(n7818), .ZN(n7817) );
  INV_X1 U10366 ( .A(n8801), .ZN(n7818) );
  INV_X1 U10367 ( .A(n7823), .ZN(n7819) );
  NAND2_X1 U10368 ( .A1(n7822), .A2(n7821), .ZN(n7820) );
  NAND2_X1 U10369 ( .A1(n7823), .A2(n8801), .ZN(n7822) );
  OAI211_X1 U10370 ( .C1(n9004), .C2(n6761), .A(n7824), .B(n7826), .ZN(
        P2_U3328) );
  NAND2_X1 U10371 ( .A1(n9004), .A2(n7825), .ZN(n7824) );
  OR2_X1 U10372 ( .A1(n9023), .A2(n7827), .ZN(n7825) );
  AOI21_X1 U10373 ( .B1(n8840), .B2(n8839), .A(n8838), .ZN(n8841) );
  OAI22_X2 U10374 ( .A1(n7858), .A2(n7856), .B1(n8825), .B2(n7855), .ZN(n8831)
         );
  INV_X1 U10375 ( .A(n8825), .ZN(n7857) );
  NAND2_X1 U10376 ( .A1(n8906), .A2(n7864), .ZN(n7860) );
  NAND3_X1 U10377 ( .A1(n7861), .A2(n7860), .A3(n7862), .ZN(n8914) );
  NAND2_X2 U10378 ( .A1(n7869), .A2(n9518), .ZN(n13629) );
  NAND2_X1 U10379 ( .A1(n9322), .A2(n7874), .ZN(n7872) );
  NAND2_X1 U10380 ( .A1(n13710), .A2(n9550), .ZN(n7890) );
  NAND2_X1 U10381 ( .A1(n7890), .A2(n9108), .ZN(n13618) );
  INV_X1 U10382 ( .A(n11770), .ZN(n7899) );
  NAND2_X1 U10383 ( .A1(n6571), .A2(n11770), .ZN(n7895) );
  OAI21_X1 U10384 ( .B1(n11770), .B2(n9289), .A(n9288), .ZN(n11842) );
  NAND2_X1 U10385 ( .A1(n9524), .A2(n9683), .ZN(n13356) );
  NAND3_X1 U10386 ( .A1(n7939), .A2(n7942), .A3(n15608), .ZN(n7940) );
  NAND2_X1 U10387 ( .A1(n14930), .A2(n14935), .ZN(n7946) );
  NAND3_X1 U10388 ( .A1(n7942), .A2(n7944), .A3(n7941), .ZN(n15215) );
  INV_X1 U10389 ( .A(n12074), .ZN(n7948) );
  INV_X1 U10390 ( .A(n7962), .ZN(n15086) );
  NAND2_X1 U10391 ( .A1(n14704), .A2(n7987), .ZN(n7986) );
  INV_X1 U10392 ( .A(n12504), .ZN(n7999) );
  INV_X1 U10393 ( .A(n6562), .ZN(n11359) );
  NAND2_X1 U10394 ( .A1(n13900), .A2(n13748), .ZN(n13787) );
  INV_X1 U10395 ( .A(n10223), .ZN(n10226) );
  NAND2_X2 U10396 ( .A1(n10523), .A2(n10522), .ZN(n10587) );
  OR2_X1 U10397 ( .A1(n14938), .A2(n14937), .ZN(n15222) );
  OR2_X1 U10398 ( .A1(n9891), .A2(n13561), .ZN(n9897) );
  CLKBUF_X1 U10399 ( .A(n9747), .Z(n13716) );
  INV_X1 U10400 ( .A(n13789), .ZN(n11633) );
  NAND2_X1 U10401 ( .A1(n12593), .A2(n12592), .ZN(n12594) );
  AOI21_X2 U10402 ( .B1(n13064), .B2(n13433), .A(n12976), .ZN(n13035) );
  NAND2_X1 U10403 ( .A1(n13269), .A2(n13279), .ZN(n13292) );
  NAND2_X1 U10404 ( .A1(n14114), .A2(n15740), .ZN(n8769) );
  AND2_X1 U10405 ( .A1(n10675), .A2(n10692), .ZN(n15180) );
  XNOR2_X1 U10406 ( .A(n8314), .B(SI_22_), .ZN(n12326) );
  AND2_X1 U10407 ( .A1(n8781), .A2(n12612), .ZN(n10014) );
  NAND2_X1 U10408 ( .A1(n8753), .A2(n9904), .ZN(n8754) );
  NAND2_X1 U10409 ( .A1(n9368), .A2(n9059), .ZN(n9062) );
  OR2_X1 U10410 ( .A1(n12328), .A2(n10887), .ZN(n10888) );
  NOR2_X1 U10411 ( .A1(n14086), .A2(n9010), .ZN(n8950) );
  INV_X1 U10412 ( .A(n8271), .ZN(n8244) );
  AND2_X1 U10413 ( .A1(n8234), .A2(n8271), .ZN(n11886) );
  NAND2_X1 U10414 ( .A1(n10670), .A2(n10669), .ZN(n10671) );
  INV_X1 U10415 ( .A(n9211), .ZN(n9531) );
  NAND2_X1 U10416 ( .A1(n11356), .A2(n12874), .ZN(n11160) );
  INV_X1 U10417 ( .A(n10259), .ZN(n15374) );
  NAND2_X1 U10418 ( .A1(n13354), .A2(n9753), .ZN(n9755) );
  NAND2_X1 U10419 ( .A1(n10668), .A2(n6553), .ZN(n10669) );
  NAND2_X1 U10420 ( .A1(n10257), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10258) );
  NAND2_X1 U10421 ( .A1(n9703), .A2(n9702), .ZN(n9870) );
  INV_X1 U10422 ( .A(n11656), .ZN(n8496) );
  AND2_X1 U10423 ( .A1(n14167), .A2(n13768), .ZN(n8010) );
  AND2_X1 U10424 ( .A1(n9896), .A2(n8014), .ZN(n8011) );
  AND2_X1 U10425 ( .A1(n12452), .A2(n15189), .ZN(n15525) );
  OR2_X1 U10426 ( .A1(n14086), .A2(n9003), .ZN(n8012) );
  OR2_X1 U10427 ( .A1(n15743), .A2(n8771), .ZN(n8013) );
  AND2_X2 U10428 ( .A1(n9926), .A2(n9925), .ZN(n15750) );
  INV_X1 U10429 ( .A(n15750), .ZN(n12591) );
  AND2_X2 U10430 ( .A1(n11617), .A2(n9925), .ZN(n15743) );
  INV_X1 U10431 ( .A(n13566), .ZN(n9690) );
  OR2_X1 U10432 ( .A1(n13553), .A2(n9895), .ZN(n8014) );
  AND2_X1 U10433 ( .A1(n14968), .A2(n12434), .ZN(n8016) );
  OR2_X1 U10434 ( .A1(n7520), .A2(n14574), .ZN(n8017) );
  AND2_X1 U10435 ( .A1(n13935), .A2(n6556), .ZN(n8018) );
  AND2_X1 U10436 ( .A1(n8078), .A2(n8077), .ZN(n8019) );
  INV_X1 U10437 ( .A(n13733), .ZN(n13726) );
  AND2_X1 U10438 ( .A1(n10703), .A2(n10702), .ZN(n8020) );
  INV_X1 U10439 ( .A(n11957), .ZN(n8149) );
  INV_X1 U10440 ( .A(n11771), .ZN(n9778) );
  AND2_X1 U10441 ( .A1(n8250), .A2(n8242), .ZN(n8023) );
  AND2_X1 U10442 ( .A1(n8239), .A2(n8228), .ZN(n8024) );
  OR2_X1 U10443 ( .A1(n8298), .A2(SI_21_), .ZN(n8025) );
  AND2_X1 U10444 ( .A1(n8987), .A2(n8978), .ZN(n8028) );
  INV_X1 U10445 ( .A(n8995), .ZN(n14408) );
  AND2_X1 U10446 ( .A1(n8074), .A2(n8073), .ZN(n8029) );
  AND2_X1 U10447 ( .A1(n9905), .A2(n9904), .ZN(n8030) );
  OR2_X1 U10448 ( .A1(n14111), .A2(n14574), .ZN(n8031) );
  OR2_X1 U10449 ( .A1(n8296), .A2(SI_20_), .ZN(n8032) );
  NOR3_X1 U10450 ( .A1(n14446), .A2(n14445), .A3(n14444), .ZN(n8033) );
  INV_X1 U10451 ( .A(n14222), .ZN(n14226) );
  NAND2_X1 U10452 ( .A1(n9174), .A2(n9584), .ZN(n10799) );
  AOI21_X1 U10453 ( .B1(n12684), .B2(n12683), .A(n12682), .ZN(n12685) );
  OAI21_X1 U10454 ( .B1(n8785), .B2(n15660), .A(n8921), .ZN(n8786) );
  INV_X1 U10455 ( .A(n8786), .ZN(n8787) );
  NAND2_X1 U10456 ( .A1(n8788), .A2(n8787), .ZN(n8789) );
  NAND2_X1 U10457 ( .A1(n8799), .A2(n8798), .ZN(n8801) );
  INV_X1 U10458 ( .A(n12736), .ZN(n12737) );
  OAI21_X1 U10459 ( .B1(n9640), .B2(n9377), .A(n6888), .ZN(n9641) );
  AND2_X1 U10460 ( .A1(n8883), .A2(n8873), .ZN(n8874) );
  INV_X1 U10461 ( .A(n12775), .ZN(n12776) );
  NOR2_X1 U10462 ( .A1(n13089), .A2(n9961), .ZN(n9689) );
  NAND2_X1 U10463 ( .A1(n9690), .A2(n9689), .ZN(n9691) );
  INV_X1 U10464 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n10216) );
  INV_X1 U10465 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n9093) );
  INV_X1 U10466 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9812) );
  INV_X1 U10467 ( .A(n15149), .ZN(n12270) );
  INV_X1 U10468 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9941) );
  AND2_X1 U10469 ( .A1(n14282), .A2(n8590), .ZN(n8589) );
  INV_X1 U10470 ( .A(n11870), .ZN(n11867) );
  INV_X1 U10471 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n15823) );
  INV_X1 U10472 ( .A(n15126), .ZN(n12281) );
  INV_X1 U10473 ( .A(n13390), .ZN(n9504) );
  AND2_X1 U10474 ( .A1(n9071), .A2(n9454), .ZN(n9072) );
  INV_X1 U10475 ( .A(n9323), .ZN(n9324) );
  INV_X1 U10476 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8037) );
  AND2_X1 U10477 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n8518) );
  INV_X1 U10478 ( .A(n11224), .ZN(n8148) );
  INV_X1 U10479 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8391) );
  AND2_X1 U10480 ( .A1(n8268), .A2(n8267), .ZN(n8269) );
  INV_X1 U10481 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n11527) );
  INV_X1 U10482 ( .A(n10218), .ZN(n9943) );
  OR2_X1 U10483 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n16119), .ZN(n10611) );
  INV_X1 U10484 ( .A(n9542), .ZN(n9127) );
  INV_X1 U10485 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9120) );
  INV_X1 U10486 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n9115) );
  NOR2_X1 U10487 ( .A1(n6620), .A2(n13503), .ZN(n13501) );
  AND2_X1 U10488 ( .A1(n10498), .A2(n15770), .ZN(n10530) );
  XNOR2_X1 U10489 ( .A(n13789), .B(n15707), .ZN(n10016) );
  INV_X1 U10490 ( .A(n10858), .ZN(n10854) );
  INV_X1 U10491 ( .A(n11925), .ZN(n11922) );
  AND2_X1 U10492 ( .A1(n13741), .A2(n13740), .ZN(n13742) );
  NAND2_X1 U10493 ( .A1(n8594), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8601) );
  INV_X1 U10494 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10873) );
  OAI21_X1 U10495 ( .B1(n9917), .B2(n13915), .A(n9916), .ZN(n9918) );
  INV_X1 U10496 ( .A(n13931), .ZN(n8764) );
  INV_X1 U10497 ( .A(n10009), .ZN(n11653) );
  AND2_X1 U10498 ( .A1(n10038), .A2(n6562), .ZN(n8951) );
  OR2_X1 U10499 ( .A1(n14339), .A2(n13945), .ZN(n8564) );
  INV_X1 U10500 ( .A(n14632), .ZN(n12518) );
  INV_X1 U10501 ( .A(n14736), .ZN(n12511) );
  XNOR2_X1 U10502 ( .A(n12712), .B(n14786), .ZN(n12877) );
  AND3_X1 U10503 ( .A1(n11893), .A2(P1_B_REG_SCAN_IN), .A3(n11786), .ZN(n10187) );
  NAND2_X1 U10504 ( .A1(n8260), .A2(SI_19_), .ZN(n8283) );
  AND2_X1 U10505 ( .A1(n10129), .A2(n10128), .ZN(n10142) );
  OR2_X1 U10506 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n10621), .ZN(n10622) );
  INV_X1 U10507 ( .A(n12953), .ZN(n12954) );
  INV_X1 U10508 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9110) );
  NAND2_X1 U10509 ( .A1(n10515), .A2(n10514), .ZN(n13088) );
  AND2_X1 U10510 ( .A1(n9560), .A2(n9144), .ZN(n12004) );
  NAND2_X2 U10511 ( .A1(n13714), .A2(n9132), .ZN(n9175) );
  INV_X1 U10512 ( .A(n13374), .ZN(n13406) );
  INV_X1 U10513 ( .A(n11052), .ZN(n10766) );
  OAI211_X1 U10514 ( .C1(n13701), .C2(n9887), .A(n9886), .B(n9885), .ZN(n9892)
         );
  AND2_X1 U10515 ( .A1(n9560), .A2(n9136), .ZN(n13336) );
  INV_X1 U10516 ( .A(n13547), .ZN(n13535) );
  INV_X1 U10517 ( .A(n13915), .ZN(n13905) );
  XNOR2_X1 U10518 ( .A(n10016), .B(n10014), .ZN(n10401) );
  AND2_X1 U10519 ( .A1(n8674), .A2(n8665), .ZN(n14150) );
  INV_X1 U10520 ( .A(n8739), .ZN(n8755) );
  OR2_X1 U10521 ( .A1(n8468), .A2(n8444), .ZN(n8451) );
  INV_X1 U10522 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n13894) );
  NAND2_X1 U10523 ( .A1(n10036), .A2(n15702), .ZN(n14398) );
  INV_X1 U10524 ( .A(n14575), .ZN(n14513) );
  AND2_X1 U10525 ( .A1(n9008), .A2(n9007), .ZN(n14326) );
  NOR2_X1 U10526 ( .A1(n9924), .A2(n8419), .ZN(n10007) );
  OR2_X1 U10527 ( .A1(n10700), .A2(n10359), .ZN(n10363) );
  INV_X1 U10528 ( .A(n15130), .ZN(n15178) );
  INV_X1 U10529 ( .A(n15599), .ZN(n15530) );
  INV_X1 U10530 ( .A(n13088), .ZN(n13096) );
  INV_X1 U10531 ( .A(n11312), .ZN(n9731) );
  INV_X1 U10532 ( .A(n13085), .ZN(n13386) );
  INV_X1 U10533 ( .A(n11845), .ZN(n11759) );
  NAND2_X1 U10534 ( .A1(n9746), .A2(n9745), .ZN(n10501) );
  INV_X1 U10535 ( .A(n13610), .ZN(n13614) );
  AND4_X1 U10536 ( .A1(n10535), .A2(n9844), .A3(n9843), .A4(n9884), .ZN(n9845)
         );
  INV_X1 U10537 ( .A(n13502), .ZN(n13552) );
  INV_X1 U10538 ( .A(n15771), .ZN(n15784) );
  NAND2_X1 U10539 ( .A1(n9764), .A2(n11382), .ZN(n15770) );
  INV_X4 U10540 ( .A(n8097), .ZN(n10885) );
  INV_X1 U10541 ( .A(n13917), .ZN(n13907) );
  INV_X1 U10542 ( .A(n13925), .ZN(n13903) );
  AND2_X1 U10543 ( .A1(n8645), .A2(n8644), .ZN(n13801) );
  AND2_X1 U10544 ( .A1(n15633), .A2(n10456), .ZN(n15651) );
  AND2_X1 U10545 ( .A1(n14285), .A2(n14086), .ZN(n14401) );
  INV_X1 U10546 ( .A(n14361), .ZN(n14312) );
  NAND2_X1 U10547 ( .A1(n12591), .A2(n12590), .ZN(n12592) );
  INV_X1 U10548 ( .A(n14574), .ZN(n8433) );
  OAI21_X1 U10549 ( .B1(n8763), .B2(n14375), .A(n13795), .ZN(n14108) );
  OAI21_X1 U10550 ( .B1(n14086), .B2(n15659), .A(n10034), .ZN(n14518) );
  NAND2_X1 U10551 ( .A1(n8950), .A2(n11491), .ZN(n15716) );
  NAND2_X1 U10552 ( .A1(n15716), .A2(n15715), .ZN(n15740) );
  AND2_X1 U10553 ( .A1(n15701), .A2(n8431), .ZN(n9925) );
  AOI21_X1 U10554 ( .B1(n8413), .B2(n11895), .A(n12119), .ZN(n15670) );
  OR2_X1 U10555 ( .A1(n12859), .A2(n10692), .ZN(n15130) );
  AND4_X1 U10556 ( .A1(n12166), .A2(n12165), .A3(n12164), .A4(n12163), .ZN(
        n14758) );
  INV_X1 U10557 ( .A(n15814), .ZN(n15483) );
  OR2_X1 U10558 ( .A1(n15478), .A2(n12912), .ZN(n15817) );
  INV_X1 U10559 ( .A(n15815), .ZN(n15812) );
  INV_X1 U10560 ( .A(n15538), .ZN(n15517) );
  XOR2_X1 U10561 ( .A(n14770), .B(n15230), .Z(n14955) );
  OAI21_X1 U10562 ( .B1(n10349), .B2(P1_D_REG_0__SCAN_IN), .A(n10348), .ZN(
        n15202) );
  AND2_X1 U10563 ( .A1(n12674), .A2(n10355), .ZN(n15558) );
  INV_X1 U10564 ( .A(n15561), .ZN(n15588) );
  INV_X1 U10565 ( .A(n15558), .ZN(n15552) );
  NAND2_X1 U10566 ( .A1(n10188), .A2(n10376), .ZN(n11131) );
  XNOR2_X1 U10567 ( .A(n9946), .B(n15963), .ZN(n10185) );
  AND2_X1 U10568 ( .A1(n9998), .A2(n9997), .ZN(n15751) );
  INV_X1 U10569 ( .A(n13102), .ZN(n13081) );
  INV_X1 U10570 ( .A(n13536), .ZN(n13111) );
  INV_X1 U10571 ( .A(n13332), .ZN(n13210) );
  INV_X1 U10572 ( .A(n13318), .ZN(n13283) );
  NAND2_X1 U10573 ( .A1(n13553), .A2(n9890), .ZN(n13561) );
  INV_X1 U10574 ( .A(n13400), .ZN(n11912) );
  INV_X1 U10575 ( .A(n13622), .ZN(n13565) );
  NAND2_X1 U10576 ( .A1(n15804), .A2(n15755), .ZN(n13617) );
  INV_X1 U10577 ( .A(n15804), .ZN(n15801) );
  OR2_X1 U10578 ( .A1(n15788), .A2(n9876), .ZN(n13699) );
  INV_X2 U10579 ( .A(n15788), .ZN(n15786) );
  NAND2_X1 U10580 ( .A1(n10082), .A2(n10081), .ZN(n10116) );
  INV_X1 U10581 ( .A(SI_26_), .ZN(n12055) );
  INV_X1 U10582 ( .A(SI_16_), .ZN(n10307) );
  NAND2_X1 U10583 ( .A1(n10040), .A2(n10039), .ZN(n13855) );
  INV_X1 U10584 ( .A(n13923), .ZN(n13912) );
  INV_X1 U10585 ( .A(n9917), .ZN(n13930) );
  INV_X1 U10586 ( .A(n12655), .ZN(n13937) );
  INV_X1 U10587 ( .A(n15644), .ZN(n15624) );
  OR2_X1 U10588 ( .A1(n10455), .A2(n8399), .ZN(n15623) );
  NAND2_X1 U10589 ( .A1(n14285), .A2(n11623), .ZN(n14399) );
  NAND2_X1 U10590 ( .A1(n14285), .A2(n11621), .ZN(n14361) );
  NAND2_X1 U10591 ( .A1(n15750), .A2(n14518), .ZN(n14514) );
  INV_X1 U10592 ( .A(n14274), .ZN(n14555) );
  NAND2_X1 U10593 ( .A1(n15743), .A2(n14518), .ZN(n14574) );
  INV_X1 U10594 ( .A(n15743), .ZN(n15741) );
  OR2_X1 U10595 ( .A1(n10005), .A2(n15699), .ZN(n15697) );
  NAND2_X1 U10596 ( .A1(n8405), .A2(n8403), .ZN(n11788) );
  INV_X1 U10597 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10644) );
  INV_X1 U10598 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10194) );
  OR2_X1 U10599 ( .A1(n14737), .A2(n15130), .ZN(n14706) );
  INV_X1 U10600 ( .A(n14753), .ZN(n14742) );
  INV_X1 U10601 ( .A(n14740), .ZN(n14765) );
  INV_X1 U10602 ( .A(n14990), .ZN(n14771) );
  INV_X1 U10603 ( .A(n15131), .ZN(n14777) );
  OR2_X1 U10604 ( .A1(n15478), .A2(n10692), .ZN(n15814) );
  OR2_X1 U10605 ( .A1(n15478), .A2(n10244), .ZN(n15815) );
  INV_X1 U10606 ( .A(n15097), .ZN(n15512) );
  OR2_X1 U10607 ( .A1(n15525), .A2(n11320), .ZN(n15195) );
  AND2_X1 U10608 ( .A1(n15500), .A2(n11147), .ZN(n15122) );
  INV_X2 U10609 ( .A(n15620), .ZN(n15622) );
  OR3_X1 U10610 ( .A1(n15328), .A2(n15327), .A3(n15326), .ZN(n15362) );
  AND3_X1 U10611 ( .A1(n15579), .A2(n15578), .A3(n15577), .ZN(n15616) );
  INV_X2 U10612 ( .A(n15606), .ZN(n15608) );
  INV_X1 U10613 ( .A(n15527), .ZN(n15526) );
  OR2_X1 U10614 ( .A1(n10189), .A2(n11131), .ZN(n15527) );
  INV_X1 U10615 ( .A(n12911), .ZN(n12915) );
  INV_X1 U10616 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11107) );
  INV_X1 U10617 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10316) );
  AND2_X1 U10618 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10430), .ZN(P2_U3947) );
  OAI21_X1 U10619 ( .B1(n12589), .B2(n15741), .A(n8772), .ZN(P2_U3495) );
  INV_X1 U10620 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8432) );
  INV_X1 U10621 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10053) );
  INV_X2 U10622 ( .A(P1_RD_REG_SCAN_IN), .ZN(n8035) );
  INV_X2 U10623 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9028) );
  AND2_X1 U10624 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8038) );
  INV_X1 U10625 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10051) );
  NAND2_X1 U10626 ( .A1(n8050), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8039) );
  INV_X1 U10627 ( .A(SI_1_), .ZN(n10101) );
  OAI211_X1 U10628 ( .C1(n8050), .C2(n10051), .A(n8039), .B(n10101), .ZN(n8040) );
  NAND2_X1 U10629 ( .A1(n8106), .A2(n8040), .ZN(n8043) );
  NAND2_X1 U10630 ( .A1(n8050), .A2(n9030), .ZN(n8041) );
  OAI211_X1 U10631 ( .C1(P2_DATAO_REG_1__SCAN_IN), .C2(n8050), .A(n8041), .B(
        SI_1_), .ZN(n8042) );
  INV_X1 U10632 ( .A(n8044), .ZN(n8045) );
  NAND2_X1 U10633 ( .A1(n8045), .A2(SI_2_), .ZN(n8046) );
  MUX2_X1 U10634 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8050), .Z(n8049) );
  XNOR2_X1 U10635 ( .A(n8049), .B(SI_4_), .ZN(n8136) );
  NOR2_X1 U10636 ( .A1(n8124), .A2(SI_3_), .ZN(n8047) );
  NOR2_X1 U10637 ( .A1(n8136), .A2(n8047), .ZN(n8048) );
  NAND2_X1 U10638 ( .A1(n8049), .A2(SI_4_), .ZN(n8140) );
  INV_X4 U10639 ( .A(n8097), .ZN(n12325) );
  NAND2_X1 U10640 ( .A1(n8142), .A2(SI_5_), .ZN(n8153) );
  NAND3_X1 U10641 ( .A1(n8141), .A2(n8140), .A3(n8153), .ZN(n8053) );
  XNOR2_X1 U10642 ( .A(n8054), .B(SI_6_), .ZN(n8155) );
  NOR2_X1 U10643 ( .A1(n8142), .A2(SI_5_), .ZN(n8051) );
  NOR2_X1 U10644 ( .A1(n8155), .A2(n8051), .ZN(n8052) );
  NAND2_X1 U10645 ( .A1(n8053), .A2(n8052), .ZN(n8056) );
  NAND2_X1 U10646 ( .A1(n8054), .A2(SI_6_), .ZN(n8055) );
  MUX2_X1 U10647 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n10885), .Z(n8058) );
  XNOR2_X1 U10648 ( .A(n8058), .B(SI_7_), .ZN(n8160) );
  INV_X1 U10649 ( .A(n8160), .ZN(n8057) );
  NAND2_X1 U10650 ( .A1(n8161), .A2(n8057), .ZN(n8060) );
  NAND2_X1 U10651 ( .A1(n8058), .A2(SI_7_), .ZN(n8059) );
  INV_X1 U10652 ( .A(n8166), .ZN(n8061) );
  MUX2_X1 U10653 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n12325), .Z(n8064) );
  INV_X1 U10654 ( .A(n8174), .ZN(n8063) );
  MUX2_X1 U10655 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10885), .Z(n8066) );
  XNOR2_X1 U10656 ( .A(n8066), .B(SI_10_), .ZN(n8184) );
  INV_X1 U10657 ( .A(n8184), .ZN(n8065) );
  NAND2_X1 U10658 ( .A1(n8066), .A2(SI_10_), .ZN(n8067) );
  MUX2_X1 U10659 ( .A(n10201), .B(n10194), .S(n8050), .Z(n8068) );
  INV_X1 U10660 ( .A(n8068), .ZN(n8069) );
  NAND2_X1 U10661 ( .A1(n8069), .A2(SI_11_), .ZN(n8070) );
  NAND2_X1 U10662 ( .A1(n8071), .A2(n8070), .ZN(n8189) );
  MUX2_X1 U10663 ( .A(n10316), .B(n10309), .S(n12325), .Z(n8075) );
  INV_X1 U10664 ( .A(n8075), .ZN(n8076) );
  NAND2_X1 U10665 ( .A1(n8076), .A2(SI_13_), .ZN(n8077) );
  MUX2_X1 U10666 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n12325), .Z(n8220) );
  INV_X1 U10667 ( .A(n8220), .ZN(n8079) );
  NOR2_X1 U10668 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), 
        .ZN(n8083) );
  NAND4_X1 U10669 ( .A1(n8086), .A2(n8383), .A3(n8417), .A4(n8401), .ZN(n8091)
         );
  INV_X1 U10670 ( .A(n8091), .ZN(n8087) );
  XNOR2_X1 U10671 ( .A(P2_IR_REG_31__SCAN_IN), .B(P2_IR_REG_27__SCAN_IN), .ZN(
        n8088) );
  NAND2_X1 U10672 ( .A1(n8090), .A2(n8089), .ZN(n8092) );
  NAND2_X2 U10673 ( .A1(n8111), .A2(n10885), .ZN(n8121) );
  INV_X2 U10674 ( .A(n8121), .ZN(n8264) );
  NAND2_X1 U10675 ( .A1(n12244), .A2(n8264), .ZN(n8105) );
  INV_X1 U10676 ( .A(n8099), .ZN(n8100) );
  NAND2_X1 U10677 ( .A1(n8214), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8103) );
  XNOR2_X1 U10678 ( .A(n8103), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11292) );
  AOI22_X1 U10679 ( .A1(n8235), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8274), 
        .B2(n11292), .ZN(n8104) );
  INV_X1 U10680 ( .A(n14481), .ZN(n14325) );
  XNOR2_X1 U10681 ( .A(n8106), .B(n10101), .ZN(n8108) );
  INV_X1 U10682 ( .A(n8109), .ZN(n8115) );
  OR2_X1 U10683 ( .A1(n8111), .A2(n10433), .ZN(n8110) );
  INV_X1 U10684 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8112) );
  XNOR2_X1 U10685 ( .A(n9159), .B(n9028), .ZN(n14596) );
  MUX2_X1 U10686 ( .A(n8112), .B(n14596), .S(n8111), .Z(n15660) );
  XNOR2_X1 U10687 ( .A(n8113), .B(n8114), .ZN(n10689) );
  NAND2_X1 U10688 ( .A1(n8115), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8116) );
  MUX2_X1 U10689 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8116), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n8118) );
  NAND2_X1 U10690 ( .A1(n8118), .A2(n8117), .ZN(n13964) );
  OAI211_X2 U10691 ( .C1(n8121), .C2(n10689), .A(n8120), .B(n8119), .ZN(n11934) );
  NAND2_X1 U10692 ( .A1(n8117), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8122) );
  MUX2_X1 U10693 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8122), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8123) );
  OR2_X1 U10694 ( .A1(n8117), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n8128) );
  NAND2_X1 U10695 ( .A1(n8123), .A2(n8128), .ZN(n15642) );
  XNOR2_X1 U10696 ( .A(n8124), .B(SI_3_), .ZN(n8132) );
  NAND2_X1 U10697 ( .A1(n8264), .A2(n10886), .ZN(n8126) );
  OR2_X1 U10698 ( .A1(n8376), .A2(n10056), .ZN(n8125) );
  OAI211_X1 U10699 ( .C1(n10428), .C2(n15642), .A(n8126), .B(n8125), .ZN(n8465) );
  NAND2_X1 U10700 ( .A1(n8128), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8127) );
  MUX2_X1 U10701 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8127), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8131) );
  INV_X1 U10702 ( .A(n8128), .ZN(n8130) );
  NAND2_X1 U10703 ( .A1(n8130), .A2(n8129), .ZN(n8143) );
  NAND2_X1 U10704 ( .A1(n8131), .A2(n8143), .ZN(n13977) );
  INV_X1 U10705 ( .A(n8132), .ZN(n8133) );
  NAND2_X1 U10706 ( .A1(n8135), .A2(n8134), .ZN(n8137) );
  XNOR2_X1 U10707 ( .A(n8137), .B(n8136), .ZN(n10899) );
  NAND2_X1 U10708 ( .A1(n10899), .A2(n8264), .ZN(n8139) );
  OR2_X1 U10709 ( .A1(n8376), .A2(n10067), .ZN(n8138) );
  NAND2_X1 U10710 ( .A1(n8141), .A2(n8140), .ZN(n8152) );
  XNOR2_X1 U10711 ( .A(n8142), .B(SI_5_), .ZN(n8150) );
  XNOR2_X1 U10712 ( .A(n8152), .B(n8150), .ZN(n11019) );
  NAND2_X1 U10713 ( .A1(n11019), .A2(n8264), .ZN(n8147) );
  NAND2_X1 U10714 ( .A1(n8143), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8144) );
  MUX2_X1 U10715 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8144), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n8145) );
  AND2_X1 U10716 ( .A1(n8145), .A2(n8098), .ZN(n13990) );
  AOI22_X1 U10717 ( .A1(n8235), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8274), .B2(
        n13990), .ZN(n8146) );
  NAND2_X1 U10718 ( .A1(n8147), .A2(n8146), .ZN(n11224) );
  INV_X1 U10719 ( .A(n8150), .ZN(n8151) );
  NAND2_X1 U10720 ( .A1(n8152), .A2(n8151), .ZN(n8154) );
  NAND2_X1 U10721 ( .A1(n8154), .A2(n8153), .ZN(n8156) );
  NAND2_X1 U10722 ( .A1(n11189), .A2(n8264), .ZN(n8159) );
  NAND2_X1 U10723 ( .A1(n8098), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8157) );
  XNOR2_X1 U10724 ( .A(n8157), .B(P2_IR_REG_6__SCAN_IN), .ZN(n14004) );
  AOI22_X1 U10725 ( .A1(n8235), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8274), .B2(
        n14004), .ZN(n8158) );
  NAND2_X1 U10726 ( .A1(n8159), .A2(n8158), .ZN(n11661) );
  XNOR2_X1 U10727 ( .A(n8161), .B(n8160), .ZN(n11439) );
  NAND2_X1 U10728 ( .A1(n11439), .A2(n8264), .ZN(n8165) );
  INV_X1 U10729 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8162) );
  NAND2_X1 U10730 ( .A1(n7349), .A2(n8162), .ZN(n8168) );
  NAND2_X1 U10731 ( .A1(n8168), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8163) );
  XNOR2_X1 U10732 ( .A(n8163), .B(P2_IR_REG_7__SCAN_IN), .ZN(n14020) );
  AOI22_X1 U10733 ( .A1(n8235), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8274), .B2(
        n14020), .ZN(n8164) );
  XNOR2_X1 U10734 ( .A(n8167), .B(n8166), .ZN(n11510) );
  NAND2_X1 U10735 ( .A1(n11510), .A2(n8264), .ZN(n8173) );
  NAND2_X1 U10736 ( .A1(n8170), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8169) );
  MUX2_X1 U10737 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8169), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n8171) );
  NAND2_X1 U10738 ( .A1(n8171), .A2(n8177), .ZN(n14033) );
  INV_X1 U10739 ( .A(n14033), .ZN(n14029) );
  AOI22_X1 U10740 ( .A1(n8235), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n14029), 
        .B2(n8274), .ZN(n8172) );
  INV_X1 U10741 ( .A(n14519), .ZN(n11696) );
  XNOR2_X1 U10742 ( .A(n8175), .B(n8174), .ZN(n11515) );
  NAND2_X1 U10743 ( .A1(n11515), .A2(n8264), .ZN(n8183) );
  NAND2_X1 U10744 ( .A1(n8177), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8176) );
  MUX2_X1 U10745 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8176), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n8180) );
  INV_X1 U10746 ( .A(n8177), .ZN(n8179) );
  INV_X1 U10747 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8178) );
  NAND2_X1 U10748 ( .A1(n8179), .A2(n8178), .ZN(n8191) );
  NAND2_X1 U10749 ( .A1(n8180), .A2(n8191), .ZN(n10484) );
  OAI22_X1 U10750 ( .A1(n10484), .A2(n10428), .B1(n8376), .B2(n10168), .ZN(
        n8181) );
  INV_X1 U10751 ( .A(n8181), .ZN(n8182) );
  XNOR2_X1 U10752 ( .A(n8185), .B(n8184), .ZN(n11493) );
  NAND2_X1 U10753 ( .A1(n11493), .A2(n8264), .ZN(n8188) );
  NAND2_X1 U10754 ( .A1(n8191), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8186) );
  XNOR2_X1 U10755 ( .A(n8186), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10724) );
  AOI22_X1 U10756 ( .A1(n10724), .A2(n8274), .B1(n8235), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n8187) );
  INV_X1 U10757 ( .A(n14367), .ZN(n14504) );
  OAI21_X1 U10758 ( .B1(n8191), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8192) );
  XNOR2_X1 U10759 ( .A(n8192), .B(P2_IR_REG_11__SCAN_IN), .ZN(n14052) );
  AOI22_X1 U10760 ( .A1(n14052), .A2(n8274), .B1(n8235), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8193) );
  XNOR2_X1 U10761 ( .A(n8194), .B(n8029), .ZN(n12070) );
  NAND2_X1 U10762 ( .A1(n12070), .A2(n8264), .ZN(n8201) );
  INV_X1 U10763 ( .A(n8195), .ZN(n8196) );
  NAND2_X1 U10764 ( .A1(n8196), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8197) );
  MUX2_X1 U10765 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8197), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8199) );
  INV_X1 U10766 ( .A(n8198), .ZN(n8203) );
  AOI22_X1 U10767 ( .A1(n8235), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8274), 
        .B2(n10495), .ZN(n8200) );
  XNOR2_X1 U10768 ( .A(n8202), .B(n8019), .ZN(n12153) );
  NAND2_X1 U10769 ( .A1(n12153), .A2(n8264), .ZN(n8207) );
  NAND2_X1 U10770 ( .A1(n8203), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8204) );
  MUX2_X1 U10771 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8204), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8205) );
  NAND2_X1 U10772 ( .A1(n8205), .A2(n8214), .ZN(n10876) );
  INV_X1 U10773 ( .A(n10876), .ZN(n10843) );
  AOI22_X1 U10774 ( .A1(n8235), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8274), 
        .B2(n10843), .ZN(n8206) );
  INV_X1 U10775 ( .A(n8219), .ZN(n8209) );
  NAND2_X1 U10776 ( .A1(n8209), .A2(SI_14_), .ZN(n8210) );
  NOR2_X1 U10777 ( .A1(n8211), .A2(SI_15_), .ZN(n8221) );
  INV_X1 U10778 ( .A(n8221), .ZN(n8212) );
  NAND2_X1 U10779 ( .A1(n8222), .A2(n8212), .ZN(n8213) );
  NAND2_X1 U10780 ( .A1(n12250), .A2(n8264), .ZN(n8217) );
  NAND2_X1 U10781 ( .A1(n8229), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8215) );
  XNOR2_X1 U10782 ( .A(n8215), .B(P2_IR_REG_15__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U10783 ( .A1(n8235), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8274), 
        .B2(n11830), .ZN(n8216) );
  NAND2_X1 U10784 ( .A1(n8220), .A2(SI_14_), .ZN(n8218) );
  NOR2_X1 U10785 ( .A1(n8220), .A2(SI_14_), .ZN(n8223) );
  AOI21_X1 U10786 ( .B1(n8223), .B2(n8222), .A(n8221), .ZN(n8224) );
  MUX2_X1 U10787 ( .A(n10545), .B(n15888), .S(n10885), .Z(n8226) );
  INV_X1 U10788 ( .A(n8226), .ZN(n8227) );
  NAND2_X1 U10789 ( .A1(n8227), .A2(SI_16_), .ZN(n8228) );
  XNOR2_X1 U10790 ( .A(n8238), .B(n8024), .ZN(n12261) );
  NAND2_X1 U10791 ( .A1(n12261), .A2(n8264), .ZN(n8237) );
  INV_X1 U10792 ( .A(n8233), .ZN(n8230) );
  NAND2_X1 U10793 ( .A1(n8230), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8231) );
  MUX2_X1 U10794 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8231), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n8234) );
  INV_X1 U10795 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8232) );
  AOI22_X1 U10796 ( .A1(n11886), .A2(n8274), .B1(n8235), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n8236) );
  MUX2_X1 U10797 ( .A(n16042), .B(n10644), .S(n12325), .Z(n8240) );
  INV_X1 U10798 ( .A(n8240), .ZN(n8241) );
  NAND2_X1 U10799 ( .A1(n8241), .A2(SI_17_), .ZN(n8242) );
  NAND2_X1 U10800 ( .A1(n12272), .A2(n8264), .ZN(n8248) );
  NAND2_X1 U10801 ( .A1(n8271), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8243) );
  MUX2_X1 U10802 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8243), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8245) );
  NAND2_X1 U10803 ( .A1(n8244), .A2(n8265), .ZN(n8251) );
  NAND2_X1 U10804 ( .A1(n8245), .A2(n8251), .ZN(n11836) );
  OAI22_X1 U10805 ( .A1(n11836), .A2(n10428), .B1(n8376), .B2(n10644), .ZN(
        n8246) );
  INV_X1 U10806 ( .A(n8246), .ZN(n8247) );
  MUX2_X1 U10807 ( .A(n11107), .B(n15896), .S(n10885), .Z(n8277) );
  XNOR2_X1 U10808 ( .A(n8256), .B(n8277), .ZN(n12282) );
  NAND2_X1 U10809 ( .A1(n12282), .A2(n8264), .ZN(n8255) );
  NAND2_X1 U10810 ( .A1(n8251), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8252) );
  XNOR2_X1 U10811 ( .A(n8252), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14067) );
  NOR2_X1 U10812 ( .A1(n8376), .A2(n15896), .ZN(n8253) );
  AOI21_X1 U10813 ( .B1(n14067), .B2(n8274), .A(n8253), .ZN(n8254) );
  INV_X1 U10814 ( .A(n8277), .ZN(n8280) );
  NAND2_X1 U10815 ( .A1(n8256), .A2(n8280), .ZN(n8259) );
  INV_X1 U10816 ( .A(n8279), .ZN(n8257) );
  NAND2_X1 U10817 ( .A1(n8257), .A2(SI_18_), .ZN(n8258) );
  NAND2_X1 U10818 ( .A1(n8259), .A2(n8258), .ZN(n8263) );
  INV_X1 U10819 ( .A(n8260), .ZN(n8261) );
  NAND2_X1 U10820 ( .A1(n8261), .A2(n10630), .ZN(n8281) );
  NAND2_X1 U10821 ( .A1(n8283), .A2(n8281), .ZN(n8262) );
  NAND2_X1 U10822 ( .A1(n12293), .A2(n8264), .ZN(n8276) );
  XNOR2_X1 U10823 ( .A(P2_IR_REG_19__SCAN_IN), .B(P2_IR_REG_31__SCAN_IN), .ZN(
        n8268) );
  INV_X1 U10824 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8266) );
  NAND3_X1 U10825 ( .A1(n8266), .A2(n8265), .A3(P2_IR_REG_19__SCAN_IN), .ZN(
        n8267) );
  INV_X1 U10826 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n15836) );
  NOR2_X1 U10827 ( .A1(n8376), .A2(n15836), .ZN(n8273) );
  AOI21_X1 U10828 ( .B1(n8775), .B2(n8274), .A(n8273), .ZN(n8275) );
  OAI21_X1 U10829 ( .B1(n8277), .B2(n10549), .A(n8283), .ZN(n8278) );
  INV_X1 U10830 ( .A(n8281), .ZN(n8282) );
  XNOR2_X1 U10831 ( .A(n8301), .B(SI_20_), .ZN(n8289) );
  MUX2_X1 U10832 ( .A(n11281), .B(n11284), .S(n12325), .Z(n8297) );
  XNOR2_X1 U10833 ( .A(n8289), .B(n8297), .ZN(n12301) );
  NAND2_X1 U10834 ( .A1(n12301), .A2(n8264), .ZN(n8288) );
  OR2_X1 U10835 ( .A1(n8376), .A2(n11284), .ZN(n8287) );
  INV_X1 U10836 ( .A(n8297), .ZN(n8296) );
  NAND2_X1 U10837 ( .A1(n8289), .A2(n8296), .ZN(n8291) );
  OR2_X1 U10838 ( .A1(n8301), .A2(n11250), .ZN(n8290) );
  NAND2_X1 U10839 ( .A1(n8291), .A2(n8290), .ZN(n8293) );
  XNOR2_X1 U10840 ( .A(n8298), .B(SI_21_), .ZN(n8292) );
  NAND2_X1 U10841 ( .A1(n12312), .A2(n8264), .ZN(n8295) );
  INV_X1 U10842 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n15958) );
  OR2_X1 U10843 ( .A1(n8376), .A2(n15958), .ZN(n8294) );
  NOR2_X1 U10844 ( .A1(n8297), .A2(n11250), .ZN(n8299) );
  AOI22_X1 U10845 ( .A1(n8299), .A2(n8025), .B1(n8298), .B2(SI_21_), .ZN(n8300) );
  MUX2_X1 U10846 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n10885), .Z(n8315) );
  XNOR2_X1 U10847 ( .A(n12326), .B(n8315), .ZN(n11490) );
  NAND2_X1 U10848 ( .A1(n11490), .A2(n8264), .ZN(n8303) );
  INV_X1 U10849 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n15835) );
  OR2_X1 U10850 ( .A1(n8376), .A2(n15835), .ZN(n8302) );
  INV_X1 U10851 ( .A(n12326), .ZN(n8304) );
  NAND2_X1 U10852 ( .A1(n8304), .A2(n8315), .ZN(n8306) );
  NAND2_X1 U10853 ( .A1(n8314), .A2(SI_22_), .ZN(n8305) );
  XNOR2_X1 U10854 ( .A(n8317), .B(SI_23_), .ZN(n8307) );
  NAND2_X1 U10855 ( .A1(n12340), .A2(n8264), .ZN(n8310) );
  INV_X1 U10856 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11743) );
  OR2_X1 U10857 ( .A1(n8376), .A2(n11743), .ZN(n8309) );
  INV_X1 U10858 ( .A(n8317), .ZN(n8311) );
  NAND2_X1 U10859 ( .A1(n8311), .A2(n11314), .ZN(n8318) );
  OAI21_X1 U10860 ( .B1(SI_22_), .B2(n8315), .A(n8318), .ZN(n8312) );
  INV_X1 U10861 ( .A(n8312), .ZN(n8313) );
  INV_X1 U10862 ( .A(n8315), .ZN(n8316) );
  INV_X1 U10863 ( .A(SI_22_), .ZN(n9469) );
  NOR2_X1 U10864 ( .A1(n8316), .A2(n9469), .ZN(n8319) );
  AOI22_X1 U10865 ( .A1(n8319), .A2(n8318), .B1(n8317), .B2(SI_23_), .ZN(n8320) );
  INV_X1 U10866 ( .A(n8325), .ZN(n8321) );
  NAND2_X1 U10867 ( .A1(n12360), .A2(n8264), .ZN(n8323) );
  INV_X1 U10868 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11790) );
  OR2_X1 U10869 ( .A1(n8376), .A2(n11790), .ZN(n8322) );
  NAND2_X1 U10870 ( .A1(n8326), .A2(SI_24_), .ZN(n8327) );
  MUX2_X1 U10871 ( .A(n11894), .B(n11898), .S(n12325), .Z(n8329) );
  INV_X1 U10872 ( .A(SI_25_), .ZN(n11891) );
  INV_X1 U10873 ( .A(n8329), .ZN(n8330) );
  NAND2_X1 U10874 ( .A1(n8330), .A2(SI_25_), .ZN(n8331) );
  NAND2_X1 U10875 ( .A1(n8336), .A2(n8331), .ZN(n8334) );
  XNOR2_X1 U10876 ( .A(n8335), .B(n8334), .ZN(n12350) );
  NAND2_X1 U10877 ( .A1(n12350), .A2(n8264), .ZN(n8333) );
  OR2_X1 U10878 ( .A1(n8376), .A2(n11898), .ZN(n8332) );
  INV_X1 U10879 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n12586) );
  XNOR2_X1 U10880 ( .A(n8340), .B(SI_26_), .ZN(n8337) );
  NAND2_X1 U10881 ( .A1(n12372), .A2(n8264), .ZN(n8339) );
  OR2_X1 U10882 ( .A1(n8376), .A2(n16023), .ZN(n8338) );
  NAND2_X1 U10883 ( .A1(n8343), .A2(n8342), .ZN(n8349) );
  INV_X1 U10884 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15380) );
  INV_X1 U10885 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12239) );
  MUX2_X1 U10886 ( .A(n15380), .B(n12239), .S(n10885), .Z(n8347) );
  XNOR2_X1 U10887 ( .A(n8347), .B(SI_27_), .ZN(n8344) );
  NAND2_X1 U10888 ( .A1(n12394), .A2(n8264), .ZN(n8346) );
  OR2_X1 U10889 ( .A1(n8376), .A2(n12239), .ZN(n8345) );
  INV_X1 U10890 ( .A(n8347), .ZN(n8350) );
  NOR2_X1 U10891 ( .A1(n8350), .A2(SI_27_), .ZN(n8348) );
  NAND2_X1 U10892 ( .A1(n8350), .A2(SI_27_), .ZN(n8351) );
  MUX2_X1 U10893 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n12325), .Z(n8354) );
  XNOR2_X1 U10894 ( .A(n8354), .B(SI_28_), .ZN(n8355) );
  NAND2_X1 U10895 ( .A1(n12461), .A2(n8264), .ZN(n8353) );
  INV_X1 U10896 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9085) );
  OR2_X1 U10897 ( .A1(n8376), .A2(n9085), .ZN(n8352) );
  INV_X1 U10898 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15376) );
  INV_X1 U10899 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14589) );
  XNOR2_X1 U10900 ( .A(n8361), .B(SI_29_), .ZN(n8359) );
  NAND2_X1 U10901 ( .A1(n14586), .A2(n8264), .ZN(n8358) );
  OR2_X1 U10902 ( .A1(n8376), .A2(n14589), .ZN(n8357) );
  NAND2_X1 U10903 ( .A1(n8360), .A2(n8359), .ZN(n8363) );
  INV_X1 U10904 ( .A(SI_29_), .ZN(n12241) );
  NAND2_X1 U10905 ( .A1(n8361), .A2(n12241), .ZN(n8362) );
  INV_X1 U10906 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n15371) );
  INV_X1 U10907 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12595) );
  MUX2_X1 U10908 ( .A(n15371), .B(n12595), .S(n12325), .Z(n8369) );
  XNOR2_X1 U10909 ( .A(n8369), .B(SI_30_), .ZN(n8367) );
  NAND2_X1 U10910 ( .A1(n12811), .A2(n8264), .ZN(n8365) );
  OR2_X1 U10911 ( .A1(n8376), .A2(n12595), .ZN(n8364) );
  INV_X1 U10912 ( .A(n8366), .ZN(n8368) );
  NAND2_X1 U10913 ( .A1(n8368), .A2(n8367), .ZN(n8372) );
  INV_X1 U10914 ( .A(n8369), .ZN(n8370) );
  NAND2_X1 U10915 ( .A1(n8370), .A2(SI_30_), .ZN(n8371) );
  XNOR2_X1 U10916 ( .A(n8373), .B(SI_31_), .ZN(n8374) );
  NAND2_X1 U10917 ( .A1(n14579), .A2(n8264), .ZN(n8378) );
  INV_X1 U10918 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n14582) );
  OR2_X1 U10919 ( .A1(n8376), .A2(n14582), .ZN(n8377) );
  XNOR2_X1 U10920 ( .A(n14092), .B(n8995), .ZN(n8389) );
  NAND2_X1 U10921 ( .A1(n8382), .A2(n8383), .ZN(n8380) );
  NAND2_X1 U10922 ( .A1(n8380), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8379) );
  MUX2_X1 U10923 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8379), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n8381) );
  INV_X1 U10924 ( .A(n8382), .ZN(n8387) );
  NAND2_X2 U10925 ( .A1(n11491), .A2(n11359), .ZN(n15659) );
  OR2_X4 U10926 ( .A1(n15659), .A2(n9010), .ZN(n14338) );
  NAND2_X1 U10927 ( .A1(n8393), .A2(n8391), .ZN(n14580) );
  XNOR2_X2 U10928 ( .A(n8392), .B(n14581), .ZN(n8395) );
  XNOR2_X2 U10929 ( .A(n8394), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8436) );
  INV_X1 U10930 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n15880) );
  NAND2_X2 U10931 ( .A1(n8395), .A2(n14587), .ZN(n8468) );
  NAND2_X1 U10932 ( .A1(n8757), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8397) );
  NAND2_X1 U10933 ( .A1(n8756), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8396) );
  OAI211_X1 U10934 ( .C1(n8944), .C2(n15880), .A(n8397), .B(n8396), .ZN(n13927) );
  INV_X1 U10935 ( .A(n11491), .ZN(n8782) );
  NAND2_X1 U10936 ( .A1(n10427), .A2(n8398), .ZN(n13917) );
  INV_X1 U10937 ( .A(P2_B_REG_SCAN_IN), .ZN(n15938) );
  NOR2_X1 U10938 ( .A1(n8399), .A2(n15938), .ZN(n8400) );
  NOR2_X1 U10939 ( .A1(n13917), .A2(n8400), .ZN(n9915) );
  AND2_X1 U10940 ( .A1(n13927), .A2(n9915), .ZN(n14089) );
  NOR2_X1 U10941 ( .A1(n14088), .A2(n14089), .ZN(n14406) );
  OAI21_X1 U10942 ( .B1(n8416), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8402) );
  MUX2_X1 U10943 ( .A(n8402), .B(P2_IR_REG_31__SCAN_IN), .S(n8401), .Z(n8403)
         );
  NAND2_X1 U10944 ( .A1(n8405), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8404) );
  MUX2_X1 U10945 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8404), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8406) );
  NAND2_X1 U10946 ( .A1(n8408), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8407) );
  MUX2_X1 U10947 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8407), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8412) );
  INV_X1 U10948 ( .A(n8408), .ZN(n8410) );
  INV_X1 U10949 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8409) );
  NAND2_X1 U10950 ( .A1(n8410), .A2(n8409), .ZN(n8411) );
  INV_X1 U10951 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15698) );
  NAND2_X1 U10952 ( .A1(n15670), .A2(n15698), .ZN(n8415) );
  NAND2_X1 U10953 ( .A1(n11788), .A2(n12119), .ZN(n8414) );
  NAND2_X1 U10954 ( .A1(n8415), .A2(n8414), .ZN(n10005) );
  NAND2_X1 U10955 ( .A1(n14086), .A2(n11283), .ZN(n10038) );
  NAND2_X1 U10956 ( .A1(n8416), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8418) );
  NAND2_X1 U10957 ( .A1(n10426), .A2(n9929), .ZN(n8419) );
  INV_X1 U10958 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15700) );
  NAND2_X1 U10959 ( .A1(n15670), .A2(n15700), .ZN(n8421) );
  NAND2_X1 U10960 ( .A1(n12119), .A2(n11895), .ZN(n8420) );
  NOR4_X1 U10961 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n8425) );
  NOR4_X1 U10962 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8424) );
  INV_X1 U10963 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15936) );
  INV_X1 U10964 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n15983) );
  INV_X1 U10965 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n16091) );
  INV_X1 U10966 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n16004) );
  NAND4_X1 U10967 ( .A1(n15936), .A2(n15983), .A3(n16091), .A4(n16004), .ZN(
        n8422) );
  NOR2_X1 U10968 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n8422), .ZN(n15871) );
  NOR4_X1 U10969 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n8423) );
  NAND4_X1 U10970 ( .A1(n8425), .A2(n8424), .A3(n15871), .A4(n8423), .ZN(n8430) );
  NOR4_X1 U10971 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n8428) );
  NOR4_X1 U10972 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n8427) );
  NOR4_X1 U10973 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n8426) );
  INV_X1 U10974 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n15674) );
  NAND4_X1 U10975 ( .A1(n8428), .A2(n8427), .A3(n8426), .A4(n15674), .ZN(n8429) );
  OAI21_X1 U10976 ( .B1(n8430), .B2(n8429), .A(n15670), .ZN(n10004) );
  AND2_X1 U10977 ( .A1(n10004), .A2(n10035), .ZN(n8431) );
  MUX2_X1 U10978 ( .A(n8432), .B(n14406), .S(n15743), .Z(n8435) );
  NAND2_X1 U10979 ( .A1(n8995), .A2(n8433), .ZN(n8434) );
  NAND2_X1 U10980 ( .A1(n8435), .A2(n8434), .ZN(P2_U3498) );
  INV_X1 U10981 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8749) );
  INV_X1 U10982 ( .A(n8455), .ZN(n8676) );
  NAND2_X1 U10983 ( .A1(n8676), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8443) );
  INV_X1 U10984 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11977) );
  NAND2_X4 U10985 ( .A1(n8437), .A2(n8436), .ZN(n8739) );
  INV_X1 U10986 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8438) );
  INV_X1 U10987 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n8439) );
  NAND4_X4 U10988 ( .A1(n8443), .A2(n8442), .A3(n8441), .A4(n8440), .ZN(n8781)
         );
  INV_X1 U10989 ( .A(n8691), .ZN(n8452) );
  INV_X1 U10990 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n8444) );
  INV_X1 U10991 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n8445) );
  OR2_X1 U10992 ( .A1(n8455), .A2(n8445), .ZN(n8450) );
  INV_X1 U10993 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n8446) );
  OR2_X1 U10994 ( .A1(n8739), .A2(n8446), .ZN(n8449) );
  INV_X1 U10995 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n8447) );
  INV_X1 U10996 ( .A(n15660), .ZN(n10558) );
  NAND2_X1 U10997 ( .A1(n11968), .A2(n8453), .ZN(n10575) );
  NAND2_X1 U10998 ( .A1(n8757), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8459) );
  INV_X1 U10999 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n13958) );
  OR2_X1 U11000 ( .A1(n8739), .A2(n13958), .ZN(n8458) );
  INV_X1 U11001 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n8454) );
  OR2_X1 U11002 ( .A1(n8944), .A2(n8454), .ZN(n8457) );
  INV_X1 U11003 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10435) );
  OR2_X1 U11004 ( .A1(n8945), .A2(n10435), .ZN(n8456) );
  OR2_X1 U11005 ( .A1(n13956), .A2(n11934), .ZN(n8460) );
  NAND2_X1 U11006 ( .A1(n10576), .A2(n8460), .ZN(n11704) );
  NAND2_X1 U11007 ( .A1(n8757), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8464) );
  OR2_X1 U11008 ( .A1(n8739), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8463) );
  INV_X1 U11009 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10417) );
  INV_X1 U11010 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11714) );
  OR2_X1 U11011 ( .A1(n8945), .A2(n11714), .ZN(n8461) );
  INV_X1 U11012 ( .A(n8465), .ZN(n15717) );
  XNOR2_X1 U11013 ( .A(n13955), .B(n15717), .ZN(n9011) );
  NAND2_X1 U11014 ( .A1(n11704), .A2(n9011), .ZN(n8467) );
  OR2_X1 U11015 ( .A1(n13955), .A2(n11717), .ZN(n8466) );
  NAND2_X1 U11016 ( .A1(n8756), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8474) );
  INV_X1 U11017 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n8469) );
  OR2_X1 U11018 ( .A1(n8468), .A2(n8469), .ZN(n8473) );
  XNOR2_X1 U11019 ( .A(P2_REG3_REG_3__SCAN_IN), .B(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n11624) );
  OR2_X1 U11020 ( .A1(n8739), .A2(n11624), .ZN(n8472) );
  INV_X1 U11021 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n8470) );
  OR2_X1 U11022 ( .A1(n8944), .A2(n8470), .ZN(n8471) );
  XNOR2_X1 U11023 ( .A(n13954), .B(n11625), .ZN(n10790) );
  OR2_X1 U11024 ( .A1(n13954), .A2(n10851), .ZN(n8475) );
  NAND2_X1 U11025 ( .A1(n8756), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8484) );
  INV_X1 U11026 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n8476) );
  OR2_X1 U11027 ( .A1(n8468), .A2(n8476), .ZN(n8483) );
  NAND3_X1 U11028 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n8489) );
  INV_X1 U11029 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8478) );
  NAND2_X1 U11030 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n8477) );
  NAND2_X1 U11031 ( .A1(n8478), .A2(n8477), .ZN(n8479) );
  NAND2_X1 U11032 ( .A1(n8489), .A2(n8479), .ZN(n11956) );
  OR2_X1 U11033 ( .A1(n8739), .A2(n11956), .ZN(n8482) );
  INV_X1 U11034 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n8480) );
  OR2_X1 U11035 ( .A1(n8944), .A2(n8480), .ZN(n8481) );
  NAND4_X1 U11036 ( .A1(n8484), .A2(n8483), .A3(n8482), .A4(n8481), .ZN(n13953) );
  NAND2_X1 U11037 ( .A1(n11224), .A2(n13953), .ZN(n8485) );
  OR2_X1 U11038 ( .A1(n11224), .A2(n13953), .ZN(n8486) );
  NAND2_X1 U11039 ( .A1(n8757), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8495) );
  INV_X1 U11040 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10444) );
  OR2_X1 U11041 ( .A1(n8945), .A2(n10444), .ZN(n8494) );
  INV_X1 U11042 ( .A(n8489), .ZN(n8487) );
  NAND2_X1 U11043 ( .A1(n8487), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8504) );
  INV_X1 U11044 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U11045 ( .A1(n8489), .A2(n8488), .ZN(n8490) );
  NAND2_X1 U11046 ( .A1(n8504), .A2(n8490), .ZN(n11663) );
  OR2_X1 U11047 ( .A1(n8739), .A2(n11663), .ZN(n8493) );
  INV_X1 U11048 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n8491) );
  OR2_X1 U11049 ( .A1(n8944), .A2(n8491), .ZN(n8492) );
  NAND4_X1 U11050 ( .A1(n8495), .A2(n8494), .A3(n8493), .A4(n8492), .ZN(n13952) );
  XNOR2_X1 U11051 ( .A(n11661), .B(n13952), .ZN(n11656) );
  NAND2_X1 U11052 ( .A1(n8757), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8501) );
  INV_X1 U11053 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n16075) );
  OR2_X1 U11054 ( .A1(n8455), .A2(n16075), .ZN(n8500) );
  INV_X1 U11055 ( .A(n8504), .ZN(n8497) );
  INV_X1 U11056 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8516) );
  XNOR2_X1 U11057 ( .A(n8517), .B(n8516), .ZN(n11695) );
  OR2_X1 U11058 ( .A1(n8739), .A2(n11695), .ZN(n8499) );
  INV_X1 U11059 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11693) );
  OR2_X1 U11060 ( .A1(n8945), .A2(n11693), .ZN(n8498) );
  NAND4_X1 U11061 ( .A1(n8501), .A2(n8500), .A3(n8499), .A4(n8498), .ZN(n13950) );
  NAND2_X1 U11062 ( .A1(n8757), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8509) );
  INV_X1 U11063 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n8502) );
  OR2_X1 U11064 ( .A1(n8944), .A2(n8502), .ZN(n8508) );
  INV_X1 U11065 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8503) );
  NAND2_X1 U11066 ( .A1(n8504), .A2(n8503), .ZN(n8505) );
  NAND2_X1 U11067 ( .A1(n8517), .A2(n8505), .ZN(n11989) );
  OR2_X1 U11068 ( .A1(n8739), .A2(n11989), .ZN(n8507) );
  INV_X1 U11069 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11996) );
  OR2_X1 U11070 ( .A1(n8945), .A2(n11996), .ZN(n8506) );
  NAND4_X1 U11071 ( .A1(n8509), .A2(n8508), .A3(n8507), .A4(n8506), .ZN(n13951) );
  NAND2_X1 U11072 ( .A1(n14519), .A2(n13950), .ZN(n8510) );
  NAND2_X1 U11073 ( .A1(n8511), .A2(n8510), .ZN(n8512) );
  AND2_X1 U11074 ( .A1(n11661), .A2(n13952), .ZN(n11681) );
  INV_X1 U11075 ( .A(n8512), .ZN(n14384) );
  NOR2_X1 U11076 ( .A1(n11683), .A2(n13951), .ZN(n8513) );
  OR2_X1 U11077 ( .A1(n11688), .A2(n8513), .ZN(n14385) );
  NAND2_X1 U11078 ( .A1(n8756), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8524) );
  INV_X1 U11079 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8514) );
  OR2_X1 U11080 ( .A1(n8468), .A2(n8514), .ZN(n8523) );
  INV_X1 U11081 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8515) );
  OAI21_X1 U11082 ( .B1(n8517), .B2(n8516), .A(n8515), .ZN(n8520) );
  INV_X1 U11083 ( .A(n8517), .ZN(n8519) );
  NAND2_X1 U11084 ( .A1(n8520), .A2(n8530), .ZN(n14397) );
  OR2_X1 U11085 ( .A1(n8739), .A2(n14397), .ZN(n8522) );
  INV_X1 U11086 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n14512) );
  OR2_X1 U11087 ( .A1(n8944), .A2(n14512), .ZN(n8521) );
  NAND4_X1 U11088 ( .A1(n8524), .A2(n8523), .A3(n8522), .A4(n8521), .ZN(n13949) );
  INV_X1 U11089 ( .A(n13949), .ZN(n11645) );
  NAND2_X1 U11090 ( .A1(n14575), .A2(n11645), .ZN(n14373) );
  NAND2_X1 U11091 ( .A1(n8707), .A2(n14373), .ZN(n14387) );
  INV_X1 U11092 ( .A(n14387), .ZN(n14391) );
  AOI21_X1 U11093 ( .B1(n14384), .B2(n14385), .A(n14391), .ZN(n8525) );
  NAND2_X1 U11094 ( .A1(n14575), .A2(n13949), .ZN(n8526) );
  NAND2_X1 U11095 ( .A1(n8757), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8536) );
  INV_X1 U11096 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8527) );
  OR2_X1 U11097 ( .A1(n8945), .A2(n8527), .ZN(n8535) );
  INV_X1 U11098 ( .A(n8530), .ZN(n8528) );
  INV_X1 U11099 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8529) );
  NAND2_X1 U11100 ( .A1(n8530), .A2(n8529), .ZN(n8531) );
  NAND2_X1 U11101 ( .A1(n8541), .A2(n8531), .ZN(n14365) );
  OR2_X1 U11102 ( .A1(n8739), .A2(n14365), .ZN(n8534) );
  INV_X1 U11103 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8532) );
  OR2_X1 U11104 ( .A1(n8944), .A2(n8532), .ZN(n8533) );
  NAND4_X1 U11105 ( .A1(n8536), .A2(n8535), .A3(n8534), .A4(n8533), .ZN(n13948) );
  INV_X1 U11106 ( .A(n13948), .ZN(n11728) );
  NAND2_X1 U11107 ( .A1(n14367), .A2(n11728), .ZN(n11730) );
  OR2_X1 U11108 ( .A1(n14367), .A2(n11728), .ZN(n8537) );
  NAND2_X1 U11109 ( .A1(n11730), .A2(n8537), .ZN(n14374) );
  NAND2_X1 U11110 ( .A1(n14367), .A2(n13948), .ZN(n8538) );
  NAND2_X1 U11111 ( .A1(n8756), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8546) );
  INV_X1 U11112 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14568) );
  OR2_X1 U11113 ( .A1(n8468), .A2(n14568), .ZN(n8545) );
  NAND2_X1 U11114 ( .A1(n8541), .A2(n8540), .ZN(n8542) );
  NAND2_X1 U11115 ( .A1(n8550), .A2(n8542), .ZN(n13885) );
  OR2_X1 U11116 ( .A1(n8739), .A2(n13885), .ZN(n8544) );
  INV_X1 U11117 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n14501) );
  OR2_X1 U11118 ( .A1(n8944), .A2(n14501), .ZN(n8543) );
  NOR2_X1 U11119 ( .A1(n14570), .A2(n13812), .ZN(n8548) );
  NAND2_X1 U11120 ( .A1(n14570), .A2(n13812), .ZN(n8547) );
  NAND2_X1 U11121 ( .A1(n8757), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8555) );
  INV_X1 U11122 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n14352) );
  OR2_X1 U11123 ( .A1(n8945), .A2(n14352), .ZN(n8554) );
  NAND2_X1 U11124 ( .A1(n8550), .A2(n8549), .ZN(n8551) );
  NAND2_X1 U11125 ( .A1(n8558), .A2(n8551), .ZN(n14351) );
  OR2_X1 U11126 ( .A1(n8739), .A2(n14351), .ZN(n8553) );
  INV_X1 U11127 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10839) );
  OR2_X1 U11128 ( .A1(n8944), .A2(n10839), .ZN(n8552) );
  NAND4_X1 U11129 ( .A1(n8555), .A2(n8554), .A3(n8553), .A4(n8552), .ZN(n13946) );
  NOR2_X1 U11130 ( .A1(n14357), .A2(n13946), .ZN(n8557) );
  NAND2_X1 U11131 ( .A1(n14357), .A2(n13946), .ZN(n8556) );
  NAND2_X1 U11132 ( .A1(n8756), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8563) );
  INV_X1 U11133 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n15879) );
  OR2_X1 U11134 ( .A1(n8468), .A2(n15879), .ZN(n8562) );
  INV_X1 U11135 ( .A(n8567), .ZN(n8568) );
  NAND2_X1 U11136 ( .A1(n8558), .A2(n10873), .ZN(n8559) );
  NAND2_X1 U11137 ( .A1(n8568), .A2(n8559), .ZN(n14340) );
  OR2_X1 U11138 ( .A1(n8739), .A2(n14340), .ZN(n8561) );
  INV_X1 U11139 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n14489) );
  OR2_X1 U11140 ( .A1(n8944), .A2(n14489), .ZN(n8560) );
  NAND4_X1 U11141 ( .A1(n8563), .A2(n8562), .A3(n8561), .A4(n8560), .ZN(n13945) );
  AND2_X1 U11142 ( .A1(n14339), .A2(n13945), .ZN(n8565) );
  NAND2_X1 U11143 ( .A1(n8756), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8573) );
  INV_X1 U11144 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8566) );
  OR2_X1 U11145 ( .A1(n8468), .A2(n8566), .ZN(n8572) );
  INV_X1 U11146 ( .A(n8582), .ZN(n8580) );
  INV_X1 U11147 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n15922) );
  NAND2_X1 U11148 ( .A1(n8568), .A2(n15922), .ZN(n8569) );
  NAND2_X1 U11149 ( .A1(n8580), .A2(n8569), .ZN(n14322) );
  OR2_X1 U11150 ( .A1(n8739), .A2(n14322), .ZN(n8571) );
  INV_X1 U11151 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10845) );
  OR2_X1 U11152 ( .A1(n8944), .A2(n10845), .ZN(n8570) );
  NAND4_X1 U11153 ( .A1(n8573), .A2(n8572), .A3(n8571), .A4(n8570), .ZN(n13944) );
  OR2_X1 U11154 ( .A1(n14481), .A2(n13944), .ZN(n9008) );
  INV_X1 U11155 ( .A(n9008), .ZN(n8574) );
  NAND2_X1 U11156 ( .A1(n14481), .A2(n13944), .ZN(n9007) );
  NAND2_X1 U11157 ( .A1(n8756), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8578) );
  INV_X1 U11158 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14558) );
  OR2_X1 U11159 ( .A1(n8468), .A2(n14558), .ZN(n8577) );
  INV_X1 U11160 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11289) );
  XNOR2_X1 U11161 ( .A(n8580), .B(n11289), .ZN(n14307) );
  OR2_X1 U11162 ( .A1(n8739), .A2(n14307), .ZN(n8576) );
  INV_X1 U11163 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14478) );
  OR2_X1 U11164 ( .A1(n8944), .A2(n14478), .ZN(n8575) );
  NAND4_X1 U11165 ( .A1(n8578), .A2(n8577), .A3(n8576), .A4(n8575), .ZN(n13943) );
  OR2_X1 U11166 ( .A1(n14306), .A2(n13943), .ZN(n14282) );
  INV_X1 U11167 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8579) );
  OAI21_X1 U11168 ( .B1(n8580), .B2(n11289), .A(n8579), .ZN(n8583) );
  AND2_X1 U11169 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n8581) );
  INV_X1 U11170 ( .A(n8594), .ZN(n8595) );
  AND2_X1 U11171 ( .A1(n8583), .A2(n8595), .ZN(n14292) );
  NAND2_X1 U11172 ( .A1(n8755), .A2(n14292), .ZN(n8588) );
  INV_X1 U11173 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8584) );
  OR2_X1 U11174 ( .A1(n8468), .A2(n8584), .ZN(n8587) );
  INV_X1 U11175 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11822) );
  OR2_X1 U11176 ( .A1(n8944), .A2(n11822), .ZN(n8586) );
  INV_X1 U11177 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n14284) );
  OR2_X1 U11178 ( .A1(n8945), .A2(n14284), .ZN(n8585) );
  NAND4_X1 U11179 ( .A1(n8588), .A2(n8587), .A3(n8586), .A4(n8585), .ZN(n13942) );
  NAND3_X1 U11180 ( .A1(n14306), .A2(n13943), .A3(n8590), .ZN(n8592) );
  NAND2_X1 U11181 ( .A1(n14469), .A2(n13942), .ZN(n8591) );
  AND2_X1 U11182 ( .A1(n8592), .A2(n8591), .ZN(n8593) );
  INV_X1 U11183 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n15845) );
  NAND2_X1 U11184 ( .A1(n8595), .A2(n15845), .ZN(n8596) );
  NAND2_X1 U11185 ( .A1(n8601), .A2(n8596), .ZN(n13837) );
  NOR2_X1 U11186 ( .A1(n13837), .A2(n8739), .ZN(n8600) );
  INV_X1 U11187 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14467) );
  NOR2_X1 U11188 ( .A1(n8944), .A2(n14467), .ZN(n8599) );
  INV_X1 U11189 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11837) );
  NAND2_X1 U11190 ( .A1(n8757), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8597) );
  OAI21_X1 U11191 ( .B1(n11837), .B2(n8945), .A(n8597), .ZN(n8598) );
  INV_X1 U11192 ( .A(n13941), .ZN(n13892) );
  XNOR2_X1 U11193 ( .A(n14274), .B(n13892), .ZN(n14272) );
  NAND2_X1 U11194 ( .A1(n8601), .A2(n13894), .ZN(n8602) );
  AND2_X1 U11195 ( .A1(n8610), .A2(n8602), .ZN(n14258) );
  NAND2_X1 U11196 ( .A1(n14258), .A2(n8755), .ZN(n8605) );
  AOI22_X1 U11197 ( .A1(n8756), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8757), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U11198 ( .A1(n8676), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8603) );
  XNOR2_X1 U11199 ( .A(n14460), .B(n13940), .ZN(n14264) );
  INV_X1 U11200 ( .A(n14264), .ZN(n8606) );
  NAND2_X1 U11201 ( .A1(n14260), .A2(n12639), .ZN(n8607) );
  INV_X1 U11202 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8609) );
  NAND2_X1 U11203 ( .A1(n8610), .A2(n8609), .ZN(n8611) );
  NAND2_X1 U11204 ( .A1(n8619), .A2(n8611), .ZN(n14247) );
  OR2_X1 U11205 ( .A1(n14247), .A2(n8739), .ZN(n8617) );
  INV_X1 U11206 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8614) );
  NAND2_X1 U11207 ( .A1(n8757), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8613) );
  NAND2_X1 U11208 ( .A1(n8756), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8612) );
  OAI211_X1 U11209 ( .C1(n8944), .C2(n8614), .A(n8613), .B(n8612), .ZN(n8615)
         );
  INV_X1 U11210 ( .A(n8615), .ZN(n8616) );
  NAND2_X1 U11211 ( .A1(n14456), .A2(n13939), .ZN(n9013) );
  INV_X1 U11212 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13854) );
  NAND2_X1 U11213 ( .A1(n8619), .A2(n13854), .ZN(n8620) );
  AND2_X1 U11214 ( .A1(n8630), .A2(n8620), .ZN(n14232) );
  NAND2_X1 U11215 ( .A1(n14232), .A2(n8755), .ZN(n8626) );
  INV_X1 U11216 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8623) );
  NAND2_X1 U11217 ( .A1(n8756), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8622) );
  NAND2_X1 U11218 ( .A1(n8757), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8621) );
  OAI211_X1 U11219 ( .C1(n8623), .C2(n8944), .A(n8622), .B(n8621), .ZN(n8624)
         );
  INV_X1 U11220 ( .A(n8624), .ZN(n8625) );
  NAND2_X1 U11221 ( .A1(n8626), .A2(n8625), .ZN(n13938) );
  NAND2_X1 U11222 ( .A1(n14451), .A2(n13938), .ZN(n8627) );
  INV_X1 U11223 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U11224 ( .A1(n8630), .A2(n8629), .ZN(n8631) );
  NAND2_X1 U11225 ( .A1(n8639), .A2(n8631), .ZN(n14209) );
  OR2_X1 U11226 ( .A1(n14209), .A2(n8739), .ZN(n8636) );
  INV_X1 U11227 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n14447) );
  NAND2_X1 U11228 ( .A1(n8757), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8633) );
  NAND2_X1 U11229 ( .A1(n8756), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8632) );
  OAI211_X1 U11230 ( .C1(n14447), .C2(n8944), .A(n8633), .B(n8632), .ZN(n8634)
         );
  INV_X1 U11231 ( .A(n8634), .ZN(n8635) );
  XNOR2_X1 U11232 ( .A(n14214), .B(n12655), .ZN(n9016) );
  INV_X1 U11233 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U11234 ( .A1(n8639), .A2(n8638), .ZN(n8640) );
  NAND2_X1 U11235 ( .A1(n8647), .A2(n8640), .ZN(n14198) );
  OR2_X1 U11236 ( .A1(n14198), .A2(n8739), .ZN(n8645) );
  INV_X1 U11237 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n14441) );
  NAND2_X1 U11238 ( .A1(n8757), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8642) );
  NAND2_X1 U11239 ( .A1(n8756), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8641) );
  OAI211_X1 U11240 ( .C1(n14441), .C2(n8944), .A(n8642), .B(n8641), .ZN(n8643)
         );
  INV_X1 U11241 ( .A(n8643), .ZN(n8644) );
  NAND2_X1 U11242 ( .A1(n14194), .A2(n13801), .ZN(n8725) );
  NAND2_X1 U11243 ( .A1(n14157), .A2(n8725), .ZN(n9015) );
  OR2_X1 U11244 ( .A1(n14545), .A2(n13801), .ZN(n8646) );
  INV_X1 U11245 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n16033) );
  OR2_X2 U11246 ( .A1(n8647), .A2(n16033), .ZN(n8664) );
  NAND2_X1 U11247 ( .A1(n8647), .A2(n16033), .ZN(n8648) );
  NAND2_X1 U11248 ( .A1(n8664), .A2(n8648), .ZN(n14181) );
  OR2_X1 U11249 ( .A1(n14181), .A2(n8739), .ZN(n8654) );
  INV_X1 U11250 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U11251 ( .A1(n8757), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8650) );
  NAND2_X1 U11252 ( .A1(n8756), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8649) );
  OAI211_X1 U11253 ( .C1(n8944), .C2(n8651), .A(n8650), .B(n8649), .ZN(n8652)
         );
  INV_X1 U11254 ( .A(n8652), .ZN(n8653) );
  INV_X1 U11255 ( .A(n14175), .ZN(n8655) );
  XNOR2_X1 U11256 ( .A(n8664), .B(P2_REG3_REG_24__SCAN_IN), .ZN(n14168) );
  NAND2_X1 U11257 ( .A1(n14168), .A2(n8755), .ZN(n8661) );
  INV_X1 U11258 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U11259 ( .A1(n8676), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8657) );
  NAND2_X1 U11260 ( .A1(n8757), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8656) );
  OAI211_X1 U11261 ( .C1(n8945), .C2(n8658), .A(n8657), .B(n8656), .ZN(n8659)
         );
  INV_X1 U11262 ( .A(n8659), .ZN(n8660) );
  AND2_X2 U11263 ( .A1(n8661), .A2(n8660), .ZN(n13768) );
  INV_X2 U11264 ( .A(n13768), .ZN(n13934) );
  XNOR2_X1 U11265 ( .A(n14167), .B(n13934), .ZN(n14163) );
  NAND2_X1 U11266 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n8662) );
  INV_X1 U11267 ( .A(n8673), .ZN(n8674) );
  INV_X1 U11268 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13846) );
  INV_X1 U11269 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8663) );
  OAI21_X1 U11270 ( .B1(n8664), .B2(n13846), .A(n8663), .ZN(n8665) );
  NAND2_X1 U11271 ( .A1(n14150), .A2(n8755), .ZN(n8670) );
  INV_X1 U11272 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14423) );
  NAND2_X1 U11273 ( .A1(n8756), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U11274 ( .A1(n8757), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8666) );
  OAI211_X1 U11275 ( .C1(n14423), .C2(n8944), .A(n8667), .B(n8666), .ZN(n8668)
         );
  INV_X1 U11276 ( .A(n8668), .ZN(n8669) );
  INV_X1 U11277 ( .A(n13933), .ZN(n8671) );
  NOR2_X1 U11278 ( .A1(n14534), .A2(n8671), .ZN(n8672) );
  INV_X1 U11279 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n15965) );
  NAND2_X1 U11280 ( .A1(n8674), .A2(n15965), .ZN(n8675) );
  NAND2_X1 U11281 ( .A1(n8734), .A2(n8675), .ZN(n14132) );
  OR2_X1 U11282 ( .A1(n14132), .A2(n8739), .ZN(n8681) );
  INV_X1 U11283 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n14131) );
  NAND2_X1 U11284 ( .A1(n8676), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8678) );
  NAND2_X1 U11285 ( .A1(n8757), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8677) );
  OAI211_X1 U11286 ( .C1(n8945), .C2(n14131), .A(n8678), .B(n8677), .ZN(n8679)
         );
  INV_X1 U11287 ( .A(n8679), .ZN(n8680) );
  INV_X1 U11288 ( .A(n13932), .ZN(n8746) );
  XNOR2_X1 U11289 ( .A(n8734), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n14120) );
  NAND2_X1 U11290 ( .A1(n14120), .A2(n8755), .ZN(n8686) );
  INV_X1 U11291 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n16101) );
  NAND2_X1 U11292 ( .A1(n8757), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8683) );
  NAND2_X1 U11293 ( .A1(n8756), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8682) );
  OAI211_X1 U11294 ( .C1(n8944), .C2(n16101), .A(n8683), .B(n8682), .ZN(n8684)
         );
  INV_X1 U11295 ( .A(n8684), .ZN(n8685) );
  INV_X1 U11296 ( .A(n14128), .ZN(n8690) );
  INV_X1 U11297 ( .A(n8767), .ZN(n8689) );
  AOI211_X1 U11298 ( .C1(n13752), .C2(n8690), .A(n14338), .B(n8689), .ZN(
        n14119) );
  NOR2_X1 U11299 ( .A1(n8788), .A2(n15660), .ZN(n11974) );
  NAND2_X1 U11300 ( .A1(n8691), .A2(n11974), .ZN(n11973) );
  OR2_X1 U11301 ( .A1(n8781), .A2(n15707), .ZN(n8692) );
  NOR2_X1 U11302 ( .A1(n13956), .A2(n10584), .ZN(n11705) );
  INV_X1 U11303 ( .A(n9011), .ZN(n11708) );
  NAND2_X1 U11304 ( .A1(n13956), .A2(n10584), .ZN(n8693) );
  OAI211_X1 U11305 ( .C1(n11707), .C2(n11705), .A(n11708), .B(n8693), .ZN(
        n8695) );
  OR2_X1 U11306 ( .A1(n13955), .A2(n15717), .ZN(n8694) );
  NAND2_X1 U11307 ( .A1(n8695), .A2(n8694), .ZN(n10793) );
  INV_X1 U11308 ( .A(n10790), .ZN(n10792) );
  NAND2_X1 U11309 ( .A1(n10793), .A2(n10792), .ZN(n8697) );
  OR2_X1 U11310 ( .A1(n11625), .A2(n13954), .ZN(n8696) );
  NAND2_X1 U11311 ( .A1(n8697), .A2(n8696), .ZN(n11961) );
  XNOR2_X1 U11312 ( .A(n8148), .B(n13953), .ZN(n11955) );
  INV_X1 U11313 ( .A(n11955), .ZN(n11962) );
  NAND2_X1 U11314 ( .A1(n11961), .A2(n11962), .ZN(n8700) );
  INV_X1 U11315 ( .A(n13953), .ZN(n8698) );
  NAND2_X1 U11316 ( .A1(n8698), .A2(n11224), .ZN(n8699) );
  NAND2_X1 U11317 ( .A1(n8700), .A2(n8699), .ZN(n11655) );
  INV_X1 U11318 ( .A(n13952), .ZN(n11387) );
  NAND2_X1 U11319 ( .A1(n11661), .A2(n11387), .ZN(n8701) );
  INV_X1 U11320 ( .A(n13951), .ZN(n11644) );
  AND2_X1 U11321 ( .A1(n11683), .A2(n11644), .ZN(n8704) );
  OR2_X1 U11322 ( .A1(n11683), .A2(n11644), .ZN(n8703) );
  INV_X1 U11323 ( .A(n14371), .ZN(n8706) );
  INV_X1 U11324 ( .A(n14374), .ZN(n14363) );
  XNOR2_X1 U11325 ( .A(n13887), .B(n13812), .ZN(n11731) );
  INV_X1 U11326 ( .A(n11731), .ZN(n11726) );
  INV_X1 U11327 ( .A(n13812), .ZN(n13947) );
  OR2_X1 U11328 ( .A1(n14570), .A2(n13947), .ZN(n8709) );
  INV_X1 U11329 ( .A(n13946), .ZN(n13864) );
  OR2_X1 U11330 ( .A1(n14357), .A2(n13864), .ZN(n8710) );
  INV_X1 U11331 ( .A(n13945), .ZN(n8712) );
  AND2_X1 U11332 ( .A1(n14339), .A2(n8712), .ZN(n8711) );
  OR2_X1 U11333 ( .A1(n14339), .A2(n8712), .ZN(n8713) );
  INV_X1 U11334 ( .A(n13944), .ZN(n13916) );
  NOR2_X1 U11335 ( .A1(n14481), .A2(n13916), .ZN(n8714) );
  INV_X1 U11336 ( .A(n13943), .ZN(n8716) );
  AND2_X1 U11337 ( .A1(n14306), .A2(n8716), .ZN(n8715) );
  OR2_X1 U11338 ( .A1(n14306), .A2(n8716), .ZN(n8717) );
  INV_X1 U11339 ( .A(n13942), .ZN(n13918) );
  OR2_X1 U11340 ( .A1(n14274), .A2(n13892), .ZN(n8718) );
  AND2_X1 U11341 ( .A1(n14260), .A2(n13940), .ZN(n8719) );
  NOR2_X1 U11342 ( .A1(n14251), .A2(n13939), .ZN(n8721) );
  NAND2_X1 U11343 ( .A1(n14251), .A2(n13939), .ZN(n8720) );
  INV_X1 U11344 ( .A(n13938), .ZN(n8911) );
  NAND2_X1 U11345 ( .A1(n14451), .A2(n8911), .ZN(n8723) );
  OR2_X1 U11346 ( .A1(n14451), .A2(n8911), .ZN(n8722) );
  NAND2_X1 U11347 ( .A1(n14548), .A2(n13937), .ZN(n8724) );
  NAND2_X1 U11348 ( .A1(n14182), .A2(n13731), .ZN(n14158) );
  INV_X1 U11349 ( .A(n14157), .ZN(n8727) );
  AOI21_X1 U11350 ( .B1(n13731), .B2(n14157), .A(n14182), .ZN(n8726) );
  INV_X1 U11351 ( .A(n14163), .ZN(n14159) );
  AOI211_X1 U11352 ( .C1(n8727), .C2(n13935), .A(n8726), .B(n14159), .ZN(n8728) );
  XNOR2_X1 U11353 ( .A(n14146), .B(n13933), .ZN(n14142) );
  INV_X1 U11354 ( .A(n14142), .ZN(n8730) );
  XNOR2_X1 U11355 ( .A(n14130), .B(n13932), .ZN(n14136) );
  XNOR2_X1 U11356 ( .A(n8752), .B(n8765), .ZN(n8748) );
  NAND2_X1 U11357 ( .A1(n6562), .A2(n9010), .ZN(n8731) );
  OAI21_X2 U11358 ( .B1(n14086), .B2(n11491), .A(n8731), .ZN(n15662) );
  INV_X1 U11359 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8733) );
  INV_X1 U11360 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8732) );
  OAI21_X1 U11361 ( .B1(n8734), .B2(n8733), .A(n8732), .ZN(n8738) );
  INV_X1 U11362 ( .A(n8734), .ZN(n8736) );
  AND2_X1 U11363 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n8735) );
  INV_X1 U11364 ( .A(n14101), .ZN(n8737) );
  NAND2_X1 U11365 ( .A1(n8738), .A2(n8737), .ZN(n13793) );
  OR2_X1 U11366 ( .A1(n13793), .A2(n8739), .ZN(n8744) );
  INV_X1 U11367 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n12590) );
  NAND2_X1 U11368 ( .A1(n8756), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8741) );
  NAND2_X1 U11369 ( .A1(n8757), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8740) );
  OAI211_X1 U11370 ( .C1(n12590), .C2(n8944), .A(n8741), .B(n8740), .ZN(n8742)
         );
  INV_X1 U11371 ( .A(n8742), .ZN(n8743) );
  INV_X1 U11372 ( .A(n8398), .ZN(n8745) );
  OAI22_X1 U11373 ( .A1(n9917), .A2(n13917), .B1(n8746), .B2(n13915), .ZN(
        n8747) );
  INV_X1 U11374 ( .A(n8747), .ZN(n13750) );
  MUX2_X1 U11375 ( .A(n8749), .B(n14413), .S(n15743), .Z(n8751) );
  NAND2_X1 U11376 ( .A1(n13752), .A2(n8433), .ZN(n8750) );
  NAND2_X1 U11377 ( .A1(n8751), .A2(n8750), .ZN(P2_U3494) );
  INV_X1 U11378 ( .A(n9906), .ZN(n8753) );
  NAND2_X1 U11379 ( .A1(n13752), .A2(n8764), .ZN(n9904) );
  NAND2_X1 U11380 ( .A1(n13797), .A2(n9917), .ZN(n9905) );
  XNOR2_X1 U11381 ( .A(n8754), .B(n9900), .ZN(n8763) );
  NAND2_X1 U11382 ( .A1(n14101), .A2(n8755), .ZN(n8762) );
  INV_X1 U11383 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9928) );
  NAND2_X1 U11384 ( .A1(n8756), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8759) );
  NAND2_X1 U11385 ( .A1(n8757), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8758) );
  OAI211_X1 U11386 ( .C1(n8944), .C2(n9928), .A(n8759), .B(n8758), .ZN(n8760)
         );
  INV_X1 U11387 ( .A(n8760), .ZN(n8761) );
  NAND2_X1 U11388 ( .A1(n8762), .A2(n8761), .ZN(n13929) );
  AOI22_X1 U11389 ( .A1(n13931), .A2(n13905), .B1(n13929), .B2(n13907), .ZN(
        n13795) );
  XNOR2_X1 U11390 ( .A(n9901), .B(n7168), .ZN(n14114) );
  INV_X1 U11391 ( .A(n9903), .ZN(n8766) );
  AOI211_X1 U11392 ( .C1(n13797), .C2(n8767), .A(n14338), .B(n8766), .ZN(
        n14113) );
  NAND2_X1 U11393 ( .A1(n8769), .A2(n8768), .ZN(n8770) );
  INV_X1 U11394 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8771) );
  INV_X1 U11395 ( .A(n8773), .ZN(n8774) );
  OAI22_X1 U11396 ( .A1(n14545), .A2(n8997), .B1(n13801), .B2(n8960), .ZN(
        n8924) );
  OAI22_X1 U11397 ( .A1(n14260), .A2(n8960), .B1(n12639), .B2(n8997), .ZN(
        n8904) );
  INV_X1 U11398 ( .A(n8904), .ZN(n8908) );
  NAND2_X1 U11399 ( .A1(n8921), .A2(n7528), .ZN(n8778) );
  NAND2_X1 U11400 ( .A1(n8781), .A2(n8776), .ZN(n8777) );
  NAND2_X1 U11401 ( .A1(n8778), .A2(n8777), .ZN(n8793) );
  NOR2_X1 U11402 ( .A1(n8921), .A2(n8779), .ZN(n8780) );
  NAND2_X1 U11403 ( .A1(n8793), .A2(n8794), .ZN(n8792) );
  NAND2_X1 U11404 ( .A1(n8788), .A2(n15660), .ZN(n8784) );
  OAI21_X1 U11405 ( .B1(n10011), .B2(n8782), .A(n10009), .ZN(n8785) );
  NAND3_X1 U11406 ( .A1(n8784), .A2(n8785), .A3(n8783), .ZN(n8790) );
  NAND2_X1 U11407 ( .A1(n8790), .A2(n8789), .ZN(n8791) );
  INV_X1 U11408 ( .A(n8793), .ZN(n8796) );
  INV_X1 U11409 ( .A(n8794), .ZN(n8795) );
  NAND2_X1 U11410 ( .A1(n8796), .A2(n8795), .ZN(n8797) );
  NAND2_X1 U11411 ( .A1(n8961), .A2(n13956), .ZN(n8799) );
  NAND2_X1 U11412 ( .A1(n6561), .A2(n11934), .ZN(n8798) );
  AOI22_X1 U11413 ( .A1(n8961), .A2(n11934), .B1(n6561), .B2(n13956), .ZN(
        n8800) );
  NAND2_X1 U11414 ( .A1(n8961), .A2(n11717), .ZN(n8803) );
  NAND2_X1 U11415 ( .A1(n13955), .A2(n8776), .ZN(n8802) );
  NAND2_X1 U11416 ( .A1(n8803), .A2(n8802), .ZN(n8805) );
  AOI22_X1 U11417 ( .A1(n8961), .A2(n13955), .B1(n8776), .B2(n11717), .ZN(
        n8804) );
  NOR2_X1 U11418 ( .A1(n8806), .A2(n8805), .ZN(n8807) );
  NAND2_X1 U11419 ( .A1(n8961), .A2(n13954), .ZN(n8810) );
  NAND2_X1 U11420 ( .A1(n8997), .A2(n10851), .ZN(n8809) );
  NAND2_X1 U11421 ( .A1(n8810), .A2(n8809), .ZN(n8812) );
  AOI22_X1 U11422 ( .A1(n8961), .A2(n10851), .B1(n8997), .B2(n13954), .ZN(
        n8811) );
  AOI21_X1 U11423 ( .B1(n8813), .B2(n8812), .A(n8811), .ZN(n8815) );
  NOR2_X1 U11424 ( .A1(n8813), .A2(n8812), .ZN(n8814) );
  NAND2_X1 U11425 ( .A1(n8961), .A2(n11224), .ZN(n8817) );
  NAND2_X1 U11426 ( .A1(n13953), .A2(n8997), .ZN(n8816) );
  NAND2_X1 U11427 ( .A1(n8817), .A2(n8816), .ZN(n8819) );
  AOI22_X1 U11428 ( .A1(n8961), .A2(n13953), .B1(n8997), .B2(n11224), .ZN(
        n8818) );
  NAND2_X1 U11429 ( .A1(n8961), .A2(n13952), .ZN(n8822) );
  NAND2_X1 U11430 ( .A1(n11661), .A2(n8997), .ZN(n8821) );
  NAND2_X1 U11431 ( .A1(n8822), .A2(n8821), .ZN(n8825) );
  NAND2_X1 U11432 ( .A1(n8961), .A2(n11661), .ZN(n8823) );
  OAI21_X1 U11433 ( .B1(n11387), .B2(n8961), .A(n8823), .ZN(n8824) );
  NAND2_X1 U11434 ( .A1(n8960), .A2(n11683), .ZN(n8827) );
  NAND2_X1 U11435 ( .A1(n13951), .A2(n8997), .ZN(n8826) );
  NAND2_X1 U11436 ( .A1(n8827), .A2(n8826), .ZN(n8830) );
  AOI22_X1 U11437 ( .A1(n13951), .A2(n8961), .B1(n11683), .B2(n8997), .ZN(
        n8828) );
  AOI21_X1 U11438 ( .B1(n8831), .B2(n8830), .A(n8828), .ZN(n8829) );
  NOR2_X1 U11439 ( .A1(n8831), .A2(n8830), .ZN(n8832) );
  AOI22_X1 U11440 ( .A1(n14519), .A2(n8997), .B1(n13950), .B2(n8961), .ZN(
        n8835) );
  NAND2_X1 U11441 ( .A1(n14519), .A2(n8961), .ZN(n8833) );
  OAI21_X1 U11442 ( .B1(n11388), .B2(n8960), .A(n8833), .ZN(n8834) );
  INV_X1 U11443 ( .A(n8840), .ZN(n8843) );
  NAND2_X1 U11444 ( .A1(n14575), .A2(n8960), .ZN(n8837) );
  NAND2_X1 U11445 ( .A1(n13949), .A2(n8997), .ZN(n8836) );
  NAND2_X1 U11446 ( .A1(n8837), .A2(n8836), .ZN(n8839) );
  INV_X1 U11447 ( .A(n8839), .ZN(n8842) );
  AOI22_X1 U11448 ( .A1(n14575), .A2(n8997), .B1(n13949), .B2(n8960), .ZN(
        n8838) );
  AOI22_X1 U11449 ( .A1(n14367), .A2(n8997), .B1(n13948), .B2(n8960), .ZN(
        n8845) );
  OAI22_X1 U11450 ( .A1(n14504), .A2(n8997), .B1(n11728), .B2(n8960), .ZN(
        n8844) );
  AOI22_X1 U11451 ( .A1(n13887), .A2(n8960), .B1(n8997), .B2(n13947), .ZN(
        n8851) );
  OAI22_X1 U11452 ( .A1(n14570), .A2(n8960), .B1(n13812), .B2(n8997), .ZN(
        n8850) );
  AND2_X1 U11453 ( .A1(n13946), .A2(n8997), .ZN(n8847) );
  AOI21_X1 U11454 ( .B1(n14357), .B2(n8960), .A(n8847), .ZN(n8872) );
  NAND2_X1 U11455 ( .A1(n14357), .A2(n8997), .ZN(n8849) );
  NAND2_X1 U11456 ( .A1(n8960), .A2(n13946), .ZN(n8848) );
  NAND2_X1 U11457 ( .A1(n8849), .A2(n8848), .ZN(n8871) );
  OAI22_X1 U11458 ( .A1(n8872), .A2(n8871), .B1(n8851), .B2(n8850), .ZN(n8875)
         );
  AND2_X1 U11459 ( .A1(n13941), .A2(n8997), .ZN(n8852) );
  AOI21_X1 U11460 ( .B1(n14274), .B2(n8960), .A(n8852), .ZN(n8893) );
  NAND2_X1 U11461 ( .A1(n14274), .A2(n8997), .ZN(n8854) );
  NAND2_X1 U11462 ( .A1(n8960), .A2(n13941), .ZN(n8853) );
  NAND2_X1 U11463 ( .A1(n8854), .A2(n8853), .ZN(n8891) );
  NAND2_X1 U11464 ( .A1(n8893), .A2(n8891), .ZN(n8859) );
  AND2_X1 U11465 ( .A1(n13942), .A2(n8997), .ZN(n8855) );
  AOI21_X1 U11466 ( .B1(n14469), .B2(n8960), .A(n8855), .ZN(n8888) );
  NAND2_X1 U11467 ( .A1(n14469), .A2(n8997), .ZN(n8857) );
  NAND2_X1 U11468 ( .A1(n8960), .A2(n13942), .ZN(n8856) );
  NAND2_X1 U11469 ( .A1(n8857), .A2(n8856), .ZN(n8887) );
  NAND2_X1 U11470 ( .A1(n8888), .A2(n8887), .ZN(n8858) );
  NAND2_X1 U11471 ( .A1(n8859), .A2(n8858), .ZN(n8886) );
  AND2_X1 U11472 ( .A1(n13943), .A2(n8997), .ZN(n8860) );
  AOI21_X1 U11473 ( .B1(n14306), .B2(n8960), .A(n8860), .ZN(n8885) );
  NAND2_X1 U11474 ( .A1(n14306), .A2(n8997), .ZN(n8862) );
  NAND2_X1 U11475 ( .A1(n8960), .A2(n13943), .ZN(n8861) );
  NAND2_X1 U11476 ( .A1(n8862), .A2(n8861), .ZN(n8884) );
  AND2_X1 U11477 ( .A1(n8885), .A2(n8884), .ZN(n8863) );
  OR2_X1 U11478 ( .A1(n8886), .A2(n8863), .ZN(n8878) );
  AND2_X1 U11479 ( .A1(n13944), .A2(n8997), .ZN(n8864) );
  AOI21_X1 U11480 ( .B1(n14481), .B2(n8960), .A(n8864), .ZN(n8877) );
  NAND2_X1 U11481 ( .A1(n14481), .A2(n8997), .ZN(n8866) );
  NAND2_X1 U11482 ( .A1(n8960), .A2(n13944), .ZN(n8865) );
  NAND2_X1 U11483 ( .A1(n8866), .A2(n8865), .ZN(n8876) );
  AND2_X1 U11484 ( .A1(n8877), .A2(n8876), .ZN(n8867) );
  NOR2_X1 U11485 ( .A1(n8878), .A2(n8867), .ZN(n8883) );
  AND2_X1 U11486 ( .A1(n13945), .A2(n8997), .ZN(n8868) );
  AOI21_X1 U11487 ( .B1(n14339), .B2(n8960), .A(n8868), .ZN(n8880) );
  NAND2_X1 U11488 ( .A1(n14339), .A2(n8997), .ZN(n8870) );
  NAND2_X1 U11489 ( .A1(n8960), .A2(n13945), .ZN(n8869) );
  NAND2_X1 U11490 ( .A1(n8870), .A2(n8869), .ZN(n8879) );
  AOI22_X1 U11491 ( .A1(n8880), .A2(n8879), .B1(n8872), .B2(n8871), .ZN(n8873)
         );
  OR3_X1 U11492 ( .A1(n8878), .A2(n8877), .A3(n8876), .ZN(n8902) );
  INV_X1 U11493 ( .A(n8879), .ZN(n8882) );
  INV_X1 U11494 ( .A(n8880), .ZN(n8881) );
  NAND3_X1 U11495 ( .A1(n8883), .A2(n8882), .A3(n8881), .ZN(n8901) );
  OR3_X1 U11496 ( .A1(n8886), .A2(n8885), .A3(n8884), .ZN(n8899) );
  INV_X1 U11497 ( .A(n8887), .ZN(n8890) );
  INV_X1 U11498 ( .A(n8888), .ZN(n8889) );
  NAND2_X1 U11499 ( .A1(n8890), .A2(n8889), .ZN(n8892) );
  NAND3_X1 U11500 ( .A1(n8892), .A2(n14555), .A3(n13892), .ZN(n8897) );
  INV_X1 U11501 ( .A(n8891), .ZN(n8896) );
  INV_X1 U11502 ( .A(n8892), .ZN(n8895) );
  INV_X1 U11503 ( .A(n8893), .ZN(n8894) );
  AOI22_X1 U11504 ( .A1(n8897), .A2(n8896), .B1(n8895), .B2(n8894), .ZN(n8898)
         );
  AND2_X1 U11505 ( .A1(n8899), .A2(n8898), .ZN(n8900) );
  INV_X1 U11506 ( .A(n8905), .ZN(n8907) );
  AOI22_X1 U11507 ( .A1(n14460), .A2(n8960), .B1(n8997), .B2(n13940), .ZN(
        n8903) );
  AOI21_X1 U11508 ( .B1(n8905), .B2(n8904), .A(n8903), .ZN(n8906) );
  OAI22_X1 U11509 ( .A1(n14251), .A2(n8997), .B1(n13893), .B2(n8960), .ZN(
        n8909) );
  OAI22_X1 U11510 ( .A1(n14251), .A2(n8960), .B1(n13893), .B2(n8997), .ZN(
        n8910) );
  AOI22_X1 U11511 ( .A1(n14451), .A2(n8997), .B1(n13938), .B2(n8960), .ZN(
        n8913) );
  INV_X1 U11512 ( .A(n14451), .ZN(n13856) );
  OAI22_X1 U11513 ( .A1(n13856), .A2(n8997), .B1(n8911), .B2(n8960), .ZN(n8912) );
  OAI21_X1 U11514 ( .B1(n8914), .B2(n8913), .A(n8912), .ZN(n8916) );
  NAND2_X1 U11515 ( .A1(n8914), .A2(n8913), .ZN(n8915) );
  NAND2_X1 U11516 ( .A1(n8916), .A2(n8915), .ZN(n8917) );
  OAI22_X1 U11517 ( .A1(n14548), .A2(n8997), .B1(n12655), .B2(n8960), .ZN(
        n8918) );
  OAI22_X1 U11518 ( .A1(n14548), .A2(n8960), .B1(n12655), .B2(n8997), .ZN(
        n8920) );
  INV_X1 U11519 ( .A(n8918), .ZN(n8919) );
  OAI22_X1 U11520 ( .A1(n14545), .A2(n8960), .B1(n13801), .B2(n8997), .ZN(
        n8922) );
  INV_X1 U11521 ( .A(n8922), .ZN(n8923) );
  AOI22_X1 U11522 ( .A1(n14182), .A2(n8960), .B1(n8997), .B2(n13935), .ZN(
        n8925) );
  NOR2_X1 U11523 ( .A1(n8926), .A2(n8925), .ZN(n8929) );
  AOI22_X1 U11524 ( .A1(n14182), .A2(n8997), .B1(n13935), .B2(n8960), .ZN(
        n8928) );
  NAND2_X1 U11525 ( .A1(n8926), .A2(n8925), .ZN(n8927) );
  OAI22_X1 U11526 ( .A1(n14537), .A2(n8960), .B1(n13768), .B2(n8997), .ZN(
        n8942) );
  AOI22_X1 U11527 ( .A1(n14167), .A2(n8960), .B1(n8997), .B2(n13934), .ZN(
        n8930) );
  AOI21_X1 U11528 ( .B1(n8943), .B2(n8942), .A(n8930), .ZN(n8980) );
  AND2_X1 U11529 ( .A1(n13933), .A2(n8997), .ZN(n8931) );
  AOI21_X1 U11530 ( .B1(n14146), .B2(n8960), .A(n8931), .ZN(n8964) );
  NAND2_X1 U11531 ( .A1(n14146), .A2(n8997), .ZN(n8933) );
  NAND2_X1 U11532 ( .A1(n13933), .A2(n8960), .ZN(n8932) );
  NAND2_X1 U11533 ( .A1(n8933), .A2(n8932), .ZN(n8963) );
  AND2_X1 U11534 ( .A1(n13931), .A2(n8960), .ZN(n8934) );
  AOI21_X1 U11535 ( .B1(n13752), .B2(n8997), .A(n8934), .ZN(n8974) );
  NAND2_X1 U11536 ( .A1(n13752), .A2(n8960), .ZN(n8936) );
  NAND2_X1 U11537 ( .A1(n13931), .A2(n8997), .ZN(n8935) );
  NAND2_X1 U11538 ( .A1(n8936), .A2(n8935), .ZN(n8973) );
  NAND2_X1 U11539 ( .A1(n8974), .A2(n8973), .ZN(n8962) );
  AND2_X1 U11540 ( .A1(n13932), .A2(n8960), .ZN(n8937) );
  AOI21_X1 U11541 ( .B1(n14130), .B2(n8997), .A(n8937), .ZN(n8968) );
  NAND2_X1 U11542 ( .A1(n14130), .A2(n8960), .ZN(n8939) );
  NAND2_X1 U11543 ( .A1(n13932), .A2(n8997), .ZN(n8938) );
  NAND2_X1 U11544 ( .A1(n8939), .A2(n8938), .ZN(n8967) );
  NAND2_X1 U11545 ( .A1(n8968), .A2(n8967), .ZN(n8972) );
  OAI211_X1 U11546 ( .C1(n8964), .C2(n8963), .A(n8962), .B(n8972), .ZN(n8940)
         );
  INV_X1 U11547 ( .A(n8940), .ZN(n8941) );
  OAI21_X1 U11548 ( .B1(n8943), .B2(n8942), .A(n8941), .ZN(n8979) );
  INV_X1 U11549 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n14411) );
  OR2_X1 U11550 ( .A1(n8944), .A2(n14411), .ZN(n8948) );
  INV_X1 U11551 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n14094) );
  OR2_X1 U11552 ( .A1(n8945), .A2(n14094), .ZN(n8947) );
  INV_X1 U11553 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14524) );
  OR2_X1 U11554 ( .A1(n8468), .A2(n14524), .ZN(n8946) );
  AND3_X1 U11555 ( .A1(n8948), .A2(n8947), .A3(n8946), .ZN(n8949) );
  OAI22_X1 U11556 ( .A1(n14526), .A2(n8997), .B1(n8949), .B2(n8960), .ZN(n8991) );
  INV_X1 U11557 ( .A(n14526), .ZN(n14097) );
  INV_X1 U11558 ( .A(n8949), .ZN(n13928) );
  INV_X1 U11559 ( .A(n8950), .ZN(n15665) );
  NAND2_X1 U11560 ( .A1(n8960), .A2(n13927), .ZN(n8952) );
  OAI211_X1 U11561 ( .C1(n15665), .C2(n11491), .A(n8952), .B(n8951), .ZN(n8953) );
  AOI22_X1 U11562 ( .A1(n14097), .A2(n8997), .B1(n13928), .B2(n8953), .ZN(
        n8992) );
  AND2_X1 U11563 ( .A1(n13929), .A2(n8960), .ZN(n8954) );
  AOI21_X1 U11564 ( .B1(n9922), .B2(n8997), .A(n8954), .ZN(n8986) );
  NAND2_X1 U11565 ( .A1(n9922), .A2(n8960), .ZN(n8956) );
  NAND2_X1 U11566 ( .A1(n13929), .A2(n8997), .ZN(n8955) );
  NAND2_X1 U11567 ( .A1(n8956), .A2(n8955), .ZN(n8985) );
  OAI22_X1 U11568 ( .A1(n8991), .A2(n8992), .B1(n8986), .B2(n8985), .ZN(n8959)
         );
  INV_X1 U11569 ( .A(n13927), .ZN(n8957) );
  NAND2_X1 U11570 ( .A1(n8995), .A2(n8957), .ZN(n8998) );
  OR2_X1 U11571 ( .A1(n8995), .A2(n8957), .ZN(n8958) );
  NAND2_X1 U11572 ( .A1(n8959), .A2(n9021), .ZN(n8987) );
  AOI22_X1 U11573 ( .A1(n13797), .A2(n8960), .B1(n8997), .B2(n13930), .ZN(
        n8982) );
  OAI22_X1 U11574 ( .A1(n14111), .A2(n8960), .B1(n9917), .B2(n8997), .ZN(n8981) );
  INV_X1 U11575 ( .A(n8962), .ZN(n8976) );
  INV_X1 U11576 ( .A(n8963), .ZN(n8966) );
  INV_X1 U11577 ( .A(n8964), .ZN(n8965) );
  NOR2_X1 U11578 ( .A1(n8966), .A2(n8965), .ZN(n8971) );
  INV_X1 U11579 ( .A(n8967), .ZN(n8970) );
  INV_X1 U11580 ( .A(n8968), .ZN(n8969) );
  AOI22_X1 U11581 ( .A1(n8972), .A2(n8971), .B1(n8970), .B2(n8969), .ZN(n8975)
         );
  OAI22_X1 U11582 ( .A1(n8976), .A2(n8975), .B1(n8974), .B2(n8973), .ZN(n8977)
         );
  AOI21_X1 U11583 ( .B1(n8982), .B2(n8981), .A(n8977), .ZN(n8978) );
  OAI21_X1 U11584 ( .B1(n8980), .B2(n8979), .A(n8028), .ZN(n8994) );
  INV_X1 U11585 ( .A(n8981), .ZN(n8984) );
  INV_X1 U11586 ( .A(n8982), .ZN(n8983) );
  AOI22_X1 U11587 ( .A1(n8986), .A2(n8985), .B1(n8984), .B2(n8983), .ZN(n8989)
         );
  INV_X1 U11588 ( .A(n8987), .ZN(n8988) );
  AOI21_X1 U11589 ( .B1(n9021), .B2(n8989), .A(n8988), .ZN(n8990) );
  AOI21_X1 U11590 ( .B1(n8992), .B2(n8991), .A(n8990), .ZN(n8993) );
  NAND2_X1 U11591 ( .A1(n8994), .A2(n8993), .ZN(n9001) );
  NAND2_X1 U11592 ( .A1(n8997), .A2(n13927), .ZN(n8996) );
  OAI22_X1 U11593 ( .A1(n8998), .A2(n8997), .B1(n8996), .B2(n8995), .ZN(n8999)
         );
  INV_X1 U11594 ( .A(n8999), .ZN(n9000) );
  NAND2_X1 U11595 ( .A1(n9001), .A2(n9000), .ZN(n9004) );
  OAI21_X1 U11596 ( .B1(n6562), .B2(n11283), .A(n14086), .ZN(n9002) );
  MUX2_X1 U11597 ( .A(n11359), .B(n11491), .S(n11283), .Z(n9003) );
  INV_X1 U11598 ( .A(n10426), .ZN(n9005) );
  AND2_X1 U11599 ( .A1(n9005), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9026) );
  INV_X1 U11600 ( .A(n13929), .ZN(n9006) );
  XOR2_X1 U11601 ( .A(n14306), .B(n13943), .Z(n14298) );
  XNOR2_X1 U11602 ( .A(n14469), .B(n13942), .ZN(n14287) );
  OR2_X1 U11603 ( .A1(n8788), .A2(n10558), .ZN(n9009) );
  NAND2_X1 U11604 ( .A1(n11969), .A2(n9009), .ZN(n15661) );
  XNOR2_X1 U11605 ( .A(n11683), .B(n13951), .ZN(n11992) );
  XNOR2_X1 U11606 ( .A(n14339), .B(n13945), .ZN(n14332) );
  XNOR2_X1 U11607 ( .A(n14357), .B(n13946), .ZN(n14348) );
  NAND2_X1 U11608 ( .A1(n9014), .A2(n9013), .ZN(n14240) );
  NOR4_X1 U11609 ( .A1(n14175), .A2(n9017), .A3(n9016), .A4(n9015), .ZN(n9018)
         );
  XNOR2_X1 U11610 ( .A(n14097), .B(n13928), .ZN(n9020) );
  INV_X1 U11611 ( .A(n9026), .ZN(n11741) );
  NOR3_X1 U11612 ( .A1(n9022), .A2(n6562), .A3(n11741), .ZN(n9023) );
  NOR4_X1 U11613 ( .A1(n10038), .A2(n15699), .A3(n13915), .A4(n8399), .ZN(
        n9025) );
  AOI211_X1 U11614 ( .C1(n9026), .C2(n11491), .A(n15938), .B(n9025), .ZN(n9027) );
  INV_X1 U11615 ( .A(n9161), .ZN(n9029) );
  NAND2_X1 U11616 ( .A1(n9030), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9031) );
  NAND2_X1 U11617 ( .A1(n9163), .A2(n9031), .ZN(n9154) );
  NAND2_X1 U11618 ( .A1(n10053), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9033) );
  NAND2_X1 U11619 ( .A1(n10095), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n9032) );
  AND2_X1 U11620 ( .A1(n9033), .A2(n9032), .ZN(n9153) );
  NAND2_X1 U11621 ( .A1(n10890), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n9034) );
  NAND2_X1 U11622 ( .A1(n16025), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n9036) );
  NAND2_X1 U11623 ( .A1(n10076), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n9038) );
  NAND2_X1 U11624 ( .A1(n10087), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9040) );
  NAND2_X1 U11625 ( .A1(n10124), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n9041) );
  NAND2_X1 U11626 ( .A1(n9042), .A2(n9041), .ZN(n9244) );
  NAND2_X1 U11627 ( .A1(n10121), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n9043) );
  NAND2_X1 U11628 ( .A1(n10174), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9046) );
  NAND2_X1 U11629 ( .A1(n10168), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n9045) );
  NAND2_X1 U11630 ( .A1(n10179), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U11631 ( .A1(n16097), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U11632 ( .A1(n10201), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9049) );
  XNOR2_X1 U11633 ( .A(n9052), .B(P1_DATAO_REG_12__SCAN_IN), .ZN(n9321) );
  INV_X1 U11634 ( .A(n9321), .ZN(n9051) );
  NAND2_X1 U11635 ( .A1(n9052), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9053) );
  NAND2_X1 U11636 ( .A1(n10554), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9056) );
  NAND2_X1 U11637 ( .A1(n10309), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n9054) );
  AND2_X1 U11638 ( .A1(n9056), .A2(n9054), .ZN(n9055) );
  AND2_X1 U11639 ( .A1(n10316), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9057) );
  INV_X1 U11640 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U11641 ( .A1(n9057), .A2(n9056), .B1(P1_DATAO_REG_14__SCAN_IN), 
        .B2(n10553), .ZN(n9058) );
  XNOR2_X1 U11642 ( .A(n10641), .B(P2_DATAO_REG_15__SCAN_IN), .ZN(n9367) );
  INV_X1 U11643 ( .A(n9367), .ZN(n9059) );
  INV_X1 U11644 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9060) );
  NAND2_X1 U11645 ( .A1(n9060), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9061) );
  XNOR2_X1 U11646 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n9380) );
  NAND2_X1 U11647 ( .A1(n10545), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9063) );
  XNOR2_X1 U11648 ( .A(n10644), .B(P2_DATAO_REG_17__SCAN_IN), .ZN(n9399) );
  INV_X1 U11649 ( .A(n9399), .ZN(n9064) );
  NAND2_X1 U11650 ( .A1(n16042), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n9065) );
  XNOR2_X1 U11651 ( .A(n15896), .B(P2_DATAO_REG_18__SCAN_IN), .ZN(n9411) );
  INV_X1 U11652 ( .A(n9411), .ZN(n9066) );
  NAND2_X1 U11653 ( .A1(n11107), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9067) );
  XNOR2_X1 U11654 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .ZN(n9422) );
  INV_X1 U11655 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11145) );
  NAND2_X1 U11656 ( .A1(n11145), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9069) );
  INV_X1 U11657 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16016) );
  NAND2_X1 U11658 ( .A1(n16016), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9455) );
  OAI21_X1 U11659 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(n11284), .A(n9455), 
        .ZN(n9070) );
  NAND3_X1 U11660 ( .A1(n9455), .A2(P2_DATAO_REG_20__SCAN_IN), .A3(n11284), 
        .ZN(n9071) );
  NAND2_X1 U11661 ( .A1(n15958), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9454) );
  NAND2_X1 U11662 ( .A1(n15835), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9075) );
  INV_X1 U11663 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9073) );
  NAND2_X1 U11664 ( .A1(n9073), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9074) );
  NAND2_X1 U11665 ( .A1(n11743), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9077) );
  INV_X1 U11666 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n15918) );
  NAND2_X1 U11667 ( .A1(n15918), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9076) );
  AND2_X1 U11668 ( .A1(n9077), .A2(n9076), .ZN(n9480) );
  INV_X1 U11669 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11787) );
  AND2_X1 U11670 ( .A1(n11894), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9080) );
  NAND2_X1 U11671 ( .A1(n11898), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9081) );
  AND2_X1 U11672 ( .A1(n16023), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9082) );
  NAND2_X1 U11673 ( .A1(n12586), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9083) );
  NAND2_X1 U11674 ( .A1(n12239), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9084) );
  INV_X1 U11675 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12462) );
  XNOR2_X1 U11676 ( .A(n14589), .B(P2_DATAO_REG_29__SCAN_IN), .ZN(n9548) );
  INV_X1 U11677 ( .A(n9548), .ZN(n9086) );
  NAND2_X1 U11678 ( .A1(n9549), .A2(n9086), .ZN(n9088) );
  NAND2_X1 U11679 ( .A1(n15376), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9087) );
  NAND2_X1 U11680 ( .A1(n9088), .A2(n9087), .ZN(n9138) );
  XNOR2_X1 U11681 ( .A(n12595), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n9137) );
  NAND2_X1 U11682 ( .A1(n12595), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9089) );
  OAI21_X1 U11683 ( .B1(n9138), .B2(n9137), .A(n9089), .ZN(n9091) );
  XNOR2_X1 U11684 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n9090) );
  XNOR2_X1 U11685 ( .A(n9091), .B(n9090), .ZN(n13710) );
  NOR2_X2 U11686 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n9092) );
  NAND4_X1 U11687 ( .A1(n9092), .A2(n9812), .A3(n7627), .A4(n9729), .ZN(n9095)
         );
  NOR2_X2 U11688 ( .A1(n9095), .A2(n9323), .ZN(n9736) );
  NOR2_X1 U11689 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), 
        .ZN(n9097) );
  NOR2_X1 U11690 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), 
        .ZN(n9096) );
  INV_X1 U11691 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9384) );
  NOR2_X1 U11692 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), 
        .ZN(n9100) );
  NAND2_X4 U11693 ( .A1(n6559), .A2(n10885), .ZN(n9202) );
  INV_X1 U11694 ( .A(SI_31_), .ZN(n13705) );
  OR2_X1 U11695 ( .A1(n9202), .A2(n13705), .ZN(n9108) );
  INV_X1 U11696 ( .A(n9212), .ZN(n9111) );
  INV_X1 U11697 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n9118) );
  INV_X1 U11698 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n9121) );
  INV_X1 U11699 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n9123) );
  INV_X1 U11700 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n16003) );
  INV_X1 U11701 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n15924) );
  NAND2_X1 U11702 ( .A1(n16003), .A2(n15924), .ZN(n9125) );
  INV_X1 U11703 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n9126) );
  NAND2_X2 U11704 ( .A1(n9131), .A2(n9132), .ZN(n9177) );
  INV_X1 U11705 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n13621) );
  NAND2_X1 U11706 ( .A1(n9554), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n9134) );
  INV_X1 U11707 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n16010) );
  OR2_X1 U11708 ( .A1(n9175), .A2(n16010), .ZN(n9133) );
  OAI211_X1 U11709 ( .C1(n9211), .C2(n13621), .A(n9134), .B(n9133), .ZN(n9135)
         );
  INV_X1 U11710 ( .A(n9135), .ZN(n9136) );
  XNOR2_X1 U11711 ( .A(n9138), .B(n9137), .ZN(n13712) );
  NAND2_X1 U11712 ( .A1(n13712), .A2(n9550), .ZN(n9140) );
  INV_X1 U11713 ( .A(SI_30_), .ZN(n16017) );
  OR2_X1 U11714 ( .A1(n9202), .A2(n16017), .ZN(n9139) );
  INV_X1 U11715 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n13625) );
  NAND2_X1 U11716 ( .A1(n9554), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9142) );
  NAND2_X1 U11717 ( .A1(n9553), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9141) );
  OAI211_X1 U11718 ( .C1(n13625), .C2(n9211), .A(n9142), .B(n9141), .ZN(n9143)
         );
  INV_X1 U11719 ( .A(n9143), .ZN(n9144) );
  NAND2_X1 U11720 ( .A1(n13622), .A2(n12004), .ZN(n9145) );
  NAND2_X1 U11721 ( .A1(n9554), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9150) );
  INV_X1 U11722 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15791) );
  OR2_X1 U11723 ( .A1(n9175), .A2(n15791), .ZN(n9149) );
  INV_X1 U11724 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n9146) );
  OR2_X1 U11725 ( .A1(n9211), .A2(n9146), .ZN(n9148) );
  INV_X1 U11726 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10767) );
  OR2_X1 U11727 ( .A1(n9177), .A2(n10767), .ZN(n9147) );
  INV_X1 U11728 ( .A(n9980), .ZN(n9151) );
  INV_X1 U11729 ( .A(n10106), .ZN(n10755) );
  OR2_X1 U11730 ( .A1(n9202), .A2(SI_2_), .ZN(n9156) );
  OAI21_X1 U11731 ( .B1(n9154), .B2(n9153), .A(n9152), .ZN(n10103) );
  OR2_X1 U11732 ( .A1(n9256), .A2(n10103), .ZN(n9155) );
  OAI211_X1 U11733 ( .C1(n10755), .C2(n8022), .A(n9156), .B(n9155), .ZN(n9767)
         );
  INV_X1 U11734 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11062) );
  INV_X1 U11735 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n9157) );
  INV_X1 U11736 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10713) );
  INV_X1 U11737 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n15964) );
  NAND2_X1 U11738 ( .A1(n15964), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9158) );
  AND2_X1 U11739 ( .A1(n9161), .A2(n9158), .ZN(n9160) );
  OAI21_X1 U11740 ( .B1(n10885), .B2(n9160), .A(n9159), .ZN(n13725) );
  MUX2_X1 U11741 ( .A(P3_IR_REG_0__SCAN_IN), .B(n13725), .S(n8022), .Z(n9766)
         );
  INV_X1 U11742 ( .A(n11055), .ZN(n9172) );
  OR2_X1 U11743 ( .A1(n9202), .A2(n10101), .ZN(n9167) );
  NAND2_X1 U11744 ( .A1(n9162), .A2(n9161), .ZN(n9164) );
  AND2_X1 U11745 ( .A1(n9163), .A2(n9164), .ZN(n10102) );
  OR2_X1 U11746 ( .A1(n9256), .A2(n10102), .ZN(n9166) );
  INV_X1 U11747 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15789) );
  OR2_X1 U11748 ( .A1(n9175), .A2(n15789), .ZN(n9171) );
  INV_X1 U11749 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n9168) );
  INV_X1 U11750 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11089) );
  OR2_X1 U11751 ( .A1(n9177), .A2(n11089), .ZN(n9169) );
  NAND2_X1 U11752 ( .A1(n9172), .A2(n9708), .ZN(n10526) );
  INV_X2 U11753 ( .A(n11046), .ZN(n9173) );
  NAND2_X1 U11754 ( .A1(n9585), .A2(n10758), .ZN(n9174) );
  OR2_X1 U11755 ( .A1(n13120), .A2(n9767), .ZN(n9584) );
  NAND2_X1 U11756 ( .A1(n9554), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9181) );
  INV_X1 U11757 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15793) );
  OR2_X1 U11758 ( .A1(n9175), .A2(n15793), .ZN(n9180) );
  INV_X1 U11759 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n9176) );
  OR2_X1 U11760 ( .A1(n9211), .A2(n9176), .ZN(n9179) );
  OR2_X1 U11761 ( .A1(n9177), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n9178) );
  NAND4_X1 U11762 ( .A1(n9181), .A2(n9180), .A3(n9179), .A4(n9178), .ZN(n11241) );
  OR2_X1 U11763 ( .A1(n9202), .A2(SI_3_), .ZN(n9188) );
  OR2_X1 U11764 ( .A1(n9184), .A2(n9183), .ZN(n9185) );
  NAND2_X1 U11765 ( .A1(n9186), .A2(n9185), .ZN(n10060) );
  OR2_X1 U11766 ( .A1(n9256), .A2(n10060), .ZN(n9187) );
  OAI211_X1 U11767 ( .C1(n10739), .C2(n8022), .A(n9188), .B(n9187), .ZN(n10810) );
  NAND2_X1 U11768 ( .A1(n11241), .A2(n10810), .ZN(n9595) );
  NAND2_X1 U11769 ( .A1(n9594), .A2(n9595), .ZN(n10802) );
  INV_X1 U11770 ( .A(n10802), .ZN(n10800) );
  NAND2_X1 U11771 ( .A1(n10799), .A2(n10800), .ZN(n9189) );
  NAND2_X1 U11772 ( .A1(n9189), .A2(n9594), .ZN(n11234) );
  NAND2_X1 U11773 ( .A1(n9554), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9195) );
  INV_X1 U11774 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15795) );
  OR2_X1 U11775 ( .A1(n9175), .A2(n15795), .ZN(n9194) );
  NAND2_X1 U11776 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9190) );
  AND2_X1 U11777 ( .A1(n9212), .A2(n9190), .ZN(n11237) );
  OR2_X1 U11778 ( .A1(n9177), .A2(n11237), .ZN(n9193) );
  INV_X1 U11779 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n9191) );
  OR2_X1 U11780 ( .A1(n9211), .A2(n9191), .ZN(n9192) );
  NAND4_X1 U11781 ( .A1(n9195), .A2(n9194), .A3(n9193), .A4(n9192), .ZN(n13119) );
  NAND2_X1 U11782 ( .A1(n9198), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9197) );
  MUX2_X1 U11783 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9197), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n9201) );
  INV_X1 U11784 ( .A(n10991), .ZN(n9209) );
  OR2_X1 U11785 ( .A1(n9202), .A2(SI_4_), .ZN(n9208) );
  OR2_X1 U11786 ( .A1(n9204), .A2(n9203), .ZN(n9205) );
  NAND2_X1 U11787 ( .A1(n9206), .A2(n9205), .ZN(n10057) );
  OR2_X1 U11788 ( .A1(n9256), .A2(n10057), .ZN(n9207) );
  OAI211_X1 U11789 ( .C1(n9209), .C2(n8022), .A(n9208), .B(n9207), .ZN(n11236)
         );
  OR2_X1 U11790 ( .A1(n13119), .A2(n11236), .ZN(n9599) );
  NAND2_X1 U11791 ( .A1(n13119), .A2(n11236), .ZN(n9598) );
  NAND2_X1 U11792 ( .A1(n9599), .A2(n9598), .ZN(n11240) );
  INV_X1 U11793 ( .A(n11240), .ZN(n11235) );
  NAND2_X1 U11794 ( .A1(n11234), .A2(n11235), .ZN(n9210) );
  NAND2_X1 U11795 ( .A1(n9210), .A2(n9599), .ZN(n11360) );
  NAND2_X1 U11796 ( .A1(n9531), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9217) );
  INV_X1 U11797 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15797) );
  OR2_X1 U11798 ( .A1(n9175), .A2(n15797), .ZN(n9216) );
  INV_X1 U11799 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15939) );
  OR2_X1 U11800 ( .A1(n9436), .A2(n15939), .ZN(n9215) );
  NAND2_X1 U11801 ( .A1(n9212), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n9213) );
  AND2_X1 U11802 ( .A1(n9226), .A2(n9213), .ZN(n11362) );
  OR2_X1 U11803 ( .A1(n9177), .A2(n11362), .ZN(n9214) );
  NAND4_X1 U11804 ( .A1(n9217), .A2(n9216), .A3(n9215), .A4(n9214), .ZN(n13118) );
  OR2_X1 U11805 ( .A1(n9219), .A2(n9218), .ZN(n9220) );
  NAND2_X1 U11806 ( .A1(n9221), .A2(n9220), .ZN(n10112) );
  OR2_X1 U11807 ( .A1(n9256), .A2(n10112), .ZN(n9225) );
  OR2_X1 U11808 ( .A1(n9202), .A2(SI_5_), .ZN(n9224) );
  NAND2_X1 U11809 ( .A1(n9232), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9222) );
  XNOR2_X1 U11810 ( .A(n9222), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10779) );
  OR2_X1 U11811 ( .A1(n8022), .A2(n10779), .ZN(n9223) );
  NAND2_X1 U11812 ( .A1(n13118), .A2(n15769), .ZN(n9605) );
  NAND2_X1 U11813 ( .A1(n9603), .A2(n9605), .ZN(n11361) );
  NAND2_X1 U11814 ( .A1(n9531), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9231) );
  INV_X1 U11815 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15799) );
  OR2_X1 U11816 ( .A1(n9175), .A2(n15799), .ZN(n9230) );
  INV_X1 U11817 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n16060) );
  OR2_X1 U11818 ( .A1(n9436), .A2(n16060), .ZN(n9229) );
  NAND2_X1 U11819 ( .A1(n9226), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9227) );
  AND2_X1 U11820 ( .A1(n9238), .A2(n9227), .ZN(n11412) );
  OR2_X1 U11821 ( .A1(n9177), .A2(n11412), .ZN(n9228) );
  INV_X2 U11822 ( .A(n8022), .ZN(n9428) );
  NAND2_X1 U11823 ( .A1(n9246), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9233) );
  XNOR2_X1 U11824 ( .A(n9233), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10952) );
  AOI22_X1 U11825 ( .A1(n9429), .A2(SI_6_), .B1(n9428), .B2(n10952), .ZN(n9237) );
  XNOR2_X1 U11826 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n9234) );
  XNOR2_X1 U11827 ( .A(n9235), .B(n9234), .ZN(n10064) );
  NAND2_X1 U11828 ( .A1(n10064), .A2(n9550), .ZN(n9236) );
  NAND2_X1 U11829 ( .A1(n13117), .A2(n11411), .ZN(n9607) );
  NAND2_X1 U11830 ( .A1(n9609), .A2(n9607), .ZN(n11402) );
  INV_X1 U11831 ( .A(n11402), .ZN(n11399) );
  NAND2_X1 U11832 ( .A1(n9531), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9243) );
  INV_X1 U11833 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15802) );
  OR2_X1 U11834 ( .A1(n9175), .A2(n15802), .ZN(n9242) );
  NAND2_X1 U11835 ( .A1(n9238), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9239) );
  AND2_X1 U11836 ( .A1(n9263), .A2(n9239), .ZN(n11469) );
  OR2_X1 U11837 ( .A1(n9177), .A2(n11469), .ZN(n9241) );
  INV_X1 U11838 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11426) );
  OR2_X1 U11839 ( .A1(n9436), .A2(n11426), .ZN(n9240) );
  NAND4_X1 U11840 ( .A1(n9243), .A2(n9242), .A3(n9241), .A4(n9240), .ZN(n13116) );
  XNOR2_X1 U11841 ( .A(n9245), .B(n9244), .ZN(n10080) );
  NAND2_X1 U11842 ( .A1(n10080), .A2(n9550), .ZN(n9251) );
  INV_X1 U11843 ( .A(SI_7_), .ZN(n10079) );
  INV_X1 U11844 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9247) );
  NAND2_X1 U11845 ( .A1(n9257), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9249) );
  INV_X1 U11846 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9248) );
  XNOR2_X1 U11847 ( .A(n9249), .B(n9248), .ZN(n10965) );
  AOI22_X1 U11848 ( .A1(n9429), .A2(n10079), .B1(n9428), .B2(n10965), .ZN(
        n9250) );
  NAND2_X1 U11849 ( .A1(n9251), .A2(n9250), .ZN(n11427) );
  NAND2_X1 U11850 ( .A1(n13116), .A2(n11427), .ZN(n9611) );
  OR2_X1 U11851 ( .A1(n9253), .A2(n9252), .ZN(n9254) );
  NAND2_X1 U11852 ( .A1(n9255), .A2(n9254), .ZN(n10078) );
  OR2_X1 U11853 ( .A1(n10078), .A2(n9256), .ZN(n9262) );
  NAND2_X1 U11854 ( .A1(n9259), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9258) );
  MUX2_X1 U11855 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9258), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n9260) );
  INV_X1 U11856 ( .A(n11568), .ZN(n11560) );
  AOI22_X1 U11857 ( .A1(n9428), .A2(n11560), .B1(n9429), .B2(SI_8_), .ZN(n9261) );
  NAND2_X1 U11858 ( .A1(n9554), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9269) );
  INV_X1 U11859 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11559) );
  OR2_X1 U11860 ( .A1(n9175), .A2(n11559), .ZN(n9268) );
  NAND2_X1 U11861 ( .A1(n9263), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9264) );
  AND2_X1 U11862 ( .A1(n9281), .A2(n9264), .ZN(n11763) );
  OR2_X1 U11863 ( .A1(n9177), .A2(n11763), .ZN(n9267) );
  INV_X1 U11864 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n9265) );
  OR2_X1 U11865 ( .A1(n9211), .A2(n9265), .ZN(n9266) );
  NAND4_X1 U11866 ( .A1(n9269), .A2(n9268), .A3(n9267), .A4(n9266), .ZN(n13114) );
  NAND2_X1 U11867 ( .A1(n11720), .A2(n13114), .ZN(n9615) );
  INV_X1 U11868 ( .A(n13114), .ZN(n9776) );
  NAND2_X1 U11869 ( .A1(n11767), .A2(n9776), .ZN(n9616) );
  NAND2_X1 U11870 ( .A1(n11371), .A2(n9775), .ZN(n9270) );
  NAND2_X1 U11871 ( .A1(n9270), .A2(n9616), .ZN(n11770) );
  OR2_X1 U11872 ( .A1(n9272), .A2(n9271), .ZN(n9273) );
  NAND2_X1 U11873 ( .A1(n9274), .A2(n9273), .ZN(n10108) );
  NAND2_X1 U11874 ( .A1(n10108), .A2(n9550), .ZN(n9280) );
  NAND2_X1 U11875 ( .A1(n9276), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9275) );
  MUX2_X1 U11876 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9275), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n9278) );
  INV_X1 U11877 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9277) );
  NAND2_X1 U11878 ( .A1(n9278), .A2(n9308), .ZN(n11569) );
  INV_X1 U11879 ( .A(SI_9_), .ZN(n10107) );
  AOI22_X1 U11880 ( .A1(n11569), .A2(n9428), .B1(n9429), .B2(n10107), .ZN(
        n9279) );
  NAND2_X1 U11881 ( .A1(n9554), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n9287) );
  INV_X1 U11882 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11983) );
  OR2_X1 U11883 ( .A1(n9175), .A2(n11983), .ZN(n9286) );
  NAND2_X1 U11884 ( .A1(n9281), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n9282) );
  AND2_X1 U11885 ( .A1(n9299), .A2(n9282), .ZN(n11794) );
  OR2_X1 U11886 ( .A1(n9177), .A2(n11794), .ZN(n9285) );
  INV_X1 U11887 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n9283) );
  OR2_X1 U11888 ( .A1(n9211), .A2(n9283), .ZN(n9284) );
  NOR2_X1 U11889 ( .A1(n11985), .A2(n11759), .ZN(n9289) );
  NAND2_X1 U11890 ( .A1(n11985), .A2(n11759), .ZN(n9288) );
  OR2_X1 U11891 ( .A1(n9291), .A2(n9290), .ZN(n9292) );
  NAND2_X1 U11892 ( .A1(n9293), .A2(n9292), .ZN(n10111) );
  NAND2_X1 U11893 ( .A1(n10111), .A2(n9550), .ZN(n9298) );
  NAND2_X1 U11894 ( .A1(n9308), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9295) );
  INV_X1 U11895 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9294) );
  NOR2_X1 U11896 ( .A1(n9202), .A2(SI_10_), .ZN(n9296) );
  AOI21_X1 U11897 ( .B1(n13124), .B2(n9428), .A(n9296), .ZN(n9297) );
  NAND2_X1 U11898 ( .A1(n9554), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n9305) );
  INV_X1 U11899 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n13133) );
  OR2_X1 U11900 ( .A1(n9175), .A2(n13133), .ZN(n9304) );
  NAND2_X1 U11901 ( .A1(n9299), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9300) );
  AND2_X1 U11902 ( .A1(n9314), .A2(n9300), .ZN(n11907) );
  OR2_X1 U11903 ( .A1(n9177), .A2(n11907), .ZN(n9303) );
  INV_X1 U11904 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n9301) );
  OR2_X1 U11905 ( .A1(n9211), .A2(n9301), .ZN(n9302) );
  NAND4_X1 U11906 ( .A1(n9305), .A2(n9304), .A3(n9303), .A4(n9302), .ZN(n13113) );
  OR2_X1 U11907 ( .A1(n12053), .A2(n13113), .ZN(n9620) );
  NAND2_X1 U11908 ( .A1(n12053), .A2(n13113), .ZN(n9621) );
  NAND2_X1 U11909 ( .A1(n9620), .A2(n9621), .ZN(n9780) );
  XNOR2_X1 U11910 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9306) );
  XNOR2_X1 U11911 ( .A(n9307), .B(n9306), .ZN(n10167) );
  NAND2_X1 U11912 ( .A1(n10167), .A2(n9550), .ZN(n9313) );
  OAI21_X1 U11913 ( .B1(n9308), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9310) );
  INV_X1 U11914 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9309) );
  NOR2_X1 U11915 ( .A1(n9202), .A2(SI_11_), .ZN(n9311) );
  AOI21_X1 U11916 ( .B1(n13153), .B2(n9428), .A(n9311), .ZN(n9312) );
  NAND2_X1 U11917 ( .A1(n9313), .A2(n9312), .ZN(n12003) );
  NAND2_X1 U11918 ( .A1(n9314), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9315) );
  AND2_X1 U11919 ( .A1(n9332), .A2(n9315), .ZN(n11900) );
  OR2_X1 U11920 ( .A1(n9177), .A2(n11900), .ZN(n9320) );
  INV_X1 U11921 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n13136) );
  OR2_X1 U11922 ( .A1(n9175), .A2(n13136), .ZN(n9319) );
  INV_X1 U11923 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n9316) );
  OR2_X1 U11924 ( .A1(n9211), .A2(n9316), .ZN(n9318) );
  INV_X1 U11925 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11899) );
  OR2_X1 U11926 ( .A1(n9436), .A2(n11899), .ZN(n9317) );
  NAND4_X1 U11927 ( .A1(n9320), .A2(n9319), .A3(n9318), .A4(n9317), .ZN(n13112) );
  NAND2_X1 U11928 ( .A1(n12003), .A2(n13112), .ZN(n9625) );
  NAND2_X1 U11929 ( .A1(n9624), .A2(n9625), .ZN(n11782) );
  XNOR2_X1 U11930 ( .A(n9322), .B(n9321), .ZN(n10182) );
  NAND2_X1 U11931 ( .A1(n10182), .A2(n9550), .ZN(n9331) );
  NAND2_X1 U11932 ( .A1(n9328), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9327) );
  MUX2_X1 U11933 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9327), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n9329) );
  AND2_X1 U11934 ( .A1(n9570), .A2(n9329), .ZN(n13171) );
  AOI22_X1 U11935 ( .A1(n9429), .A2(SI_12_), .B1(n9428), .B2(n13171), .ZN(
        n9330) );
  NAND2_X1 U11936 ( .A1(n9332), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9333) );
  NAND2_X1 U11937 ( .A1(n9343), .A2(n9333), .ZN(n12110) );
  NAND2_X1 U11938 ( .A1(n9547), .A2(n12110), .ZN(n9338) );
  INV_X1 U11939 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n13162) );
  OR2_X1 U11940 ( .A1(n9436), .A2(n13162), .ZN(n9337) );
  INV_X1 U11941 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n15909) );
  OR2_X1 U11942 ( .A1(n9175), .A2(n15909), .ZN(n9336) );
  INV_X1 U11943 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n9334) );
  OR2_X1 U11944 ( .A1(n9211), .A2(n9334), .ZN(n9335) );
  OR2_X1 U11945 ( .A1(n12113), .A2(n13059), .ZN(n9628) );
  NAND2_X1 U11946 ( .A1(n12113), .A2(n13059), .ZN(n9629) );
  NAND2_X1 U11947 ( .A1(n9628), .A2(n9629), .ZN(n12103) );
  XNOR2_X1 U11948 ( .A(n9349), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10282) );
  NAND2_X1 U11949 ( .A1(n10282), .A2(n9550), .ZN(n9342) );
  NAND2_X1 U11950 ( .A1(n9570), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9339) );
  MUX2_X1 U11951 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9339), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n9340) );
  INV_X1 U11952 ( .A(n9424), .ZN(n9355) );
  NAND2_X1 U11953 ( .A1(n9340), .A2(n9355), .ZN(n13207) );
  AOI22_X1 U11954 ( .A1(n9429), .A2(n10281), .B1(n9428), .B2(n13207), .ZN(
        n9341) );
  NAND2_X1 U11955 ( .A1(n9343), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9344) );
  NAND2_X1 U11956 ( .A1(n9361), .A2(n9344), .ZN(n13556) );
  NAND2_X1 U11957 ( .A1(n9547), .A2(n13556), .ZN(n9348) );
  INV_X1 U11958 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13554) );
  OR2_X1 U11959 ( .A1(n9436), .A2(n13554), .ZN(n9347) );
  INV_X1 U11960 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n13613) );
  OR2_X1 U11961 ( .A1(n9175), .A2(n13613), .ZN(n9346) );
  INV_X1 U11962 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n15873) );
  OR2_X1 U11963 ( .A1(n9211), .A2(n15873), .ZN(n9345) );
  NOR2_X1 U11964 ( .A1(n13555), .A2(n12106), .ZN(n9633) );
  NAND2_X1 U11965 ( .A1(n13555), .A2(n12106), .ZN(n9637) );
  NAND2_X1 U11966 ( .A1(n9349), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9352) );
  NAND2_X1 U11967 ( .A1(n9350), .A2(n10316), .ZN(n9351) );
  NAND2_X1 U11968 ( .A1(n9352), .A2(n9351), .ZN(n9354) );
  XNOR2_X1 U11969 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n9353) );
  XNOR2_X1 U11970 ( .A(n9354), .B(n9353), .ZN(n10305) );
  NAND2_X1 U11971 ( .A1(n10305), .A2(n9550), .ZN(n9360) );
  INV_X1 U11972 ( .A(SI_14_), .ZN(n10304) );
  NAND2_X1 U11973 ( .A1(n9355), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9356) );
  MUX2_X1 U11974 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9356), .S(
        P3_IR_REG_14__SCAN_IN), .Z(n9358) );
  INV_X1 U11975 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9357) );
  NAND2_X1 U11976 ( .A1(n9424), .A2(n9357), .ZN(n9383) );
  NAND2_X1 U11977 ( .A1(n9358), .A2(n9383), .ZN(n13202) );
  AOI22_X1 U11978 ( .A1(n9429), .A2(n10304), .B1(n9428), .B2(n13202), .ZN(
        n9359) );
  NAND2_X1 U11979 ( .A1(n9361), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9362) );
  NAND2_X1 U11980 ( .A1(n9372), .A2(n9362), .ZN(n13528) );
  NAND2_X1 U11981 ( .A1(n13528), .A2(n9547), .ZN(n9366) );
  NAND2_X1 U11982 ( .A1(n9554), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9365) );
  NAND2_X1 U11983 ( .A1(n9553), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9364) );
  NAND2_X1 U11984 ( .A1(n9531), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9363) );
  NAND4_X1 U11985 ( .A1(n9366), .A2(n9365), .A3(n9364), .A4(n9363), .ZN(n13548) );
  NAND2_X1 U11986 ( .A1(n13689), .A2(n13548), .ZN(n9639) );
  INV_X1 U11987 ( .A(n9639), .ZN(n9377) );
  XNOR2_X1 U11988 ( .A(n9368), .B(n9367), .ZN(n10283) );
  NAND2_X1 U11989 ( .A1(n10283), .A2(n9550), .ZN(n9371) );
  NAND2_X1 U11990 ( .A1(n9383), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9369) );
  XNOR2_X1 U11991 ( .A(n9369), .B(P3_IR_REG_15__SCAN_IN), .ZN(n13256) );
  AOI22_X1 U11992 ( .A1(n9429), .A2(SI_15_), .B1(n9428), .B2(n13256), .ZN(
        n9370) );
  NAND2_X1 U11993 ( .A1(n9372), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9373) );
  NAND2_X1 U11994 ( .A1(n9395), .A2(n9373), .ZN(n13513) );
  NAND2_X1 U11995 ( .A1(n13513), .A2(n9547), .ZN(n9376) );
  AOI22_X1 U11996 ( .A1(n9553), .A2(P3_REG1_REG_15__SCAN_IN), .B1(n9554), .B2(
        P3_REG2_REG_15__SCAN_IN), .ZN(n9375) );
  NAND2_X1 U11997 ( .A1(n9531), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9374) );
  NAND2_X1 U11998 ( .A1(n13685), .A2(n13536), .ZN(n9643) );
  INV_X1 U11999 ( .A(n9643), .ZN(n9378) );
  AOI21_X1 U12000 ( .B1(n13511), .B2(n9638), .A(n9378), .ZN(n9379) );
  INV_X1 U12001 ( .A(n9380), .ZN(n9381) );
  XNOR2_X1 U12002 ( .A(n9382), .B(n9381), .ZN(n10306) );
  NAND2_X1 U12003 ( .A1(n10306), .A2(n9550), .ZN(n9393) );
  INV_X1 U12004 ( .A(n9383), .ZN(n9385) );
  AND2_X1 U12005 ( .A1(n9385), .A2(n9384), .ZN(n9389) );
  INV_X1 U12006 ( .A(n9389), .ZN(n9386) );
  NAND2_X1 U12007 ( .A1(n9386), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9387) );
  MUX2_X1 U12008 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9387), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n9390) );
  INV_X1 U12009 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n9388) );
  NAND2_X1 U12010 ( .A1(n9389), .A2(n9388), .ZN(n9413) );
  NAND2_X1 U12011 ( .A1(n9390), .A2(n9413), .ZN(n13257) );
  OAI22_X1 U12012 ( .A1(n13257), .A2(n8022), .B1(n9202), .B2(n10307), .ZN(
        n9391) );
  INV_X1 U12013 ( .A(n9391), .ZN(n9392) );
  INV_X1 U12014 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13678) );
  INV_X1 U12015 ( .A(n9394), .ZN(n9404) );
  NAND2_X1 U12016 ( .A1(n9395), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9396) );
  NAND2_X1 U12017 ( .A1(n9404), .A2(n9396), .ZN(n13508) );
  NAND2_X1 U12018 ( .A1(n13508), .A2(n9547), .ZN(n9398) );
  AOI22_X1 U12019 ( .A1(n9553), .A2(P3_REG1_REG_16__SCAN_IN), .B1(n9554), .B2(
        P3_REG2_REG_16__SCAN_IN), .ZN(n9397) );
  OAI211_X1 U12020 ( .C1(n9211), .C2(n13678), .A(n9398), .B(n9397), .ZN(n13519) );
  INV_X1 U12021 ( .A(n13519), .ZN(n13489) );
  OR2_X1 U12022 ( .A1(n13679), .A2(n13489), .ZN(n9581) );
  NAND2_X1 U12023 ( .A1(n13679), .A2(n13489), .ZN(n9645) );
  NAND2_X1 U12024 ( .A1(n9581), .A2(n9645), .ZN(n13499) );
  INV_X1 U12025 ( .A(n13499), .ZN(n13503) );
  XNOR2_X1 U12026 ( .A(n9400), .B(n9399), .ZN(n10394) );
  NAND2_X1 U12027 ( .A1(n10394), .A2(n9550), .ZN(n9403) );
  NAND2_X1 U12028 ( .A1(n9413), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9401) );
  XNOR2_X1 U12029 ( .A(n9401), .B(P3_IR_REG_17__SCAN_IN), .ZN(n13301) );
  AOI22_X1 U12030 ( .A1(n13301), .A2(n9428), .B1(SI_17_), .B2(n9429), .ZN(
        n9402) );
  NAND2_X1 U12031 ( .A1(n9404), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9405) );
  NAND2_X1 U12032 ( .A1(n9417), .A2(n9405), .ZN(n13495) );
  NAND2_X1 U12033 ( .A1(n13495), .A2(n9547), .ZN(n9410) );
  INV_X1 U12034 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13671) );
  NAND2_X1 U12035 ( .A1(n9554), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n9407) );
  NAND2_X1 U12036 ( .A1(n9553), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9406) );
  OAI211_X1 U12037 ( .C1(n13671), .C2(n9211), .A(n9407), .B(n9406), .ZN(n9408)
         );
  INV_X1 U12038 ( .A(n9408), .ZN(n9409) );
  OR2_X1 U12039 ( .A1(n13672), .A2(n13504), .ZN(n9648) );
  NAND2_X1 U12040 ( .A1(n13672), .A2(n13504), .ZN(n9652) );
  NAND2_X1 U12041 ( .A1(n9648), .A2(n9652), .ZN(n13487) );
  INV_X1 U12042 ( .A(n13487), .ZN(n13485) );
  XNOR2_X1 U12043 ( .A(n9412), .B(n9411), .ZN(n10548) );
  NAND2_X1 U12044 ( .A1(n10548), .A2(n9550), .ZN(n9416) );
  OAI21_X1 U12045 ( .B1(n9413), .B2(P3_IR_REG_17__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9414) );
  XNOR2_X1 U12046 ( .A(n9414), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13302) );
  AOI22_X1 U12047 ( .A1(n13302), .A2(n9428), .B1(SI_18_), .B2(n9429), .ZN(
        n9415) );
  NAND2_X1 U12048 ( .A1(n9417), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9418) );
  NAND2_X1 U12049 ( .A1(n9432), .A2(n9418), .ZN(n13477) );
  INV_X1 U12050 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n16057) );
  NAND2_X1 U12051 ( .A1(n9554), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9420) );
  NAND2_X1 U12052 ( .A1(n9553), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9419) );
  OAI211_X1 U12053 ( .C1(n16057), .C2(n9211), .A(n9420), .B(n9419), .ZN(n9421)
         );
  NAND2_X1 U12054 ( .A1(n13597), .A2(n13490), .ZN(n9655) );
  XNOR2_X1 U12055 ( .A(n9423), .B(n9422), .ZN(n10629) );
  NAND2_X1 U12056 ( .A1(n10629), .A2(n9550), .ZN(n9431) );
  NAND2_X1 U12057 ( .A1(n9424), .A2(n9569), .ZN(n9426) );
  NAND2_X1 U12058 ( .A1(n9426), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9425) );
  MUX2_X1 U12059 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9425), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n9427) );
  AOI22_X1 U12060 ( .A1(n9429), .A2(n10630), .B1(n9428), .B2(n10631), .ZN(
        n9430) );
  NAND2_X2 U12061 ( .A1(n9431), .A2(n9430), .ZN(n13593) );
  NAND2_X1 U12062 ( .A1(n9432), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U12063 ( .A1(n9442), .A2(n9433), .ZN(n13466) );
  NAND2_X1 U12064 ( .A1(n13466), .A2(n9547), .ZN(n9439) );
  INV_X1 U12065 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n15877) );
  NAND2_X1 U12066 ( .A1(n9531), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9435) );
  NAND2_X1 U12067 ( .A1(n9553), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9434) );
  OAI211_X1 U12068 ( .C1(n9436), .C2(n15877), .A(n9435), .B(n9434), .ZN(n9437)
         );
  INV_X1 U12069 ( .A(n9437), .ZN(n9438) );
  NAND2_X1 U12070 ( .A1(n13593), .A2(n13108), .ZN(n9705) );
  XNOR2_X1 U12071 ( .A(n9450), .B(n11281), .ZN(n11248) );
  NAND2_X1 U12072 ( .A1(n11248), .A2(n9550), .ZN(n9441) );
  OR2_X1 U12073 ( .A1(n9202), .A2(n11250), .ZN(n9440) );
  NAND2_X2 U12074 ( .A1(n9441), .A2(n9440), .ZN(n13590) );
  NAND2_X1 U12075 ( .A1(n9442), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9443) );
  NAND2_X1 U12076 ( .A1(n9460), .A2(n9443), .ZN(n13451) );
  NAND2_X1 U12077 ( .A1(n13451), .A2(n9547), .ZN(n9449) );
  INV_X1 U12078 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n9446) );
  NAND2_X1 U12079 ( .A1(n9554), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9445) );
  NAND2_X1 U12080 ( .A1(n9553), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9444) );
  OAI211_X1 U12081 ( .C1(n9446), .C2(n9211), .A(n9445), .B(n9444), .ZN(n9447)
         );
  INV_X1 U12082 ( .A(n9447), .ZN(n9448) );
  OR2_X2 U12083 ( .A1(n13590), .A2(n13460), .ZN(n9659) );
  NAND2_X1 U12084 ( .A1(n13590), .A2(n13460), .ZN(n9660) );
  NAND2_X1 U12085 ( .A1(n9659), .A2(n9660), .ZN(n13445) );
  NAND2_X1 U12086 ( .A1(n9451), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9452) );
  NAND2_X1 U12087 ( .A1(n9453), .A2(n9452), .ZN(n9457) );
  NAND2_X1 U12088 ( .A1(n9455), .A2(n9454), .ZN(n9456) );
  XNOR2_X1 U12089 ( .A(n9457), .B(n9456), .ZN(n11379) );
  NAND2_X1 U12090 ( .A1(n11379), .A2(n9550), .ZN(n9459) );
  INV_X1 U12091 ( .A(SI_21_), .ZN(n11380) );
  OR2_X1 U12092 ( .A1(n9202), .A2(n11380), .ZN(n9458) );
  NAND2_X1 U12093 ( .A1(n9460), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9461) );
  NAND2_X1 U12094 ( .A1(n9472), .A2(n9461), .ZN(n13435) );
  INV_X1 U12095 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13654) );
  NAND2_X1 U12096 ( .A1(n9554), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9463) );
  NAND2_X1 U12097 ( .A1(n9553), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9462) );
  OAI211_X1 U12098 ( .C1(n13654), .C2(n9211), .A(n9463), .B(n9462), .ZN(n9464)
         );
  NAND2_X1 U12099 ( .A1(n13434), .A2(n13446), .ZN(n9664) );
  OR2_X1 U12100 ( .A1(n9466), .A2(n9465), .ZN(n9467) );
  NAND2_X1 U12101 ( .A1(n9468), .A2(n9467), .ZN(n11109) );
  NAND2_X1 U12102 ( .A1(n11109), .A2(n9550), .ZN(n9471) );
  OR2_X1 U12103 ( .A1(n9202), .A2(n9469), .ZN(n9470) );
  NAND2_X1 U12104 ( .A1(n9472), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9473) );
  NAND2_X1 U12105 ( .A1(n9486), .A2(n9473), .ZN(n13424) );
  NAND2_X1 U12106 ( .A1(n13424), .A2(n9547), .ZN(n9478) );
  INV_X1 U12107 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13648) );
  NAND2_X1 U12108 ( .A1(n9553), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9475) );
  NAND2_X1 U12109 ( .A1(n9554), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n9474) );
  OAI211_X1 U12110 ( .C1(n13648), .C2(n9211), .A(n9475), .B(n9474), .ZN(n9476)
         );
  INV_X1 U12111 ( .A(n9476), .ZN(n9477) );
  NAND2_X1 U12112 ( .A1(n13649), .A2(n13433), .ZN(n9667) );
  NAND2_X1 U12113 ( .A1(n9479), .A2(n9666), .ZN(n13408) );
  OR2_X1 U12114 ( .A1(n9481), .A2(n9480), .ZN(n9482) );
  NAND2_X1 U12115 ( .A1(n9483), .A2(n9482), .ZN(n11311) );
  NAND2_X1 U12116 ( .A1(n11311), .A2(n9550), .ZN(n9485) );
  OR2_X1 U12117 ( .A1(n9202), .A2(n11314), .ZN(n9484) );
  NAND2_X1 U12118 ( .A1(n9486), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9487) );
  NAND2_X1 U12119 ( .A1(n9497), .A2(n9487), .ZN(n13411) );
  NAND2_X1 U12120 ( .A1(n13411), .A2(n9547), .ZN(n9492) );
  INV_X1 U12121 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n15999) );
  NAND2_X1 U12122 ( .A1(n9553), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9489) );
  NAND2_X1 U12123 ( .A1(n9554), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9488) );
  OAI211_X1 U12124 ( .C1(n15999), .C2(n9211), .A(n9489), .B(n9488), .ZN(n9490)
         );
  INV_X1 U12125 ( .A(n9490), .ZN(n9491) );
  NAND2_X1 U12126 ( .A1(n13580), .A2(n13069), .ZN(n9493) );
  NAND2_X1 U12127 ( .A1(n9674), .A2(n9493), .ZN(n13404) );
  XNOR2_X1 U12128 ( .A(n9494), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n11700) );
  NAND2_X1 U12129 ( .A1(n11700), .A2(n9550), .ZN(n9496) );
  OR2_X1 U12130 ( .A1(n9202), .A2(n11701), .ZN(n9495) );
  NAND2_X1 U12131 ( .A1(n9497), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9498) );
  NAND2_X1 U12132 ( .A1(n9509), .A2(n9498), .ZN(n13397) );
  NAND2_X1 U12133 ( .A1(n13397), .A2(n9547), .ZN(n9503) );
  INV_X1 U12134 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13641) );
  NAND2_X1 U12135 ( .A1(n9554), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9500) );
  NAND2_X1 U12136 ( .A1(n9553), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9499) );
  OAI211_X1 U12137 ( .C1(n13641), .C2(n9211), .A(n9500), .B(n9499), .ZN(n9501)
         );
  INV_X1 U12138 ( .A(n9501), .ZN(n9502) );
  NAND2_X1 U12139 ( .A1(n13396), .A2(n13406), .ZN(n9672) );
  XNOR2_X1 U12140 ( .A(n11898), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n9505) );
  XNOR2_X1 U12141 ( .A(n9506), .B(n9505), .ZN(n11889) );
  NAND2_X1 U12142 ( .A1(n11889), .A2(n9550), .ZN(n9508) );
  OR2_X1 U12143 ( .A1(n9202), .A2(n11891), .ZN(n9507) );
  NAND2_X2 U12144 ( .A1(n9508), .A2(n9507), .ZN(n13636) );
  NAND2_X1 U12145 ( .A1(n9509), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9510) );
  NAND2_X1 U12146 ( .A1(n9529), .A2(n9510), .ZN(n13379) );
  NAND2_X1 U12147 ( .A1(n13379), .A2(n9547), .ZN(n9515) );
  INV_X1 U12148 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13634) );
  NAND2_X1 U12149 ( .A1(n9554), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9512) );
  NAND2_X1 U12150 ( .A1(n9553), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9511) );
  OAI211_X1 U12151 ( .C1(n13634), .C2(n9211), .A(n9512), .B(n9511), .ZN(n9513)
         );
  INV_X1 U12152 ( .A(n9513), .ZN(n9514) );
  OR2_X1 U12153 ( .A1(n13636), .A2(n13085), .ZN(n9679) );
  NAND2_X1 U12154 ( .A1(n13636), .A2(n13085), .ZN(n9680) );
  AND2_X2 U12155 ( .A1(n9679), .A2(n9680), .ZN(n13370) );
  XNOR2_X1 U12156 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .ZN(n9516) );
  XNOR2_X1 U12157 ( .A(n9517), .B(n9516), .ZN(n12054) );
  OR2_X1 U12158 ( .A1(n9202), .A2(n12055), .ZN(n9518) );
  XNOR2_X1 U12159 ( .A(n9529), .B(P3_REG3_REG_26__SCAN_IN), .ZN(n13366) );
  NAND2_X1 U12160 ( .A1(n13366), .A2(n9547), .ZN(n9523) );
  INV_X1 U12161 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13628) );
  NAND2_X1 U12162 ( .A1(n9553), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9520) );
  NAND2_X1 U12163 ( .A1(n9554), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9519) );
  OAI211_X1 U12164 ( .C1(n9211), .C2(n13628), .A(n9520), .B(n9519), .ZN(n9521)
         );
  INV_X1 U12165 ( .A(n9521), .ZN(n9522) );
  NAND2_X1 U12166 ( .A1(n13362), .A2(n9684), .ZN(n9524) );
  XNOR2_X1 U12167 ( .A(n12239), .B(P2_DATAO_REG_27__SCAN_IN), .ZN(n9525) );
  XNOR2_X1 U12168 ( .A(n9526), .B(n9525), .ZN(n13719) );
  NAND2_X1 U12169 ( .A1(n13719), .A2(n9550), .ZN(n9528) );
  INV_X1 U12170 ( .A(SI_27_), .ZN(n13722) );
  OR2_X1 U12171 ( .A1(n9202), .A2(n13722), .ZN(n9527) );
  OAI21_X1 U12172 ( .B1(n9529), .B2(P3_REG3_REG_26__SCAN_IN), .A(
        P3_REG3_REG_27__SCAN_IN), .ZN(n9530) );
  NAND2_X1 U12173 ( .A1(n9530), .A2(n9542), .ZN(n13357) );
  NAND2_X1 U12174 ( .A1(n13357), .A2(n9547), .ZN(n9536) );
  INV_X1 U12175 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n16073) );
  NAND2_X1 U12176 ( .A1(n9531), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9533) );
  NAND2_X1 U12177 ( .A1(n9554), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9532) );
  OAI211_X1 U12178 ( .C1(n9175), .C2(n16073), .A(n9533), .B(n9532), .ZN(n9534)
         );
  INV_X1 U12179 ( .A(n9534), .ZN(n9535) );
  NAND2_X1 U12180 ( .A1(n13566), .A2(n13089), .ZN(n9753) );
  OR2_X1 U12181 ( .A1(n13566), .A2(n13089), .ZN(n9537) );
  AND2_X2 U12182 ( .A1(n9753), .A2(n9537), .ZN(n13355) );
  XNOR2_X1 U12183 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .ZN(n9538) );
  XNOR2_X1 U12184 ( .A(n9539), .B(n9538), .ZN(n13715) );
  NAND2_X1 U12185 ( .A1(n13715), .A2(n9550), .ZN(n9541) );
  INV_X1 U12186 ( .A(SI_28_), .ZN(n13718) );
  OR2_X1 U12187 ( .A1(n9202), .A2(n13718), .ZN(n9540) );
  NAND2_X1 U12188 ( .A1(n9542), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9543) );
  NAND2_X1 U12189 ( .A1(n9893), .A2(n9543), .ZN(n13343) );
  INV_X1 U12190 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n16000) );
  NAND2_X1 U12191 ( .A1(n9553), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9545) );
  NAND2_X1 U12192 ( .A1(n9554), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9544) );
  OAI211_X1 U12193 ( .C1(n9211), .C2(n16000), .A(n9545), .B(n9544), .ZN(n9546)
         );
  AND2_X1 U12194 ( .A1(n9694), .A2(n9753), .ZN(n9696) );
  XNOR2_X1 U12195 ( .A(n9549), .B(n9548), .ZN(n12240) );
  NAND2_X1 U12196 ( .A1(n12240), .A2(n9550), .ZN(n9552) );
  OR2_X1 U12197 ( .A1(n9202), .A2(n12241), .ZN(n9551) );
  INV_X1 U12198 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9557) );
  NAND2_X1 U12199 ( .A1(n9553), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9556) );
  NAND2_X1 U12200 ( .A1(n9554), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9555) );
  OAI211_X1 U12201 ( .C1(n9211), .C2(n9557), .A(n9556), .B(n9555), .ZN(n9558)
         );
  INV_X1 U12202 ( .A(n9558), .ZN(n9559) );
  NAND2_X1 U12203 ( .A1(n9894), .A2(n12999), .ZN(n9702) );
  NAND2_X1 U12204 ( .A1(n9702), .A2(n10631), .ZN(n9561) );
  AOI21_X1 U12205 ( .B1(n13336), .B2(n13622), .A(n9561), .ZN(n9562) );
  INV_X1 U12206 ( .A(n9563), .ZN(n9565) );
  INV_X1 U12207 ( .A(n13336), .ZN(n12049) );
  NAND3_X1 U12208 ( .A1(n9718), .A2(n13324), .A3(n12049), .ZN(n9566) );
  OAI21_X1 U12209 ( .B1(n13618), .B2(n10631), .A(n9566), .ZN(n9564) );
  OAI21_X1 U12210 ( .B1(n9565), .B2(n9701), .A(n9564), .ZN(n9580) );
  INV_X1 U12211 ( .A(n13618), .ZN(n13339) );
  AOI211_X1 U12212 ( .C1(n12049), .C2(n9718), .A(n13324), .B(n13339), .ZN(
        n9578) );
  AOI211_X1 U12213 ( .C1(n13565), .C2(n9702), .A(n10631), .B(n13618), .ZN(
        n9577) );
  NOR2_X1 U12214 ( .A1(n9566), .A2(n9702), .ZN(n9576) );
  NAND2_X1 U12215 ( .A1(n9569), .A2(n9568), .ZN(n9735) );
  INV_X1 U12216 ( .A(n9574), .ZN(n9571) );
  INV_X1 U12217 ( .A(n11251), .ZN(n9762) );
  NAND2_X1 U12218 ( .A1(n9571), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9572) );
  MUX2_X1 U12219 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9572), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n9575) );
  NAND2_X1 U12220 ( .A1(n9762), .A2(n10521), .ZN(n9805) );
  NOR4_X1 U12221 ( .A1(n9578), .A2(n9577), .A3(n9576), .A4(n9805), .ZN(n9579)
         );
  INV_X1 U12222 ( .A(n9581), .ZN(n9647) );
  NAND2_X1 U12223 ( .A1(n9582), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9583) );
  NAND2_X2 U12224 ( .A1(n11110), .A2(n10521), .ZN(n9855) );
  NAND2_X1 U12225 ( .A1(n9594), .A2(n9584), .ZN(n9588) );
  NAND2_X1 U12226 ( .A1(n13122), .A2(n10715), .ZN(n9707) );
  AND3_X1 U12227 ( .A1(n9708), .A2(n9707), .A3(n11110), .ZN(n9589) );
  NAND2_X1 U12228 ( .A1(n13120), .A2(n9767), .ZN(n9586) );
  OAI211_X1 U12229 ( .C1(n9592), .C2(n9589), .A(n9595), .B(n9586), .ZN(n9587)
         );
  INV_X1 U12230 ( .A(n9589), .ZN(n9590) );
  NAND2_X1 U12231 ( .A1(n9590), .A2(n9707), .ZN(n9591) );
  MUX2_X1 U12232 ( .A(n11055), .B(n9591), .S(n10521), .Z(n9593) );
  MUX2_X1 U12233 ( .A(n9595), .B(n9594), .S(n9961), .Z(n9596) );
  INV_X1 U12234 ( .A(n9598), .ZN(n9601) );
  INV_X1 U12235 ( .A(n9599), .ZN(n9600) );
  MUX2_X1 U12236 ( .A(n9601), .B(n9600), .S(n9961), .Z(n9602) );
  AND2_X1 U12237 ( .A1(n9609), .A2(n9603), .ZN(n9604) );
  AOI21_X1 U12238 ( .B1(n9607), .B2(n9605), .A(n9961), .ZN(n9606) );
  AOI21_X1 U12239 ( .B1(n9608), .B2(n9607), .A(n9606), .ZN(n9614) );
  OAI21_X1 U12240 ( .B1(n9961), .B2(n9609), .A(n11464), .ZN(n9613) );
  MUX2_X1 U12241 ( .A(n9611), .B(n9610), .S(n9961), .Z(n9612) );
  OAI211_X1 U12242 ( .C1(n9614), .C2(n9613), .A(n9775), .B(n9612), .ZN(n9618)
         );
  XNOR2_X1 U12243 ( .A(n11985), .B(n11845), .ZN(n11771) );
  MUX2_X1 U12244 ( .A(n9616), .B(n9615), .S(n9961), .Z(n9617) );
  INV_X1 U12245 ( .A(n11782), .ZN(n11779) );
  INV_X1 U12246 ( .A(n11985), .ZN(n11796) );
  MUX2_X1 U12247 ( .A(n11759), .B(n11796), .S(n9961), .Z(n9619) );
  OR2_X1 U12248 ( .A1(n11985), .A2(n11845), .ZN(n9779) );
  NAND3_X1 U12249 ( .A1(n11843), .A2(n9619), .A3(n9779), .ZN(n9623) );
  MUX2_X1 U12250 ( .A(n9621), .B(n9620), .S(n9961), .Z(n9622) );
  NAND2_X1 U12251 ( .A1(n9629), .A2(n9624), .ZN(n9627) );
  NAND2_X1 U12252 ( .A1(n9628), .A2(n9625), .ZN(n9626) );
  MUX2_X1 U12253 ( .A(n9627), .B(n9626), .S(n9961), .Z(n9631) );
  MUX2_X1 U12254 ( .A(n9629), .B(n9628), .S(n9855), .Z(n9630) );
  OR2_X1 U12255 ( .A1(n9633), .A2(n7933), .ZN(n13544) );
  NAND2_X1 U12256 ( .A1(n9633), .A2(n9855), .ZN(n9634) );
  NAND2_X1 U12257 ( .A1(n13530), .A2(n9634), .ZN(n9635) );
  AOI22_X1 U12258 ( .A1(n9640), .A2(n9637), .B1(n9961), .B2(n13511), .ZN(n9642) );
  NAND2_X1 U12259 ( .A1(n9638), .A2(n9643), .ZN(n13515) );
  AOI21_X1 U12260 ( .B1(n9645), .B2(n9643), .A(n9855), .ZN(n9644) );
  AOI21_X1 U12261 ( .B1(n9647), .B2(n9961), .A(n9646), .ZN(n9653) );
  INV_X1 U12262 ( .A(n9648), .ZN(n9651) );
  INV_X1 U12263 ( .A(n9649), .ZN(n9650) );
  AOI211_X1 U12264 ( .C1(n9651), .C2(n9655), .A(n9855), .B(n9650), .ZN(n9654)
         );
  INV_X1 U12265 ( .A(n9654), .ZN(n9657) );
  NAND3_X1 U12266 ( .A1(n9706), .A2(n9855), .A3(n9655), .ZN(n9656) );
  MUX2_X1 U12267 ( .A(n9705), .B(n9706), .S(n9961), .Z(n9658) );
  NAND2_X1 U12268 ( .A1(n13441), .A2(n9658), .ZN(n9662) );
  MUX2_X1 U12269 ( .A(n9660), .B(n9659), .S(n9961), .Z(n9661) );
  MUX2_X1 U12270 ( .A(n9664), .B(n9663), .S(n9855), .Z(n9665) );
  MUX2_X1 U12271 ( .A(n9667), .B(n9666), .S(n9961), .Z(n9668) );
  NAND3_X1 U12272 ( .A1(n9669), .A2(n13407), .A3(n9668), .ZN(n9671) );
  NAND3_X1 U12273 ( .A1(n13580), .A2(n13069), .A3(n9961), .ZN(n9670) );
  AOI21_X1 U12274 ( .B1(n9671), .B2(n9670), .A(n13390), .ZN(n9678) );
  INV_X1 U12275 ( .A(n9672), .ZN(n9676) );
  OAI21_X1 U12276 ( .B1(n9676), .B2(n9674), .A(n9673), .ZN(n9675) );
  MUX2_X1 U12277 ( .A(n9676), .B(n9675), .S(n9855), .Z(n9677) );
  OAI21_X1 U12278 ( .B1(n9678), .B2(n9677), .A(n13370), .ZN(n9682) );
  MUX2_X1 U12279 ( .A(n9680), .B(n9679), .S(n9855), .Z(n9681) );
  INV_X1 U12280 ( .A(n9683), .ZN(n9686) );
  INV_X1 U12281 ( .A(n9684), .ZN(n9685) );
  INV_X1 U12282 ( .A(n9702), .ZN(n9698) );
  AOI21_X1 U12283 ( .B1(n9698), .B2(n9718), .A(n9701), .ZN(n9699) );
  AND2_X1 U12284 ( .A1(n13618), .A2(n13336), .ZN(n9717) );
  AOI21_X2 U12285 ( .B1(n9700), .B2(n9699), .A(n9717), .ZN(n9725) );
  NAND2_X1 U12286 ( .A1(n11251), .A2(n10631), .ZN(n9856) );
  NAND2_X1 U12287 ( .A1(n11251), .A2(n13324), .ZN(n11052) );
  INV_X1 U12288 ( .A(n9701), .ZN(n9721) );
  INV_X1 U12289 ( .A(n13417), .ZN(n13418) );
  NAND2_X1 U12290 ( .A1(n9706), .A2(n9705), .ZN(n13458) );
  INV_X1 U12291 ( .A(n11464), .ZN(n11420) );
  INV_X1 U12292 ( .A(n9775), .ZN(n11373) );
  AND2_X1 U12293 ( .A1(n11055), .A2(n9707), .ZN(n10564) );
  NOR3_X1 U12294 ( .A1(n11056), .A2(n11240), .A3(n11361), .ZN(n9709) );
  NAND4_X1 U12295 ( .A1(n10564), .A2(n9585), .A3(n10800), .A4(n9709), .ZN(
        n9710) );
  NOR4_X1 U12296 ( .A1(n11420), .A2(n11373), .A3(n9710), .A4(n11402), .ZN(
        n9711) );
  NAND4_X1 U12297 ( .A1(n9711), .A2(n11771), .A3(n11843), .A4(n11779), .ZN(
        n9712) );
  NOR4_X1 U12298 ( .A1(n13499), .A2(n13515), .A3(n12103), .A4(n9712), .ZN(
        n9713) );
  NAND4_X1 U12299 ( .A1(n13530), .A2(n7443), .A3(n13485), .A4(n9713), .ZN(
        n9714) );
  NOR4_X1 U12300 ( .A1(n13418), .A2(n13473), .A3(n13458), .A4(n9714), .ZN(
        n9715) );
  NAND4_X1 U12301 ( .A1(n13407), .A2(n13441), .A3(n13431), .A4(n9715), .ZN(
        n9716) );
  INV_X1 U12302 ( .A(n9717), .ZN(n9719) );
  NAND4_X1 U12303 ( .A1(n9721), .A2(n9720), .A3(n9719), .A4(n9718), .ZN(n9722)
         );
  XNOR2_X1 U12304 ( .A(n9722), .B(n13324), .ZN(n9723) );
  NOR2_X1 U12305 ( .A1(n11251), .A2(n10521), .ZN(n10520) );
  NAND2_X1 U12306 ( .A1(n9723), .A2(n10520), .ZN(n9724) );
  INV_X1 U12307 ( .A(n9732), .ZN(n9728) );
  NAND2_X1 U12308 ( .A1(n9728), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9730) );
  OR2_X1 U12309 ( .A1(n10500), .A2(P3_U3151), .ZN(n11312) );
  NAND2_X1 U12310 ( .A1(n9732), .A2(n16100), .ZN(n9809) );
  NAND2_X1 U12311 ( .A1(n9809), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9733) );
  INV_X1 U12312 ( .A(n9735), .ZN(n9738) );
  INV_X1 U12313 ( .A(n11703), .ZN(n9746) );
  NAND2_X1 U12314 ( .A1(n9743), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9740) );
  MUX2_X1 U12315 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9740), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n9741) );
  NAND2_X1 U12316 ( .A1(n9815), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9742) );
  MUX2_X1 U12317 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9742), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9744) );
  NOR2_X1 U12318 ( .A1(n12057), .A2(n11892), .ZN(n9745) );
  INV_X1 U12319 ( .A(n9856), .ZN(n9760) );
  NAND2_X1 U12320 ( .A1(n10535), .A2(n9760), .ZN(n10513) );
  INV_X1 U12321 ( .A(n13716), .ZN(n9995) );
  INV_X1 U12322 ( .A(n13724), .ZN(n13328) );
  NAND2_X1 U12323 ( .A1(n9995), .A2(n13328), .ZN(n9992) );
  NAND2_X1 U12324 ( .A1(n8022), .A2(n9992), .ZN(n9765) );
  INV_X1 U12325 ( .A(n9765), .ZN(n9749) );
  NOR2_X1 U12326 ( .A1(n10513), .A2(n13533), .ZN(n10512) );
  NAND2_X1 U12327 ( .A1(n10512), .A2(n9995), .ZN(n9750) );
  OAI211_X1 U12328 ( .C1(n11110), .C2(n11312), .A(n9750), .B(P3_B_REG_SCAN_IN), 
        .ZN(n9751) );
  NAND2_X1 U12329 ( .A1(n9752), .A2(n9751), .ZN(P3_U3296) );
  INV_X1 U12330 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n9846) );
  NAND2_X1 U12331 ( .A1(n11251), .A2(n11110), .ZN(n9756) );
  NAND2_X1 U12332 ( .A1(n9756), .A2(n13324), .ZN(n9757) );
  NAND2_X1 U12333 ( .A1(n9757), .A2(n11382), .ZN(n9759) );
  NAND2_X1 U12334 ( .A1(n11251), .A2(n11382), .ZN(n9758) );
  NAND2_X1 U12335 ( .A1(n9758), .A2(n9764), .ZN(n9828) );
  NAND2_X1 U12336 ( .A1(n9759), .A2(n9828), .ZN(n10498) );
  NAND2_X1 U12337 ( .A1(n10530), .A2(n9760), .ZN(n9763) );
  AND2_X1 U12338 ( .A1(n10631), .A2(n11110), .ZN(n9761) );
  NAND2_X1 U12339 ( .A1(n9762), .A2(n9761), .ZN(n9827) );
  NAND2_X1 U12340 ( .A1(n10766), .A2(n9764), .ZN(n15771) );
  NAND2_X1 U12341 ( .A1(n13394), .A2(n15771), .ZN(n15755) );
  NAND2_X1 U12342 ( .A1(n13122), .A2(n9766), .ZN(n11048) );
  INV_X1 U12343 ( .A(n9767), .ZN(n10765) );
  OR2_X1 U12344 ( .A1(n13120), .A2(n10765), .ZN(n10803) );
  AND2_X1 U12345 ( .A1(n10802), .A2(n10803), .ZN(n9768) );
  NAND2_X1 U12346 ( .A1(n10804), .A2(n9768), .ZN(n10801) );
  INV_X1 U12347 ( .A(n10810), .ZN(n10599) );
  NAND2_X1 U12348 ( .A1(n11241), .A2(n10599), .ZN(n9769) );
  NAND2_X1 U12349 ( .A1(n10801), .A2(n9769), .ZN(n11239) );
  NAND2_X1 U12350 ( .A1(n11239), .A2(n11240), .ZN(n9771) );
  INV_X1 U12351 ( .A(n11236), .ZN(n10999) );
  NAND2_X1 U12352 ( .A1(n13119), .A2(n10999), .ZN(n9770) );
  NAND2_X1 U12353 ( .A1(n9771), .A2(n9770), .ZN(n11363) );
  INV_X1 U12354 ( .A(n11411), .ZN(n9772) );
  NAND2_X1 U12355 ( .A1(n13117), .A2(n9772), .ZN(n11418) );
  NAND2_X1 U12356 ( .A1(n11361), .A2(n11418), .ZN(n9774) );
  OR2_X1 U12357 ( .A1(n13118), .A2(n11269), .ZN(n11403) );
  NAND2_X1 U12358 ( .A1(n11402), .A2(n11403), .ZN(n11405) );
  AOI21_X1 U12359 ( .B1(n11418), .B2(n11405), .A(n11464), .ZN(n9773) );
  INV_X1 U12360 ( .A(n11427), .ZN(n11472) );
  NAND2_X1 U12361 ( .A1(n11720), .A2(n9776), .ZN(n9777) );
  INV_X1 U12362 ( .A(n13113), .ZN(n11604) );
  OR2_X1 U12363 ( .A1(n12053), .A2(n11604), .ZN(n9781) );
  NAND2_X1 U12364 ( .A1(n9782), .A2(n9781), .ZN(n11778) );
  NAND2_X1 U12365 ( .A1(n11778), .A2(n11782), .ZN(n9784) );
  INV_X1 U12366 ( .A(n13112), .ZN(n11949) );
  OR2_X1 U12367 ( .A1(n12003), .A2(n11949), .ZN(n9783) );
  NAND2_X1 U12368 ( .A1(n9784), .A2(n9783), .ZN(n12105) );
  NAND2_X1 U12369 ( .A1(n12113), .A2(n13550), .ZN(n9785) );
  NOR2_X1 U12370 ( .A1(n13555), .A2(n13534), .ZN(n9788) );
  NAND2_X1 U12371 ( .A1(n13555), .A2(n13534), .ZN(n9787) );
  INV_X1 U12372 ( .A(n13548), .ZN(n13100) );
  OR2_X1 U12373 ( .A1(n13689), .A2(n13100), .ZN(n13516) );
  NAND2_X1 U12374 ( .A1(n13685), .A2(n13111), .ZN(n9789) );
  AND2_X1 U12375 ( .A1(n13679), .A2(n13519), .ZN(n13488) );
  INV_X1 U12376 ( .A(n13504), .ZN(n13110) );
  AND2_X1 U12377 ( .A1(n13672), .A2(n13110), .ZN(n9790) );
  AOI21_X1 U12378 ( .B1(n13487), .B2(n13488), .A(n9790), .ZN(n13471) );
  NAND2_X1 U12379 ( .A1(n13487), .A2(n13499), .ZN(n13472) );
  NAND3_X1 U12380 ( .A1(n13471), .A2(n13473), .A3(n13472), .ZN(n9792) );
  INV_X1 U12381 ( .A(n13490), .ZN(n13109) );
  OR2_X1 U12382 ( .A1(n13597), .A2(n13109), .ZN(n9791) );
  AND2_X1 U12383 ( .A1(n9792), .A2(n9791), .ZN(n9793) );
  OR2_X1 U12384 ( .A1(n13593), .A2(n13476), .ZN(n9794) );
  NAND2_X1 U12385 ( .A1(n13457), .A2(n9794), .ZN(n13444) );
  NAND2_X1 U12386 ( .A1(n13444), .A2(n13445), .ZN(n13443) );
  NAND2_X1 U12387 ( .A1(n13590), .A2(n13107), .ZN(n9795) );
  INV_X1 U12388 ( .A(n13446), .ZN(n13420) );
  OR2_X1 U12389 ( .A1(n13434), .A2(n13420), .ZN(n9796) );
  INV_X1 U12390 ( .A(n13649), .ZN(n9797) );
  NAND2_X1 U12391 ( .A1(n13580), .A2(n13421), .ZN(n13387) );
  INV_X1 U12392 ( .A(n13387), .ZN(n9799) );
  AND2_X1 U12393 ( .A1(n13396), .A2(n13374), .ZN(n9798) );
  NOR2_X1 U12394 ( .A1(n9799), .A2(n9798), .ZN(n9800) );
  OR2_X1 U12395 ( .A1(n13396), .A2(n13374), .ZN(n9801) );
  INV_X1 U12396 ( .A(n13629), .ZN(n9802) );
  NAND2_X1 U12397 ( .A1(n13324), .A2(n11110), .ZN(n9849) );
  NAND2_X1 U12398 ( .A1(n9803), .A2(n13549), .ZN(n9807) );
  INV_X1 U12399 ( .A(n9809), .ZN(n9808) );
  NAND3_X1 U12400 ( .A1(n9808), .A2(P3_B_REG_SCAN_IN), .A3(n9815), .ZN(n9820)
         );
  INV_X1 U12401 ( .A(P3_B_REG_SCAN_IN), .ZN(n9864) );
  NAND4_X1 U12402 ( .A1(n9809), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_IR_REG_24__SCAN_IN), .A4(n9864), .ZN(n9819) );
  XNOR2_X1 U12403 ( .A(n9811), .B(P3_IR_REG_24__SCAN_IN), .ZN(n9810) );
  NAND3_X1 U12404 ( .A1(n9815), .A2(P3_B_REG_SCAN_IN), .A3(n9810), .ZN(n9814)
         );
  NAND3_X1 U12405 ( .A1(n9812), .A2(n9864), .A3(n9811), .ZN(n9813) );
  OAI211_X1 U12406 ( .C1(n9815), .C2(P3_B_REG_SCAN_IN), .A(n9814), .B(n9813), 
        .ZN(n9816) );
  INV_X1 U12407 ( .A(n9816), .ZN(n9817) );
  NAND3_X1 U12408 ( .A1(n9820), .A2(n9819), .A3(n9818), .ZN(n9822) );
  NAND2_X1 U12409 ( .A1(n11703), .A2(n12057), .ZN(n9823) );
  NAND2_X1 U12410 ( .A1(n12057), .A2(n11892), .ZN(n9825) );
  NAND2_X1 U12411 ( .A1(n13703), .A2(n13701), .ZN(n9847) );
  INV_X1 U12412 ( .A(n13701), .ZN(n9830) );
  NAND2_X1 U12413 ( .A1(n9824), .A2(n9830), .ZN(n9852) );
  NAND2_X1 U12414 ( .A1(n9827), .A2(n9855), .ZN(n9882) );
  NAND2_X1 U12415 ( .A1(n9856), .A2(n9961), .ZN(n10499) );
  NAND2_X1 U12416 ( .A1(n9882), .A2(n10499), .ZN(n9881) );
  NAND2_X1 U12417 ( .A1(n9881), .A2(n13701), .ZN(n9844) );
  NAND3_X1 U12418 ( .A1(n9828), .A2(n9849), .A3(n9856), .ZN(n9829) );
  NAND2_X1 U12419 ( .A1(n9829), .A2(n9855), .ZN(n9831) );
  NAND2_X1 U12420 ( .A1(n9831), .A2(n9830), .ZN(n9843) );
  NOR2_X1 U12421 ( .A1(P3_D_REG_5__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .ZN(
        n9835) );
  NOR4_X1 U12422 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9834) );
  NOR4_X1 U12423 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_29__SCAN_IN), .ZN(n9833) );
  NOR4_X1 U12424 ( .A1(P3_D_REG_10__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9832) );
  NAND4_X1 U12425 ( .A1(n9835), .A2(n9834), .A3(n9833), .A4(n9832), .ZN(n9841)
         );
  NOR4_X1 U12426 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n9839) );
  NOR4_X1 U12427 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n9838) );
  NOR4_X1 U12428 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9837) );
  NOR4_X1 U12429 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n9836) );
  NAND4_X1 U12430 ( .A1(n9839), .A2(n9838), .A3(n9837), .A4(n9836), .ZN(n9840)
         );
  NOR2_X1 U12431 ( .A1(n9841), .A2(n9840), .ZN(n9842) );
  INV_X1 U12432 ( .A(n9847), .ZN(n9848) );
  INV_X1 U12433 ( .A(n9849), .ZN(n9850) );
  NAND2_X1 U12434 ( .A1(n10520), .A2(n9850), .ZN(n10531) );
  INV_X1 U12435 ( .A(n10498), .ZN(n9853) );
  INV_X1 U12436 ( .A(n9884), .ZN(n9851) );
  OAI22_X1 U12437 ( .A1(n10534), .A2(n10531), .B1(n9853), .B2(n10532), .ZN(
        n9854) );
  NAND2_X1 U12438 ( .A1(n9854), .A2(n10535), .ZN(n9860) );
  INV_X1 U12439 ( .A(n10534), .ZN(n9858) );
  NOR2_X1 U12440 ( .A1(n9856), .A2(n9855), .ZN(n9857) );
  AND2_X1 U12441 ( .A1(n10535), .A2(n9857), .ZN(n10507) );
  NAND2_X1 U12442 ( .A1(n9858), .A2(n10507), .ZN(n9859) );
  XNOR2_X1 U12443 ( .A(n9863), .B(n9870), .ZN(n9868) );
  OAI21_X1 U12444 ( .B1(n9864), .B2(n13716), .A(n13547), .ZN(n13335) );
  OAI21_X1 U12445 ( .B1(n9868), .B2(n13502), .A(n9867), .ZN(n9889) );
  MUX2_X1 U12446 ( .A(P3_REG1_REG_29__SCAN_IN), .B(n9889), .S(n15804), .Z(
        n9869) );
  INV_X1 U12447 ( .A(n9869), .ZN(n9874) );
  XNOR2_X1 U12448 ( .A(n9871), .B(n9870), .ZN(n9891) );
  INV_X1 U12449 ( .A(n9894), .ZN(n9877) );
  OAI22_X1 U12450 ( .A1(n9891), .A2(n13617), .B1(n9877), .B2(n13610), .ZN(
        n9872) );
  INV_X1 U12451 ( .A(n9872), .ZN(n9873) );
  NAND2_X1 U12452 ( .A1(n9874), .A2(n9873), .ZN(P3_U3488) );
  MUX2_X1 U12453 ( .A(P3_REG0_REG_29__SCAN_IN), .B(n9889), .S(n15786), .Z(
        n9875) );
  INV_X1 U12454 ( .A(n9875), .ZN(n9880) );
  INV_X1 U12455 ( .A(n15755), .ZN(n9876) );
  OAI22_X1 U12456 ( .A1(n9891), .A2(n13699), .B1(n9877), .B2(n13688), .ZN(
        n9878) );
  INV_X1 U12457 ( .A(n9878), .ZN(n9879) );
  NAND2_X1 U12458 ( .A1(n9880), .A2(n9879), .ZN(P3_U3456) );
  INV_X1 U12459 ( .A(n9881), .ZN(n9887) );
  NAND2_X1 U12460 ( .A1(n13701), .A2(n9882), .ZN(n9883) );
  AND3_X1 U12461 ( .A1(n10535), .A2(n9884), .A3(n9883), .ZN(n9885) );
  NOR2_X1 U12462 ( .A1(n11052), .A2(n15770), .ZN(n9888) );
  NAND2_X2 U12463 ( .A1(n9892), .A2(n13479), .ZN(n13553) );
  NAND2_X1 U12464 ( .A1(n9889), .A2(n13553), .ZN(n9898) );
  NAND2_X1 U12465 ( .A1(n10766), .A2(n10521), .ZN(n10759) );
  NAND2_X1 U12466 ( .A1(n13394), .A2(n10759), .ZN(n9890) );
  NOR2_X1 U12467 ( .A1(n9892), .A2(n10766), .ZN(n11429) );
  NOR2_X1 U12468 ( .A1(n9893), .A2(n13479), .ZN(n13337) );
  AOI21_X1 U12469 ( .B1(n9894), .B2(n13558), .A(n13337), .ZN(n9896) );
  INV_X1 U12470 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n9895) );
  NAND3_X1 U12471 ( .A1(n9898), .A2(n9897), .A3(n8011), .ZN(P3_U3204) );
  INV_X1 U12472 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9921) );
  XNOR2_X1 U12473 ( .A(n9902), .B(n9910), .ZN(n14099) );
  NAND3_X1 U12474 ( .A1(n8753), .A2(n7165), .A3(n8030), .ZN(n9914) );
  NAND3_X1 U12475 ( .A1(n9906), .A2(n9910), .A3(n9907), .ZN(n9913) );
  INV_X1 U12476 ( .A(n9907), .ZN(n9909) );
  OAI21_X1 U12477 ( .B1(n9909), .B2(n8030), .A(n9910), .ZN(n9908) );
  OAI21_X1 U12478 ( .B1(n9910), .B2(n9909), .A(n9908), .ZN(n9911) );
  NAND3_X1 U12479 ( .A1(n9914), .A2(n9913), .A3(n9912), .ZN(n9920) );
  NAND2_X1 U12480 ( .A1(n13928), .A2(n9915), .ZN(n9916) );
  INV_X1 U12481 ( .A(n9918), .ZN(n9919) );
  NAND2_X1 U12482 ( .A1(n9920), .A2(n9919), .ZN(n14105) );
  MUX2_X1 U12483 ( .A(n9921), .B(n9927), .S(n15743), .Z(n9923) );
  NAND2_X1 U12484 ( .A1(n9923), .A2(n8017), .ZN(P2_U3496) );
  NOR2_X1 U12485 ( .A1(n15697), .A2(n9924), .ZN(n9926) );
  INV_X1 U12486 ( .A(n9929), .ZN(n9930) );
  INV_X2 U12487 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9931) );
  NOR2_X2 U12488 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n10195) );
  INV_X2 U12489 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10570) );
  INV_X2 U12490 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10310) );
  NAND4_X1 U12491 ( .A1(n10570), .A2(n10310), .A3(n10196), .A4(n10096), .ZN(
        n9936) );
  NAND2_X1 U12492 ( .A1(n10205), .A2(n10208), .ZN(n9938) );
  NAND2_X1 U12493 ( .A1(n9940), .A2(n9943), .ZN(n9949) );
  INV_X1 U12494 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9947) );
  XNOR2_X1 U12495 ( .A(n9948), .B(n9947), .ZN(n11893) );
  NAND2_X1 U12496 ( .A1(n9949), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9950) );
  MUX2_X1 U12497 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9950), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9952) );
  OR3_X4 U12498 ( .A1(n10185), .A2(n11893), .A3(n11786), .ZN(n10376) );
  NOR2_X1 U12499 ( .A1(n10191), .A2(n10376), .ZN(P1_U4016) );
  INV_X1 U12500 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10371) );
  NOR2_X1 U12501 ( .A1(n10371), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11065) );
  NAND2_X1 U12502 ( .A1(n11065), .A2(n9953), .ZN(n9954) );
  OAI21_X1 U12503 ( .B1(n11102), .B2(n11065), .A(n9954), .ZN(n11092) );
  INV_X1 U12504 ( .A(n9954), .ZN(n9955) );
  NAND2_X1 U12505 ( .A1(n9956), .A2(n10739), .ZN(n9957) );
  XNOR2_X1 U12506 ( .A(n10991), .B(P3_REG1_REG_4__SCAN_IN), .ZN(n10985) );
  XNOR2_X1 U12507 ( .A(n10952), .B(n15799), .ZN(n9959) );
  INV_X1 U12508 ( .A(n10948), .ZN(n9965) );
  NAND3_X1 U12509 ( .A1(n10778), .A2(n9959), .A3(n6999), .ZN(n9964) );
  INV_X1 U12510 ( .A(n10535), .ZN(n9960) );
  NAND2_X1 U12511 ( .A1(n9960), .A2(n11312), .ZN(n9998) );
  NAND2_X1 U12512 ( .A1(n9961), .A2(n10500), .ZN(n9962) );
  NAND2_X1 U12513 ( .A1(n9962), .A2(n8022), .ZN(n9997) );
  INV_X1 U12514 ( .A(n9997), .ZN(n9963) );
  AND2_X1 U12515 ( .A1(n9998), .A2(n9963), .ZN(n9996) );
  INV_X1 U12516 ( .A(n13313), .ZN(n13190) );
  AOI21_X1 U12517 ( .B1(n9965), .B2(n9964), .A(n13190), .ZN(n10003) );
  INV_X1 U12518 ( .A(n11102), .ZN(n9968) );
  MUX2_X1 U12519 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n13724), .Z(n9966) );
  INV_X1 U12520 ( .A(n9966), .ZN(n9967) );
  XNOR2_X1 U12521 ( .A(n9966), .B(n11102), .ZN(n11095) );
  MUX2_X1 U12522 ( .A(n10713), .B(n10371), .S(n13724), .Z(n11059) );
  NAND2_X1 U12523 ( .A1(n11059), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11094) );
  NOR2_X1 U12524 ( .A1(n11095), .A2(n11094), .ZN(n11093) );
  MUX2_X1 U12525 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n13724), .Z(n9969) );
  XNOR2_X1 U12526 ( .A(n9969), .B(n10739), .ZN(n10730) );
  INV_X1 U12527 ( .A(n9969), .ZN(n9970) );
  MUX2_X1 U12528 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13724), .Z(n9971) );
  XNOR2_X1 U12529 ( .A(n9971), .B(n10991), .ZN(n10975) );
  MUX2_X1 U12530 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n13724), .Z(n9972) );
  INV_X1 U12531 ( .A(n10779), .ZN(n10115) );
  NAND2_X1 U12532 ( .A1(n9972), .A2(n10115), .ZN(n10774) );
  INV_X1 U12533 ( .A(n9972), .ZN(n9973) );
  NAND2_X1 U12534 ( .A1(n9973), .A2(n10779), .ZN(n10776) );
  MUX2_X1 U12535 ( .A(n16060), .B(n15799), .S(n13724), .Z(n9974) );
  NAND2_X1 U12536 ( .A1(n9974), .A2(n10952), .ZN(n10962) );
  INV_X1 U12537 ( .A(n9974), .ZN(n9975) );
  INV_X1 U12538 ( .A(n10952), .ZN(n10949) );
  NAND2_X1 U12539 ( .A1(n9975), .A2(n10949), .ZN(n9976) );
  NAND2_X1 U12540 ( .A1(n10962), .A2(n9976), .ZN(n9977) );
  INV_X1 U12541 ( .A(n10970), .ZN(n9979) );
  NAND3_X1 U12542 ( .A1(n10772), .A2(n10776), .A3(n9977), .ZN(n9978) );
  AND2_X1 U12543 ( .A1(P3_U3897), .A2(n13716), .ZN(n13332) );
  AOI21_X1 U12544 ( .B1(n9979), .B2(n9978), .A(n13210), .ZN(n10002) );
  NOR2_X1 U12545 ( .A1(n10713), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9981) );
  NAND2_X1 U12546 ( .A1(n9980), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9982) );
  OAI21_X1 U12547 ( .B1(n11102), .B2(n9981), .A(n9982), .ZN(n11086) );
  INV_X1 U12548 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11054) );
  OR2_X1 U12549 ( .A1(n11086), .A2(n11054), .ZN(n11087) );
  NAND2_X1 U12550 ( .A1(n11087), .A2(n9982), .ZN(n10748) );
  INV_X1 U12551 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10770) );
  NAND2_X1 U12552 ( .A1(n10748), .A2(n10749), .ZN(n10747) );
  NAND2_X1 U12553 ( .A1(n10106), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9983) );
  NAND2_X1 U12554 ( .A1(n10747), .A2(n9983), .ZN(n9984) );
  INV_X1 U12555 ( .A(n10739), .ZN(n10063) );
  NAND2_X1 U12556 ( .A1(n9984), .A2(n10063), .ZN(n10978) );
  INV_X1 U12557 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10809) );
  INV_X1 U12558 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n9985) );
  XNOR2_X1 U12559 ( .A(n10991), .B(n9985), .ZN(n10977) );
  NAND2_X1 U12560 ( .A1(n10991), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9986) );
  NAND2_X1 U12561 ( .A1(n10982), .A2(n9986), .ZN(n9987) );
  XNOR2_X1 U12562 ( .A(n10952), .B(P3_REG2_REG_6__SCAN_IN), .ZN(n9989) );
  NAND2_X1 U12563 ( .A1(n9988), .A2(n9989), .ZN(n10954) );
  INV_X1 U12564 ( .A(n9989), .ZN(n9991) );
  NAND3_X1 U12565 ( .A1(n10783), .A2(n9991), .A3(n9990), .ZN(n9994) );
  INV_X1 U12566 ( .A(n9992), .ZN(n9993) );
  AOI21_X1 U12567 ( .B1(n10954), .B2(n9994), .A(n13283), .ZN(n10001) );
  MUX2_X1 U12568 ( .A(n9996), .B(P3_U3897), .S(n9995), .Z(n13323) );
  INV_X1 U12569 ( .A(n13323), .ZN(n13295) );
  AND2_X1 U12570 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n11396) );
  AOI21_X1 U12571 ( .B1(n15751), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11396), .ZN(
        n9999) );
  OAI21_X1 U12572 ( .B1(n13295), .B2(n10949), .A(n9999), .ZN(n10000) );
  OR4_X1 U12573 ( .A1(n10003), .A2(n10002), .A3(n10001), .A4(n10000), .ZN(
        P3_U3188) );
  INV_X1 U12574 ( .A(n10004), .ZN(n10028) );
  OR2_X1 U12575 ( .A1(n10005), .A2(n10028), .ZN(n10006) );
  OAI21_X1 U12576 ( .B1(n10006), .B2(n15701), .A(n10035), .ZN(n10008) );
  NAND2_X1 U12577 ( .A1(n10008), .A2(n10007), .ZN(n10397) );
  MUX2_X1 U12578 ( .A(n13859), .B(P2_U3088), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n10043) );
  NAND2_X4 U12579 ( .A1(n15715), .A2(n11653), .ZN(n13789) );
  INV_X1 U12580 ( .A(n10022), .ZN(n14293) );
  OR2_X1 U12581 ( .A1(n11969), .A2(n14293), .ZN(n10013) );
  NAND2_X1 U12582 ( .A1(n11633), .A2(n15660), .ZN(n10012) );
  INV_X1 U12583 ( .A(n10014), .ZN(n10015) );
  NAND2_X1 U12584 ( .A1(n10016), .A2(n10015), .ZN(n10017) );
  XNOR2_X1 U12585 ( .A(n13789), .B(n11934), .ZN(n10018) );
  NAND2_X1 U12586 ( .A1(n13956), .A2(n12612), .ZN(n10019) );
  XNOR2_X1 U12587 ( .A(n10018), .B(n10019), .ZN(n10410) );
  INV_X1 U12588 ( .A(n10018), .ZN(n10020) );
  NAND2_X1 U12589 ( .A1(n10020), .A2(n10019), .ZN(n10021) );
  XNOR2_X1 U12590 ( .A(n13789), .B(n11717), .ZN(n10023) );
  AND2_X1 U12591 ( .A1(n13955), .A2(n12612), .ZN(n10024) );
  NAND2_X1 U12592 ( .A1(n10023), .A2(n10024), .ZN(n10852) );
  INV_X1 U12593 ( .A(n10023), .ZN(n10026) );
  INV_X1 U12594 ( .A(n10024), .ZN(n10025) );
  NAND2_X1 U12595 ( .A1(n10026), .A2(n10025), .ZN(n10027) );
  NAND2_X1 U12596 ( .A1(n10852), .A2(n10027), .ZN(n10032) );
  NOR2_X1 U12597 ( .A1(n14518), .A2(n10427), .ZN(n10029) );
  INV_X1 U12598 ( .A(n10853), .ZN(n10031) );
  AOI211_X1 U12599 ( .C1(n10033), .C2(n10032), .A(n13925), .B(n10031), .ZN(
        n10042) );
  INV_X1 U12600 ( .A(n10034), .ZN(n11623) );
  NAND2_X1 U12601 ( .A1(n10040), .A2(n11623), .ZN(n10037) );
  AOI22_X1 U12602 ( .A1(n13905), .A2(n13956), .B1(n13954), .B2(n13907), .ZN(
        n11710) );
  INV_X1 U12603 ( .A(n10038), .ZN(n10039) );
  OAI22_X1 U12604 ( .A1(n13912), .A2(n15717), .B1(n11710), .B2(n13855), .ZN(
        n10041) );
  OR3_X1 U12605 ( .A1(n10043), .A2(n10042), .A3(n10041), .ZN(P2_U3190) );
  INV_X1 U12606 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n11063) );
  AOI21_X1 U12607 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n11063), .A(n7196), .ZN(
        n10045) );
  INV_X1 U12608 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10044) );
  NOR2_X1 U12609 ( .A1(n10045), .A2(n10044), .ZN(n16127) );
  AOI21_X1 U12610 ( .B1(n10045), .B2(n10044), .A(n16127), .ZN(SUB_1596_U53) );
  INV_X1 U12611 ( .A(SI_0_), .ZN(n10046) );
  OAI21_X1 U12612 ( .B1(n10885), .B2(n10046), .A(n15964), .ZN(n10047) );
  NAND2_X1 U12613 ( .A1(n10048), .A2(n10047), .ZN(n10351) );
  MUX2_X1 U12614 ( .A(n10351), .B(n6932), .S(P1_STATE_REG_SCAN_IN), .Z(n10049)
         );
  INV_X1 U12615 ( .A(n10049), .ZN(P1_U3355) );
  AND2_X1 U12616 ( .A1(n10052), .A2(P1_U3086), .ZN(n11744) );
  INV_X2 U12617 ( .A(n11744), .ZN(n15379) );
  OAI222_X1 U12618 ( .A1(n10666), .A2(P1_U3086), .B1(n15379), .B2(n10663), 
        .C1(n10051), .C2(n15370), .ZN(P1_U3354) );
  AND2_X1 U12619 ( .A1(n10052), .A2(P2_U3088), .ZN(n14592) );
  INV_X2 U12620 ( .A(n14592), .ZN(n14590) );
  NAND2_X1 U12621 ( .A1(n10885), .A2(P2_U3088), .ZN(n14594) );
  OAI222_X1 U12622 ( .A1(n14590), .A2(n10053), .B1(n14594), .B2(n10689), .C1(
        P2_U3088), .C2(n13964), .ZN(P2_U3325) );
  INV_X1 U12623 ( .A(n10886), .ZN(n10055) );
  NAND2_X1 U12624 ( .A1(n10093), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10054) );
  OAI222_X1 U12625 ( .A1(n15370), .A2(n10890), .B1(n15379), .B2(n10055), .C1(
        P1_U3086), .C2(n10887), .ZN(P1_U3352) );
  OAI222_X1 U12626 ( .A1(n14590), .A2(n10056), .B1(n14594), .B2(n10055), .C1(
        P2_U3088), .C2(n15642), .ZN(P2_U3324) );
  NOR2_X1 U12627 ( .A1(n10885), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13709) );
  INV_X2 U12628 ( .A(n13709), .ZN(n13721) );
  INV_X1 U12629 ( .A(n10057), .ZN(n10059) );
  INV_X1 U12630 ( .A(SI_4_), .ZN(n10058) );
  OAI222_X1 U12631 ( .A1(n10991), .A2(P3_U3151), .B1(n13721), .B2(n10059), 
        .C1(n10058), .C2(n13723), .ZN(P3_U3291) );
  INV_X1 U12632 ( .A(n10060), .ZN(n10062) );
  INV_X1 U12633 ( .A(SI_3_), .ZN(n10061) );
  OAI222_X1 U12634 ( .A1(n10063), .A2(P3_U3151), .B1(n13721), .B2(n10062), 
        .C1(n10061), .C2(n13723), .ZN(P3_U3292) );
  INV_X1 U12635 ( .A(n10064), .ZN(n10066) );
  INV_X1 U12636 ( .A(SI_6_), .ZN(n10065) );
  OAI222_X1 U12637 ( .A1(n10949), .A2(P3_U3151), .B1(n13721), .B2(n10066), 
        .C1(n10065), .C2(n13723), .ZN(P3_U3289) );
  INV_X1 U12638 ( .A(n10899), .ZN(n10091) );
  OAI222_X1 U12639 ( .A1(n14590), .A2(n10067), .B1(n14594), .B2(n10091), .C1(
        P2_U3088), .C2(n13977), .ZN(P2_U3323) );
  INV_X1 U12640 ( .A(n11019), .ZN(n10075) );
  INV_X1 U12641 ( .A(n13990), .ZN(n10068) );
  OAI222_X1 U12642 ( .A1(n14590), .A2(n10069), .B1(n14594), .B2(n10075), .C1(
        P2_U3088), .C2(n10068), .ZN(P2_U3322) );
  INV_X1 U12643 ( .A(n10088), .ZN(n10071) );
  NAND2_X1 U12644 ( .A1(n10071), .A2(n10070), .ZN(n10073) );
  NAND2_X1 U12645 ( .A1(n10073), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10072) );
  MUX2_X1 U12646 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10072), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n10074) );
  AND2_X1 U12647 ( .A1(n10074), .A2(n10543), .ZN(n11020) );
  OAI222_X1 U12648 ( .A1(n15370), .A2(n10076), .B1(n15379), .B2(n10075), .C1(
        P1_U3086), .C2(n7500), .ZN(P1_U3350) );
  INV_X1 U12649 ( .A(SI_8_), .ZN(n10077) );
  OAI222_X1 U12650 ( .A1(n13721), .A2(n10078), .B1(n13723), .B2(n10077), .C1(
        n11568), .C2(P3_U3151), .ZN(P3_U3287) );
  OAI222_X1 U12651 ( .A1(n13721), .A2(n10080), .B1(n13723), .B2(n10079), .C1(
        n10965), .C2(P3_U3151), .ZN(P3_U3288) );
  AND2_X1 U12652 ( .A1(n10116), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12653 ( .A1(n10116), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12654 ( .A1(n10116), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12655 ( .A1(n10116), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12656 ( .A1(n10116), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12657 ( .A1(n10116), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12658 ( .A1(n10116), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12659 ( .A1(n10116), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12660 ( .A1(n10116), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12661 ( .A1(n10116), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12662 ( .A1(n10116), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12663 ( .A1(n10116), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12664 ( .A1(n10116), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12665 ( .A1(n10116), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12666 ( .A1(n10116), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12667 ( .A1(n10116), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12668 ( .A1(n10116), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12669 ( .A1(n10116), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12670 ( .A1(n10116), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12671 ( .A1(n10116), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12672 ( .A1(n10116), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12673 ( .A1(n10116), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12674 ( .A1(n10116), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12675 ( .A1(n10116), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  INV_X1 U12676 ( .A(n11189), .ZN(n10086) );
  INV_X1 U12677 ( .A(n14004), .ZN(n10083) );
  OAI222_X1 U12678 ( .A1(n14590), .A2(n10084), .B1(n14594), .B2(n10086), .C1(
        P2_U3088), .C2(n10083), .ZN(P2_U3321) );
  INV_X1 U12679 ( .A(n15370), .ZN(n15367) );
  NAND2_X1 U12680 ( .A1(n10543), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10085) );
  XNOR2_X1 U12681 ( .A(n10085), .B(P1_IR_REG_6__SCAN_IN), .ZN(n11190) );
  INV_X1 U12682 ( .A(n11190), .ZN(n10288) );
  OAI222_X1 U12683 ( .A1(n15370), .A2(n10087), .B1(n15379), .B2(n10086), .C1(
        P1_U3086), .C2(n10288), .ZN(P1_U3349) );
  INV_X1 U12684 ( .A(n10898), .ZN(n10090) );
  OAI222_X1 U12685 ( .A1(n15370), .A2(n16025), .B1(n15379), .B2(n10091), .C1(
        P1_U3086), .C2(n10090), .ZN(P1_U3351) );
  NAND2_X1 U12686 ( .A1(n10094), .A2(n10093), .ZN(n10694) );
  OAI222_X1 U12687 ( .A1(n15370), .A2(n10095), .B1(n15379), .B2(n10689), .C1(
        P1_U3086), .C2(n10694), .ZN(P1_U3353) );
  INV_X1 U12688 ( .A(n11439), .ZN(n10123) );
  INV_X1 U12689 ( .A(n10543), .ZN(n10097) );
  NAND2_X1 U12690 ( .A1(n10097), .A2(n10096), .ZN(n10118) );
  NAND2_X1 U12691 ( .A1(n10118), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10098) );
  XNOR2_X1 U12692 ( .A(n10098), .B(P1_IR_REG_7__SCAN_IN), .ZN(n11440) );
  INV_X1 U12693 ( .A(n11440), .ZN(n10099) );
  OAI222_X1 U12694 ( .A1(n15370), .A2(n10100), .B1(n15379), .B2(n10123), .C1(
        P1_U3086), .C2(n10099), .ZN(P1_U3348) );
  OAI222_X1 U12695 ( .A1(n11102), .A2(P3_U3151), .B1(n13721), .B2(n10102), 
        .C1(n10101), .C2(n13723), .ZN(P3_U3294) );
  INV_X1 U12696 ( .A(n10103), .ZN(n10105) );
  INV_X1 U12697 ( .A(SI_2_), .ZN(n10104) );
  OAI222_X1 U12698 ( .A1(n10106), .A2(P3_U3151), .B1(n13721), .B2(n10105), 
        .C1(n10104), .C2(n13723), .ZN(P3_U3293) );
  OAI222_X1 U12699 ( .A1(n13721), .A2(n10108), .B1(n13723), .B2(n10107), .C1(
        n11569), .C2(P3_U3151), .ZN(P3_U3286) );
  INV_X1 U12700 ( .A(n14594), .ZN(n11740) );
  INV_X1 U12701 ( .A(n11740), .ZN(n11897) );
  NOR2_X1 U12702 ( .A1(n10433), .A2(P2_U3088), .ZN(n15632) );
  AOI21_X1 U12703 ( .B1(n14592), .B2(P1_DATAO_REG_1__SCAN_IN), .A(n15632), 
        .ZN(n10109) );
  OAI21_X1 U12704 ( .B1(n10663), .B2(n11897), .A(n10109), .ZN(P2_U3326) );
  INV_X1 U12705 ( .A(SI_10_), .ZN(n10110) );
  OAI222_X1 U12706 ( .A1(n13721), .A2(n10111), .B1(n13723), .B2(n10110), .C1(
        n13124), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X1 U12707 ( .A(n10112), .ZN(n10114) );
  INV_X1 U12708 ( .A(SI_5_), .ZN(n10113) );
  OAI222_X1 U12709 ( .A1(n10115), .A2(P3_U3151), .B1(n13721), .B2(n10114), 
        .C1(n10113), .C2(n13723), .ZN(P3_U3290) );
  INV_X1 U12710 ( .A(n10116), .ZN(n10117) );
  INV_X1 U12711 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n16077) );
  NOR2_X1 U12712 ( .A1(n10117), .A2(n16077), .ZN(P3_U3260) );
  INV_X1 U12713 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n15954) );
  NOR2_X1 U12714 ( .A1(n10117), .A2(n15954), .ZN(P3_U3243) );
  INV_X1 U12715 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n15955) );
  NOR2_X1 U12716 ( .A1(n10117), .A2(n15955), .ZN(P3_U3255) );
  INV_X1 U12717 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n15907) );
  NOR2_X1 U12718 ( .A1(n10117), .A2(n15907), .ZN(P3_U3241) );
  INV_X1 U12719 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n16047) );
  NOR2_X1 U12720 ( .A1(n10117), .A2(n16047), .ZN(P3_U3240) );
  INV_X1 U12721 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n16043) );
  NOR2_X1 U12722 ( .A1(n10117), .A2(n16043), .ZN(P3_U3251) );
  INV_X1 U12723 ( .A(n11510), .ZN(n10120) );
  NAND2_X1 U12724 ( .A1(n10198), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10170) );
  XNOR2_X1 U12725 ( .A(n10170), .B(P1_IR_REG_8__SCAN_IN), .ZN(n11511) );
  INV_X1 U12726 ( .A(n11511), .ZN(n10653) );
  OAI222_X1 U12727 ( .A1(n15370), .A2(n10119), .B1(n15379), .B2(n10120), .C1(
        P1_U3086), .C2(n10653), .ZN(P1_U3347) );
  OAI222_X1 U12728 ( .A1(n14590), .A2(n10121), .B1(n14594), .B2(n10120), .C1(
        P2_U3088), .C2(n14033), .ZN(P2_U3319) );
  INV_X1 U12729 ( .A(n14020), .ZN(n10122) );
  OAI222_X1 U12730 ( .A1(n14590), .A2(n10124), .B1(n11897), .B2(n10123), .C1(
        P2_U3088), .C2(n10122), .ZN(P2_U3320) );
  NAND2_X1 U12731 ( .A1(n10147), .A2(n10125), .ZN(n10143) );
  NAND2_X1 U12732 ( .A1(n10126), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n10129) );
  NAND2_X1 U12733 ( .A1(n10127), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n10128) );
  NAND2_X1 U12734 ( .A1(n10143), .A2(n10142), .ZN(n10141) );
  NAND2_X1 U12735 ( .A1(n10141), .A2(n10129), .ZN(n10130) );
  OAI21_X1 U12736 ( .B1(n10132), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n10133), .ZN(
        n10135) );
  NAND2_X1 U12737 ( .A1(n10137), .A2(n10133), .ZN(n10134) );
  NAND2_X1 U12738 ( .A1(n10134), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n10605) );
  NAND2_X1 U12739 ( .A1(n10135), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n10136) );
  INV_X1 U12740 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10138) );
  NAND2_X1 U12741 ( .A1(n10140), .A2(n10139), .ZN(n10154) );
  OAI21_X1 U12742 ( .B1(n10143), .B2(n10142), .A(n10141), .ZN(n10152) );
  NAND2_X1 U12743 ( .A1(n10145), .A2(n10144), .ZN(n10146) );
  NAND2_X1 U12744 ( .A1(n10147), .A2(n10146), .ZN(n10148) );
  NAND2_X1 U12745 ( .A1(n10148), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n10150) );
  XOR2_X1 U12746 ( .A(n10148), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n16126) );
  NAND2_X1 U12747 ( .A1(n16127), .A2(n16126), .ZN(n10149) );
  NAND2_X1 U12748 ( .A1(n10150), .A2(n10149), .ZN(n10151) );
  NAND2_X1 U12749 ( .A1(n10152), .A2(n10151), .ZN(n15467) );
  INV_X1 U12750 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15469) );
  NAND2_X1 U12751 ( .A1(n15467), .A2(n15469), .ZN(n10153) );
  AND2_X1 U12752 ( .A1(n15468), .A2(n10153), .ZN(n10155) );
  NAND2_X1 U12753 ( .A1(n10154), .A2(n10155), .ZN(n16122) );
  INV_X1 U12754 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n16124) );
  NAND2_X1 U12755 ( .A1(n16122), .A2(n16124), .ZN(n10158) );
  INV_X1 U12756 ( .A(n10154), .ZN(n10157) );
  INV_X1 U12757 ( .A(n10155), .ZN(n10156) );
  NAND2_X1 U12758 ( .A1(n10157), .A2(n10156), .ZN(n16123) );
  AND2_X1 U12759 ( .A1(n10158), .A2(n16123), .ZN(n15383) );
  INV_X1 U12760 ( .A(n10162), .ZN(n10163) );
  INV_X1 U12761 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n13984) );
  OAI21_X1 U12762 ( .B1(n6760), .B2(n13984), .A(n10604), .ZN(SUB_1596_U58) );
  OAI222_X1 U12763 ( .A1(n13721), .A2(n10167), .B1(n13723), .B2(n10166), .C1(
        n13153), .C2(P3_U3151), .ZN(P3_U3284) );
  INV_X1 U12764 ( .A(n11515), .ZN(n10173) );
  OAI222_X1 U12765 ( .A1(n14590), .A2(n10168), .B1(n14594), .B2(n10173), .C1(
        P2_U3088), .C2(n10484), .ZN(P2_U3318) );
  INV_X1 U12766 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n10169) );
  NAND2_X1 U12767 ( .A1(n10170), .A2(n10169), .ZN(n10171) );
  NAND2_X1 U12768 ( .A1(n10171), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10176) );
  XNOR2_X1 U12769 ( .A(n10176), .B(P1_IR_REG_9__SCAN_IN), .ZN(n14842) );
  INV_X1 U12770 ( .A(n14842), .ZN(n10172) );
  OAI222_X1 U12771 ( .A1(n15370), .A2(n10174), .B1(n15379), .B2(n10173), .C1(
        P1_U3086), .C2(n10172), .ZN(P1_U3346) );
  INV_X1 U12772 ( .A(n11493), .ZN(n10181) );
  INV_X1 U12773 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10175) );
  NAND2_X1 U12774 ( .A1(n10176), .A2(n10175), .ZN(n10177) );
  NAND2_X1 U12775 ( .A1(n10177), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10178) );
  XNOR2_X1 U12776 ( .A(n10178), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11494) );
  INV_X1 U12777 ( .A(n11494), .ZN(n10822) );
  OAI222_X1 U12778 ( .A1(n15370), .A2(n10179), .B1(n15379), .B2(n10181), .C1(
        P1_U3086), .C2(n10822), .ZN(P1_U3345) );
  INV_X1 U12779 ( .A(n10724), .ZN(n10180) );
  OAI222_X1 U12780 ( .A1(n14590), .A2(n16097), .B1(n14594), .B2(n10181), .C1(
        P2_U3088), .C2(n10180), .ZN(P2_U3317) );
  INV_X1 U12781 ( .A(n10182), .ZN(n10184) );
  INV_X1 U12782 ( .A(n13171), .ZN(n13183) );
  OAI222_X1 U12783 ( .A1(n13721), .A2(n10184), .B1(n13723), .B2(n10183), .C1(
        n13183), .C2(P3_U3151), .ZN(P3_U3283) );
  NOR2_X1 U12784 ( .A1(n11786), .A2(P1_B_REG_SCAN_IN), .ZN(n10186) );
  INV_X1 U12785 ( .A(n10349), .ZN(n10189) );
  INV_X1 U12786 ( .A(n10191), .ZN(n10188) );
  NAND2_X1 U12787 ( .A1(n12588), .A2(n11786), .ZN(n10348) );
  OAI22_X1 U12788 ( .A1(n15526), .A2(P1_D_REG_0__SCAN_IN), .B1(n10191), .B2(
        n10348), .ZN(n10190) );
  INV_X1 U12789 ( .A(n10190), .ZN(P1_U3445) );
  NAND2_X1 U12790 ( .A1(n12588), .A2(n11893), .ZN(n10336) );
  OAI22_X1 U12791 ( .A1(n15526), .A2(P1_D_REG_1__SCAN_IN), .B1(n10191), .B2(
        n10336), .ZN(n10192) );
  INV_X1 U12792 ( .A(n10192), .ZN(P1_U3446) );
  INV_X1 U12793 ( .A(n12007), .ZN(n10200) );
  INV_X1 U12794 ( .A(n14052), .ZN(n10193) );
  OAI222_X1 U12795 ( .A1(n14590), .A2(n10194), .B1(n14594), .B2(n10200), .C1(
        P2_U3088), .C2(n10193), .ZN(P2_U3316) );
  NAND2_X1 U12796 ( .A1(n10195), .A2(n10196), .ZN(n10197) );
  NAND2_X1 U12797 ( .A1(n10572), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10199) );
  XNOR2_X1 U12798 ( .A(n10199), .B(P1_IR_REG_11__SCAN_IN), .ZN(n12008) );
  INV_X1 U12799 ( .A(n12008), .ZN(n11114) );
  OAI222_X1 U12800 ( .A1(n15370), .A2(n10201), .B1(n15379), .B2(n10200), .C1(
        P1_U3086), .C2(n11114), .ZN(P1_U3344) );
  AND2_X1 U12801 ( .A1(n10333), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12911) );
  NAND2_X1 U12802 ( .A1(n11131), .A2(n12915), .ZN(n10231) );
  NAND2_X1 U12803 ( .A1(n10205), .A2(n10204), .ZN(n10206) );
  INV_X1 U12804 ( .A(n10206), .ZN(n10207) );
  AND2_X1 U12805 ( .A1(n10207), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n10210) );
  XNOR2_X1 U12806 ( .A(n10208), .B(P1_IR_REG_31__SCAN_IN), .ZN(n10209) );
  NOR2_X1 U12807 ( .A1(n10210), .A2(n10209), .ZN(n10211) );
  AOI21_X1 U12808 ( .B1(n9937), .B2(n10212), .A(n10211), .ZN(n10215) );
  AND2_X1 U12809 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .ZN(n10213) );
  NAND2_X1 U12810 ( .A1(n10330), .A2(n10213), .ZN(n10214) );
  INV_X1 U12811 ( .A(n12673), .ZN(n15381) );
  NAND2_X1 U12812 ( .A1(n10354), .A2(n15381), .ZN(n12859) );
  OR2_X1 U12813 ( .A1(n12859), .A2(n10333), .ZN(n10227) );
  INV_X1 U12814 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10221) );
  AND2_X1 U12815 ( .A1(n12328), .A2(n10227), .ZN(n10230) );
  INV_X1 U12816 ( .A(n10230), .ZN(n10228) );
  NOR2_X1 U12817 ( .A1(n15475), .A2(n14791), .ZN(P1_U3085) );
  INV_X1 U12818 ( .A(n12070), .ZN(n10287) );
  XNOR2_X1 U12819 ( .A(n10311), .B(P1_IR_REG_12__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U12820 ( .A1(n12071), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n15367), .ZN(n10229) );
  OAI21_X1 U12821 ( .B1(n10287), .B2(n15379), .A(n10229), .ZN(P1_U3343) );
  NAND2_X1 U12822 ( .A1(n10231), .A2(n10230), .ZN(n15478) );
  INV_X1 U12823 ( .A(n15817), .ZN(n15486) );
  XOR2_X1 U12824 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n11020), .Z(n10235) );
  INV_X1 U12825 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n15996) );
  AND2_X1 U12826 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14801) );
  INV_X1 U12827 ( .A(n10666), .ZN(n14796) );
  NAND2_X1 U12828 ( .A1(n14796), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10232) );
  NAND2_X1 U12829 ( .A1(n14800), .A2(n10232), .ZN(n14809) );
  INV_X1 U12830 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n15610) );
  MUX2_X1 U12831 ( .A(n15610), .B(P1_REG1_REG_2__SCAN_IN), .S(n10694), .Z(
        n14810) );
  NAND2_X1 U12832 ( .A1(n14809), .A2(n14810), .ZN(n14808) );
  INV_X1 U12833 ( .A(n10694), .ZN(n14814) );
  NAND2_X1 U12834 ( .A1(n14814), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n10233) );
  NAND2_X1 U12835 ( .A1(n14808), .A2(n10233), .ZN(n14820) );
  INV_X1 U12836 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n16062) );
  MUX2_X1 U12837 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n16062), .S(n14828), .Z(
        n14821) );
  NAND2_X1 U12838 ( .A1(n14820), .A2(n14821), .ZN(n14819) );
  NAND2_X1 U12839 ( .A1(n14828), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10234) );
  NAND2_X1 U12840 ( .A1(n14819), .A2(n10234), .ZN(n10469) );
  INV_X1 U12841 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n15613) );
  MUX2_X1 U12842 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n15613), .S(n10898), .Z(
        n10470) );
  OAI21_X1 U12843 ( .B1(n10235), .B2(n6568), .A(n10267), .ZN(n10249) );
  INV_X1 U12844 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n11140) );
  AND2_X1 U12845 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10236) );
  NAND2_X1 U12846 ( .A1(n14799), .A2(n10236), .ZN(n14798) );
  NAND2_X1 U12847 ( .A1(n14796), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10237) );
  NAND2_X1 U12848 ( .A1(n14798), .A2(n10237), .ZN(n14806) );
  INV_X1 U12849 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10238) );
  MUX2_X1 U12850 ( .A(n10238), .B(P1_REG2_REG_2__SCAN_IN), .S(n10694), .Z(
        n14807) );
  NAND2_X1 U12851 ( .A1(n14806), .A2(n14807), .ZN(n14825) );
  NAND2_X1 U12852 ( .A1(n14814), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14824) );
  NAND2_X1 U12853 ( .A1(n14825), .A2(n14824), .ZN(n10240) );
  INV_X1 U12854 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n14822) );
  MUX2_X1 U12855 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n14822), .S(n14828), .Z(
        n10239) );
  NAND2_X1 U12856 ( .A1(n10240), .A2(n10239), .ZN(n14827) );
  NAND2_X1 U12857 ( .A1(n14828), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n10241) );
  NAND2_X1 U12858 ( .A1(n14827), .A2(n10241), .ZN(n10468) );
  INV_X1 U12859 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10242) );
  MUX2_X1 U12860 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10242), .S(n10898), .Z(
        n10467) );
  AOI22_X1 U12861 ( .A1(n10468), .A2(n10467), .B1(n10898), .B2(
        P1_REG2_REG_4__SCAN_IN), .ZN(n10247) );
  INV_X1 U12862 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10243) );
  MUX2_X1 U12863 ( .A(n10243), .B(P1_REG2_REG_5__SCAN_IN), .S(n11020), .Z(
        n10246) );
  INV_X1 U12864 ( .A(n10273), .ZN(n10245) );
  NAND2_X1 U12865 ( .A1(n10692), .A2(n12912), .ZN(n10244) );
  AOI211_X1 U12866 ( .C1(n10247), .C2(n10246), .A(n10245), .B(n15815), .ZN(
        n10248) );
  AOI21_X1 U12867 ( .B1(n15486), .B2(n10249), .A(n10248), .ZN(n10252) );
  NAND2_X1 U12868 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n11039) );
  INV_X1 U12869 ( .A(n11039), .ZN(n10250) );
  AOI21_X1 U12870 ( .B1(n15475), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10250), .ZN(
        n10251) );
  OAI211_X1 U12871 ( .C1(n7500), .C2(n15814), .A(n10252), .B(n10251), .ZN(
        P1_U3248) );
  NAND2_X1 U12872 ( .A1(n11031), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10263) );
  NAND2_X1 U12873 ( .A1(n10902), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10262) );
  NAND2_X1 U12874 ( .A1(n12157), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n10261) );
  AND3_X1 U12875 ( .A1(n10263), .A2(n10262), .A3(n10261), .ZN(n10265) );
  NAND2_X1 U12876 ( .A1(n11032), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n10264) );
  NAND2_X1 U12877 ( .A1(n14791), .A2(n10356), .ZN(n10266) );
  OAI21_X1 U12878 ( .B1(n14791), .B2(n9028), .A(n10266), .ZN(P1_U3560) );
  XNOR2_X1 U12879 ( .A(n11190), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n10269) );
  AOI211_X1 U12880 ( .C1(n10269), .C2(n10268), .A(n10294), .B(n15817), .ZN(
        n10280) );
  NAND2_X1 U12881 ( .A1(n11020), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10272) );
  INV_X1 U12882 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10270) );
  MUX2_X1 U12883 ( .A(n10270), .B(P1_REG2_REG_6__SCAN_IN), .S(n11190), .Z(
        n10271) );
  INV_X1 U12884 ( .A(n10323), .ZN(n10275) );
  NAND3_X1 U12885 ( .A1(n10273), .A2(n10272), .A3(n10271), .ZN(n10274) );
  NAND3_X1 U12886 ( .A1(n15812), .A2(n10275), .A3(n10274), .ZN(n10278) );
  NOR2_X1 U12887 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11028), .ZN(n10276) );
  AOI21_X1 U12888 ( .B1(n15475), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10276), .ZN(
        n10277) );
  OAI211_X1 U12889 ( .C1(n15814), .C2(n10288), .A(n10278), .B(n10277), .ZN(
        n10279) );
  OR2_X1 U12890 ( .A1(n10280), .A2(n10279), .ZN(P1_U3249) );
  OAI222_X1 U12891 ( .A1(n13721), .A2(n10282), .B1(n13723), .B2(n10281), .C1(
        n13207), .C2(P3_U3151), .ZN(P3_U3282) );
  INV_X1 U12892 ( .A(n10283), .ZN(n10285) );
  INV_X1 U12893 ( .A(SI_15_), .ZN(n10284) );
  INV_X1 U12894 ( .A(n13256), .ZN(n13235) );
  OAI222_X1 U12895 ( .A1(n13721), .A2(n10285), .B1(n13723), .B2(n10284), .C1(
        n13235), .C2(P3_U3151), .ZN(P3_U3280) );
  INV_X1 U12896 ( .A(n10495), .ZN(n10840) );
  OAI222_X1 U12897 ( .A1(P2_U3088), .A2(n10840), .B1(n11897), .B2(n10287), 
        .C1(n10286), .C2(n14590), .ZN(P2_U3315) );
  NOR2_X1 U12898 ( .A1(n10288), .A2(n10270), .ZN(n10322) );
  INV_X1 U12899 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10289) );
  MUX2_X1 U12900 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10289), .S(n11440), .Z(
        n10321) );
  NAND2_X1 U12901 ( .A1(n11440), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10292) );
  INV_X1 U12902 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10290) );
  MUX2_X1 U12903 ( .A(n10290), .B(P1_REG2_REG_8__SCAN_IN), .S(n11511), .Z(
        n10291) );
  NAND3_X1 U12904 ( .A1(n10320), .A2(n10292), .A3(n10291), .ZN(n10293) );
  NAND2_X1 U12905 ( .A1(n15812), .A2(n10293), .ZN(n10302) );
  INV_X1 U12906 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n15824) );
  XNOR2_X1 U12907 ( .A(n11511), .B(n15824), .ZN(n10296) );
  XNOR2_X1 U12908 ( .A(n11440), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n10318) );
  OAI21_X1 U12909 ( .B1(n10296), .B2(n10295), .A(n10649), .ZN(n10297) );
  NAND2_X1 U12910 ( .A1(n10297), .A2(n15486), .ZN(n10301) );
  NAND2_X1 U12911 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11874) );
  INV_X1 U12912 ( .A(n11874), .ZN(n10299) );
  NOR2_X1 U12913 ( .A1(n15814), .A2(n10653), .ZN(n10298) );
  AOI211_X1 U12914 ( .C1(n15475), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10299), .B(
        n10298), .ZN(n10300) );
  OAI211_X1 U12915 ( .C1(n14848), .C2(n10302), .A(n10301), .B(n10300), .ZN(
        P1_U3251) );
  INV_X1 U12916 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n15952) );
  NAND2_X1 U12917 ( .A1(n13115), .A2(n13548), .ZN(n10303) );
  OAI21_X1 U12918 ( .B1(P3_U3897), .B2(n15952), .A(n10303), .ZN(P3_U3505) );
  OAI222_X1 U12919 ( .A1(n13721), .A2(n10305), .B1(n13723), .B2(n10304), .C1(
        n13202), .C2(P3_U3151), .ZN(P3_U3281) );
  INV_X1 U12920 ( .A(n10306), .ZN(n10308) );
  OAI222_X1 U12921 ( .A1(n13721), .A2(n10308), .B1(n13723), .B2(n10307), .C1(
        n13257), .C2(P3_U3151), .ZN(P3_U3279) );
  INV_X1 U12922 ( .A(n12153), .ZN(n10315) );
  OAI222_X1 U12923 ( .A1(P2_U3088), .A2(n10876), .B1(n11897), .B2(n10315), 
        .C1(n10309), .C2(n14590), .ZN(P2_U3314) );
  NAND2_X1 U12924 ( .A1(n10311), .A2(n10310), .ZN(n10312) );
  NAND2_X1 U12925 ( .A1(n10312), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10313) );
  NAND2_X1 U12926 ( .A1(n10313), .A2(n10570), .ZN(n10551) );
  OR2_X1 U12927 ( .A1(n10313), .A2(n10570), .ZN(n10314) );
  INV_X1 U12928 ( .A(n14859), .ZN(n11487) );
  OAI222_X1 U12929 ( .A1(n15370), .A2(n10316), .B1(n15379), .B2(n10315), .C1(
        n11487), .C2(P1_U3086), .ZN(P1_U3342) );
  AOI211_X1 U12930 ( .C1(n10319), .C2(n10318), .A(n15817), .B(n10317), .ZN(
        n10329) );
  INV_X1 U12931 ( .A(n10320), .ZN(n10325) );
  NOR3_X1 U12932 ( .A1(n10323), .A2(n10322), .A3(n10321), .ZN(n10324) );
  NOR3_X1 U12933 ( .A1(n15815), .A2(n10325), .A3(n10324), .ZN(n10328) );
  INV_X1 U12934 ( .A(n15475), .ZN(n15821) );
  INV_X1 U12935 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10616) );
  NAND2_X1 U12936 ( .A1(n15483), .A2(n11440), .ZN(n10326) );
  NAND2_X1 U12937 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11458) );
  OAI211_X1 U12938 ( .C1(n15821), .C2(n10616), .A(n10326), .B(n11458), .ZN(
        n10327) );
  OR3_X1 U12939 ( .A1(n10329), .A2(n10328), .A3(n10327), .ZN(P1_U3250) );
  NAND2_X1 U12940 ( .A1(n10330), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10331) );
  INV_X1 U12941 ( .A(n9940), .ZN(n11105) );
  AND2_X1 U12942 ( .A1(n11280), .A2(n15819), .ZN(n10385) );
  INV_X1 U12943 ( .A(n10333), .ZN(n10334) );
  OAI211_X1 U12944 ( .C1(n12859), .C2(n10385), .A(n10376), .B(n10334), .ZN(
        n10915) );
  NAND2_X1 U12945 ( .A1(n11280), .A2(n12673), .ZN(n12858) );
  INV_X1 U12946 ( .A(n12858), .ZN(n10335) );
  NAND2_X2 U12947 ( .A1(n10335), .A2(n12917), .ZN(n15538) );
  OAI21_X1 U12948 ( .B1(n10349), .B2(P1_D_REG_1__SCAN_IN), .A(n10336), .ZN(
        n10375) );
  NOR4_X1 U12949 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n10337) );
  INV_X1 U12950 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n16084) );
  INV_X1 U12951 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15980) );
  NAND3_X1 U12952 ( .A1(n10337), .A2(n16084), .A3(n15980), .ZN(n10343) );
  NOR4_X1 U12953 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n10341) );
  NOR4_X1 U12954 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n10340) );
  NOR4_X1 U12955 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n10339) );
  NOR4_X1 U12956 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n10338) );
  NAND4_X1 U12957 ( .A1(n10341), .A2(n10340), .A3(n10339), .A4(n10338), .ZN(
        n10342) );
  NOR4_X1 U12958 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n10343), .A4(n10342), .ZN(n10345) );
  INV_X1 U12959 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n16039) );
  INV_X1 U12960 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n16034) );
  INV_X1 U12961 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15894) );
  INV_X1 U12962 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15893) );
  NAND4_X1 U12963 ( .A1(n16039), .A2(n16034), .A3(n15894), .A4(n15893), .ZN(
        n10344) );
  NOR3_X1 U12964 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        n10344), .ZN(n15837) );
  AND2_X1 U12965 ( .A1(n10345), .A2(n15837), .ZN(n10346) );
  NOR2_X1 U12966 ( .A1(n10349), .A2(n10346), .ZN(n10374) );
  INV_X1 U12967 ( .A(n10374), .ZN(n10347) );
  NAND4_X1 U12968 ( .A1(n12913), .A2(n11130), .A3(n10375), .A4(n10347), .ZN(
        n15203) );
  INV_X1 U12969 ( .A(n15202), .ZN(n10350) );
  INV_X1 U12970 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10366) );
  NAND2_X1 U12971 ( .A1(n12917), .A2(n12673), .ZN(n10386) );
  MUX2_X1 U12972 ( .A(n6932), .B(n10351), .S(n6555), .Z(n11317) );
  NOR2_X1 U12973 ( .A1(n12673), .A2(n12672), .ZN(n10352) );
  OR2_X2 U12974 ( .A1(n12683), .A2(n10352), .ZN(n11860) );
  NAND2_X1 U12975 ( .A1(n12683), .A2(n15381), .ZN(n10353) );
  NAND2_X1 U12976 ( .A1(n11860), .A2(n10353), .ZN(n11320) );
  OR2_X1 U12977 ( .A1(n12858), .A2(n15819), .ZN(n15565) );
  NAND2_X1 U12978 ( .A1(n10354), .A2(n12675), .ZN(n12674) );
  OR2_X1 U12979 ( .A1(n12673), .A2(n15819), .ZN(n10355) );
  INV_X1 U12980 ( .A(n12679), .ZN(n10358) );
  NAND2_X1 U12981 ( .A1(n10356), .A2(n11317), .ZN(n10357) );
  INV_X1 U12982 ( .A(n12684), .ZN(n12869) );
  OAI21_X1 U12983 ( .B1(n15561), .B2(n15552), .A(n12869), .ZN(n10364) );
  INV_X1 U12984 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10359) );
  NAND2_X1 U12985 ( .A1(n10902), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10362) );
  NAND2_X1 U12986 ( .A1(n12157), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n10361) );
  NAND2_X1 U12987 ( .A1(n11031), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10360) );
  NAND2_X1 U12988 ( .A1(n14792), .A2(n15178), .ZN(n11316) );
  OAI211_X1 U12989 ( .C1(n10386), .C2(n11317), .A(n10364), .B(n11316), .ZN(
        n15341) );
  NAND2_X1 U12990 ( .A1(n15341), .A2(n15608), .ZN(n10365) );
  OAI21_X1 U12991 ( .B1(n15608), .B2(n10366), .A(n10365), .ZN(P1_U3459) );
  INV_X1 U12992 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n15903) );
  NAND2_X1 U12993 ( .A1(P3_U3897), .A2(n11241), .ZN(n10367) );
  OAI21_X1 U12994 ( .B1(n13115), .B2(n15903), .A(n10367), .ZN(P3_U3494) );
  INV_X1 U12995 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n15904) );
  NAND2_X1 U12996 ( .A1(n11759), .A2(P3_U3897), .ZN(n10368) );
  OAI21_X1 U12997 ( .B1(n13115), .B2(n15904), .A(n10368), .ZN(P3_U3500) );
  INV_X1 U12998 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n15997) );
  NAND2_X1 U12999 ( .A1(n12106), .A2(P3_U3897), .ZN(n10369) );
  OAI21_X1 U13000 ( .B1(P3_U3897), .B2(n15997), .A(n10369), .ZN(P3_U3504) );
  NOR2_X1 U13001 ( .A1(n10530), .A2(n13552), .ZN(n10370) );
  OAI22_X1 U13002 ( .A1(n10564), .A2(n10370), .B1(n7429), .B2(n13535), .ZN(
        n10711) );
  INV_X1 U13003 ( .A(n10711), .ZN(n10372) );
  MUX2_X1 U13004 ( .A(n10372), .B(n10371), .S(n15801), .Z(n10373) );
  OAI21_X1 U13005 ( .B1(n10715), .B2(n13610), .A(n10373), .ZN(P3_U3459) );
  INV_X1 U13006 ( .A(n14792), .ZN(n11134) );
  OR2_X1 U13007 ( .A1(n10375), .A2(n10374), .ZN(n11127) );
  NOR2_X1 U13008 ( .A1(n11127), .A2(n15202), .ZN(n10389) );
  NAND2_X1 U13009 ( .A1(n10389), .A2(n12913), .ZN(n14737) );
  INV_X1 U13010 ( .A(n12683), .ZN(n11132) );
  NAND2_X1 U13011 ( .A1(n10910), .A2(n10356), .ZN(n10378) );
  INV_X1 U13012 ( .A(n10376), .ZN(n10380) );
  NAND2_X2 U13013 ( .A1(n10376), .A2(n12683), .ZN(n10379) );
  NAND2_X1 U13014 ( .A1(n10356), .A2(n12552), .ZN(n10382) );
  NAND2_X1 U13015 ( .A1(n10380), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10381) );
  OAI211_X1 U13016 ( .C1(n14638), .C2(n11317), .A(n10382), .B(n10381), .ZN(
        n10672) );
  INV_X1 U13017 ( .A(n10673), .ZN(n10383) );
  OAI21_X1 U13018 ( .B1(n10384), .B2(n10672), .A(n10383), .ZN(n10462) );
  NAND2_X1 U13019 ( .A1(n15599), .A2(n12859), .ZN(n10387) );
  NOR2_X1 U13020 ( .A1(n11131), .A2(n10387), .ZN(n10388) );
  INV_X1 U13021 ( .A(n10389), .ZN(n10390) );
  NAND2_X1 U13022 ( .A1(n10390), .A2(n11130), .ZN(n10917) );
  NAND2_X1 U13023 ( .A1(n10917), .A2(n12913), .ZN(n10706) );
  AOI22_X1 U13024 ( .A1(n10462), .A2(n14753), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n10706), .ZN(n10393) );
  INV_X1 U13025 ( .A(n11131), .ZN(n10391) );
  AND2_X1 U13026 ( .A1(n10917), .A2(n10391), .ZN(n11042) );
  NAND2_X1 U13027 ( .A1(n14740), .A2(n6937), .ZN(n10392) );
  OAI211_X1 U13028 ( .C1(n11134), .C2(n14706), .A(n10393), .B(n10392), .ZN(
        P1_U3232) );
  INV_X1 U13029 ( .A(n10394), .ZN(n10396) );
  INV_X1 U13030 ( .A(n13301), .ZN(n13279) );
  OAI222_X1 U13031 ( .A1(n13721), .A2(n10396), .B1(n13723), .B2(n10395), .C1(
        n13279), .C2(P3_U3151), .ZN(P3_U3278) );
  OR2_X1 U13032 ( .A1(n10397), .A2(P2_U3088), .ZN(n10561) );
  INV_X1 U13033 ( .A(n10561), .ZN(n10414) );
  INV_X1 U13034 ( .A(n8788), .ZN(n10399) );
  INV_X1 U13035 ( .A(n13956), .ZN(n10398) );
  OAI22_X1 U13036 ( .A1(n10399), .A2(n13915), .B1(n10398), .B2(n13917), .ZN(
        n11975) );
  AOI22_X1 U13037 ( .A1(n13919), .A2(n11975), .B1(n13923), .B2(n7528), .ZN(
        n10405) );
  OAI21_X1 U13038 ( .B1(n10402), .B2(n10401), .A(n10400), .ZN(n10403) );
  NAND2_X1 U13039 ( .A1(n13903), .A2(n10403), .ZN(n10404) );
  OAI211_X1 U13040 ( .C1(n10414), .C2(n8438), .A(n10405), .B(n10404), .ZN(
        P2_U3194) );
  INV_X1 U13041 ( .A(n8781), .ZN(n10407) );
  INV_X1 U13042 ( .A(n13955), .ZN(n10406) );
  OAI22_X1 U13043 ( .A1(n10407), .A2(n13915), .B1(n10406), .B2(n13917), .ZN(
        n10579) );
  AOI22_X1 U13044 ( .A1(n13919), .A2(n10579), .B1(n13923), .B2(n11934), .ZN(
        n10413) );
  OAI21_X1 U13045 ( .B1(n10410), .B2(n10409), .A(n10408), .ZN(n10411) );
  NAND2_X1 U13046 ( .A1(n13903), .A2(n10411), .ZN(n10412) );
  OAI211_X1 U13047 ( .C1(n10414), .C2(n13958), .A(n10413), .B(n10412), .ZN(
        P2_U3209) );
  XNOR2_X1 U13048 ( .A(n10484), .B(n14512), .ZN(n10425) );
  INV_X1 U13049 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10415) );
  NAND2_X1 U13050 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15630) );
  OAI22_X1 U13051 ( .A1(n15631), .A2(n15630), .B1(n10433), .B2(n10415), .ZN(
        n13962) );
  MUX2_X1 U13052 ( .A(n8454), .B(P2_REG1_REG_2__SCAN_IN), .S(n13964), .Z(
        n13963) );
  NAND2_X1 U13053 ( .A1(n13962), .A2(n13963), .ZN(n13961) );
  INV_X1 U13054 ( .A(n13964), .ZN(n13960) );
  NAND2_X1 U13055 ( .A1(n13960), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10416) );
  NAND2_X1 U13056 ( .A1(n13961), .A2(n10416), .ZN(n15645) );
  MUX2_X1 U13057 ( .A(n10417), .B(P2_REG1_REG_3__SCAN_IN), .S(n15642), .Z(
        n15646) );
  NAND2_X1 U13058 ( .A1(n15645), .A2(n15646), .ZN(n15643) );
  OR2_X1 U13059 ( .A1(n15642), .A2(n10417), .ZN(n10418) );
  NAND2_X1 U13060 ( .A1(n15643), .A2(n10418), .ZN(n13975) );
  MUX2_X1 U13061 ( .A(n8470), .B(P2_REG1_REG_4__SCAN_IN), .S(n13977), .Z(
        n13976) );
  NAND2_X1 U13062 ( .A1(n13975), .A2(n13976), .ZN(n13974) );
  INV_X1 U13063 ( .A(n13977), .ZN(n10441) );
  NAND2_X1 U13064 ( .A1(n10441), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10419) );
  NAND2_X1 U13065 ( .A1(n13974), .A2(n10419), .ZN(n13988) );
  MUX2_X1 U13066 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n8480), .S(n13990), .Z(
        n13989) );
  NAND2_X1 U13067 ( .A1(n13988), .A2(n13989), .ZN(n13987) );
  NAND2_X1 U13068 ( .A1(n13990), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10420) );
  NAND2_X1 U13069 ( .A1(n13987), .A2(n10420), .ZN(n14002) );
  MUX2_X1 U13070 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n8491), .S(n14004), .Z(
        n14003) );
  NAND2_X1 U13071 ( .A1(n14002), .A2(n14003), .ZN(n14001) );
  NAND2_X1 U13072 ( .A1(n14004), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10421) );
  MUX2_X1 U13073 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n8502), .S(n14020), .Z(
        n14014) );
  XNOR2_X1 U13074 ( .A(n14033), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n14031) );
  NAND2_X1 U13075 ( .A1(n14029), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10422) );
  NAND2_X1 U13076 ( .A1(n14030), .A2(n10422), .ZN(n10424) );
  INV_X1 U13077 ( .A(n10477), .ZN(n10423) );
  AOI21_X1 U13078 ( .B1(n10425), .B2(n10424), .A(n10423), .ZN(n10461) );
  NAND2_X1 U13079 ( .A1(n10427), .A2(n10426), .ZN(n10429) );
  NAND2_X1 U13080 ( .A1(n10429), .A2(n10428), .ZN(n10432) );
  INV_X1 U13081 ( .A(n10430), .ZN(n10431) );
  NAND2_X1 U13082 ( .A1(n10432), .A2(n10431), .ZN(n15633) );
  NOR2_X1 U13083 ( .A1(n8398), .A2(P2_U3088), .ZN(n14591) );
  AND2_X1 U13084 ( .A1(n15633), .A2(n14591), .ZN(n10454) );
  MUX2_X1 U13085 ( .A(n11977), .B(P2_REG2_REG_1__SCAN_IN), .S(n10433), .Z(
        n15637) );
  AND2_X1 U13086 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n15638) );
  NAND2_X1 U13087 ( .A1(n15637), .A2(n15638), .ZN(n15636) );
  INV_X1 U13088 ( .A(n10433), .ZN(n10434) );
  NAND2_X1 U13089 ( .A1(n10434), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n13965) );
  NAND2_X1 U13090 ( .A1(n15636), .A2(n13965), .ZN(n10437) );
  MUX2_X1 U13091 ( .A(n10435), .B(P2_REG2_REG_2__SCAN_IN), .S(n13964), .Z(
        n10436) );
  NAND2_X1 U13092 ( .A1(n10437), .A2(n10436), .ZN(n13968) );
  NAND2_X1 U13093 ( .A1(n13960), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10438) );
  NAND2_X1 U13094 ( .A1(n13968), .A2(n10438), .ZN(n15654) );
  MUX2_X1 U13095 ( .A(n11714), .B(P2_REG2_REG_3__SCAN_IN), .S(n15642), .Z(
        n15655) );
  NAND2_X1 U13096 ( .A1(n15654), .A2(n15655), .ZN(n15652) );
  OR2_X1 U13097 ( .A1(n15642), .A2(n11714), .ZN(n13978) );
  NAND2_X1 U13098 ( .A1(n15652), .A2(n13978), .ZN(n10440) );
  INV_X1 U13099 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11629) );
  MUX2_X1 U13100 ( .A(n11629), .B(P2_REG2_REG_4__SCAN_IN), .S(n13977), .Z(
        n10439) );
  NAND2_X1 U13101 ( .A1(n10440), .A2(n10439), .ZN(n13993) );
  NAND2_X1 U13102 ( .A1(n10441), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n13992) );
  NAND2_X1 U13103 ( .A1(n13993), .A2(n13992), .ZN(n10443) );
  INV_X1 U13104 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11965) );
  MUX2_X1 U13105 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11965), .S(n13990), .Z(
        n10442) );
  NAND2_X1 U13106 ( .A1(n10443), .A2(n10442), .ZN(n14007) );
  NAND2_X1 U13107 ( .A1(n13990), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n14006) );
  NAND2_X1 U13108 ( .A1(n14007), .A2(n14006), .ZN(n10446) );
  MUX2_X1 U13109 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10444), .S(n14004), .Z(
        n10445) );
  NAND2_X1 U13110 ( .A1(n10446), .A2(n10445), .ZN(n14017) );
  NAND2_X1 U13111 ( .A1(n14004), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n14016) );
  NAND2_X1 U13112 ( .A1(n14017), .A2(n14016), .ZN(n10448) );
  MUX2_X1 U13113 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11996), .S(n14020), .Z(
        n10447) );
  NAND2_X1 U13114 ( .A1(n10448), .A2(n10447), .ZN(n14036) );
  NAND2_X1 U13115 ( .A1(n14020), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n14035) );
  NAND2_X1 U13116 ( .A1(n14036), .A2(n14035), .ZN(n10450) );
  MUX2_X1 U13117 ( .A(n11693), .B(P2_REG2_REG_8__SCAN_IN), .S(n14033), .Z(
        n10449) );
  NAND2_X1 U13118 ( .A1(n10450), .A2(n10449), .ZN(n14038) );
  NAND2_X1 U13119 ( .A1(n14029), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10451) );
  AND2_X1 U13120 ( .A1(n14038), .A2(n10451), .ZN(n10453) );
  INV_X1 U13121 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10483) );
  MUX2_X1 U13122 ( .A(n10483), .B(P2_REG2_REG_9__SCAN_IN), .S(n10484), .Z(
        n10452) );
  NAND2_X1 U13123 ( .A1(n10453), .A2(n10452), .ZN(n10486) );
  OAI21_X1 U13124 ( .B1(n10453), .B2(n10452), .A(n10486), .ZN(n10459) );
  INV_X1 U13125 ( .A(n10454), .ZN(n10455) );
  INV_X1 U13126 ( .A(n15623), .ZN(n15653) );
  AND2_X1 U13127 ( .A1(n8398), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10456) );
  INV_X1 U13128 ( .A(n15651), .ZN(n14082) );
  OR2_X1 U13129 ( .A1(n15633), .A2(P2_U3088), .ZN(n15658) );
  INV_X1 U13130 ( .A(n15658), .ZN(n15629) );
  AND2_X1 U13131 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n11928) );
  AOI21_X1 U13132 ( .B1(n15629), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n11928), .ZN(
        n10457) );
  OAI21_X1 U13133 ( .B1(n10484), .B2(n14082), .A(n10457), .ZN(n10458) );
  AOI21_X1 U13134 ( .B1(n10459), .B2(n15653), .A(n10458), .ZN(n10460) );
  OAI21_X1 U13135 ( .B1(n10461), .B2(n15624), .A(n10460), .ZN(P2_U3223) );
  NAND2_X1 U13136 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14797) );
  MUX2_X1 U13137 ( .A(n14797), .B(n10462), .S(n6762), .Z(n10465) );
  OAI21_X1 U13138 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n6762), .A(n10692), .ZN(
        n15471) );
  NAND2_X1 U13139 ( .A1(n15471), .A2(n6932), .ZN(n10464) );
  OAI211_X1 U13140 ( .C1(n10465), .C2(n10463), .A(n14791), .B(n10464), .ZN(
        n14818) );
  INV_X1 U13141 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10466) );
  NAND2_X1 U13142 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10929) );
  OAI21_X1 U13143 ( .B1(n15821), .B2(n10466), .A(n10929), .ZN(n10474) );
  XNOR2_X1 U13144 ( .A(n10468), .B(n10467), .ZN(n10472) );
  OAI21_X1 U13145 ( .B1(n10470), .B2(n10469), .A(n7303), .ZN(n10471) );
  OAI22_X1 U13146 ( .A1(n15815), .A2(n10472), .B1(n15817), .B2(n10471), .ZN(
        n10473) );
  AOI211_X1 U13147 ( .C1(n10898), .C2(n15483), .A(n10474), .B(n10473), .ZN(
        n10475) );
  NAND2_X1 U13148 ( .A1(n14818), .A2(n10475), .ZN(P1_U3247) );
  XNOR2_X1 U13149 ( .A(n10495), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n10482) );
  NAND2_X1 U13150 ( .A1(n10484), .A2(n14512), .ZN(n10476) );
  XNOR2_X1 U13151 ( .A(n10724), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n10719) );
  NAND2_X1 U13152 ( .A1(n10724), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10478) );
  XNOR2_X1 U13153 ( .A(n14052), .B(n14501), .ZN(n14043) );
  NAND2_X1 U13154 ( .A1(n14044), .A2(n14043), .ZN(n14042) );
  NAND2_X1 U13155 ( .A1(n14052), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10479) );
  NAND2_X1 U13156 ( .A1(n14042), .A2(n10479), .ZN(n10481) );
  INV_X1 U13157 ( .A(n10842), .ZN(n10480) );
  AOI21_X1 U13158 ( .B1(n10482), .B2(n10481), .A(n10480), .ZN(n10497) );
  INV_X1 U13159 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n12192) );
  NAND2_X1 U13160 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n13816)
         );
  OAI21_X1 U13161 ( .B1(n15658), .B2(n12192), .A(n13816), .ZN(n10494) );
  NAND2_X1 U13162 ( .A1(n10484), .A2(n10483), .ZN(n10485) );
  NAND2_X1 U13163 ( .A1(n10486), .A2(n10485), .ZN(n10723) );
  MUX2_X1 U13164 ( .A(n8527), .B(P2_REG2_REG_10__SCAN_IN), .S(n10724), .Z(
        n10722) );
  OR2_X1 U13165 ( .A1(n10723), .A2(n10722), .ZN(n10720) );
  NAND2_X1 U13166 ( .A1(n10724), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10487) );
  AND2_X1 U13167 ( .A1(n10720), .A2(n10487), .ZN(n14047) );
  INV_X1 U13168 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n16086) );
  MUX2_X1 U13169 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n16086), .S(n14052), .Z(
        n14046) );
  NAND2_X1 U13170 ( .A1(n14047), .A2(n14046), .ZN(n14045) );
  OR2_X1 U13171 ( .A1(n14052), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10490) );
  NAND2_X1 U13172 ( .A1(n14045), .A2(n10490), .ZN(n10488) );
  MUX2_X1 U13173 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n14352), .S(n10495), .Z(
        n10489) );
  NAND2_X1 U13174 ( .A1(n10488), .A2(n10489), .ZN(n10834) );
  INV_X1 U13175 ( .A(n10489), .ZN(n10491) );
  NAND3_X1 U13176 ( .A1(n14045), .A2(n10491), .A3(n10490), .ZN(n10492) );
  AOI21_X1 U13177 ( .B1(n10834), .B2(n10492), .A(n15623), .ZN(n10493) );
  AOI211_X1 U13178 ( .C1(n15651), .C2(n10495), .A(n10494), .B(n10493), .ZN(
        n10496) );
  OAI21_X1 U13179 ( .B1(n10497), .B2(n15624), .A(n10496), .ZN(P2_U3226) );
  NAND2_X1 U13180 ( .A1(n10534), .A2(n10498), .ZN(n10505) );
  INV_X1 U13181 ( .A(n10531), .ZN(n10503) );
  NAND3_X1 U13182 ( .A1(n10501), .A2(n10500), .A3(n10499), .ZN(n10502) );
  AOI21_X1 U13183 ( .B1(n10532), .B2(n10503), .A(n10502), .ZN(n10504) );
  NAND2_X1 U13184 ( .A1(n10505), .A2(n10504), .ZN(n10506) );
  NAND2_X1 U13185 ( .A1(n10506), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10509) );
  NAND2_X1 U13186 ( .A1(n10507), .A2(n10532), .ZN(n10508) );
  NOR2_X1 U13187 ( .A1(n13095), .A2(P3_U3151), .ZN(n10639) );
  NAND2_X1 U13188 ( .A1(n10535), .A2(n13598), .ZN(n10510) );
  OR2_X1 U13189 ( .A1(n10534), .A2(n10510), .ZN(n10511) );
  INV_X1 U13190 ( .A(n10532), .ZN(n10514) );
  NOR2_X1 U13191 ( .A1(n10513), .A2(n13535), .ZN(n10515) );
  INV_X1 U13192 ( .A(n13120), .ZN(n10596) );
  OAI22_X1 U13193 ( .A1(n13099), .A2(n10516), .B1(n13088), .B2(n10596), .ZN(
        n10517) );
  AOI21_X1 U13194 ( .B1(n9173), .B2(n13102), .A(n10517), .ZN(n10539) );
  NAND2_X1 U13195 ( .A1(n13121), .A2(n9173), .ZN(n10518) );
  NAND2_X1 U13196 ( .A1(n13703), .A2(n10520), .ZN(n10523) );
  OAI21_X1 U13197 ( .B1(n10521), .B2(n10631), .A(n11251), .ZN(n10522) );
  NAND2_X1 U13198 ( .A1(n12995), .A2(n11048), .ZN(n10525) );
  NAND2_X1 U13199 ( .A1(n10526), .A2(n10525), .ZN(n10527) );
  NAND3_X1 U13200 ( .A1(n11056), .A2(n7247), .A3(n11055), .ZN(n10528) );
  OAI211_X1 U13201 ( .C1(n10529), .C2(n11048), .A(n10590), .B(n10528), .ZN(
        n10537) );
  INV_X1 U13202 ( .A(n10530), .ZN(n10533) );
  OAI22_X1 U13203 ( .A1(n10534), .A2(n10533), .B1(n10532), .B2(n10531), .ZN(
        n10536) );
  INV_X1 U13204 ( .A(n13104), .ZN(n11608) );
  NAND2_X1 U13205 ( .A1(n10537), .A2(n11608), .ZN(n10538) );
  OAI211_X1 U13206 ( .C1(n10639), .C2(n11089), .A(n10539), .B(n10538), .ZN(
        P3_U3162) );
  BUF_X1 U13207 ( .A(n10540), .Z(n10541) );
  INV_X1 U13208 ( .A(n10541), .ZN(n10542) );
  OAI21_X1 U13209 ( .B1(n10543), .B2(n10542), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n10544) );
  XNOR2_X1 U13210 ( .A(n10544), .B(P1_IR_REG_16__SCAN_IN), .ZN(n14887) );
  INV_X1 U13211 ( .A(n14887), .ZN(n14881) );
  INV_X1 U13212 ( .A(n12261), .ZN(n10546) );
  OAI222_X1 U13213 ( .A1(P1_U3086), .A2(n14881), .B1(n15379), .B2(n10546), 
        .C1(n10545), .C2(n15370), .ZN(P1_U3339) );
  INV_X1 U13214 ( .A(n11886), .ZN(n10547) );
  OAI222_X1 U13215 ( .A1(P2_U3088), .A2(n10547), .B1(n11897), .B2(n10546), 
        .C1(n15888), .C2(n14590), .ZN(P2_U3311) );
  INV_X1 U13216 ( .A(n10548), .ZN(n10550) );
  INV_X1 U13217 ( .A(n13302), .ZN(n13326) );
  OAI222_X1 U13218 ( .A1(n13721), .A2(n10550), .B1(n13723), .B2(n10549), .C1(
        n13326), .C2(P3_U3151), .ZN(P3_U3277) );
  INV_X1 U13219 ( .A(n12244), .ZN(n10555) );
  NAND2_X1 U13220 ( .A1(n10551), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10552) );
  INV_X1 U13221 ( .A(n14868), .ZN(n14873) );
  OAI222_X1 U13222 ( .A1(n15370), .A2(n10553), .B1(n15379), .B2(n10555), .C1(
        n14873), .C2(P1_U3086), .ZN(P1_U3341) );
  INV_X1 U13223 ( .A(n11292), .ZN(n10837) );
  OAI222_X1 U13224 ( .A1(P2_U3088), .A2(n10837), .B1(n11897), .B2(n10555), 
        .C1(n10554), .C2(n14590), .ZN(P2_U3313) );
  NAND2_X1 U13225 ( .A1(n8781), .A2(n13907), .ZN(n15663) );
  NAND2_X1 U13226 ( .A1(n8788), .A2(n6556), .ZN(n10557) );
  INV_X1 U13227 ( .A(n10557), .ZN(n10556) );
  NAND2_X1 U13228 ( .A1(n13903), .A2(n10556), .ZN(n10560) );
  AOI21_X1 U13229 ( .B1(n13903), .B2(n10557), .A(n13923), .ZN(n10559) );
  MUX2_X1 U13230 ( .A(n10560), .B(n10559), .S(n10558), .Z(n10563) );
  NAND2_X1 U13231 ( .A1(n10561), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n10562) );
  OAI211_X1 U13232 ( .C1(n13855), .C2(n15663), .A(n10563), .B(n10562), .ZN(
        P2_U3204) );
  INV_X1 U13233 ( .A(n10564), .ZN(n10566) );
  OAI22_X1 U13234 ( .A1(n13081), .A2(n10715), .B1(n7429), .B2(n13088), .ZN(
        n10565) );
  AOI21_X1 U13235 ( .B1(n11608), .B2(n10566), .A(n10565), .ZN(n10567) );
  OAI21_X1 U13236 ( .B1(n10639), .B2(n11062), .A(n10567), .ZN(P3_U3172) );
  INV_X1 U13237 ( .A(n12250), .ZN(n10640) );
  INV_X1 U13238 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n10569) );
  INV_X1 U13239 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10568) );
  NAND4_X1 U13240 ( .A1(n10570), .A2(n10310), .A3(n10569), .A4(n10568), .ZN(
        n10571) );
  OAI21_X1 U13241 ( .B1(n10572), .B2(n10571), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n10573) );
  XNOR2_X1 U13242 ( .A(n10573), .B(P1_IR_REG_15__SCAN_IN), .ZN(n15484) );
  AOI22_X1 U13243 ( .A1(n15484), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n15367), .ZN(n10574) );
  OAI21_X1 U13244 ( .B1(n10640), .B2(n15379), .A(n10574), .ZN(P1_U3340) );
  OAI21_X1 U13245 ( .B1(n10575), .B2(n10577), .A(n10576), .ZN(n11938) );
  INV_X1 U13246 ( .A(n11970), .ZN(n10578) );
  OAI211_X1 U13247 ( .C1(n10578), .C2(n10584), .A(n14470), .B(n11716), .ZN(
        n11936) );
  INV_X1 U13248 ( .A(n11936), .ZN(n10582) );
  XNOR2_X1 U13249 ( .A(n11707), .B(n11706), .ZN(n10580) );
  AOI21_X1 U13250 ( .B1(n10580), .B2(n15662), .A(n10579), .ZN(n11940) );
  INV_X1 U13251 ( .A(n11940), .ZN(n10581) );
  AOI211_X1 U13252 ( .C1(n15740), .C2(n11938), .A(n10582), .B(n10581), .ZN(
        n10648) );
  INV_X1 U13253 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10583) );
  OAI22_X1 U13254 ( .A1(n14574), .A2(n10584), .B1(n15743), .B2(n10583), .ZN(
        n10585) );
  INV_X1 U13255 ( .A(n10585), .ZN(n10586) );
  OAI21_X1 U13256 ( .B1(n10648), .B2(n15741), .A(n10586), .ZN(P2_U3436) );
  XNOR2_X1 U13257 ( .A(n12947), .B(n9173), .ZN(n10588) );
  NAND2_X1 U13258 ( .A1(n10588), .A2(n7429), .ZN(n10589) );
  XNOR2_X1 U13259 ( .A(n10587), .B(n10765), .ZN(n10591) );
  XNOR2_X1 U13260 ( .A(n10591), .B(n13120), .ZN(n10634) );
  NAND2_X1 U13261 ( .A1(n10591), .A2(n10596), .ZN(n10592) );
  XNOR2_X1 U13262 ( .A(n10587), .B(n10599), .ZN(n10995) );
  XNOR2_X1 U13263 ( .A(n10995), .B(n11241), .ZN(n10593) );
  AOI21_X1 U13264 ( .B1(n10632), .B2(n10592), .A(n10593), .ZN(n10602) );
  AND2_X1 U13265 ( .A1(n10593), .A2(n10592), .ZN(n10594) );
  NAND2_X1 U13266 ( .A1(n10998), .A2(n11608), .ZN(n10601) );
  INV_X1 U13267 ( .A(n13119), .ZN(n11275) );
  OAI22_X1 U13268 ( .A1(n13099), .A2(n10596), .B1(n13088), .B2(n11275), .ZN(
        n10598) );
  MUX2_X1 U13269 ( .A(n13095), .B(P3_U3151), .S(P3_REG3_REG_3__SCAN_IN), .Z(
        n10597) );
  AOI211_X1 U13270 ( .C1(n10599), .C2(n13102), .A(n10598), .B(n10597), .ZN(
        n10600) );
  OAI21_X1 U13271 ( .B1(n10602), .B2(n10601), .A(n10600), .ZN(P3_U3158) );
  NAND2_X1 U13272 ( .A1(n10606), .A2(n10605), .ZN(n10612) );
  XNOR2_X1 U13273 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n10607) );
  XNOR2_X1 U13274 ( .A(n10612), .B(n10607), .ZN(n15386) );
  INV_X1 U13275 ( .A(n10608), .ZN(n10609) );
  NAND2_X1 U13276 ( .A1(n10609), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10610) );
  INV_X1 U13277 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n10614) );
  NAND2_X1 U13278 ( .A1(n10612), .A2(n10611), .ZN(n10613) );
  INV_X1 U13279 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n10615) );
  XNOR2_X1 U13280 ( .A(n10621), .B(n10615), .ZN(n10620) );
  XNOR2_X1 U13281 ( .A(n10620), .B(n10616), .ZN(n15388) );
  NAND2_X1 U13282 ( .A1(n10617), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n10618) );
  NAND2_X1 U13283 ( .A1(n10620), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n10623) );
  INV_X1 U13284 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n10624) );
  NAND2_X1 U13285 ( .A1(n10624), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n10942) );
  INV_X1 U13286 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10625) );
  NAND2_X1 U13287 ( .A1(n10625), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n10626) );
  AND2_X1 U13288 ( .A1(n10942), .A2(n10626), .ZN(n10940) );
  XNOR2_X1 U13289 ( .A(n10941), .B(n10940), .ZN(n10936) );
  INV_X1 U13290 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14026) );
  XNOR2_X1 U13291 ( .A(n10935), .B(n14026), .ZN(SUB_1596_U55) );
  NOR2_X1 U13292 ( .A1(n15786), .A2(n9157), .ZN(n10627) );
  AOI21_X1 U13293 ( .B1(n15786), .B2(n10711), .A(n10627), .ZN(n10628) );
  OAI21_X1 U13294 ( .B1(n10715), .B2(n13688), .A(n10628), .ZN(P3_U3390) );
  OAI222_X1 U13295 ( .A1(P3_U3151), .A2(n10631), .B1(n13723), .B2(n10630), 
        .C1(n13721), .C2(n10629), .ZN(P3_U3276) );
  OAI21_X1 U13296 ( .B1(n10634), .B2(n10633), .A(n10632), .ZN(n10635) );
  NAND2_X1 U13297 ( .A1(n10635), .A2(n11608), .ZN(n10638) );
  INV_X1 U13298 ( .A(n11241), .ZN(n11006) );
  OAI22_X1 U13299 ( .A1(n13099), .A2(n7429), .B1(n13088), .B2(n11006), .ZN(
        n10636) );
  AOI21_X1 U13300 ( .B1(n10765), .B2(n13102), .A(n10636), .ZN(n10637) );
  OAI211_X1 U13301 ( .C1(n10639), .C2(n10767), .A(n10638), .B(n10637), .ZN(
        P3_U3177) );
  INV_X1 U13302 ( .A(n11830), .ZN(n11295) );
  OAI222_X1 U13303 ( .A1(n14590), .A2(n10641), .B1(n11897), .B2(n10640), .C1(
        P2_U3088), .C2(n11295), .ZN(P2_U3312) );
  NAND2_X1 U13304 ( .A1(n10642), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10643) );
  XNOR2_X1 U13305 ( .A(n10643), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14902) );
  INV_X1 U13306 ( .A(n14902), .ZN(n14907) );
  INV_X1 U13307 ( .A(n12272), .ZN(n10645) );
  OAI222_X1 U13308 ( .A1(P1_U3086), .A2(n14907), .B1(n15379), .B2(n10645), 
        .C1(n16042), .C2(n15370), .ZN(P1_U3338) );
  OAI222_X1 U13309 ( .A1(P2_U3088), .A2(n11836), .B1(n11897), .B2(n10645), 
        .C1(n10644), .C2(n14590), .ZN(P2_U3310) );
  INV_X1 U13310 ( .A(n14514), .ZN(n10646) );
  AOI22_X1 U13311 ( .A1(n10646), .A2(n11934), .B1(n12591), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n10647) );
  OAI21_X1 U13312 ( .B1(n10648), .B2(n12591), .A(n10647), .ZN(P2_U3501) );
  XNOR2_X1 U13313 ( .A(n11494), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n10652) );
  OAI21_X1 U13314 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n11511), .A(n10649), .ZN(
        n14836) );
  INV_X1 U13315 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10650) );
  MUX2_X1 U13316 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10650), .S(n14842), .Z(
        n14837) );
  NAND2_X1 U13317 ( .A1(n14836), .A2(n14837), .ZN(n14835) );
  AOI211_X1 U13318 ( .C1(n10652), .C2(n10651), .A(n15817), .B(n10818), .ZN(
        n10662) );
  NOR2_X1 U13319 ( .A1(n10653), .A2(n10290), .ZN(n14843) );
  INV_X1 U13320 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10654) );
  MUX2_X1 U13321 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10654), .S(n14842), .Z(
        n10655) );
  OAI21_X1 U13322 ( .B1(n14848), .B2(n14843), .A(n10655), .ZN(n14846) );
  NAND2_X1 U13323 ( .A1(n14842), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10657) );
  INV_X1 U13324 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10821) );
  MUX2_X1 U13325 ( .A(n10821), .B(P1_REG2_REG_10__SCAN_IN), .S(n11494), .Z(
        n10656) );
  AND3_X1 U13326 ( .A1(n14846), .A2(n10657), .A3(n10656), .ZN(n10658) );
  NOR3_X1 U13327 ( .A1(n10826), .A2(n10658), .A3(n15815), .ZN(n10661) );
  NAND2_X1 U13328 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n12213)
         );
  NAND2_X1 U13329 ( .A1(n15475), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n10659) );
  OAI211_X1 U13330 ( .C1(n15814), .C2(n10822), .A(n12213), .B(n10659), .ZN(
        n10660) );
  OR3_X1 U13331 ( .A1(n10662), .A2(n10661), .A3(n10660), .ZN(P1_U3253) );
  INV_X1 U13332 ( .A(n10663), .ZN(n10664) );
  NAND2_X1 U13333 ( .A1(n11018), .A2(n10664), .ZN(n10667) );
  AND2_X1 U13334 ( .A1(n10885), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n10665) );
  INV_X1 U13335 ( .A(n11133), .ZN(n10668) );
  XNOR2_X1 U13336 ( .A(n10671), .B(n11860), .ZN(n10686) );
  XNOR2_X1 U13337 ( .A(n10685), .B(n10686), .ZN(n10687) );
  INV_X1 U13338 ( .A(n10672), .ZN(n10674) );
  XOR2_X1 U13339 ( .A(n10687), .B(n10688), .Z(n10684) );
  INV_X1 U13340 ( .A(n10356), .ZN(n11138) );
  INV_X1 U13341 ( .A(n12859), .ZN(n10675) );
  INV_X1 U13342 ( .A(n14706), .ZN(n14720) );
  NAND2_X1 U13343 ( .A1(n12157), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n10677) );
  NAND2_X1 U13344 ( .A1(n10902), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n10676) );
  AND2_X1 U13345 ( .A1(n10677), .A2(n10676), .ZN(n10680) );
  NAND2_X1 U13346 ( .A1(n11031), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n10679) );
  NAND2_X1 U13347 ( .A1(n11032), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n10678) );
  AOI22_X1 U13348 ( .A1(n14720), .A2(n14790), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n10706), .ZN(n10681) );
  OAI21_X1 U13349 ( .B1(n11138), .B2(n14715), .A(n10681), .ZN(n10682) );
  AOI21_X1 U13350 ( .B1(n14740), .B2(n10668), .A(n10682), .ZN(n10683) );
  OAI21_X1 U13351 ( .B1(n10684), .B2(n14742), .A(n10683), .ZN(P1_U3222) );
  OAI22_X1 U13352 ( .A1(n10688), .A2(n10687), .B1(n10686), .B2(n10685), .ZN(
        n10884) );
  INV_X1 U13353 ( .A(n10689), .ZN(n10690) );
  NAND2_X1 U13354 ( .A1(n11018), .A2(n10690), .ZN(n10697) );
  AND2_X1 U13355 ( .A1(n12325), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n10691) );
  OAI21_X1 U13356 ( .B1(n10692), .B2(n12912), .A(n10691), .ZN(n10693) );
  OAI21_X1 U13357 ( .B1(n12328), .B2(n10694), .A(n10693), .ZN(n10695) );
  INV_X1 U13358 ( .A(n10695), .ZN(n10696) );
  NAND2_X2 U13359 ( .A1(n10697), .A2(n10696), .ZN(n12691) );
  AOI22_X1 U13360 ( .A1(n6553), .A2(n12691), .B1(n14790), .B2(n12552), .ZN(
        n10698) );
  XNOR2_X1 U13361 ( .A(n10698), .B(n11860), .ZN(n10881) );
  INV_X1 U13362 ( .A(n14790), .ZN(n11353) );
  INV_X1 U13363 ( .A(n12691), .ZN(n15537) );
  XNOR2_X1 U13364 ( .A(n10881), .B(n10880), .ZN(n10883) );
  XOR2_X1 U13365 ( .A(n10884), .B(n10883), .Z(n10710) );
  OR2_X1 U13366 ( .A1(n11447), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10705) );
  INV_X1 U13367 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10701) );
  NAND2_X1 U13368 ( .A1(n10902), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n10702) );
  INV_X1 U13369 ( .A(n14715), .ZN(n14627) );
  AOI22_X1 U13370 ( .A1(n14627), .A2(n14792), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10706), .ZN(n10707) );
  OAI21_X1 U13371 ( .B1(n11153), .B2(n14706), .A(n10707), .ZN(n10708) );
  AOI21_X1 U13372 ( .B1(n14740), .B2(n12691), .A(n10708), .ZN(n10709) );
  OAI21_X1 U13373 ( .B1(n10710), .B2(n14742), .A(n10709), .ZN(P1_U3237) );
  AOI21_X1 U13374 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n13557), .A(n10711), .ZN(
        n10712) );
  MUX2_X1 U13375 ( .A(n10713), .B(n10712), .S(n13553), .Z(n10714) );
  OAI21_X1 U13376 ( .B1(n13456), .B2(n10715), .A(n10714), .ZN(P3_U3233) );
  INV_X1 U13377 ( .A(n10716), .ZN(n10717) );
  AOI211_X1 U13378 ( .C1(n10719), .C2(n10718), .A(n15624), .B(n10717), .ZN(
        n10728) );
  INV_X1 U13379 ( .A(n10720), .ZN(n10721) );
  AOI211_X1 U13380 ( .C1(n10723), .C2(n10722), .A(n15623), .B(n10721), .ZN(
        n10727) );
  INV_X1 U13381 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n11668) );
  NAND2_X1 U13382 ( .A1(n15651), .A2(n10724), .ZN(n10725) );
  NAND2_X1 U13383 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n12033)
         );
  OAI211_X1 U13384 ( .C1(n15658), .C2(n11668), .A(n10725), .B(n12033), .ZN(
        n10726) );
  OR3_X1 U13385 ( .A1(n10728), .A2(n10727), .A3(n10726), .ZN(P2_U3224) );
  XOR2_X1 U13386 ( .A(n10730), .B(n10729), .Z(n10741) );
  INV_X1 U13387 ( .A(n10980), .ZN(n10731) );
  AOI21_X1 U13388 ( .B1(n10809), .B2(n10732), .A(n10731), .ZN(n10737) );
  AOI22_X1 U13389 ( .A1(n15751), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n10736) );
  OAI21_X1 U13390 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(n10733), .A(n10986), .ZN(
        n10734) );
  NAND2_X1 U13391 ( .A1(n13313), .A2(n10734), .ZN(n10735) );
  OAI211_X1 U13392 ( .C1(n13283), .C2(n10737), .A(n10736), .B(n10735), .ZN(
        n10738) );
  AOI21_X1 U13393 ( .B1(n10739), .B2(n13323), .A(n10738), .ZN(n10740) );
  OAI21_X1 U13394 ( .B1(n10741), .B2(n13210), .A(n10740), .ZN(P3_U3185) );
  XOR2_X1 U13395 ( .A(n10743), .B(n10742), .Z(n10757) );
  AOI21_X1 U13396 ( .B1(n10746), .B2(n10745), .A(n10744), .ZN(n10753) );
  AOI22_X1 U13397 ( .A1(n15751), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10752) );
  OAI21_X1 U13398 ( .B1(n10749), .B2(n10748), .A(n10747), .ZN(n10750) );
  NAND2_X1 U13399 ( .A1(n13318), .A2(n10750), .ZN(n10751) );
  OAI211_X1 U13400 ( .C1(n13190), .C2(n10753), .A(n10752), .B(n10751), .ZN(
        n10754) );
  AOI21_X1 U13401 ( .B1(n10755), .B2(n13323), .A(n10754), .ZN(n10756) );
  OAI21_X1 U13402 ( .B1(n10757), .B2(n13210), .A(n10756), .ZN(P3_U3184) );
  XNOR2_X1 U13403 ( .A(n10758), .B(n10760), .ZN(n15756) );
  OAI21_X1 U13404 ( .B1(n10761), .B2(n10760), .A(n10804), .ZN(n10763) );
  OAI22_X1 U13405 ( .A1(n7429), .A2(n13533), .B1(n11006), .B2(n13535), .ZN(
        n10762) );
  AOI21_X1 U13406 ( .B1(n10763), .B2(n13552), .A(n10762), .ZN(n10764) );
  OAI21_X1 U13407 ( .B1(n15756), .B2(n13394), .A(n10764), .ZN(n15758) );
  NAND2_X1 U13408 ( .A1(n10765), .A2(n13598), .ZN(n15757) );
  OAI22_X1 U13409 ( .A1(n13479), .A2(n10767), .B1(n10766), .B2(n15757), .ZN(
        n10768) );
  NOR2_X1 U13410 ( .A1(n15758), .A2(n10768), .ZN(n10769) );
  MUX2_X1 U13411 ( .A(n10770), .B(n10769), .S(n13553), .Z(n10771) );
  OAI21_X1 U13412 ( .B1(n15756), .B2(n11912), .A(n10771), .ZN(P3_U3231) );
  INV_X1 U13413 ( .A(n10772), .ZN(n10777) );
  AOI21_X1 U13414 ( .B1(n10776), .B2(n10774), .A(n10773), .ZN(n10775) );
  AOI21_X1 U13415 ( .B1(n10777), .B2(n10776), .A(n10775), .ZN(n10787) );
  OAI21_X1 U13416 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n6756), .A(n10778), .ZN(
        n10780) );
  AOI22_X1 U13417 ( .A1(n10780), .A2(n13313), .B1(n10779), .B2(n13323), .ZN(
        n10786) );
  AND2_X1 U13418 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11277) );
  NAND2_X1 U13419 ( .A1(n10781), .A2(n15939), .ZN(n10782) );
  AOI21_X1 U13420 ( .B1(n10783), .B2(n10782), .A(n13283), .ZN(n10784) );
  AOI211_X1 U13421 ( .C1(n15751), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n11277), .B(
        n10784), .ZN(n10785) );
  OAI211_X1 U13422 ( .C1(n10787), .C2(n13210), .A(n10786), .B(n10785), .ZN(
        P3_U3187) );
  OAI21_X1 U13423 ( .B1(n10788), .B2(n10790), .A(n10789), .ZN(n10791) );
  INV_X1 U13424 ( .A(n10791), .ZN(n11632) );
  XNOR2_X1 U13425 ( .A(n10792), .B(n10793), .ZN(n10796) );
  NAND2_X1 U13426 ( .A1(n13953), .A2(n13907), .ZN(n10795) );
  NAND2_X1 U13427 ( .A1(n13955), .A2(n13905), .ZN(n10794) );
  NAND2_X1 U13428 ( .A1(n10795), .A2(n10794), .ZN(n10859) );
  AOI21_X1 U13429 ( .B1(n10796), .B2(n15662), .A(n10859), .ZN(n11628) );
  OAI211_X1 U13430 ( .C1(n11715), .C2(n11625), .A(n14470), .B(n11957), .ZN(
        n11622) );
  OAI211_X1 U13431 ( .C1(n11632), .C2(n14484), .A(n11628), .B(n11622), .ZN(
        n10816) );
  OAI22_X1 U13432 ( .A1(n14574), .A2(n11625), .B1(n15743), .B2(n8469), .ZN(
        n10797) );
  AOI21_X1 U13433 ( .B1(n10816), .B2(n15743), .A(n10797), .ZN(n10798) );
  INV_X1 U13434 ( .A(n10798), .ZN(P2_U3442) );
  XNOR2_X1 U13435 ( .A(n10800), .B(n10799), .ZN(n15764) );
  INV_X1 U13436 ( .A(n15764), .ZN(n10814) );
  INV_X1 U13437 ( .A(n13394), .ZN(n11425) );
  NAND2_X1 U13438 ( .A1(n10801), .A2(n13552), .ZN(n10807) );
  AOI21_X1 U13439 ( .B1(n10804), .B2(n10803), .A(n10802), .ZN(n10806) );
  AOI22_X1 U13440 ( .A1(n13549), .A2(n13120), .B1(n13119), .B2(n13547), .ZN(
        n10805) );
  OAI21_X1 U13441 ( .B1(n10807), .B2(n10806), .A(n10805), .ZN(n10808) );
  AOI21_X1 U13442 ( .B1(n15764), .B2(n11425), .A(n10808), .ZN(n15761) );
  MUX2_X1 U13443 ( .A(n10809), .B(n15761), .S(n13553), .Z(n10813) );
  NOR2_X1 U13444 ( .A1(n10810), .A2(n15770), .ZN(n15763) );
  AOI22_X1 U13445 ( .A1(n11429), .A2(n15763), .B1(n13557), .B2(n10811), .ZN(
        n10812) );
  OAI211_X1 U13446 ( .C1(n10814), .C2(n11912), .A(n10813), .B(n10812), .ZN(
        P3_U3230) );
  OAI22_X1 U13447 ( .A1(n14514), .A2(n11625), .B1(n15750), .B2(n8470), .ZN(
        n10815) );
  AOI21_X1 U13448 ( .B1(n10816), .B2(n15750), .A(n10815), .ZN(n10817) );
  INV_X1 U13449 ( .A(n10817), .ZN(P2_U3503) );
  XOR2_X1 U13450 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n12008), .Z(n10820) );
  OAI21_X1 U13451 ( .B1(n10820), .B2(n10819), .A(n11118), .ZN(n10831) );
  INV_X1 U13452 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11115) );
  MUX2_X1 U13453 ( .A(n11115), .B(P1_REG2_REG_11__SCAN_IN), .S(n12008), .Z(
        n10823) );
  NAND2_X1 U13454 ( .A1(n6748), .A2(n10823), .ZN(n10825) );
  MUX2_X1 U13455 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n11115), .S(n12008), .Z(
        n10824) );
  OAI211_X1 U13456 ( .C1(n10826), .C2(n10825), .A(n11113), .B(n15812), .ZN(
        n10829) );
  NAND2_X1 U13457 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n12144)
         );
  INV_X1 U13458 ( .A(n12144), .ZN(n10827) );
  AOI21_X1 U13459 ( .B1(n15475), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n10827), 
        .ZN(n10828) );
  OAI211_X1 U13460 ( .C1(n15814), .C2(n11114), .A(n10829), .B(n10828), .ZN(
        n10830) );
  AOI21_X1 U13461 ( .B1(n10831), .B2(n15486), .A(n10830), .ZN(n10832) );
  INV_X1 U13462 ( .A(n10832), .ZN(P1_U3254) );
  NAND2_X1 U13463 ( .A1(n10840), .A2(n14352), .ZN(n10833) );
  NAND2_X1 U13464 ( .A1(n10834), .A2(n10833), .ZN(n10872) );
  INV_X1 U13465 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10835) );
  MUX2_X1 U13466 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n10835), .S(n10876), .Z(
        n10871) );
  NAND2_X1 U13467 ( .A1(n10843), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10836) );
  NAND2_X1 U13468 ( .A1(n10869), .A2(n10836), .ZN(n11286) );
  XNOR2_X1 U13469 ( .A(n11286), .B(n10837), .ZN(n11285) );
  XNOR2_X1 U13470 ( .A(n11285), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n10850) );
  NOR2_X1 U13471 ( .A1(n15922), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13761) );
  NOR2_X1 U13472 ( .A1(n14082), .A2(n10837), .ZN(n10838) );
  AOI211_X1 U13473 ( .C1(P2_ADDR_REG_14__SCAN_IN), .C2(n15629), .A(n13761), 
        .B(n10838), .ZN(n10849) );
  NAND2_X1 U13474 ( .A1(n10840), .A2(n10839), .ZN(n10841) );
  XNOR2_X1 U13475 ( .A(n10876), .B(n14489), .ZN(n10868) );
  NAND2_X1 U13476 ( .A1(n10843), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10844) );
  XNOR2_X1 U13477 ( .A(n11292), .B(n10845), .ZN(n10846) );
  NAND2_X1 U13478 ( .A1(n10847), .A2(n10846), .ZN(n11294) );
  OAI211_X1 U13479 ( .C1(n10847), .C2(n10846), .A(n11294), .B(n15644), .ZN(
        n10848) );
  OAI211_X1 U13480 ( .C1(n10850), .C2(n15623), .A(n10849), .B(n10848), .ZN(
        P2_U3228) );
  XNOR2_X1 U13481 ( .A(n13789), .B(n10851), .ZN(n11220) );
  AND2_X1 U13482 ( .A1(n13954), .A2(n6556), .ZN(n11221) );
  XNOR2_X1 U13483 ( .A(n11220), .B(n11221), .ZN(n10858) );
  INV_X1 U13484 ( .A(n10857), .ZN(n10855) );
  INV_X1 U13485 ( .A(n11228), .ZN(n10856) );
  AOI21_X1 U13486 ( .B1(n10858), .B2(n10857), .A(n10856), .ZN(n10864) );
  INV_X1 U13487 ( .A(n11624), .ZN(n10862) );
  AOI22_X1 U13488 ( .A1(n13919), .A2(n10859), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10860) );
  OAI21_X1 U13489 ( .B1(n11625), .B2(n13912), .A(n10860), .ZN(n10861) );
  AOI21_X1 U13490 ( .B1(n10862), .B2(n13859), .A(n10861), .ZN(n10863) );
  OAI21_X1 U13491 ( .B1(n10864), .B2(n13925), .A(n10863), .ZN(P2_U3202) );
  INV_X1 U13492 ( .A(n10865), .ZN(n10866) );
  AOI211_X1 U13493 ( .C1(n10868), .C2(n10867), .A(n15624), .B(n10866), .ZN(
        n10879) );
  INV_X1 U13494 ( .A(n10869), .ZN(n10870) );
  AOI211_X1 U13495 ( .C1(n10872), .C2(n10871), .A(n15623), .B(n10870), .ZN(
        n10878) );
  NOR2_X1 U13496 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10873), .ZN(n10874) );
  AOI21_X1 U13497 ( .B1(n15629), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n10874), 
        .ZN(n10875) );
  OAI21_X1 U13498 ( .B1(n10876), .B2(n14082), .A(n10875), .ZN(n10877) );
  OR3_X1 U13499 ( .A1(n10879), .A2(n10878), .A3(n10877), .ZN(P2_U3227) );
  INV_X1 U13500 ( .A(n10880), .ZN(n10882) );
  AOI21_X2 U13501 ( .B1(n10884), .B2(n10883), .A(n6629), .ZN(n14622) );
  NAND2_X1 U13502 ( .A1(n11018), .A2(n10886), .ZN(n10889) );
  INV_X1 U13503 ( .A(n14828), .ZN(n10887) );
  OAI22_X1 U13504 ( .A1(n14636), .A2(n11153), .B1(n15548), .B2(n12463), .ZN(
        n10893) );
  OAI22_X1 U13505 ( .A1(n11153), .A2(n12463), .B1(n15548), .B2(n14638), .ZN(
        n10891) );
  XNOR2_X1 U13506 ( .A(n10891), .B(n11860), .ZN(n10892) );
  XOR2_X1 U13507 ( .A(n10893), .B(n10892), .Z(n14621) );
  NAND2_X1 U13508 ( .A1(n14622), .A2(n14621), .ZN(n11017) );
  INV_X1 U13509 ( .A(n14620), .ZN(n10896) );
  INV_X1 U13510 ( .A(n10892), .ZN(n10895) );
  INV_X1 U13511 ( .A(n10893), .ZN(n10894) );
  NOR2_X1 U13512 ( .A1(n10895), .A2(n10894), .ZN(n11011) );
  NOR2_X1 U13513 ( .A1(n10896), .A2(n11011), .ZN(n10914) );
  AOI22_X1 U13514 ( .A1(n12855), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n12294), 
        .B2(n10898), .ZN(n10901) );
  NAND2_X1 U13515 ( .A1(n10899), .A2(n12393), .ZN(n10900) );
  NAND2_X1 U13516 ( .A1(n6553), .A2(n12699), .ZN(n10908) );
  NAND2_X1 U13517 ( .A1(n10902), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10906) );
  OAI21_X1 U13518 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n10921), .ZN(n11340) );
  OR2_X1 U13519 ( .A1(n11447), .A2(n11340), .ZN(n10905) );
  NAND2_X1 U13520 ( .A1(n11451), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10904) );
  NAND2_X1 U13521 ( .A1(n12410), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n10903) );
  NAND2_X1 U13522 ( .A1(n14788), .A2(n12552), .ZN(n10907) );
  NAND2_X1 U13523 ( .A1(n10908), .A2(n10907), .ZN(n10909) );
  XNOR2_X1 U13524 ( .A(n10909), .B(n11860), .ZN(n11012) );
  NAND2_X1 U13525 ( .A1(n12572), .A2(n14788), .ZN(n10912) );
  NAND2_X1 U13526 ( .A1(n6554), .A2(n12699), .ZN(n10911) );
  NAND2_X1 U13527 ( .A1(n10912), .A2(n10911), .ZN(n11013) );
  XNOR2_X1 U13528 ( .A(n11012), .B(n11013), .ZN(n10913) );
  XNOR2_X1 U13529 ( .A(n10914), .B(n10913), .ZN(n10934) );
  INV_X1 U13530 ( .A(n11340), .ZN(n10931) );
  INV_X1 U13531 ( .A(n10915), .ZN(n10916) );
  NAND2_X1 U13532 ( .A1(n10917), .A2(n10916), .ZN(n10918) );
  NAND2_X1 U13533 ( .A1(n14789), .A2(n15180), .ZN(n10928) );
  NAND2_X1 U13534 ( .A1(n11451), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n10926) );
  INV_X1 U13535 ( .A(n10921), .ZN(n10919) );
  INV_X1 U13536 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10920) );
  NAND2_X1 U13537 ( .A1(n10921), .A2(n10920), .ZN(n10922) );
  NAND2_X1 U13538 ( .A1(n11029), .A2(n10922), .ZN(n11167) );
  OR2_X1 U13539 ( .A1(n11447), .A2(n11167), .ZN(n10925) );
  NAND2_X1 U13540 ( .A1(n10902), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10924) );
  NAND2_X1 U13541 ( .A1(n11032), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n10923) );
  NAND2_X1 U13542 ( .A1(n14787), .A2(n15178), .ZN(n10927) );
  AND2_X1 U13543 ( .A1(n10928), .A2(n10927), .ZN(n11339) );
  OAI21_X1 U13544 ( .B1(n14737), .B2(n11339), .A(n10929), .ZN(n10930) );
  AOI21_X1 U13545 ( .B1(n10931), .B2(n14690), .A(n10930), .ZN(n10933) );
  AND2_X1 U13546 ( .A1(n15530), .A2(n12699), .ZN(n15554) );
  NAND2_X1 U13547 ( .A1(n11042), .A2(n15554), .ZN(n10932) );
  OAI211_X1 U13548 ( .C1(n10934), .C2(n14742), .A(n10933), .B(n10932), .ZN(
        P1_U3230) );
  INV_X1 U13549 ( .A(n10936), .ZN(n10937) );
  OR2_X1 U13550 ( .A1(n10938), .A2(n10937), .ZN(n10939) );
  NAND2_X1 U13551 ( .A1(n10941), .A2(n10940), .ZN(n10943) );
  XNOR2_X1 U13552 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10944) );
  XNOR2_X1 U13553 ( .A(n11304), .B(n10944), .ZN(n10945) );
  NAND2_X1 U13554 ( .A1(n10946), .A2(n10945), .ZN(n11302) );
  NAND2_X1 U13555 ( .A1(n11301), .A2(n11302), .ZN(n10947) );
  XNOR2_X1 U13556 ( .A(n10947), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(SUB_1596_U54)
         );
  INV_X1 U13557 ( .A(n10965), .ZN(n10963) );
  AOI21_X1 U13558 ( .B1(n15802), .B2(n10951), .A(n6739), .ZN(n10974) );
  OR2_X1 U13559 ( .A1(n10952), .A2(n16060), .ZN(n10953) );
  NAND2_X1 U13560 ( .A1(n10954), .A2(n10953), .ZN(n10955) );
  NAND2_X1 U13561 ( .A1(n10956), .A2(n11426), .ZN(n10957) );
  NAND2_X1 U13562 ( .A1(n11074), .A2(n10957), .ZN(n10958) );
  NAND2_X1 U13563 ( .A1(n10958), .A2(n13318), .ZN(n10960) );
  AND2_X1 U13564 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11465) );
  AOI21_X1 U13565 ( .B1(n15751), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11465), .ZN(
        n10959) );
  OAI211_X1 U13566 ( .C1(n13295), .C2(n10965), .A(n10960), .B(n10959), .ZN(
        n10961) );
  INV_X1 U13567 ( .A(n10961), .ZN(n10973) );
  INV_X1 U13568 ( .A(n10962), .ZN(n10969) );
  MUX2_X1 U13569 ( .A(n11426), .B(n15802), .S(n13724), .Z(n10964) );
  NAND2_X1 U13570 ( .A1(n10963), .A2(n10964), .ZN(n11069) );
  INV_X1 U13571 ( .A(n10964), .ZN(n10966) );
  NAND2_X1 U13572 ( .A1(n10966), .A2(n10965), .ZN(n10967) );
  AND2_X1 U13573 ( .A1(n11069), .A2(n10967), .ZN(n10968) );
  NOR3_X1 U13574 ( .A1(n10970), .A2(n10969), .A3(n10968), .ZN(n10971) );
  OAI21_X1 U13575 ( .B1(n6749), .B2(n10971), .A(n13332), .ZN(n10972) );
  OAI211_X1 U13576 ( .C1(n10974), .C2(n13190), .A(n10973), .B(n10972), .ZN(
        P3_U3189) );
  XNOR2_X1 U13577 ( .A(n10976), .B(n10975), .ZN(n10993) );
  AND2_X1 U13578 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n11008) );
  INV_X1 U13579 ( .A(n10977), .ZN(n10979) );
  NAND3_X1 U13580 ( .A1(n10980), .A2(n10979), .A3(n10978), .ZN(n10981) );
  AOI21_X1 U13581 ( .B1(n10982), .B2(n10981), .A(n13283), .ZN(n10983) );
  AOI211_X1 U13582 ( .C1(n15751), .C2(P3_ADDR_REG_4__SCAN_IN), .A(n11008), .B(
        n10983), .ZN(n10990) );
  AND3_X1 U13583 ( .A1(n10986), .A2(n10985), .A3(n10984), .ZN(n10987) );
  OAI21_X1 U13584 ( .B1(n10988), .B2(n10987), .A(n13313), .ZN(n10989) );
  OAI211_X1 U13585 ( .C1(n13295), .C2(n10991), .A(n10990), .B(n10989), .ZN(
        n10992) );
  AOI21_X1 U13586 ( .B1(n13332), .B2(n10993), .A(n10992), .ZN(n10994) );
  INV_X1 U13587 ( .A(n10994), .ZN(P3_U3186) );
  INV_X1 U13588 ( .A(n13095), .ZN(n11764) );
  INV_X1 U13589 ( .A(n10995), .ZN(n10996) );
  NAND2_X1 U13590 ( .A1(n10996), .A2(n11241), .ZN(n10997) );
  AND2_X2 U13591 ( .A1(n10998), .A2(n10997), .ZN(n11004) );
  XNOR2_X1 U13592 ( .A(n12947), .B(n10999), .ZN(n11000) );
  NAND2_X1 U13593 ( .A1(n11000), .A2(n11275), .ZN(n11270) );
  INV_X1 U13594 ( .A(n11000), .ZN(n11001) );
  NAND2_X1 U13595 ( .A1(n11001), .A2(n13119), .ZN(n11002) );
  AND2_X1 U13596 ( .A1(n11270), .A2(n11002), .ZN(n11003) );
  OAI21_X1 U13597 ( .B1(n11004), .B2(n11003), .A(n11271), .ZN(n11005) );
  NAND2_X1 U13598 ( .A1(n11005), .A2(n11608), .ZN(n11010) );
  OAI22_X1 U13599 ( .A1(n13081), .A2(n11236), .B1(n11006), .B2(n13099), .ZN(
        n11007) );
  AOI211_X1 U13600 ( .C1(n13096), .C2(n13118), .A(n11008), .B(n11007), .ZN(
        n11009) );
  OAI211_X1 U13601 ( .C1(n11237), .C2(n11764), .A(n11010), .B(n11009), .ZN(
        P3_U3170) );
  AOI21_X1 U13602 ( .B1(n11012), .B2(n11013), .A(n11011), .ZN(n11016) );
  INV_X1 U13603 ( .A(n11012), .ZN(n11015) );
  INV_X1 U13604 ( .A(n11013), .ZN(n11014) );
  BUF_X4 U13605 ( .A(n11018), .Z(n12393) );
  NAND2_X1 U13606 ( .A1(n11019), .A2(n12393), .ZN(n11022) );
  AOI22_X1 U13607 ( .A1(n12855), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n12294), 
        .B2(n11020), .ZN(n11021) );
  NAND2_X1 U13608 ( .A1(n11022), .A2(n11021), .ZN(n12708) );
  AOI22_X1 U13609 ( .A1(n12708), .A2(n6553), .B1(n14787), .B2(n12552), .ZN(
        n11023) );
  XOR2_X1 U13610 ( .A(n11860), .B(n11023), .Z(n11323) );
  NAND2_X1 U13611 ( .A1(n12572), .A2(n14787), .ZN(n11025) );
  NAND2_X1 U13612 ( .A1(n12708), .A2(n12552), .ZN(n11024) );
  NAND2_X1 U13613 ( .A1(n11025), .A2(n11024), .ZN(n11324) );
  XNOR2_X1 U13614 ( .A(n11323), .B(n7134), .ZN(n11026) );
  XNOR2_X1 U13615 ( .A(n11325), .B(n11026), .ZN(n11045) );
  INV_X1 U13616 ( .A(n11167), .ZN(n11041) );
  NAND2_X1 U13617 ( .A1(n14788), .A2(n15180), .ZN(n11038) );
  INV_X2 U13618 ( .A(n12161), .ZN(n12448) );
  NAND2_X1 U13619 ( .A1(n12448), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n11036) );
  INV_X1 U13620 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n11028) );
  NAND2_X1 U13621 ( .A1(n11029), .A2(n11028), .ZN(n11030) );
  NAND2_X1 U13622 ( .A1(n11199), .A2(n11030), .ZN(n11329) );
  OR2_X1 U13623 ( .A1(n11447), .A2(n11329), .ZN(n11035) );
  NAND2_X1 U13624 ( .A1(n11451), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n11034) );
  NAND2_X1 U13625 ( .A1(n12410), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n11033) );
  NAND2_X1 U13626 ( .A1(n14786), .A2(n15178), .ZN(n11037) );
  AND2_X1 U13627 ( .A1(n11038), .A2(n11037), .ZN(n11163) );
  OAI21_X1 U13628 ( .B1(n14737), .B2(n11163), .A(n11039), .ZN(n11040) );
  AOI21_X1 U13629 ( .B1(n11041), .B2(n14690), .A(n11040), .ZN(n11044) );
  AND2_X1 U13630 ( .A1(n12708), .A2(n15530), .ZN(n15568) );
  NAND2_X1 U13631 ( .A1(n11042), .A2(n15568), .ZN(n11043) );
  OAI211_X1 U13632 ( .C1(n11045), .C2(n14742), .A(n11044), .B(n11043), .ZN(
        P1_U3227) );
  NOR2_X1 U13633 ( .A1(n11046), .A2(n15770), .ZN(n15753) );
  OAI21_X1 U13634 ( .B1(n11056), .B2(n11048), .A(n11047), .ZN(n11049) );
  NAND2_X1 U13635 ( .A1(n11049), .A2(n13552), .ZN(n11051) );
  AOI22_X1 U13636 ( .A1(n13547), .A2(n13120), .B1(n13122), .B2(n13549), .ZN(
        n11050) );
  NAND2_X1 U13637 ( .A1(n11051), .A2(n11050), .ZN(n15752) );
  AOI21_X1 U13638 ( .B1(n15753), .B2(n11052), .A(n15752), .ZN(n11053) );
  MUX2_X1 U13639 ( .A(n11054), .B(n11053), .S(n13553), .Z(n11058) );
  INV_X1 U13640 ( .A(n13561), .ZN(n13360) );
  XNOR2_X1 U13641 ( .A(n11056), .B(n11055), .ZN(n15754) );
  AOI22_X1 U13642 ( .A1(n13360), .A2(n15754), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n13557), .ZN(n11057) );
  NAND2_X1 U13643 ( .A1(n11058), .A2(n11057), .ZN(P3_U3232) );
  NOR3_X1 U13644 ( .A1(n13313), .A2(n13318), .A3(n13332), .ZN(n11068) );
  INV_X1 U13645 ( .A(n11059), .ZN(n11060) );
  AOI22_X1 U13646 ( .A1(n13318), .A2(P3_REG2_REG_0__SCAN_IN), .B1(n11060), 
        .B2(n13332), .ZN(n11061) );
  MUX2_X1 U13647 ( .A(n11061), .B(n13295), .S(P3_IR_REG_0__SCAN_IN), .Z(n11067) );
  INV_X1 U13648 ( .A(n15751), .ZN(n13321) );
  OAI22_X1 U13649 ( .A1(n13321), .A2(n11063), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11062), .ZN(n11064) );
  AOI21_X1 U13650 ( .B1(n11065), .B2(n13313), .A(n11064), .ZN(n11066) );
  OAI211_X1 U13651 ( .C1(n11068), .C2(n11094), .A(n11067), .B(n11066), .ZN(
        P3_U3182) );
  MUX2_X1 U13652 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13724), .Z(n11554) );
  XNOR2_X1 U13653 ( .A(n11560), .B(n11554), .ZN(n11070) );
  OAI21_X1 U13654 ( .B1(n11071), .B2(n11070), .A(n11553), .ZN(n11084) );
  XNOR2_X1 U13655 ( .A(n11568), .B(P3_REG2_REG_8__SCAN_IN), .ZN(n11073) );
  AND3_X1 U13656 ( .A1(n11074), .A2(n11073), .A3(n11072), .ZN(n11075) );
  OAI21_X1 U13657 ( .B1(n11567), .B2(n11075), .A(n13318), .ZN(n11078) );
  NAND2_X1 U13658 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n11760) );
  INV_X1 U13659 ( .A(n11760), .ZN(n11076) );
  AOI21_X1 U13660 ( .B1(n15751), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11076), .ZN(
        n11077) );
  OAI211_X1 U13661 ( .C1(n13295), .C2(n11568), .A(n11078), .B(n11077), .ZN(
        n11083) );
  XNOR2_X1 U13662 ( .A(n11568), .B(n11559), .ZN(n11079) );
  OR3_X1 U13663 ( .A1(n11080), .A2(n6739), .A3(n11079), .ZN(n11081) );
  AOI21_X1 U13664 ( .B1(n11558), .B2(n11081), .A(n13190), .ZN(n11082) );
  AOI211_X1 U13665 ( .C1(n13332), .C2(n11084), .A(n11083), .B(n11082), .ZN(
        n11085) );
  INV_X1 U13666 ( .A(n11085), .ZN(P3_U3190) );
  INV_X1 U13667 ( .A(n11086), .ZN(n11088) );
  OAI21_X1 U13668 ( .B1(n11088), .B2(P3_REG2_REG_1__SCAN_IN), .A(n11087), .ZN(
        n11100) );
  OAI22_X1 U13669 ( .A1(n13321), .A2(n11090), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11089), .ZN(n11099) );
  AOI21_X1 U13670 ( .B1(n15789), .B2(n11092), .A(n11091), .ZN(n11097) );
  AOI21_X1 U13671 ( .B1(n11095), .B2(n11094), .A(n11093), .ZN(n11096) );
  OAI22_X1 U13672 ( .A1(n13190), .A2(n11097), .B1(n11096), .B2(n13210), .ZN(
        n11098) );
  AOI211_X1 U13673 ( .C1(n13318), .C2(n11100), .A(n11099), .B(n11098), .ZN(
        n11101) );
  OAI21_X1 U13674 ( .B1(n11102), .B2(n13295), .A(n11101), .ZN(P3_U3183) );
  INV_X1 U13675 ( .A(n14067), .ZN(n14062) );
  INV_X1 U13676 ( .A(n12282), .ZN(n11108) );
  OAI222_X1 U13677 ( .A1(P2_U3088), .A2(n14062), .B1(n11897), .B2(n11108), 
        .C1(n15896), .C2(n14590), .ZN(P2_U3309) );
  NAND2_X1 U13678 ( .A1(n11103), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11104) );
  MUX2_X1 U13679 ( .A(P1_IR_REG_31__SCAN_IN), .B(n11104), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n11106) );
  AND2_X1 U13680 ( .A1(n11106), .A2(n11105), .ZN(n15808) );
  INV_X1 U13681 ( .A(n15808), .ZN(n14911) );
  OAI222_X1 U13682 ( .A1(P1_U3086), .A2(n14911), .B1(n15379), .B2(n11108), 
        .C1(n11107), .C2(n15370), .ZN(P1_U3337) );
  INV_X1 U13683 ( .A(n11109), .ZN(n11112) );
  OAI22_X1 U13684 ( .A1(n11110), .A2(P3_U3151), .B1(SI_22_), .B2(n13723), .ZN(
        n11111) );
  AOI21_X1 U13685 ( .B1(n11112), .B2(n13709), .A(n11111), .ZN(P3_U3273) );
  INV_X1 U13686 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n12097) );
  MUX2_X1 U13687 ( .A(n12097), .B(P1_REG2_REG_12__SCAN_IN), .S(n12071), .Z(
        n11117) );
  AOI21_X1 U13688 ( .B1(n11117), .B2(n11116), .A(n11482), .ZN(n11125) );
  XOR2_X1 U13689 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n12071), .Z(n11120) );
  OAI21_X1 U13690 ( .B1(n11120), .B2(n11119), .A(n11477), .ZN(n11121) );
  NAND2_X1 U13691 ( .A1(n11121), .A2(n15486), .ZN(n11124) );
  INV_X1 U13692 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n12197) );
  NAND2_X1 U13693 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n12233)
         );
  OAI21_X1 U13694 ( .B1(n15821), .B2(n12197), .A(n12233), .ZN(n11122) );
  AOI21_X1 U13695 ( .B1(n12071), .B2(n15483), .A(n11122), .ZN(n11123) );
  OAI211_X1 U13696 ( .C1(n11125), .C2(n15815), .A(n11124), .B(n11123), .ZN(
        P1_U3255) );
  NAND2_X1 U13697 ( .A1(n10356), .A2(n6937), .ZN(n11148) );
  NAND2_X2 U13698 ( .A1(n12688), .A2(n12687), .ZN(n12870) );
  XOR2_X1 U13699 ( .A(n12870), .B(n11148), .Z(n15528) );
  AND2_X1 U13700 ( .A1(n12913), .A2(n15202), .ZN(n11129) );
  INV_X1 U13701 ( .A(n11127), .ZN(n11128) );
  NAND2_X1 U13702 ( .A1(n11129), .A2(n11128), .ZN(n12452) );
  OR2_X1 U13703 ( .A1(n11132), .A2(n15819), .ZN(n12861) );
  OR2_X1 U13704 ( .A1(n15525), .A2(n12861), .ZN(n15500) );
  NAND2_X1 U13705 ( .A1(n11133), .A2(n11317), .ZN(n11172) );
  OAI21_X1 U13706 ( .B1(n11133), .B2(n11317), .A(n11172), .ZN(n15533) );
  XNOR2_X1 U13707 ( .A(n11134), .B(n15533), .ZN(n11136) );
  INV_X1 U13708 ( .A(n12870), .ZN(n11135) );
  MUX2_X1 U13709 ( .A(n11136), .B(n11135), .S(n10356), .Z(n11137) );
  OAI222_X1 U13710 ( .A1(n15128), .A2(n11138), .B1(n15566), .B2(n15528), .C1(
        n11137), .C2(n15558), .ZN(n15534) );
  AND2_X1 U13711 ( .A1(n14790), .A2(n15178), .ZN(n15529) );
  NOR2_X1 U13712 ( .A1(n15534), .A2(n15529), .ZN(n11139) );
  MUX2_X1 U13713 ( .A(n11140), .B(n11139), .S(n15097), .Z(n11144) );
  NAND2_X1 U13714 ( .A1(n12917), .A2(n12675), .ZN(n12907) );
  OR2_X1 U13715 ( .A1(n12907), .A2(n15381), .ZN(n11141) );
  OR2_X1 U13716 ( .A1(n12452), .A2(n12672), .ZN(n15082) );
  NAND2_X1 U13717 ( .A1(n15521), .A2(n15517), .ZN(n15056) );
  INV_X1 U13718 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14793) );
  OAI22_X1 U13719 ( .A1(n15056), .A2(n15533), .B1(n14793), .B2(n15189), .ZN(
        n11142) );
  AOI21_X1 U13720 ( .B1(n15515), .B2(n10668), .A(n11142), .ZN(n11143) );
  OAI211_X1 U13721 ( .C1(n15528), .C2(n15500), .A(n11144), .B(n11143), .ZN(
        P1_U3292) );
  INV_X1 U13722 ( .A(n12293), .ZN(n11146) );
  OAI222_X1 U13723 ( .A1(n15370), .A2(n11145), .B1(n15379), .B2(n11146), .C1(
        P1_U3086), .C2(n15819), .ZN(P1_U3336) );
  OAI222_X1 U13724 ( .A1(n14590), .A2(n15836), .B1(n11897), .B2(n11146), .C1(
        n14086), .C2(P2_U3088), .ZN(P2_U3308) );
  OR2_X1 U13725 ( .A1(n15525), .A2(n15566), .ZN(n11147) );
  XNOR2_X1 U13726 ( .A(n11195), .B(n11186), .ZN(n11193) );
  NAND2_X1 U13727 ( .A1(n12870), .A2(n11148), .ZN(n11150) );
  XNOR2_X2 U13728 ( .A(n14790), .B(n12691), .ZN(n12871) );
  INV_X1 U13729 ( .A(n12871), .ZN(n11171) );
  OR2_X1 U13730 ( .A1(n14790), .A2(n12691), .ZN(n11151) );
  NAND2_X1 U13731 ( .A1(n14789), .A2(n15548), .ZN(n12697) );
  INV_X1 U13732 ( .A(n12874), .ZN(n12695) );
  NAND2_X1 U13733 ( .A1(n11348), .A2(n12695), .ZN(n11155) );
  NAND2_X1 U13734 ( .A1(n11153), .A2(n15548), .ZN(n11154) );
  NAND2_X1 U13735 ( .A1(n11345), .A2(n11344), .ZN(n11157) );
  INV_X1 U13736 ( .A(n14788), .ZN(n11352) );
  NAND2_X1 U13737 ( .A1(n11352), .A2(n7470), .ZN(n11156) );
  XNOR2_X1 U13738 ( .A(n11193), .B(n11185), .ZN(n15564) );
  INV_X1 U13739 ( .A(n11193), .ZN(n12875) );
  OR2_X1 U13740 ( .A1(n14790), .A2(n15537), .ZN(n11158) );
  NAND2_X1 U13741 ( .A1(n11159), .A2(n11158), .ZN(n11356) );
  NAND2_X1 U13742 ( .A1(n11160), .A2(n12696), .ZN(n11336) );
  NAND2_X1 U13743 ( .A1(n11336), .A2(n12872), .ZN(n11162) );
  NAND2_X1 U13744 ( .A1(n11352), .A2(n12699), .ZN(n11161) );
  NAND2_X1 U13745 ( .A1(n11162), .A2(n11161), .ZN(n11194) );
  XNOR2_X1 U13746 ( .A(n12875), .B(n11194), .ZN(n11164) );
  OAI21_X1 U13747 ( .B1(n11164), .B2(n15558), .A(n11163), .ZN(n15569) );
  INV_X1 U13748 ( .A(n15569), .ZN(n11165) );
  MUX2_X1 U13749 ( .A(n10243), .B(n11165), .S(n15097), .Z(n11170) );
  INV_X1 U13750 ( .A(n11210), .ZN(n11166) );
  AOI211_X1 U13751 ( .C1(n12708), .C2(n11337), .A(n15538), .B(n11166), .ZN(
        n15567) );
  OAI22_X1 U13752 ( .A1(n15147), .A2(n11186), .B1(n11167), .B2(n15189), .ZN(
        n11168) );
  AOI21_X1 U13753 ( .B1(n15567), .B2(n15521), .A(n11168), .ZN(n11169) );
  OAI211_X1 U13754 ( .C1(n15122), .C2(n15564), .A(n11170), .B(n11169), .ZN(
        P1_U3288) );
  INV_X1 U13755 ( .A(n15542), .ZN(n11184) );
  AND2_X1 U13756 ( .A1(n11172), .A2(n12691), .ZN(n11173) );
  OR2_X1 U13757 ( .A1(n11173), .A2(n11349), .ZN(n15539) );
  INV_X1 U13758 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n15940) );
  OAI22_X1 U13759 ( .A1(n15056), .A2(n15539), .B1(n15940), .B2(n15189), .ZN(
        n11174) );
  AOI21_X1 U13760 ( .B1(n15515), .B2(n12691), .A(n11174), .ZN(n11183) );
  XNOR2_X1 U13761 ( .A(n12871), .B(n11175), .ZN(n11178) );
  NAND2_X1 U13762 ( .A1(n14792), .A2(n15180), .ZN(n11176) );
  OAI21_X1 U13763 ( .B1(n11153), .B2(n15130), .A(n11176), .ZN(n11177) );
  AOI21_X1 U13764 ( .B1(n11178), .B2(n15552), .A(n11177), .ZN(n11180) );
  INV_X1 U13765 ( .A(n15566), .ZN(n15576) );
  NAND2_X1 U13766 ( .A1(n15542), .A2(n15576), .ZN(n11179) );
  NAND2_X1 U13767 ( .A1(n11180), .A2(n11179), .ZN(n15540) );
  MUX2_X1 U13768 ( .A(n15540), .B(P1_REG2_REG_2__SCAN_IN), .S(n15525), .Z(
        n11181) );
  INV_X1 U13769 ( .A(n11181), .ZN(n11182) );
  OAI211_X1 U13770 ( .C1(n11184), .C2(n15500), .A(n11183), .B(n11182), .ZN(
        P1_U3291) );
  NAND2_X1 U13771 ( .A1(n11185), .A2(n12875), .ZN(n11188) );
  NAND2_X1 U13772 ( .A1(n11186), .A2(n11195), .ZN(n11187) );
  NAND2_X1 U13773 ( .A1(n11188), .A2(n11187), .ZN(n11506) );
  NAND2_X1 U13774 ( .A1(n11189), .A2(n12393), .ZN(n11192) );
  AOI22_X1 U13775 ( .A1(n12855), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n12294), 
        .B2(n11190), .ZN(n11191) );
  INV_X1 U13776 ( .A(n12877), .ZN(n11505) );
  XNOR2_X1 U13777 ( .A(n11506), .B(n11505), .ZN(n15575) );
  INV_X1 U13778 ( .A(n15575), .ZN(n11216) );
  NAND2_X1 U13779 ( .A1(n11194), .A2(n11193), .ZN(n11197) );
  NAND2_X1 U13780 ( .A1(n11195), .A2(n12708), .ZN(n11196) );
  NAND2_X1 U13781 ( .A1(n11197), .A2(n11196), .ZN(n11540) );
  XNOR2_X1 U13782 ( .A(n11540), .B(n12877), .ZN(n11208) );
  NAND2_X1 U13783 ( .A1(n14787), .A2(n15180), .ZN(n11206) );
  NAND2_X1 U13784 ( .A1(n11451), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n11204) );
  NAND2_X1 U13785 ( .A1(n11199), .A2(n11198), .ZN(n11200) );
  NAND2_X1 U13786 ( .A1(n11449), .A2(n11200), .ZN(n11446) );
  OR2_X1 U13787 ( .A1(n11447), .A2(n11446), .ZN(n11203) );
  NAND2_X1 U13788 ( .A1(n12448), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n11202) );
  NAND2_X1 U13789 ( .A1(n12410), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n11201) );
  NAND4_X1 U13790 ( .A1(n11204), .A2(n11203), .A3(n11202), .A4(n11201), .ZN(
        n14785) );
  NAND2_X1 U13791 ( .A1(n14785), .A2(n15178), .ZN(n11205) );
  AND2_X1 U13792 ( .A1(n11206), .A2(n11205), .ZN(n11330) );
  INV_X1 U13793 ( .A(n11330), .ZN(n11207) );
  AOI21_X1 U13794 ( .B1(n11208), .B2(n15552), .A(n11207), .ZN(n15579) );
  INV_X1 U13795 ( .A(n15525), .ZN(n15097) );
  MUX2_X1 U13796 ( .A(n10270), .B(n15579), .S(n15097), .Z(n11215) );
  NAND2_X1 U13797 ( .A1(n11210), .A2(n12712), .ZN(n11209) );
  NAND2_X1 U13798 ( .A1(n11209), .A2(n15517), .ZN(n11211) );
  OR2_X1 U13799 ( .A1(n11211), .A2(n15519), .ZN(n15572) );
  INV_X1 U13800 ( .A(n15572), .ZN(n11213) );
  INV_X1 U13801 ( .A(n12712), .ZN(n15573) );
  OAI22_X1 U13802 ( .A1(n15147), .A2(n15573), .B1(n11329), .B2(n15189), .ZN(
        n11212) );
  AOI21_X1 U13803 ( .B1(n15521), .B2(n11213), .A(n11212), .ZN(n11214) );
  OAI211_X1 U13804 ( .C1(n15122), .C2(n11216), .A(n11215), .B(n11214), .ZN(
        P1_U3287) );
  INV_X1 U13805 ( .A(n11956), .ZN(n11232) );
  NAND2_X1 U13806 ( .A1(n13952), .A2(n13907), .ZN(n11218) );
  NAND2_X1 U13807 ( .A1(n13954), .A2(n13905), .ZN(n11217) );
  NAND2_X1 U13808 ( .A1(n11218), .A2(n11217), .ZN(n11963) );
  AOI22_X1 U13809 ( .A1(n13919), .A2(n11963), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11219) );
  OAI21_X1 U13810 ( .B1(n8148), .B2(n13912), .A(n11219), .ZN(n11231) );
  INV_X1 U13811 ( .A(n11220), .ZN(n11223) );
  INV_X1 U13812 ( .A(n11221), .ZN(n11222) );
  NAND2_X1 U13813 ( .A1(n11223), .A2(n11222), .ZN(n11226) );
  XNOR2_X1 U13814 ( .A(n11224), .B(n13789), .ZN(n11252) );
  NAND2_X1 U13815 ( .A1(n13953), .A2(n12612), .ZN(n11253) );
  XNOR2_X1 U13816 ( .A(n11252), .B(n11253), .ZN(n11225) );
  INV_X1 U13817 ( .A(n11225), .ZN(n11227) );
  NAND3_X1 U13818 ( .A1(n11228), .A2(n11227), .A3(n11226), .ZN(n11229) );
  AOI21_X1 U13819 ( .B1(n11256), .B2(n11229), .A(n13925), .ZN(n11230) );
  AOI211_X1 U13820 ( .C1(n13859), .C2(n11232), .A(n11231), .B(n11230), .ZN(
        n11233) );
  INV_X1 U13821 ( .A(n11233), .ZN(P2_U3199) );
  XNOR2_X1 U13822 ( .A(n11234), .B(n11235), .ZN(n15768) );
  INV_X1 U13823 ( .A(n11429), .ZN(n11238) );
  OR2_X1 U13824 ( .A1(n11236), .A2(n15770), .ZN(n15765) );
  OAI22_X1 U13825 ( .A1(n11238), .A2(n15765), .B1(n11237), .B2(n13479), .ZN(
        n11246) );
  XNOR2_X1 U13826 ( .A(n11239), .B(n11240), .ZN(n11244) );
  NAND2_X1 U13827 ( .A1(n15768), .A2(n11425), .ZN(n11243) );
  AOI22_X1 U13828 ( .A1(n13547), .A2(n13118), .B1(n11241), .B2(n13549), .ZN(
        n11242) );
  OAI211_X1 U13829 ( .C1(n13502), .C2(n11244), .A(n11243), .B(n11242), .ZN(
        n15766) );
  MUX2_X1 U13830 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n15766), .S(n13553), .Z(
        n11245) );
  AOI211_X1 U13831 ( .C1(n15768), .C2(n13400), .A(n11246), .B(n11245), .ZN(
        n11247) );
  INV_X1 U13832 ( .A(n11247), .ZN(P3_U3229) );
  INV_X1 U13833 ( .A(n11248), .ZN(n11249) );
  OAI222_X1 U13834 ( .A1(P3_U3151), .A2(n11251), .B1(n13723), .B2(n11250), 
        .C1(n13721), .C2(n11249), .ZN(P3_U3275) );
  INV_X1 U13835 ( .A(n11252), .ZN(n11254) );
  NAND2_X1 U13836 ( .A1(n11254), .A2(n11253), .ZN(n11255) );
  XNOR2_X1 U13837 ( .A(n11661), .B(n13789), .ZN(n11257) );
  AND2_X1 U13838 ( .A1(n13952), .A2(n12612), .ZN(n11258) );
  NAND2_X1 U13839 ( .A1(n11257), .A2(n11258), .ZN(n11383) );
  INV_X1 U13840 ( .A(n11257), .ZN(n11260) );
  INV_X1 U13841 ( .A(n11258), .ZN(n11259) );
  NAND2_X1 U13842 ( .A1(n11260), .A2(n11259), .ZN(n11261) );
  AND2_X1 U13843 ( .A1(n11383), .A2(n11261), .ZN(n11262) );
  OAI211_X1 U13844 ( .C1(n6746), .C2(n11262), .A(n11384), .B(n13903), .ZN(
        n11268) );
  INV_X1 U13845 ( .A(n11663), .ZN(n11266) );
  NAND2_X1 U13846 ( .A1(n13951), .A2(n13907), .ZN(n11264) );
  NAND2_X1 U13847 ( .A1(n13953), .A2(n13905), .ZN(n11263) );
  AND2_X1 U13848 ( .A1(n11264), .A2(n11263), .ZN(n11657) );
  NAND2_X1 U13849 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n13998) );
  OAI21_X1 U13850 ( .B1(n13855), .B2(n11657), .A(n13998), .ZN(n11265) );
  AOI21_X1 U13851 ( .B1(n11266), .B2(n13859), .A(n11265), .ZN(n11267) );
  OAI211_X1 U13852 ( .C1(n6823), .C2(n13912), .A(n11268), .B(n11267), .ZN(
        P2_U3211) );
  XNOR2_X1 U13853 ( .A(n7247), .B(n11269), .ZN(n11392) );
  XNOR2_X1 U13854 ( .A(n11392), .B(n13118), .ZN(n11273) );
  OAI21_X1 U13855 ( .B1(n11273), .B2(n11272), .A(n11586), .ZN(n11274) );
  NAND2_X1 U13856 ( .A1(n11274), .A2(n11608), .ZN(n11279) );
  OAI22_X1 U13857 ( .A1(n13081), .A2(n15769), .B1(n11275), .B2(n13099), .ZN(
        n11276) );
  AOI211_X1 U13858 ( .C1(n13096), .C2(n13117), .A(n11277), .B(n11276), .ZN(
        n11278) );
  OAI211_X1 U13859 ( .C1(n11362), .C2(n11764), .A(n11279), .B(n11278), .ZN(
        P3_U3167) );
  INV_X1 U13860 ( .A(n12301), .ZN(n11282) );
  OAI222_X1 U13861 ( .A1(n15370), .A2(n11281), .B1(n15379), .B2(n11282), .C1(
        n11280), .C2(P1_U3086), .ZN(P1_U3335) );
  OAI222_X1 U13862 ( .A1(n14590), .A2(n11284), .B1(P2_U3088), .B2(n11283), 
        .C1(n14594), .C2(n11282), .ZN(P2_U3307) );
  NAND2_X1 U13863 ( .A1(n11285), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11288) );
  NAND2_X1 U13864 ( .A1(n11286), .A2(n11292), .ZN(n11287) );
  NAND2_X1 U13865 ( .A1(n11288), .A2(n11287), .ZN(n11831) );
  XNOR2_X1 U13866 ( .A(n11831), .B(n11295), .ZN(n11829) );
  XNOR2_X1 U13867 ( .A(n11829), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n11299) );
  NOR2_X1 U13868 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11289), .ZN(n11291) );
  INV_X1 U13869 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15418) );
  NOR2_X1 U13870 ( .A1(n15658), .A2(n15418), .ZN(n11290) );
  AOI211_X1 U13871 ( .C1(n15651), .C2(n11830), .A(n11291), .B(n11290), .ZN(
        n11298) );
  NAND2_X1 U13872 ( .A1(n11292), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n11293) );
  NAND2_X1 U13873 ( .A1(n11294), .A2(n11293), .ZN(n11819) );
  XNOR2_X1 U13874 ( .A(n11819), .B(n11295), .ZN(n11296) );
  NAND2_X1 U13875 ( .A1(n11296), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n11821) );
  OAI211_X1 U13876 ( .C1(n11296), .C2(P2_REG1_REG_15__SCAN_IN), .A(n11821), 
        .B(n15644), .ZN(n11297) );
  OAI211_X1 U13877 ( .C1(n11299), .C2(n15623), .A(n11298), .B(n11297), .ZN(
        P2_U3229) );
  INV_X1 U13878 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n11300) );
  INV_X1 U13879 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14840) );
  NAND2_X1 U13880 ( .A1(n14840), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n11303) );
  NAND2_X1 U13881 ( .A1(n11304), .A2(n11303), .ZN(n11306) );
  INV_X1 U13882 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n11810) );
  NAND2_X1 U13883 ( .A1(n11810), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n11305) );
  NAND2_X1 U13884 ( .A1(n11306), .A2(n11305), .ZN(n11673) );
  XNOR2_X1 U13885 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n11307) );
  XNOR2_X1 U13886 ( .A(n11673), .B(n11307), .ZN(n11308) );
  NAND2_X1 U13887 ( .A1(n11669), .A2(n11670), .ZN(n11310) );
  XNOR2_X1 U13888 ( .A(n11310), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  NAND2_X1 U13889 ( .A1(n11311), .A2(n13709), .ZN(n11313) );
  OAI211_X1 U13890 ( .C1(n11314), .C2(n13723), .A(n11313), .B(n11312), .ZN(
        P3_U3272) );
  INV_X1 U13891 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11315) );
  OAI22_X1 U13892 ( .A1(n15525), .A2(n11316), .B1(n11315), .B2(n15189), .ZN(
        n11319) );
  AOI21_X1 U13893 ( .B1(n15056), .B2(n15147), .A(n11317), .ZN(n11318) );
  AOI211_X1 U13894 ( .C1(n15525), .C2(P1_REG2_REG_0__SCAN_IN), .A(n11319), .B(
        n11318), .ZN(n11322) );
  NAND2_X1 U13895 ( .A1(n15097), .A2(n15552), .ZN(n15104) );
  INV_X1 U13896 ( .A(n15104), .ZN(n15009) );
  OAI21_X1 U13897 ( .B1(n15009), .B2(n15101), .A(n12869), .ZN(n11321) );
  NAND2_X1 U13898 ( .A1(n11322), .A2(n11321), .ZN(P1_U3293) );
  NAND2_X1 U13899 ( .A1(n12712), .A2(n6553), .ZN(n11327) );
  NAND2_X1 U13900 ( .A1(n14786), .A2(n12552), .ZN(n11326) );
  NAND2_X1 U13901 ( .A1(n11327), .A2(n11326), .ZN(n11328) );
  XNOR2_X1 U13902 ( .A(n11328), .B(n11860), .ZN(n11435) );
  AOI22_X1 U13903 ( .A1(n6554), .A2(n12712), .B1(n12572), .B2(n14786), .ZN(
        n11436) );
  XNOR2_X1 U13904 ( .A(n11435), .B(n11436), .ZN(n11433) );
  XNOR2_X1 U13905 ( .A(n11434), .B(n11433), .ZN(n11335) );
  INV_X1 U13906 ( .A(n11329), .ZN(n11332) );
  OAI22_X1 U13907 ( .A1(n14737), .A2(n11330), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11028), .ZN(n11331) );
  AOI21_X1 U13908 ( .B1(n11332), .B2(n14690), .A(n11331), .ZN(n11334) );
  NAND2_X1 U13909 ( .A1(n14740), .A2(n12712), .ZN(n11333) );
  OAI211_X1 U13910 ( .C1(n11335), .C2(n14742), .A(n11334), .B(n11333), .ZN(
        P1_U3239) );
  XNOR2_X1 U13911 ( .A(n11344), .B(n11336), .ZN(n15559) );
  AOI21_X1 U13912 ( .B1(n11351), .B2(n12699), .A(n15538), .ZN(n11338) );
  NAND2_X1 U13913 ( .A1(n11338), .A2(n11337), .ZN(n15556) );
  INV_X1 U13914 ( .A(n15556), .ZN(n11343) );
  INV_X1 U13915 ( .A(n11339), .ZN(n15555) );
  MUX2_X1 U13916 ( .A(n15555), .B(P1_REG2_REG_4__SCAN_IN), .S(n15525), .Z(
        n11342) );
  OAI22_X1 U13917 ( .A1(n15147), .A2(n7470), .B1(n11340), .B2(n15189), .ZN(
        n11341) );
  AOI211_X1 U13918 ( .C1(n11343), .C2(n15521), .A(n11342), .B(n11341), .ZN(
        n11347) );
  XNOR2_X1 U13919 ( .A(n11345), .B(n11344), .ZN(n15562) );
  NAND2_X1 U13920 ( .A1(n15562), .A2(n15101), .ZN(n11346) );
  OAI211_X1 U13921 ( .C1(n15559), .C2(n15104), .A(n11347), .B(n11346), .ZN(
        P1_U3289) );
  XNOR2_X1 U13922 ( .A(n11348), .B(n12874), .ZN(n15549) );
  OR2_X1 U13923 ( .A1(n11349), .A2(n15548), .ZN(n11350) );
  AND3_X1 U13924 ( .A1(n11351), .A2(n15517), .A3(n11350), .ZN(n15544) );
  OAI22_X1 U13925 ( .A1(n11353), .A2(n15128), .B1(n11352), .B2(n15130), .ZN(
        n15545) );
  MUX2_X1 U13926 ( .A(n15545), .B(P1_REG2_REG_3__SCAN_IN), .S(n15525), .Z(
        n11355) );
  INV_X1 U13927 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14829) );
  OAI22_X1 U13928 ( .A1(n15147), .A2(n15548), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n15189), .ZN(n11354) );
  AOI211_X1 U13929 ( .C1(n15544), .C2(n15521), .A(n11355), .B(n11354), .ZN(
        n11358) );
  XNOR2_X1 U13930 ( .A(n11356), .B(n12874), .ZN(n15553) );
  NAND2_X1 U13931 ( .A1(n15009), .A2(n15553), .ZN(n11357) );
  OAI211_X1 U13932 ( .C1(n15122), .C2(n15549), .A(n11358), .B(n11357), .ZN(
        P1_U3290) );
  INV_X1 U13933 ( .A(n12312), .ZN(n12918) );
  OAI222_X1 U13934 ( .A1(n14590), .A2(n15958), .B1(n11897), .B2(n12918), .C1(
        n11359), .C2(P2_U3088), .ZN(P2_U3306) );
  XNOR2_X1 U13935 ( .A(n11360), .B(n11361), .ZN(n15772) );
  INV_X1 U13936 ( .A(n15772), .ZN(n11369) );
  OAI22_X1 U13937 ( .A1(n13456), .A2(n15769), .B1(n11362), .B2(n13479), .ZN(
        n11368) );
  NOR2_X1 U13938 ( .A1(n11363), .A2(n7423), .ZN(n11406) );
  AND2_X1 U13939 ( .A1(n11363), .A2(n7423), .ZN(n11364) );
  OAI21_X1 U13940 ( .B1(n11406), .B2(n11364), .A(n13552), .ZN(n11366) );
  AOI22_X1 U13941 ( .A1(n13547), .A2(n13117), .B1(n13119), .B2(n13549), .ZN(
        n11365) );
  OAI211_X1 U13942 ( .C1(n15772), .C2(n13394), .A(n11366), .B(n11365), .ZN(
        n15774) );
  MUX2_X1 U13943 ( .A(P3_REG2_REG_5__SCAN_IN), .B(n15774), .S(n13553), .Z(
        n11367) );
  AOI211_X1 U13944 ( .C1(n11369), .C2(n13400), .A(n11368), .B(n11367), .ZN(
        n11370) );
  INV_X1 U13945 ( .A(n11370), .ZN(P3_U3228) );
  XNOR2_X1 U13946 ( .A(n11371), .B(n11373), .ZN(n11377) );
  INV_X1 U13947 ( .A(n11377), .ZN(n11724) );
  OAI21_X1 U13948 ( .B1(n8009), .B2(n11373), .A(n11372), .ZN(n11375) );
  INV_X1 U13949 ( .A(n13116), .ZN(n11762) );
  OAI22_X1 U13950 ( .A1(n11762), .A2(n13533), .B1(n11845), .B2(n13535), .ZN(
        n11374) );
  AOI21_X1 U13951 ( .B1(n11375), .B2(n13552), .A(n11374), .ZN(n11376) );
  OAI21_X1 U13952 ( .B1(n11377), .B2(n13394), .A(n11376), .ZN(n11721) );
  AOI21_X1 U13953 ( .B1(n15784), .B2(n11724), .A(n11721), .ZN(n11475) );
  AOI22_X1 U13954 ( .A1(n13695), .A2(n11767), .B1(P3_REG0_REG_8__SCAN_IN), 
        .B2(n15788), .ZN(n11378) );
  OAI21_X1 U13955 ( .B1(n11475), .B2(n15788), .A(n11378), .ZN(P3_U3414) );
  INV_X1 U13956 ( .A(n11379), .ZN(n11381) );
  OAI222_X1 U13957 ( .A1(n11382), .A2(P3_U3151), .B1(n13721), .B2(n11381), 
        .C1(n11380), .C2(n13723), .ZN(P3_U3274) );
  XNOR2_X1 U13958 ( .A(n11683), .B(n13789), .ZN(n11640) );
  NAND2_X1 U13959 ( .A1(n13951), .A2(n12612), .ZN(n11638) );
  XNOR2_X1 U13960 ( .A(n11640), .B(n11638), .ZN(n11385) );
  OAI211_X1 U13961 ( .C1(n11386), .C2(n11385), .A(n11642), .B(n13903), .ZN(
        n11391) );
  OAI22_X1 U13962 ( .A1(n11388), .A2(n13917), .B1(n11387), .B2(n13915), .ZN(
        n11994) );
  AND2_X1 U13963 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n14019) );
  NOR2_X1 U13964 ( .A1(n13921), .A2(n11989), .ZN(n11389) );
  AOI211_X1 U13965 ( .C1(n13919), .C2(n11994), .A(n14019), .B(n11389), .ZN(
        n11390) );
  OAI211_X1 U13966 ( .C1(n7511), .C2(n13912), .A(n11391), .B(n11390), .ZN(
        P2_U3185) );
  INV_X1 U13967 ( .A(n13118), .ZN(n11401) );
  NAND2_X1 U13968 ( .A1(n11392), .A2(n11401), .ZN(n11582) );
  AND2_X1 U13969 ( .A1(n11586), .A2(n11582), .ZN(n11394) );
  XNOR2_X1 U13970 ( .A(n12947), .B(n11411), .ZN(n11583) );
  XOR2_X1 U13971 ( .A(n11583), .B(n13117), .Z(n11393) );
  NAND2_X1 U13972 ( .A1(n11394), .A2(n11393), .ZN(n11463) );
  OAI211_X1 U13973 ( .C1(n11394), .C2(n11393), .A(n11463), .B(n11608), .ZN(
        n11398) );
  OAI22_X1 U13974 ( .A1(n13081), .A2(n11411), .B1(n11401), .B2(n13099), .ZN(
        n11395) );
  AOI211_X1 U13975 ( .C1(n13096), .C2(n13116), .A(n11396), .B(n11395), .ZN(
        n11397) );
  OAI211_X1 U13976 ( .C1(n11412), .C2(n11764), .A(n11398), .B(n11397), .ZN(
        P3_U3179) );
  XNOR2_X1 U13977 ( .A(n11400), .B(n11399), .ZN(n15779) );
  INV_X1 U13978 ( .A(n15779), .ZN(n11416) );
  OAI22_X1 U13979 ( .A1(n11762), .A2(n13535), .B1(n11401), .B2(n13533), .ZN(
        n11410) );
  INV_X1 U13980 ( .A(n11406), .ZN(n11404) );
  AOI21_X1 U13981 ( .B1(n11404), .B2(n11403), .A(n11402), .ZN(n11408) );
  OR2_X1 U13982 ( .A1(n11406), .A2(n11405), .ZN(n11419) );
  INV_X1 U13983 ( .A(n11419), .ZN(n11407) );
  NOR3_X1 U13984 ( .A1(n11408), .A2(n11407), .A3(n13502), .ZN(n11409) );
  AOI211_X1 U13985 ( .C1(n15779), .C2(n11425), .A(n11410), .B(n11409), .ZN(
        n15776) );
  MUX2_X1 U13986 ( .A(n16060), .B(n15776), .S(n13553), .Z(n11415) );
  NOR2_X1 U13987 ( .A1(n11411), .A2(n15770), .ZN(n15778) );
  INV_X1 U13988 ( .A(n11412), .ZN(n11413) );
  AOI22_X1 U13989 ( .A1(n11429), .A2(n15778), .B1(n13557), .B2(n11413), .ZN(
        n11414) );
  OAI211_X1 U13990 ( .C1(n11416), .C2(n11912), .A(n11415), .B(n11414), .ZN(
        P3_U3227) );
  XNOR2_X1 U13991 ( .A(n11417), .B(n11464), .ZN(n15785) );
  INV_X1 U13992 ( .A(n15785), .ZN(n11432) );
  NAND2_X1 U13993 ( .A1(n11419), .A2(n11418), .ZN(n11421) );
  XNOR2_X1 U13994 ( .A(n11421), .B(n11420), .ZN(n11423) );
  AOI22_X1 U13995 ( .A1(n13549), .A2(n13117), .B1(n13114), .B2(n13547), .ZN(
        n11422) );
  OAI21_X1 U13996 ( .B1(n11423), .B2(n13502), .A(n11422), .ZN(n11424) );
  AOI21_X1 U13997 ( .B1(n15785), .B2(n11425), .A(n11424), .ZN(n15781) );
  MUX2_X1 U13998 ( .A(n11426), .B(n15781), .S(n13553), .Z(n11431) );
  NOR2_X1 U13999 ( .A1(n11427), .A2(n15770), .ZN(n15783) );
  INV_X1 U14000 ( .A(n11469), .ZN(n11428) );
  AOI22_X1 U14001 ( .A1(n11429), .A2(n15783), .B1(n13557), .B2(n11428), .ZN(
        n11430) );
  OAI211_X1 U14002 ( .C1(n11432), .C2(n11912), .A(n11431), .B(n11430), .ZN(
        P3_U3226) );
  INV_X1 U14003 ( .A(n11436), .ZN(n11437) );
  NAND2_X1 U14004 ( .A1(n11435), .A2(n11437), .ZN(n11438) );
  NAND2_X1 U14005 ( .A1(n11439), .A2(n12393), .ZN(n11442) );
  AOI22_X1 U14006 ( .A1(n12855), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n12294), 
        .B2(n11440), .ZN(n11441) );
  NAND2_X1 U14007 ( .A1(n15516), .A2(n6553), .ZN(n11444) );
  NAND2_X1 U14008 ( .A1(n14785), .A2(n6554), .ZN(n11443) );
  NAND2_X1 U14009 ( .A1(n11444), .A2(n11443), .ZN(n11445) );
  XNOR2_X1 U14010 ( .A(n11445), .B(n11860), .ZN(n11857) );
  AOI22_X1 U14011 ( .A1(n15516), .A2(n6554), .B1(n12572), .B2(n14785), .ZN(
        n11855) );
  XNOR2_X1 U14012 ( .A(n11857), .B(n11855), .ZN(n11853) );
  XNOR2_X1 U14013 ( .A(n11854), .B(n11853), .ZN(n11462) );
  INV_X1 U14014 ( .A(n11446), .ZN(n15514) );
  NAND2_X1 U14015 ( .A1(n14786), .A2(n15180), .ZN(n11457) );
  NAND2_X1 U14016 ( .A1(n11449), .A2(n11448), .ZN(n11450) );
  NAND2_X1 U14017 ( .A1(n11519), .A2(n11450), .ZN(n12059) );
  OR2_X1 U14018 ( .A1(n11447), .A2(n12059), .ZN(n11455) );
  OR2_X1 U14019 ( .A1(n12413), .A2(n15824), .ZN(n11454) );
  NAND2_X1 U14020 ( .A1(n12410), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n11453) );
  NAND2_X1 U14021 ( .A1(n12448), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n11452) );
  NAND4_X1 U14022 ( .A1(n11455), .A2(n11454), .A3(n11453), .A4(n11452), .ZN(
        n14784) );
  NAND2_X1 U14023 ( .A1(n14784), .A2(n15178), .ZN(n11456) );
  AND2_X1 U14024 ( .A1(n11457), .A2(n11456), .ZN(n15509) );
  OAI21_X1 U14025 ( .B1(n14737), .B2(n15509), .A(n11458), .ZN(n11459) );
  AOI21_X1 U14026 ( .B1(n15514), .B2(n14690), .A(n11459), .ZN(n11461) );
  NAND2_X1 U14027 ( .A1(n14740), .A2(n15516), .ZN(n11460) );
  OAI211_X1 U14028 ( .C1(n11462), .C2(n14742), .A(n11461), .B(n11460), .ZN(
        P1_U3213) );
  NAND2_X1 U14029 ( .A1(n11583), .A2(n13117), .ZN(n11587) );
  NAND2_X1 U14030 ( .A1(n11463), .A2(n11587), .ZN(n11756) );
  XNOR2_X1 U14031 ( .A(n11756), .B(n11588), .ZN(n11474) );
  INV_X1 U14032 ( .A(n13117), .ZN(n11468) );
  NAND2_X1 U14033 ( .A1(n13096), .A2(n13114), .ZN(n11467) );
  INV_X1 U14034 ( .A(n11465), .ZN(n11466) );
  OAI211_X1 U14035 ( .C1(n11468), .C2(n13099), .A(n11467), .B(n11466), .ZN(
        n11471) );
  NOR2_X1 U14036 ( .A1(n11764), .A2(n11469), .ZN(n11470) );
  AOI211_X1 U14037 ( .C1(n11472), .C2(n13102), .A(n11471), .B(n11470), .ZN(
        n11473) );
  OAI21_X1 U14038 ( .B1(n11474), .B2(n13104), .A(n11473), .ZN(P3_U3153) );
  MUX2_X1 U14039 ( .A(n11559), .B(n11475), .S(n15804), .Z(n11476) );
  OAI21_X1 U14040 ( .B1(n11720), .B2(n13610), .A(n11476), .ZN(P3_U3467) );
  XNOR2_X1 U14041 ( .A(n14859), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n11479) );
  AOI211_X1 U14042 ( .C1(n11479), .C2(n11478), .A(n15817), .B(n14853), .ZN(
        n11489) );
  NOR2_X1 U14043 ( .A1(n12071), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11481) );
  XNOR2_X1 U14044 ( .A(n14859), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n11480) );
  NOR3_X1 U14045 ( .A1(n11482), .A2(n11481), .A3(n11480), .ZN(n14862) );
  INV_X1 U14046 ( .A(n14862), .ZN(n11484) );
  OAI21_X1 U14047 ( .B1(n11482), .B2(n11481), .A(n11480), .ZN(n11483) );
  NAND3_X1 U14048 ( .A1(n11484), .A2(n15812), .A3(n11483), .ZN(n11486) );
  AND2_X1 U14049 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14719) );
  AOI21_X1 U14050 ( .B1(n15475), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n14719), 
        .ZN(n11485) );
  OAI211_X1 U14051 ( .C1(n15814), .C2(n11487), .A(n11486), .B(n11485), .ZN(
        n11488) );
  OR2_X1 U14052 ( .A1(n11489), .A2(n11488), .ZN(P1_U3256) );
  INV_X1 U14053 ( .A(n11490), .ZN(n11492) );
  OAI222_X1 U14054 ( .A1(n14590), .A2(n15835), .B1(n11897), .B2(n11492), .C1(
        n11491), .C2(P2_U3088), .ZN(P2_U3305) );
  NAND2_X1 U14055 ( .A1(n11493), .A2(n12393), .ZN(n11496) );
  AOI22_X1 U14056 ( .A1(n11494), .A2(n12294), .B1(n12855), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n11495) );
  NAND2_X1 U14057 ( .A1(n12448), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11502) );
  INV_X1 U14058 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n11497) );
  NAND2_X1 U14059 ( .A1(n11521), .A2(n11497), .ZN(n11498) );
  NAND2_X1 U14060 ( .A1(n11528), .A2(n11498), .ZN(n12216) );
  OR2_X1 U14061 ( .A1(n11447), .A2(n12216), .ZN(n11501) );
  NAND2_X1 U14062 ( .A1(n11451), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11500) );
  NAND2_X1 U14063 ( .A1(n12410), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n11499) );
  NAND4_X1 U14064 ( .A1(n11502), .A2(n11501), .A3(n11500), .A4(n11499), .ZN(
        n14782) );
  INV_X1 U14065 ( .A(n14782), .ZN(n11503) );
  OR2_X1 U14066 ( .A1(n15336), .A2(n11503), .ZN(n12014) );
  NAND2_X1 U14067 ( .A1(n15336), .A2(n11503), .ZN(n11504) );
  NAND2_X1 U14068 ( .A1(n12014), .A2(n11504), .ZN(n12882) );
  NAND2_X1 U14069 ( .A1(n11506), .A2(n11505), .ZN(n11508) );
  OR2_X1 U14070 ( .A1(n12712), .A2(n14786), .ZN(n11507) );
  XNOR2_X1 U14071 ( .A(n15516), .B(n14785), .ZN(n12878) );
  OR2_X1 U14072 ( .A1(n15516), .A2(n14785), .ZN(n11509) );
  NAND2_X1 U14073 ( .A1(n11510), .A2(n12393), .ZN(n11513) );
  AOI22_X1 U14074 ( .A1(n12855), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n12294), 
        .B2(n11511), .ZN(n11512) );
  XNOR2_X1 U14075 ( .A(n12724), .B(n14784), .ZN(n12880) );
  OR2_X1 U14076 ( .A1(n12724), .A2(n14784), .ZN(n11514) );
  NAND2_X1 U14077 ( .A1(n11515), .A2(n12393), .ZN(n11517) );
  AOI22_X1 U14078 ( .A1(n14842), .A2(n12294), .B1(n12855), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n11516) );
  NAND2_X1 U14079 ( .A1(n12448), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n11525) );
  NAND2_X1 U14080 ( .A1(n11519), .A2(n11518), .ZN(n11520) );
  NAND2_X1 U14081 ( .A1(n11521), .A2(n11520), .ZN(n12186) );
  OR2_X1 U14082 ( .A1(n11447), .A2(n12186), .ZN(n11524) );
  NAND2_X1 U14083 ( .A1(n11451), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n11523) );
  NAND2_X1 U14084 ( .A1(n12410), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n11522) );
  NAND4_X1 U14085 ( .A1(n11525), .A2(n11524), .A3(n11523), .A4(n11522), .ZN(
        n14783) );
  XNOR2_X1 U14086 ( .A(n15499), .B(n14783), .ZN(n12883) );
  OR2_X1 U14087 ( .A1(n15499), .A2(n14783), .ZN(n12090) );
  NAND2_X1 U14088 ( .A1(n12092), .A2(n12090), .ZN(n12012) );
  XOR2_X1 U14089 ( .A(n12882), .B(n12012), .Z(n15340) );
  INV_X1 U14090 ( .A(n15516), .ZN(n15582) );
  AND2_X2 U14091 ( .A1(n15519), .A2(n15582), .ZN(n12066) );
  INV_X1 U14092 ( .A(n12724), .ZN(n15592) );
  INV_X1 U14093 ( .A(n15499), .ZN(n15600) );
  XNOR2_X1 U14094 ( .A(n15501), .B(n7488), .ZN(n11526) );
  NAND2_X1 U14095 ( .A1(n11526), .A2(n15517), .ZN(n11535) );
  NAND2_X1 U14096 ( .A1(n12448), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11533) );
  OR2_X2 U14097 ( .A1(n11528), .A2(n11527), .ZN(n12081) );
  NAND2_X1 U14098 ( .A1(n11528), .A2(n11527), .ZN(n11529) );
  NAND2_X1 U14099 ( .A1(n12081), .A2(n11529), .ZN(n12023) );
  OR2_X1 U14100 ( .A1(n11447), .A2(n12023), .ZN(n11532) );
  NAND2_X1 U14101 ( .A1(n11451), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n11531) );
  NAND2_X1 U14102 ( .A1(n12410), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n11530) );
  NAND4_X1 U14103 ( .A1(n11533), .A2(n11532), .A3(n11531), .A4(n11530), .ZN(
        n14781) );
  NAND2_X1 U14104 ( .A1(n14781), .A2(n15178), .ZN(n11534) );
  NAND2_X1 U14105 ( .A1(n11535), .A2(n11534), .ZN(n15334) );
  INV_X1 U14106 ( .A(n12216), .ZN(n11537) );
  AND2_X1 U14107 ( .A1(n14783), .A2(n15180), .ZN(n15335) );
  MUX2_X1 U14108 ( .A(n15335), .B(P1_REG2_REG_10__SCAN_IN), .S(n15525), .Z(
        n11536) );
  AOI21_X1 U14109 ( .B1(n15513), .B2(n11537), .A(n11536), .ZN(n11538) );
  OAI21_X1 U14110 ( .B1(n7488), .B2(n15147), .A(n11538), .ZN(n11539) );
  AOI21_X1 U14111 ( .B1(n15334), .B2(n15521), .A(n11539), .ZN(n11552) );
  NAND2_X1 U14112 ( .A1(n11540), .A2(n12877), .ZN(n11543) );
  INV_X1 U14113 ( .A(n14786), .ZN(n11541) );
  NAND2_X1 U14114 ( .A1(n12712), .A2(n11541), .ZN(n11542) );
  NAND2_X1 U14115 ( .A1(n11543), .A2(n11542), .ZN(n15507) );
  NAND2_X1 U14116 ( .A1(n15507), .A2(n12878), .ZN(n11546) );
  INV_X1 U14117 ( .A(n14785), .ZN(n11544) );
  NAND2_X1 U14118 ( .A1(n15516), .A2(n11544), .ZN(n11545) );
  NAND2_X1 U14119 ( .A1(n11546), .A2(n11545), .ZN(n12060) );
  INV_X1 U14120 ( .A(n14784), .ZN(n11862) );
  OR2_X1 U14121 ( .A1(n12724), .A2(n11862), .ZN(n11547) );
  INV_X1 U14122 ( .A(n14783), .ZN(n12215) );
  NAND2_X1 U14123 ( .A1(n15499), .A2(n12215), .ZN(n11548) );
  NAND2_X1 U14124 ( .A1(n11550), .A2(n12882), .ZN(n15337) );
  NAND3_X1 U14125 ( .A1(n12015), .A2(n15337), .A3(n15009), .ZN(n11551) );
  OAI211_X1 U14126 ( .C1(n15340), .C2(n15195), .A(n11552), .B(n11551), .ZN(
        P1_U3283) );
  MUX2_X1 U14127 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n13724), .Z(n11555) );
  NAND2_X1 U14128 ( .A1(n11569), .A2(n11555), .ZN(n11802) );
  NOR2_X1 U14129 ( .A1(n11569), .A2(n11555), .ZN(n11800) );
  NOR2_X1 U14130 ( .A1(n11805), .A2(n11800), .ZN(n11557) );
  MUX2_X1 U14131 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13724), .Z(n13137) );
  XNOR2_X1 U14132 ( .A(n13124), .B(n13137), .ZN(n11556) );
  NOR2_X1 U14133 ( .A1(n11557), .A2(n11556), .ZN(n13138) );
  AOI21_X1 U14134 ( .B1(n11557), .B2(n11556), .A(n13138), .ZN(n11581) );
  NAND2_X1 U14135 ( .A1(n11561), .A2(n11569), .ZN(n11562) );
  INV_X1 U14136 ( .A(n11562), .ZN(n11564) );
  XNOR2_X1 U14137 ( .A(n13124), .B(n13133), .ZN(n11563) );
  INV_X1 U14138 ( .A(n13132), .ZN(n11566) );
  NOR3_X1 U14139 ( .A1(n6733), .A2(n11564), .A3(n11563), .ZN(n11565) );
  OAI21_X1 U14140 ( .B1(n11566), .B2(n11565), .A(n13313), .ZN(n11580) );
  INV_X1 U14141 ( .A(n13124), .ZN(n13140) );
  INV_X1 U14142 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n11674) );
  NAND2_X1 U14143 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n11611)
         );
  OAI21_X1 U14144 ( .B1(n13321), .B2(n11674), .A(n11611), .ZN(n11578) );
  INV_X1 U14145 ( .A(n11569), .ZN(n11807) );
  NOR2_X1 U14146 ( .A1(n11570), .A2(n11807), .ZN(n11571) );
  INV_X1 U14147 ( .A(n11571), .ZN(n11573) );
  XNOR2_X1 U14148 ( .A(n13124), .B(P3_REG2_REG_10__SCAN_IN), .ZN(n11574) );
  INV_X1 U14149 ( .A(n13123), .ZN(n11576) );
  NAND3_X1 U14150 ( .A1(n11572), .A2(n11574), .A3(n11573), .ZN(n11575) );
  AOI21_X1 U14151 ( .B1(n11576), .B2(n11575), .A(n13283), .ZN(n11577) );
  AOI211_X1 U14152 ( .C1(n13323), .C2(n13140), .A(n11578), .B(n11577), .ZN(
        n11579) );
  OAI211_X1 U14153 ( .C1(n11581), .C2(n13210), .A(n11580), .B(n11579), .ZN(
        P3_U3192) );
  XNOR2_X1 U14154 ( .A(n11985), .B(n12947), .ZN(n11602) );
  XNOR2_X1 U14155 ( .A(n11602), .B(n11759), .ZN(n11596) );
  XNOR2_X1 U14156 ( .A(n11720), .B(n12947), .ZN(n11589) );
  OAI211_X1 U14157 ( .C1(n11583), .C2(n13117), .A(n11588), .B(n11582), .ZN(
        n11584) );
  NOR2_X1 U14158 ( .A1(n11758), .A2(n11584), .ZN(n11585) );
  OAI21_X1 U14159 ( .B1(n11758), .B2(n11587), .A(n11588), .ZN(n11591) );
  OAI21_X1 U14160 ( .B1(n11758), .B2(n11762), .A(n11755), .ZN(n11590) );
  AOI22_X1 U14161 ( .A1(n11591), .A2(n11590), .B1(n11589), .B2(n13114), .ZN(
        n11592) );
  INV_X1 U14162 ( .A(n11607), .ZN(n11594) );
  AOI21_X1 U14163 ( .B1(n11596), .B2(n11595), .A(n11594), .ZN(n11601) );
  INV_X1 U14164 ( .A(n13099), .ZN(n13066) );
  NAND2_X1 U14165 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11808) );
  OAI21_X1 U14166 ( .B1(n13088), .B2(n11604), .A(n11808), .ZN(n11597) );
  AOI21_X1 U14167 ( .B1(n13066), .B2(n13114), .A(n11597), .ZN(n11598) );
  OAI21_X1 U14168 ( .B1(n11794), .B2(n11764), .A(n11598), .ZN(n11599) );
  AOI21_X1 U14169 ( .B1(n11796), .B2(n13102), .A(n11599), .ZN(n11600) );
  OAI21_X1 U14170 ( .B1(n11601), .B2(n13104), .A(n11600), .ZN(P3_U3171) );
  INV_X1 U14171 ( .A(n11602), .ZN(n11603) );
  NAND2_X1 U14172 ( .A1(n11603), .A2(n11845), .ZN(n11605) );
  AND2_X1 U14173 ( .A1(n11607), .A2(n11605), .ZN(n11610) );
  XNOR2_X1 U14174 ( .A(n11746), .B(n11604), .ZN(n11609) );
  AND2_X1 U14175 ( .A1(n11609), .A2(n11605), .ZN(n11606) );
  OAI211_X1 U14176 ( .C1(n11610), .C2(n11609), .A(n11608), .B(n11748), .ZN(
        n11615) );
  OAI21_X1 U14177 ( .B1(n13088), .B2(n11949), .A(n11611), .ZN(n11613) );
  NOR2_X1 U14178 ( .A1(n11764), .A2(n11907), .ZN(n11612) );
  AOI211_X1 U14179 ( .C1(n13066), .C2(n11759), .A(n11613), .B(n11612), .ZN(
        n11614) );
  OAI211_X1 U14180 ( .C1(n13081), .C2(n12053), .A(n11615), .B(n11614), .ZN(
        P3_U3157) );
  INV_X1 U14181 ( .A(n11616), .ZN(n11618) );
  NAND2_X1 U14182 ( .A1(n11618), .A2(n11617), .ZN(n11619) );
  NAND2_X1 U14183 ( .A1(n15715), .A2(n14086), .ZN(n11620) );
  AND2_X1 U14184 ( .A1(n13789), .A2(n11620), .ZN(n11621) );
  INV_X1 U14185 ( .A(n11622), .ZN(n11627) );
  OAI22_X1 U14186 ( .A1(n14399), .A2(n11625), .B1(n11624), .B2(n14398), .ZN(
        n11626) );
  AOI21_X1 U14187 ( .B1(n14401), .B2(n11627), .A(n11626), .ZN(n11631) );
  MUX2_X1 U14188 ( .A(n11629), .B(n11628), .S(n14285), .Z(n11630) );
  OAI211_X1 U14189 ( .C1(n14361), .C2(n11632), .A(n11631), .B(n11630), .ZN(
        P2_U3261) );
  XNOR2_X1 U14190 ( .A(n14519), .B(n12649), .ZN(n11634) );
  NAND2_X1 U14191 ( .A1(n13950), .A2(n12612), .ZN(n11635) );
  NAND2_X1 U14192 ( .A1(n11634), .A2(n11635), .ZN(n11919) );
  INV_X1 U14193 ( .A(n11634), .ZN(n11637) );
  INV_X1 U14194 ( .A(n11635), .ZN(n11636) );
  NAND2_X1 U14195 ( .A1(n11637), .A2(n11636), .ZN(n11921) );
  NAND2_X1 U14196 ( .A1(n11919), .A2(n11921), .ZN(n11643) );
  INV_X1 U14197 ( .A(n11638), .ZN(n11639) );
  NAND2_X1 U14198 ( .A1(n11640), .A2(n11639), .ZN(n11641) );
  XOR2_X1 U14199 ( .A(n11643), .B(n11920), .Z(n11649) );
  NAND2_X1 U14200 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n14025) );
  OAI22_X1 U14201 ( .A1(n11645), .A2(n13917), .B1(n11644), .B2(n13915), .ZN(
        n11691) );
  NAND2_X1 U14202 ( .A1(n13919), .A2(n11691), .ZN(n11646) );
  OAI211_X1 U14203 ( .C1(n13921), .C2(n11695), .A(n14025), .B(n11646), .ZN(
        n11647) );
  AOI21_X1 U14204 ( .B1(n14519), .B2(n13923), .A(n11647), .ZN(n11648) );
  OAI21_X1 U14205 ( .B1(n11649), .B2(n13925), .A(n11648), .ZN(P2_U3193) );
  NAND2_X1 U14206 ( .A1(n11651), .A2(n11656), .ZN(n11652) );
  NAND2_X1 U14207 ( .A1(n11650), .A2(n11652), .ZN(n15727) );
  NOR2_X1 U14208 ( .A1(n14086), .A2(n11653), .ZN(n11654) );
  AND2_X1 U14209 ( .A1(n14285), .A2(n11654), .ZN(n15667) );
  INV_X1 U14210 ( .A(n15667), .ZN(n14405) );
  XNOR2_X1 U14211 ( .A(n11655), .B(n8496), .ZN(n11659) );
  OR2_X1 U14212 ( .A1(n15727), .A2(n15715), .ZN(n11658) );
  OAI211_X1 U14213 ( .C1(n14375), .C2(n11659), .A(n11658), .B(n11657), .ZN(
        n15730) );
  MUX2_X1 U14214 ( .A(n15730), .B(P2_REG2_REG_6__SCAN_IN), .S(n6557), .Z(
        n11660) );
  INV_X1 U14215 ( .A(n11660), .ZN(n11666) );
  AOI21_X1 U14216 ( .B1(n11958), .B2(n11661), .A(n14338), .ZN(n11662) );
  AND2_X1 U14217 ( .A1(n11986), .A2(n11662), .ZN(n15728) );
  OAI22_X1 U14218 ( .A1(n14399), .A2(n6823), .B1(n11663), .B2(n14398), .ZN(
        n11664) );
  AOI21_X1 U14219 ( .B1(n14401), .B2(n15728), .A(n11664), .ZN(n11665) );
  OAI211_X1 U14220 ( .C1(n15727), .C2(n14405), .A(n11666), .B(n11665), .ZN(
        P2_U3259) );
  INV_X1 U14221 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n15921) );
  NAND2_X1 U14222 ( .A1(n13386), .A2(P3_U3897), .ZN(n11667) );
  OAI21_X1 U14223 ( .B1(n13115), .B2(n15921), .A(n11667), .ZN(P3_U3516) );
  INV_X1 U14224 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n15926) );
  NAND2_X1 U14225 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n15926), .ZN(n11672) );
  NAND2_X1 U14226 ( .A1(n11673), .A2(n11672), .ZN(n11676) );
  NAND2_X1 U14227 ( .A1(n11674), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n11675) );
  NAND2_X1 U14228 ( .A1(n11676), .A2(n11675), .ZN(n12041) );
  INV_X1 U14229 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n11677) );
  NAND2_X1 U14230 ( .A1(n11677), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n12042) );
  INV_X1 U14231 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n13131) );
  NAND2_X1 U14232 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n13131), .ZN(n12039) );
  AND2_X1 U14233 ( .A1(n12042), .A2(n12039), .ZN(n11678) );
  XNOR2_X1 U14234 ( .A(n12041), .B(n11678), .ZN(n11679) );
  NAND2_X1 U14235 ( .A1(n12037), .A2(n12038), .ZN(n11680) );
  XNOR2_X1 U14236 ( .A(n11680), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  INV_X1 U14237 ( .A(n11681), .ZN(n11682) );
  NAND2_X1 U14238 ( .A1(n11650), .A2(n11682), .ZN(n14383) );
  OAI21_X1 U14239 ( .B1(n14383), .B2(n13951), .A(n11683), .ZN(n11685) );
  NAND2_X1 U14240 ( .A1(n14383), .A2(n13951), .ZN(n11684) );
  NAND2_X1 U14241 ( .A1(n11685), .A2(n11684), .ZN(n11686) );
  XNOR2_X1 U14242 ( .A(n11686), .B(n11688), .ZN(n11692) );
  INV_X1 U14243 ( .A(n11692), .ZN(n14522) );
  INV_X1 U14244 ( .A(n15715), .ZN(n15713) );
  OR2_X1 U14245 ( .A1(n11687), .A2(n7170), .ZN(n14372) );
  NAND2_X1 U14246 ( .A1(n11687), .A2(n7170), .ZN(n11689) );
  AOI21_X1 U14247 ( .B1(n14372), .B2(n11689), .A(n14375), .ZN(n11690) );
  AOI211_X1 U14248 ( .C1(n11692), .C2(n15713), .A(n11691), .B(n11690), .ZN(
        n14521) );
  MUX2_X1 U14249 ( .A(n11693), .B(n14521), .S(n14285), .Z(n11699) );
  OAI21_X1 U14250 ( .B1(n11987), .B2(n11696), .A(n14470), .ZN(n11694) );
  NOR2_X1 U14251 ( .A1(n11694), .A2(n14396), .ZN(n14517) );
  OAI22_X1 U14252 ( .A1(n14399), .A2(n11696), .B1(n11695), .B2(n14398), .ZN(
        n11697) );
  AOI21_X1 U14253 ( .B1(n14517), .B2(n14401), .A(n11697), .ZN(n11698) );
  OAI211_X1 U14254 ( .C1(n14522), .C2(n14405), .A(n11699), .B(n11698), .ZN(
        P2_U3257) );
  INV_X1 U14255 ( .A(n11700), .ZN(n11702) );
  OAI222_X1 U14256 ( .A1(P3_U3151), .A2(n11703), .B1(n13721), .B2(n11702), 
        .C1(n11701), .C2(n13723), .ZN(P3_U3271) );
  XNOR2_X1 U14257 ( .A(n11704), .B(n11708), .ZN(n15714) );
  INV_X1 U14258 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n11712) );
  AOI21_X1 U14259 ( .B1(n11707), .B2(n11706), .A(n11705), .ZN(n11709) );
  XNOR2_X1 U14260 ( .A(n11709), .B(n11708), .ZN(n11711) );
  OAI21_X1 U14261 ( .B1(n11711), .B2(n14375), .A(n11710), .ZN(n15720) );
  AOI21_X1 U14262 ( .B1(n15666), .B2(n11712), .A(n15720), .ZN(n11713) );
  MUX2_X1 U14263 ( .A(n11714), .B(n11713), .S(n14285), .Z(n11719) );
  AOI211_X1 U14264 ( .C1(n11717), .C2(n11716), .A(n14338), .B(n11715), .ZN(
        n15718) );
  AOI22_X1 U14265 ( .A1(n14368), .A2(n11717), .B1(n14401), .B2(n15718), .ZN(
        n11718) );
  OAI211_X1 U14266 ( .C1(n14361), .C2(n15714), .A(n11719), .B(n11718), .ZN(
        P2_U3262) );
  OAI22_X1 U14267 ( .A1(n13456), .A2(n11720), .B1(n11763), .B2(n13479), .ZN(
        n11723) );
  MUX2_X1 U14268 ( .A(P3_REG2_REG_8__SCAN_IN), .B(n11721), .S(n13553), .Z(
        n11722) );
  AOI211_X1 U14269 ( .C1(n11724), .C2(n13400), .A(n11723), .B(n11722), .ZN(
        n11725) );
  INV_X1 U14270 ( .A(n11725), .ZN(P3_U3225) );
  XNOR2_X1 U14271 ( .A(n11727), .B(n11726), .ZN(n14500) );
  OAI22_X1 U14272 ( .A1(n11728), .A2(n13915), .B1(n13864), .B2(n13917), .ZN(
        n13883) );
  NAND3_X1 U14273 ( .A1(n11729), .A2(n11731), .A3(n11730), .ZN(n11732) );
  AOI21_X1 U14274 ( .B1(n11733), .B2(n11732), .A(n14375), .ZN(n11734) );
  AOI211_X1 U14275 ( .C1(n15713), .C2(n14500), .A(n13883), .B(n11734), .ZN(
        n14497) );
  INV_X1 U14276 ( .A(n8021), .ZN(n14354) );
  AOI211_X1 U14277 ( .C1(n13887), .C2(n11735), .A(n14338), .B(n14354), .ZN(
        n14499) );
  NOR2_X1 U14278 ( .A1(n14570), .A2(n14399), .ZN(n11737) );
  OAI22_X1 U14279 ( .A1(n14285), .A2(n16086), .B1(n13885), .B2(n14398), .ZN(
        n11736) );
  AOI211_X1 U14280 ( .C1(n14499), .C2(n14401), .A(n11737), .B(n11736), .ZN(
        n11739) );
  NAND2_X1 U14281 ( .A1(n14500), .A2(n15667), .ZN(n11738) );
  OAI211_X1 U14282 ( .C1(n14497), .C2(n6557), .A(n11739), .B(n11738), .ZN(
        P2_U3254) );
  NAND2_X1 U14283 ( .A1(n12340), .A2(n11740), .ZN(n11742) );
  OAI211_X1 U14284 ( .C1(n11743), .C2(n14590), .A(n11742), .B(n11741), .ZN(
        P2_U3304) );
  NAND2_X1 U14285 ( .A1(n12340), .A2(n11744), .ZN(n11745) );
  OAI211_X1 U14286 ( .C1(n15918), .C2(n15370), .A(n11745), .B(n12915), .ZN(
        P1_U3332) );
  NAND2_X1 U14287 ( .A1(n11746), .A2(n13113), .ZN(n11747) );
  XNOR2_X1 U14288 ( .A(n12003), .B(n12995), .ZN(n11943) );
  XNOR2_X1 U14289 ( .A(n11943), .B(n13112), .ZN(n11749) );
  XNOR2_X1 U14290 ( .A(n11942), .B(n11749), .ZN(n11754) );
  INV_X1 U14291 ( .A(n12003), .ZN(n11781) );
  NAND2_X1 U14292 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n13129)
         );
  OAI21_X1 U14293 ( .B1(n13088), .B2(n13059), .A(n13129), .ZN(n11750) );
  AOI21_X1 U14294 ( .B1(n13066), .B2(n13113), .A(n11750), .ZN(n11751) );
  OAI21_X1 U14295 ( .B1(n11900), .B2(n11764), .A(n11751), .ZN(n11752) );
  AOI21_X1 U14296 ( .B1(n11781), .B2(n13102), .A(n11752), .ZN(n11753) );
  OAI21_X1 U14297 ( .B1(n11754), .B2(n13104), .A(n11753), .ZN(P3_U3176) );
  MUX2_X1 U14298 ( .A(n11756), .B(n13116), .S(n11755), .Z(n11757) );
  XOR2_X1 U14299 ( .A(n11758), .B(n11757), .Z(n11769) );
  NAND2_X1 U14300 ( .A1(n13096), .A2(n11759), .ZN(n11761) );
  OAI211_X1 U14301 ( .C1(n11762), .C2(n13099), .A(n11761), .B(n11760), .ZN(
        n11766) );
  NOR2_X1 U14302 ( .A1(n11764), .A2(n11763), .ZN(n11765) );
  AOI211_X1 U14303 ( .C1(n11767), .C2(n13102), .A(n11766), .B(n11765), .ZN(
        n11768) );
  OAI21_X1 U14304 ( .B1(n11769), .B2(n13104), .A(n11768), .ZN(P3_U3161) );
  XOR2_X1 U14305 ( .A(n11771), .B(n11770), .Z(n11799) );
  INV_X1 U14306 ( .A(n11799), .ZN(n11776) );
  AOI22_X1 U14307 ( .A1(n13549), .A2(n13114), .B1(n13113), .B2(n13547), .ZN(
        n11775) );
  OAI211_X1 U14308 ( .C1(n11773), .C2(n9778), .A(n13552), .B(n11772), .ZN(
        n11774) );
  OAI211_X1 U14309 ( .C1(n11799), .C2(n13394), .A(n11775), .B(n11774), .ZN(
        n11791) );
  AOI21_X1 U14310 ( .B1(n15784), .B2(n11776), .A(n11791), .ZN(n11982) );
  AOI22_X1 U14311 ( .A1(n13695), .A2(n11796), .B1(P3_REG0_REG_9__SCAN_IN), 
        .B2(n15788), .ZN(n11777) );
  OAI21_X1 U14312 ( .B1(n11982), .B2(n15788), .A(n11777), .ZN(P3_U3417) );
  XNOR2_X1 U14313 ( .A(n11778), .B(n11779), .ZN(n11780) );
  AOI222_X1 U14314 ( .A1(n13552), .A2(n11780), .B1(n13550), .B2(n13547), .C1(
        n13113), .C2(n13549), .ZN(n11999) );
  AOI22_X1 U14315 ( .A1(n13695), .A2(n11781), .B1(P3_REG0_REG_11__SCAN_IN), 
        .B2(n15788), .ZN(n11785) );
  XNOR2_X1 U14316 ( .A(n11783), .B(n11782), .ZN(n12000) );
  INV_X1 U14317 ( .A(n13699), .ZN(n13673) );
  NAND2_X1 U14318 ( .A1(n12000), .A2(n13673), .ZN(n11784) );
  OAI211_X1 U14319 ( .C1(n11999), .C2(n15788), .A(n11785), .B(n11784), .ZN(
        P3_U3423) );
  INV_X1 U14320 ( .A(n12360), .ZN(n11789) );
  OAI222_X1 U14321 ( .A1(n15370), .A2(n11787), .B1(n15379), .B2(n11789), .C1(
        P1_U3086), .C2(n11786), .ZN(P1_U3331) );
  OAI222_X1 U14322 ( .A1(n14590), .A2(n11790), .B1(n11897), .B2(n11789), .C1(
        n11788), .C2(P2_U3088), .ZN(P2_U3303) );
  INV_X1 U14323 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11793) );
  INV_X1 U14324 ( .A(n11791), .ZN(n11792) );
  MUX2_X1 U14325 ( .A(n11793), .B(n11792), .S(n13553), .Z(n11798) );
  NOR2_X1 U14326 ( .A1(n13479), .A2(n11794), .ZN(n11795) );
  AOI21_X1 U14327 ( .B1(n13558), .B2(n11796), .A(n11795), .ZN(n11797) );
  OAI211_X1 U14328 ( .C1(n11799), .C2(n11912), .A(n11798), .B(n11797), .ZN(
        P3_U3224) );
  INV_X1 U14329 ( .A(n11800), .ZN(n11804) );
  AOI21_X1 U14330 ( .B1(n11804), .B2(n11802), .A(n11801), .ZN(n11803) );
  AOI21_X1 U14331 ( .B1(n11805), .B2(n11804), .A(n11803), .ZN(n11817) );
  OAI21_X1 U14332 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n11806), .A(n11572), .ZN(
        n11815) );
  NAND2_X1 U14333 ( .A1(n13323), .A2(n11807), .ZN(n11809) );
  OAI211_X1 U14334 ( .C1(n13321), .C2(n11810), .A(n11809), .B(n11808), .ZN(
        n11814) );
  AOI21_X1 U14335 ( .B1(n11983), .B2(n11811), .A(n6733), .ZN(n11812) );
  NOR2_X1 U14336 ( .A1(n11812), .A2(n13190), .ZN(n11813) );
  AOI211_X1 U14337 ( .C1(n13318), .C2(n11815), .A(n11814), .B(n11813), .ZN(
        n11816) );
  OAI21_X1 U14338 ( .B1(n11817), .B2(n13210), .A(n11816), .ZN(P3_U3191) );
  INV_X1 U14339 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n16012) );
  NAND2_X1 U14340 ( .A1(n9803), .A2(P3_U3897), .ZN(n11818) );
  OAI21_X1 U14341 ( .B1(n13115), .B2(n16012), .A(n11818), .ZN(P3_U3518) );
  NAND2_X1 U14342 ( .A1(n11819), .A2(n11830), .ZN(n11820) );
  NAND2_X1 U14343 ( .A1(n11821), .A2(n11820), .ZN(n11882) );
  XNOR2_X1 U14344 ( .A(n11886), .B(n11822), .ZN(n11881) );
  NAND2_X1 U14345 ( .A1(n11886), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n11823) );
  XNOR2_X1 U14346 ( .A(n11836), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n11824) );
  OAI211_X1 U14347 ( .C1(n11825), .C2(n11824), .A(n14066), .B(n15644), .ZN(
        n11828) );
  NAND2_X1 U14348 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13838)
         );
  INV_X1 U14349 ( .A(n11836), .ZN(n14065) );
  NAND2_X1 U14350 ( .A1(n15651), .A2(n14065), .ZN(n11827) );
  NAND2_X1 U14351 ( .A1(n15629), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n11826) );
  AND4_X1 U14352 ( .A1(n11828), .A2(n13838), .A3(n11827), .A4(n11826), .ZN(
        n11841) );
  NAND2_X1 U14353 ( .A1(n11829), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n11833) );
  NAND2_X1 U14354 ( .A1(n11831), .A2(n11830), .ZN(n11832) );
  NAND2_X1 U14355 ( .A1(n11833), .A2(n11832), .ZN(n11879) );
  XNOR2_X1 U14356 ( .A(n11886), .B(n14284), .ZN(n11878) );
  NAND2_X1 U14357 ( .A1(n11879), .A2(n11878), .ZN(n11835) );
  NAND2_X1 U14358 ( .A1(n11886), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11834) );
  NAND2_X1 U14359 ( .A1(n11835), .A2(n11834), .ZN(n11839) );
  MUX2_X1 U14360 ( .A(n11837), .B(P2_REG2_REG_17__SCAN_IN), .S(n11836), .Z(
        n11838) );
  NAND2_X1 U14361 ( .A1(n11839), .A2(n11838), .ZN(n14057) );
  OAI211_X1 U14362 ( .C1(n11839), .C2(n11838), .A(n14057), .B(n15653), .ZN(
        n11840) );
  NAND2_X1 U14363 ( .A1(n11841), .A2(n11840), .ZN(P2_U3231) );
  XNOR2_X1 U14364 ( .A(n11842), .B(n11843), .ZN(n11913) );
  INV_X1 U14365 ( .A(n11913), .ZN(n11849) );
  XNOR2_X1 U14366 ( .A(n11844), .B(n11843), .ZN(n11847) );
  OAI22_X1 U14367 ( .A1(n11949), .A2(n13535), .B1(n11845), .B2(n13533), .ZN(
        n11846) );
  AOI21_X1 U14368 ( .B1(n11847), .B2(n13552), .A(n11846), .ZN(n11848) );
  OAI21_X1 U14369 ( .B1(n11913), .B2(n13394), .A(n11848), .ZN(n11904) );
  AOI21_X1 U14370 ( .B1(n15784), .B2(n11849), .A(n11904), .ZN(n12051) );
  INV_X1 U14371 ( .A(n12053), .ZN(n11909) );
  AOI22_X1 U14372 ( .A1(n13695), .A2(n11909), .B1(P3_REG0_REG_10__SCAN_IN), 
        .B2(n15788), .ZN(n11850) );
  OAI21_X1 U14373 ( .B1(n12051), .B2(n15788), .A(n11850), .ZN(P3_U3420) );
  INV_X1 U14374 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n15950) );
  INV_X1 U14375 ( .A(n13352), .ZN(n11851) );
  NAND2_X1 U14376 ( .A1(n11851), .A2(P3_U3897), .ZN(n11852) );
  OAI21_X1 U14377 ( .B1(n13115), .B2(n15950), .A(n11852), .ZN(P3_U3519) );
  INV_X1 U14378 ( .A(n11855), .ZN(n11856) );
  NAND2_X1 U14379 ( .A1(n12724), .A2(n6553), .ZN(n11859) );
  NAND2_X1 U14380 ( .A1(n14784), .A2(n6554), .ZN(n11858) );
  NAND2_X1 U14381 ( .A1(n11859), .A2(n11858), .ZN(n11861) );
  XNOR2_X1 U14382 ( .A(n11861), .B(n12534), .ZN(n11865) );
  NOR2_X1 U14383 ( .A1(n14636), .A2(n11862), .ZN(n11863) );
  AOI21_X1 U14384 ( .B1(n12724), .B2(n12552), .A(n11863), .ZN(n11864) );
  NAND2_X1 U14385 ( .A1(n11865), .A2(n11864), .ZN(n12123) );
  OAI21_X1 U14386 ( .B1(n11865), .B2(n11864), .A(n12123), .ZN(n11870) );
  INV_X1 U14387 ( .A(n12124), .ZN(n11869) );
  AOI21_X1 U14388 ( .B1(n11866), .B2(n11870), .A(n11869), .ZN(n11877) );
  INV_X1 U14389 ( .A(n14737), .ZN(n14762) );
  NAND2_X1 U14390 ( .A1(n14785), .A2(n15180), .ZN(n11872) );
  NAND2_X1 U14391 ( .A1(n14783), .A2(n15178), .ZN(n11871) );
  NAND2_X1 U14392 ( .A1(n11872), .A2(n11871), .ZN(n15590) );
  NAND2_X1 U14393 ( .A1(n14762), .A2(n15590), .ZN(n11873) );
  OAI211_X1 U14394 ( .C1(n14759), .C2(n12059), .A(n11874), .B(n11873), .ZN(
        n11875) );
  AOI21_X1 U14395 ( .B1(n14740), .B2(n12724), .A(n11875), .ZN(n11876) );
  OAI21_X1 U14396 ( .B1(n11877), .B2(n14742), .A(n11876), .ZN(P1_U3221) );
  XNOR2_X1 U14397 ( .A(n11879), .B(n11878), .ZN(n11888) );
  INV_X1 U14398 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15432) );
  NAND2_X1 U14399 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13828)
         );
  OAI21_X1 U14400 ( .B1(n15658), .B2(n15432), .A(n13828), .ZN(n11885) );
  OAI211_X1 U14401 ( .C1(n11882), .C2(n11881), .A(n11880), .B(n15644), .ZN(
        n11883) );
  INV_X1 U14402 ( .A(n11883), .ZN(n11884) );
  AOI211_X1 U14403 ( .C1(n15651), .C2(n11886), .A(n11885), .B(n11884), .ZN(
        n11887) );
  OAI21_X1 U14404 ( .B1(n11888), .B2(n15623), .A(n11887), .ZN(P2_U3230) );
  INV_X1 U14405 ( .A(n11889), .ZN(n11890) );
  OAI222_X1 U14406 ( .A1(n11892), .A2(P3_U3151), .B1(n13723), .B2(n11891), 
        .C1(n13721), .C2(n11890), .ZN(P3_U3270) );
  INV_X1 U14407 ( .A(n12350), .ZN(n11896) );
  OAI222_X1 U14408 ( .A1(n15370), .A2(n11894), .B1(n15379), .B2(n11896), .C1(
        P1_U3086), .C2(n11893), .ZN(P1_U3330) );
  OAI222_X1 U14409 ( .A1(n14590), .A2(n11898), .B1(n11897), .B2(n11896), .C1(
        P2_U3088), .C2(n11895), .ZN(P2_U3302) );
  MUX2_X1 U14410 ( .A(n11899), .B(n11999), .S(n13553), .Z(n11903) );
  OAI22_X1 U14411 ( .A1(n13456), .A2(n12003), .B1(n11900), .B2(n13479), .ZN(
        n11901) );
  AOI21_X1 U14412 ( .B1(n12000), .B2(n13360), .A(n11901), .ZN(n11902) );
  NAND2_X1 U14413 ( .A1(n11903), .A2(n11902), .ZN(P3_U3222) );
  INV_X1 U14414 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11906) );
  INV_X1 U14415 ( .A(n11904), .ZN(n11905) );
  MUX2_X1 U14416 ( .A(n11906), .B(n11905), .S(n13553), .Z(n11911) );
  NOR2_X1 U14417 ( .A1(n13479), .A2(n11907), .ZN(n11908) );
  AOI21_X1 U14418 ( .B1(n13558), .B2(n11909), .A(n11908), .ZN(n11910) );
  OAI211_X1 U14419 ( .C1(n11913), .C2(n11912), .A(n11911), .B(n11910), .ZN(
        P3_U3223) );
  XNOR2_X1 U14420 ( .A(n14575), .B(n12649), .ZN(n11914) );
  NAND2_X1 U14421 ( .A1(n13949), .A2(n12612), .ZN(n11915) );
  NAND2_X1 U14422 ( .A1(n11914), .A2(n11915), .ZN(n12028) );
  INV_X1 U14423 ( .A(n11914), .ZN(n11917) );
  INV_X1 U14424 ( .A(n11915), .ZN(n11916) );
  NAND2_X1 U14425 ( .A1(n11917), .A2(n11916), .ZN(n11918) );
  NAND2_X1 U14426 ( .A1(n12028), .A2(n11918), .ZN(n11925) );
  INV_X1 U14427 ( .A(n12029), .ZN(n11923) );
  AOI21_X1 U14428 ( .B1(n11925), .B2(n11924), .A(n11923), .ZN(n11932) );
  NAND2_X1 U14429 ( .A1(n13948), .A2(n13907), .ZN(n11927) );
  NAND2_X1 U14430 ( .A1(n13950), .A2(n13905), .ZN(n11926) );
  NAND2_X1 U14431 ( .A1(n11927), .A2(n11926), .ZN(n14393) );
  AOI21_X1 U14432 ( .B1(n13919), .B2(n14393), .A(n11928), .ZN(n11929) );
  OAI21_X1 U14433 ( .B1(n14397), .B2(n13921), .A(n11929), .ZN(n11930) );
  AOI21_X1 U14434 ( .B1(n14575), .B2(n13923), .A(n11930), .ZN(n11931) );
  OAI21_X1 U14435 ( .B1(n11932), .B2(n13925), .A(n11931), .ZN(P2_U3203) );
  OAI22_X1 U14436 ( .A1(n14285), .A2(n10435), .B1(n13958), .B2(n14398), .ZN(
        n11933) );
  AOI21_X1 U14437 ( .B1(n14368), .B2(n11934), .A(n11933), .ZN(n11935) );
  OAI21_X1 U14438 ( .B1(n14370), .B2(n11936), .A(n11935), .ZN(n11937) );
  AOI21_X1 U14439 ( .B1(n14312), .B2(n11938), .A(n11937), .ZN(n11939) );
  OAI21_X1 U14440 ( .B1(n6557), .B2(n11940), .A(n11939), .ZN(P2_U3263) );
  NAND2_X1 U14441 ( .A1(n11943), .A2(n11949), .ZN(n11941) );
  NAND2_X1 U14442 ( .A1(n11942), .A2(n11941), .ZN(n11946) );
  INV_X1 U14443 ( .A(n11943), .ZN(n11944) );
  NAND2_X1 U14444 ( .A1(n11944), .A2(n13112), .ZN(n11945) );
  XNOR2_X1 U14445 ( .A(n12113), .B(n12995), .ZN(n12919) );
  XNOR2_X1 U14446 ( .A(n12919), .B(n13059), .ZN(n11947) );
  NAND2_X1 U14447 ( .A1(n13096), .A2(n12106), .ZN(n11948) );
  NAND2_X1 U14448 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n13151)
         );
  OAI211_X1 U14449 ( .C1(n11949), .C2(n13099), .A(n11948), .B(n13151), .ZN(
        n11950) );
  AOI21_X1 U14450 ( .B1(n12110), .B2(n13095), .A(n11950), .ZN(n11952) );
  NAND2_X1 U14451 ( .A1(n12113), .A2(n13102), .ZN(n11951) );
  OAI211_X1 U14452 ( .C1(n11953), .C2(n13104), .A(n11952), .B(n11951), .ZN(
        P3_U3164) );
  XNOR2_X1 U14453 ( .A(n11954), .B(n11955), .ZN(n15726) );
  OAI22_X1 U14454 ( .A1(n14399), .A2(n8148), .B1(n14398), .B2(n11956), .ZN(
        n11960) );
  OAI211_X1 U14455 ( .C1(n8149), .C2(n8148), .A(n14470), .B(n11958), .ZN(
        n15723) );
  NOR2_X1 U14456 ( .A1(n14370), .A2(n15723), .ZN(n11959) );
  AOI211_X1 U14457 ( .C1(n15726), .C2(n14312), .A(n11960), .B(n11959), .ZN(
        n11967) );
  XNOR2_X1 U14458 ( .A(n11961), .B(n11962), .ZN(n11964) );
  AOI21_X1 U14459 ( .B1(n11964), .B2(n15662), .A(n11963), .ZN(n15724) );
  MUX2_X1 U14460 ( .A(n11965), .B(n15724), .S(n14285), .Z(n11966) );
  NAND2_X1 U14461 ( .A1(n11967), .A2(n11966), .ZN(P2_U3260) );
  OAI21_X1 U14462 ( .B1(n8452), .B2(n11969), .A(n11968), .ZN(n15712) );
  OAI22_X1 U14463 ( .A1(n14399), .A2(n15707), .B1(n14398), .B2(n8438), .ZN(
        n11972) );
  OAI211_X1 U14464 ( .C1(n15707), .C2(n15660), .A(n14470), .B(n11970), .ZN(
        n15706) );
  NOR2_X1 U14465 ( .A1(n14370), .A2(n15706), .ZN(n11971) );
  AOI211_X1 U14466 ( .C1(n14312), .C2(n15712), .A(n11972), .B(n11971), .ZN(
        n11979) );
  OAI21_X1 U14467 ( .B1(n11974), .B2(n8691), .A(n11973), .ZN(n11976) );
  AOI21_X1 U14468 ( .B1(n11976), .B2(n15662), .A(n11975), .ZN(n15708) );
  MUX2_X1 U14469 ( .A(n11977), .B(n15708), .S(n14285), .Z(n11978) );
  NAND2_X1 U14470 ( .A1(n11979), .A2(n11978), .ZN(P2_U3264) );
  INV_X1 U14471 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n16026) );
  INV_X1 U14472 ( .A(n12999), .ZN(n11980) );
  NAND2_X1 U14473 ( .A1(n11980), .A2(P3_U3897), .ZN(n11981) );
  OAI21_X1 U14474 ( .B1(n13115), .B2(n16026), .A(n11981), .ZN(P3_U3520) );
  MUX2_X1 U14475 ( .A(n11983), .B(n11982), .S(n15804), .Z(n11984) );
  OAI21_X1 U14476 ( .B1(n13610), .B2(n11985), .A(n11984), .ZN(P3_U3468) );
  XNOR2_X1 U14477 ( .A(n14383), .B(n11992), .ZN(n15739) );
  INV_X1 U14478 ( .A(n11987), .ZN(n11988) );
  OAI211_X1 U14479 ( .C1(n7511), .C2(n6826), .A(n11988), .B(n14470), .ZN(
        n15735) );
  NOR2_X1 U14480 ( .A1(n15735), .A2(n14370), .ZN(n11991) );
  OAI22_X1 U14481 ( .A1(n14399), .A2(n7511), .B1(n14398), .B2(n11989), .ZN(
        n11990) );
  AOI211_X1 U14482 ( .C1(n15739), .C2(n14312), .A(n11991), .B(n11990), .ZN(
        n11998) );
  XNOR2_X1 U14483 ( .A(n11993), .B(n11992), .ZN(n11995) );
  AOI21_X1 U14484 ( .B1(n11995), .B2(n15662), .A(n11994), .ZN(n15736) );
  MUX2_X1 U14485 ( .A(n11996), .B(n15736), .S(n14285), .Z(n11997) );
  NAND2_X1 U14486 ( .A1(n11998), .A2(n11997), .ZN(P2_U3258) );
  MUX2_X1 U14487 ( .A(n13136), .B(n11999), .S(n15804), .Z(n12002) );
  INV_X1 U14488 ( .A(n13617), .ZN(n13602) );
  NAND2_X1 U14489 ( .A1(n12000), .A2(n13602), .ZN(n12001) );
  OAI211_X1 U14490 ( .C1(n13610), .C2(n12003), .A(n12002), .B(n12001), .ZN(
        P3_U3470) );
  INV_X1 U14491 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n15973) );
  INV_X1 U14492 ( .A(n12004), .ZN(n12005) );
  NAND2_X1 U14493 ( .A1(n12005), .A2(P3_U3897), .ZN(n12006) );
  OAI21_X1 U14494 ( .B1(n13115), .B2(n15973), .A(n12006), .ZN(P3_U3521) );
  NAND2_X1 U14495 ( .A1(n12007), .A2(n12393), .ZN(n12010) );
  AOI22_X1 U14496 ( .A1(n12855), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n12008), 
        .B2(n12294), .ZN(n12009) );
  INV_X1 U14497 ( .A(n14781), .ZN(n12214) );
  NAND2_X1 U14498 ( .A1(n15331), .A2(n12214), .ZN(n12011) );
  OR2_X1 U14499 ( .A1(n15336), .A2(n14782), .ZN(n12091) );
  INV_X1 U14500 ( .A(n12091), .ZN(n12093) );
  AOI21_X1 U14501 ( .B1(n12012), .B2(n12882), .A(n12093), .ZN(n12013) );
  XOR2_X1 U14502 ( .A(n12885), .B(n12013), .Z(n15333) );
  NAND2_X1 U14503 ( .A1(n12016), .A2(n12885), .ZN(n12069) );
  OAI211_X1 U14504 ( .C1(n12885), .C2(n12016), .A(n12069), .B(n15552), .ZN(
        n12021) );
  NAND2_X1 U14505 ( .A1(n12448), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n12020) );
  INV_X1 U14506 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n12080) );
  XNOR2_X1 U14507 ( .A(n12081), .B(n12080), .ZN(n12232) );
  OR2_X1 U14508 ( .A1(n11447), .A2(n12232), .ZN(n12019) );
  NAND2_X1 U14509 ( .A1(n11451), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n12018) );
  NAND2_X1 U14510 ( .A1(n12410), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n12017) );
  NAND4_X1 U14511 ( .A1(n12020), .A2(n12019), .A3(n12018), .A4(n12017), .ZN(
        n14780) );
  AOI22_X1 U14512 ( .A1(n15180), .A2(n14782), .B1(n14780), .B2(n15178), .ZN(
        n12145) );
  NAND2_X1 U14513 ( .A1(n12021), .A2(n12145), .ZN(n15329) );
  NAND2_X1 U14514 ( .A1(n15329), .A2(n15097), .ZN(n12027) );
  AOI211_X1 U14515 ( .C1(n15331), .C2(n12022), .A(n15538), .B(n12169), .ZN(
        n15330) );
  INV_X1 U14516 ( .A(n15331), .ZN(n12150) );
  INV_X1 U14517 ( .A(n12023), .ZN(n12147) );
  AOI22_X1 U14518 ( .A1(n15512), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n12147), 
        .B2(n15513), .ZN(n12024) );
  OAI21_X1 U14519 ( .B1(n12150), .B2(n15147), .A(n12024), .ZN(n12025) );
  AOI21_X1 U14520 ( .B1(n15330), .B2(n15521), .A(n12025), .ZN(n12026) );
  OAI211_X1 U14521 ( .C1(n15333), .C2(n15195), .A(n12027), .B(n12026), .ZN(
        P1_U3282) );
  XNOR2_X1 U14522 ( .A(n14367), .B(n12649), .ZN(n12596) );
  NAND2_X1 U14523 ( .A1(n13948), .A2(n12612), .ZN(n12597) );
  XNOR2_X1 U14524 ( .A(n12596), .B(n12597), .ZN(n12600) );
  XNOR2_X1 U14525 ( .A(n12601), .B(n12600), .ZN(n12036) );
  OR2_X1 U14526 ( .A1(n13812), .A2(n13917), .ZN(n12031) );
  NAND2_X1 U14527 ( .A1(n13949), .A2(n13905), .ZN(n12030) );
  NAND2_X1 U14528 ( .A1(n12031), .A2(n12030), .ZN(n14377) );
  NAND2_X1 U14529 ( .A1(n13919), .A2(n14377), .ZN(n12032) );
  OAI211_X1 U14530 ( .C1(n13921), .C2(n14365), .A(n12033), .B(n12032), .ZN(
        n12034) );
  AOI21_X1 U14531 ( .B1(n14367), .B2(n13923), .A(n12034), .ZN(n12035) );
  OAI21_X1 U14532 ( .B1(n12036), .B2(n13925), .A(n12035), .ZN(P2_U3189) );
  INV_X1 U14533 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14049) );
  INV_X1 U14534 ( .A(n12039), .ZN(n12040) );
  XNOR2_X1 U14535 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(P3_ADDR_REG_12__SCAN_IN), 
        .ZN(n12044) );
  XNOR2_X1 U14536 ( .A(n12196), .B(n12044), .ZN(n12046) );
  INV_X1 U14537 ( .A(n12046), .ZN(n12047) );
  NAND2_X1 U14538 ( .A1(n12193), .A2(n12194), .ZN(n12048) );
  XNOR2_X1 U14539 ( .A(n12048), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  INV_X1 U14540 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16061) );
  NAND2_X1 U14541 ( .A1(n12049), .A2(n13115), .ZN(n12050) );
  OAI21_X1 U14542 ( .B1(P3_U3897), .B2(n16061), .A(n12050), .ZN(P3_U3522) );
  MUX2_X1 U14543 ( .A(n13133), .B(n12051), .S(n15804), .Z(n12052) );
  OAI21_X1 U14544 ( .B1(n13610), .B2(n12053), .A(n12052), .ZN(P3_U3469) );
  INV_X1 U14545 ( .A(n12054), .ZN(n12056) );
  OAI222_X1 U14546 ( .A1(P3_U3151), .A2(n12057), .B1(n13721), .B2(n12056), 
        .C1(n12055), .C2(n13723), .ZN(P3_U3269) );
  XNOR2_X1 U14547 ( .A(n12058), .B(n12880), .ZN(n15589) );
  INV_X1 U14548 ( .A(n12059), .ZN(n12064) );
  INV_X1 U14549 ( .A(n12061), .ZN(n12062) );
  AOI211_X1 U14550 ( .C1(n12063), .C2(n12060), .A(n15558), .B(n12062), .ZN(
        n15596) );
  AOI211_X1 U14551 ( .C1(n15513), .C2(n12064), .A(n15590), .B(n15596), .ZN(
        n12065) );
  MUX2_X1 U14552 ( .A(n10290), .B(n12065), .S(n15097), .Z(n12068) );
  INV_X1 U14553 ( .A(n12066), .ZN(n15518) );
  AOI211_X1 U14554 ( .C1(n12724), .C2(n15518), .A(n15538), .B(n15502), .ZN(
        n15595) );
  AOI22_X1 U14555 ( .A1(n15595), .A2(n15521), .B1(n15515), .B2(n12724), .ZN(
        n12067) );
  OAI211_X1 U14556 ( .C1(n15195), .C2(n15589), .A(n12068), .B(n12067), .ZN(
        P1_U3285) );
  NAND2_X1 U14557 ( .A1(n12069), .A2(n12075), .ZN(n12074) );
  NAND2_X1 U14558 ( .A1(n12070), .A2(n12393), .ZN(n12073) );
  AOI22_X1 U14559 ( .A1(n12071), .A2(n12294), .B1(n12855), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n12072) );
  NAND2_X2 U14560 ( .A1(n12073), .A2(n12072), .ZN(n12745) );
  NAND3_X1 U14561 ( .A1(n12069), .A2(n12175), .A3(n12075), .ZN(n12076) );
  NAND3_X1 U14562 ( .A1(n12152), .A2(n15552), .A3(n12076), .ZN(n12089) );
  NAND2_X1 U14563 ( .A1(n14781), .A2(n15180), .ZN(n12088) );
  NAND2_X1 U14564 ( .A1(n12448), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n12086) );
  INV_X1 U14565 ( .A(n12081), .ZN(n12078) );
  INV_X1 U14566 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n12079) );
  OAI21_X1 U14567 ( .B1(n12081), .B2(n12080), .A(n12079), .ZN(n12082) );
  NAND2_X1 U14568 ( .A1(n12159), .A2(n12082), .ZN(n14717) );
  OR2_X1 U14569 ( .A1(n11447), .A2(n14717), .ZN(n12085) );
  NAND2_X1 U14570 ( .A1(n11031), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n12084) );
  NAND2_X1 U14571 ( .A1(n12410), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n12083) );
  NAND4_X1 U14572 ( .A1(n12086), .A2(n12085), .A3(n12084), .A4(n12083), .ZN(
        n15181) );
  NAND2_X1 U14573 ( .A1(n15181), .A2(n15178), .ZN(n12087) );
  AND2_X1 U14574 ( .A1(n12088), .A2(n12087), .ZN(n12234) );
  NAND2_X1 U14575 ( .A1(n12089), .A2(n12234), .ZN(n15328) );
  INV_X1 U14576 ( .A(n15328), .ZN(n12102) );
  NOR2_X1 U14577 ( .A1(n12882), .A2(n12093), .ZN(n12094) );
  NOR2_X1 U14578 ( .A1(n12885), .A2(n12094), .ZN(n12095) );
  XNOR2_X1 U14579 ( .A(n12176), .B(n12175), .ZN(n15323) );
  XNOR2_X1 U14580 ( .A(n12169), .B(n12745), .ZN(n12096) );
  NAND2_X1 U14581 ( .A1(n12096), .A2(n15517), .ZN(n15324) );
  OAI22_X1 U14582 ( .A1(n15097), .A2(n12097), .B1(n12232), .B2(n15189), .ZN(
        n12098) );
  AOI21_X1 U14583 ( .B1(n12745), .B2(n15515), .A(n12098), .ZN(n12099) );
  OAI21_X1 U14584 ( .B1(n15324), .B2(n15082), .A(n12099), .ZN(n12100) );
  AOI21_X1 U14585 ( .B1(n15323), .B2(n15101), .A(n12100), .ZN(n12101) );
  OAI21_X1 U14586 ( .B1(n12102), .B2(n15512), .A(n12101), .ZN(P1_U3281) );
  XNOR2_X1 U14587 ( .A(n12104), .B(n12103), .ZN(n12114) );
  XNOR2_X1 U14588 ( .A(n12105), .B(n6890), .ZN(n12107) );
  AOI222_X1 U14589 ( .A1(n13552), .A2(n12107), .B1(n12106), .B2(n13547), .C1(
        n13112), .C2(n13549), .ZN(n12118) );
  MUX2_X1 U14590 ( .A(n15909), .B(n12118), .S(n15804), .Z(n12109) );
  NAND2_X1 U14591 ( .A1(n12113), .A2(n13614), .ZN(n12108) );
  OAI211_X1 U14592 ( .C1(n13617), .C2(n12114), .A(n12109), .B(n12108), .ZN(
        P3_U3471) );
  MUX2_X1 U14593 ( .A(n13162), .B(n12118), .S(n13553), .Z(n12112) );
  AOI22_X1 U14594 ( .A1(n12113), .A2(n13558), .B1(n13557), .B2(n12110), .ZN(
        n12111) );
  OAI211_X1 U14595 ( .C1(n12114), .C2(n13561), .A(n12112), .B(n12111), .ZN(
        P3_U3221) );
  AOI22_X1 U14596 ( .A1(n12113), .A2(n13695), .B1(P3_REG0_REG_12__SCAN_IN), 
        .B2(n15788), .ZN(n12117) );
  INV_X1 U14597 ( .A(n12114), .ZN(n12115) );
  NAND2_X1 U14598 ( .A1(n12115), .A2(n13673), .ZN(n12116) );
  OAI211_X1 U14599 ( .C1(n12118), .C2(n15788), .A(n12117), .B(n12116), .ZN(
        P3_U3426) );
  INV_X1 U14600 ( .A(n12372), .ZN(n12587) );
  OAI222_X1 U14601 ( .A1(P2_U3088), .A2(n12119), .B1(n14594), .B2(n12587), 
        .C1(n16023), .C2(n14590), .ZN(P2_U3301) );
  NAND2_X1 U14602 ( .A1(n15331), .A2(n6553), .ZN(n12121) );
  NAND2_X1 U14603 ( .A1(n14781), .A2(n6554), .ZN(n12120) );
  NAND2_X1 U14604 ( .A1(n12121), .A2(n12120), .ZN(n12122) );
  XNOR2_X1 U14605 ( .A(n12122), .B(n11860), .ZN(n12223) );
  AOI22_X1 U14606 ( .A1(n15331), .A2(n6554), .B1(n12572), .B2(n14781), .ZN(
        n12221) );
  XNOR2_X1 U14607 ( .A(n12223), .B(n12221), .ZN(n12142) );
  NAND2_X1 U14608 ( .A1(n15499), .A2(n6554), .ZN(n12126) );
  NAND2_X1 U14609 ( .A1(n12572), .A2(n14783), .ZN(n12125) );
  NAND2_X1 U14610 ( .A1(n15499), .A2(n6553), .ZN(n12128) );
  NAND2_X1 U14611 ( .A1(n14783), .A2(n6554), .ZN(n12127) );
  NAND2_X1 U14612 ( .A1(n12128), .A2(n12127), .ZN(n12129) );
  XNOR2_X1 U14613 ( .A(n12129), .B(n12534), .ZN(n12184) );
  NAND2_X1 U14614 ( .A1(n15336), .A2(n6553), .ZN(n12131) );
  NAND2_X1 U14615 ( .A1(n14782), .A2(n6554), .ZN(n12130) );
  NAND2_X1 U14616 ( .A1(n12131), .A2(n12130), .ZN(n12132) );
  XNOR2_X1 U14617 ( .A(n12132), .B(n11860), .ZN(n12207) );
  NAND2_X1 U14618 ( .A1(n15336), .A2(n6554), .ZN(n12135) );
  NAND2_X1 U14619 ( .A1(n12572), .A2(n14782), .ZN(n12134) );
  NAND2_X1 U14620 ( .A1(n12135), .A2(n12134), .ZN(n12206) );
  NOR2_X1 U14621 ( .A1(n12207), .A2(n12206), .ZN(n12205) );
  AOI21_X1 U14622 ( .B1(n12183), .B2(n12184), .A(n12205), .ZN(n12140) );
  INV_X1 U14623 ( .A(n12184), .ZN(n12209) );
  INV_X1 U14624 ( .A(n12183), .ZN(n12208) );
  AOI21_X1 U14625 ( .B1(n12209), .B2(n12208), .A(n12206), .ZN(n12138) );
  INV_X1 U14626 ( .A(n12207), .ZN(n12137) );
  NAND3_X1 U14627 ( .A1(n12209), .A2(n12208), .A3(n12206), .ZN(n12136) );
  OAI21_X1 U14628 ( .B1(n12138), .B2(n12137), .A(n12136), .ZN(n12139) );
  OAI21_X1 U14629 ( .B1(n12142), .B2(n12141), .A(n12225), .ZN(n12143) );
  NAND2_X1 U14630 ( .A1(n12143), .A2(n14753), .ZN(n12149) );
  OAI21_X1 U14631 ( .B1(n14737), .B2(n12145), .A(n12144), .ZN(n12146) );
  AOI21_X1 U14632 ( .B1(n12147), .B2(n14690), .A(n12146), .ZN(n12148) );
  OAI211_X1 U14633 ( .C1(n12150), .C2(n14765), .A(n12149), .B(n12148), .ZN(
        P1_U3236) );
  INV_X1 U14634 ( .A(n14780), .ZN(n14716) );
  OR2_X1 U14635 ( .A1(n12745), .A2(n14716), .ZN(n12151) );
  INV_X1 U14636 ( .A(n12249), .ZN(n12156) );
  NAND2_X1 U14637 ( .A1(n12153), .A2(n12393), .ZN(n12155) );
  AOI22_X1 U14638 ( .A1(n14859), .A2(n12294), .B1(n12855), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n12154) );
  XNOR2_X1 U14639 ( .A(n15319), .B(n12754), .ZN(n12888) );
  AOI21_X1 U14640 ( .B1(n12156), .B2(n12888), .A(n15558), .ZN(n12168) );
  INV_X1 U14641 ( .A(n12888), .ZN(n12179) );
  NAND2_X1 U14642 ( .A1(n12249), .A2(n12179), .ZN(n15162) );
  OR2_X2 U14643 ( .A1(n12159), .A2(n15981), .ZN(n12254) );
  NAND2_X1 U14644 ( .A1(n12159), .A2(n15981), .ZN(n12160) );
  AND2_X1 U14645 ( .A1(n12254), .A2(n12160), .ZN(n15188) );
  NAND2_X1 U14646 ( .A1(n12158), .A2(n15188), .ZN(n12166) );
  INV_X1 U14647 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n15191) );
  OR2_X1 U14648 ( .A1(n12161), .A2(n15191), .ZN(n12165) );
  INV_X1 U14649 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14852) );
  OR2_X1 U14650 ( .A1(n12413), .A2(n14852), .ZN(n12164) );
  INV_X1 U14651 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n12162) );
  OR2_X1 U14652 ( .A1(n10700), .A2(n12162), .ZN(n12163) );
  OAI22_X1 U14653 ( .A1(n14716), .A2(n15128), .B1(n14758), .B2(n15130), .ZN(
        n12167) );
  AOI21_X1 U14654 ( .B1(n12168), .B2(n15162), .A(n12167), .ZN(n15321) );
  INV_X1 U14655 ( .A(n12745), .ZN(n15325) );
  INV_X1 U14656 ( .A(n12170), .ZN(n12172) );
  NAND2_X1 U14657 ( .A1(n12170), .A2(n14723), .ZN(n15175) );
  INV_X1 U14658 ( .A(n15175), .ZN(n12171) );
  AOI211_X1 U14659 ( .C1(n15319), .C2(n12172), .A(n15538), .B(n12171), .ZN(
        n15318) );
  INV_X1 U14660 ( .A(n14717), .ZN(n12173) );
  AOI22_X1 U14661 ( .A1(n15525), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n12173), 
        .B2(n15513), .ZN(n12174) );
  OAI21_X1 U14662 ( .B1(n14723), .B2(n15147), .A(n12174), .ZN(n12181) );
  OR2_X1 U14663 ( .A1(n12745), .A2(n14780), .ZN(n12177) );
  XNOR2_X1 U14664 ( .A(n12416), .B(n12179), .ZN(n15322) );
  NOR2_X1 U14665 ( .A1(n15322), .A2(n15195), .ZN(n12180) );
  AOI211_X1 U14666 ( .C1(n15318), .C2(n15521), .A(n12181), .B(n12180), .ZN(
        n12182) );
  OAI21_X1 U14667 ( .B1(n15321), .B2(n15512), .A(n12182), .ZN(P1_U3280) );
  XNOR2_X1 U14668 ( .A(n6614), .B(n12183), .ZN(n12210) );
  XNOR2_X1 U14669 ( .A(n12210), .B(n12184), .ZN(n12185) );
  NAND2_X1 U14670 ( .A1(n12185), .A2(n14753), .ZN(n12191) );
  INV_X1 U14671 ( .A(n12186), .ZN(n15498) );
  NAND2_X1 U14672 ( .A1(n14784), .A2(n15180), .ZN(n12188) );
  NAND2_X1 U14673 ( .A1(n14782), .A2(n15178), .ZN(n12187) );
  AND2_X1 U14674 ( .A1(n12188), .A2(n12187), .ZN(n15495) );
  NAND2_X1 U14675 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n14839) );
  OAI21_X1 U14676 ( .B1(n14737), .B2(n15495), .A(n14839), .ZN(n12189) );
  AOI21_X1 U14677 ( .B1(n15498), .B2(n14690), .A(n12189), .ZN(n12190) );
  OAI211_X1 U14678 ( .C1(n15600), .C2(n14765), .A(n12191), .B(n12190), .ZN(
        P1_U3231) );
  INV_X1 U14679 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n13152) );
  NAND2_X1 U14680 ( .A1(n13152), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n12195) );
  NAND2_X1 U14681 ( .A1(n12196), .A2(n12195), .ZN(n12199) );
  NAND2_X1 U14682 ( .A1(n12197), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n12198) );
  NAND2_X1 U14683 ( .A1(n12199), .A2(n12198), .ZN(n15394) );
  INV_X1 U14684 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n12200) );
  NAND2_X1 U14685 ( .A1(n12200), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n15395) );
  INV_X1 U14686 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n13179) );
  NAND2_X1 U14687 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n13179), .ZN(n15393) );
  NAND2_X1 U14688 ( .A1(n15395), .A2(n15393), .ZN(n12201) );
  XNOR2_X1 U14689 ( .A(n15394), .B(n12201), .ZN(n12202) );
  NAND2_X1 U14690 ( .A1(n12203), .A2(n12202), .ZN(n15391) );
  NAND2_X1 U14691 ( .A1(n15390), .A2(n15391), .ZN(n12204) );
  XNOR2_X1 U14692 ( .A(n12204), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  AOI21_X1 U14693 ( .B1(n12207), .B2(n12206), .A(n12205), .ZN(n12212) );
  AOI22_X1 U14694 ( .A1(n12210), .A2(n12209), .B1(n6614), .B2(n12208), .ZN(
        n12211) );
  XOR2_X1 U14695 ( .A(n12212), .B(n12211), .Z(n12220) );
  OAI21_X1 U14696 ( .B1(n14706), .B2(n12214), .A(n12213), .ZN(n12218) );
  OAI22_X1 U14697 ( .A1(n14759), .A2(n12216), .B1(n12215), .B2(n14715), .ZN(
        n12217) );
  AOI211_X1 U14698 ( .C1(n14740), .C2(n15336), .A(n12218), .B(n12217), .ZN(
        n12219) );
  OAI21_X1 U14699 ( .B1(n12220), .B2(n14742), .A(n12219), .ZN(P1_U3217) );
  INV_X1 U14700 ( .A(n12221), .ZN(n12222) );
  OR2_X1 U14701 ( .A1(n12223), .A2(n12222), .ZN(n12224) );
  AOI22_X1 U14702 ( .A1(n12745), .A2(n6553), .B1(n12552), .B2(n14780), .ZN(
        n12226) );
  XNOR2_X1 U14703 ( .A(n12226), .B(n11860), .ZN(n12469) );
  NOR2_X1 U14704 ( .A1(n14636), .A2(n14716), .ZN(n12227) );
  AOI21_X1 U14705 ( .B1(n12745), .B2(n12552), .A(n12227), .ZN(n12470) );
  XNOR2_X1 U14706 ( .A(n12469), .B(n12470), .ZN(n12229) );
  AOI21_X1 U14707 ( .B1(n12228), .B2(n12229), .A(n14742), .ZN(n12231) );
  INV_X1 U14708 ( .A(n12229), .ZN(n12230) );
  NAND2_X1 U14709 ( .A1(n12231), .A2(n12474), .ZN(n12238) );
  INV_X1 U14710 ( .A(n12232), .ZN(n12236) );
  OAI21_X1 U14711 ( .B1(n14737), .B2(n12234), .A(n12233), .ZN(n12235) );
  AOI21_X1 U14712 ( .B1(n12236), .B2(n14690), .A(n12235), .ZN(n12237) );
  OAI211_X1 U14713 ( .C1(n15325), .C2(n14765), .A(n12238), .B(n12237), .ZN(
        P1_U3224) );
  INV_X1 U14714 ( .A(n12394), .ZN(n15378) );
  INV_X1 U14715 ( .A(n12240), .ZN(n12243) );
  OAI222_X1 U14716 ( .A1(n13721), .A2(n12243), .B1(n12242), .B2(P3_U3151), 
        .C1(n12241), .C2(n13723), .ZN(P3_U3266) );
  AOI22_X1 U14717 ( .A1(n14868), .A2(n12294), .B1(n12855), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n12245) );
  NAND2_X1 U14718 ( .A1(n15319), .A2(n12754), .ZN(n12246) );
  NOR2_X1 U14719 ( .A1(n15319), .A2(n12754), .ZN(n15160) );
  NAND2_X1 U14720 ( .A1(n12757), .A2(n15160), .ZN(n12247) );
  AOI22_X1 U14721 ( .A1(n15484), .A2(n12294), .B1(n12855), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n12251) );
  NAND2_X1 U14722 ( .A1(n12254), .A2(n12253), .ZN(n12255) );
  NAND2_X1 U14723 ( .A1(n12265), .A2(n12255), .ZN(n15171) );
  NAND2_X1 U14724 ( .A1(n12448), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n12256) );
  OAI21_X1 U14725 ( .B1(n15171), .B2(n11447), .A(n12256), .ZN(n12260) );
  INV_X1 U14726 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n12258) );
  NAND2_X1 U14727 ( .A1(n12410), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n12257) );
  OAI21_X1 U14728 ( .B1(n12258), .B2(n12413), .A(n12257), .ZN(n12259) );
  NAND2_X1 U14729 ( .A1(n15308), .A2(n14681), .ZN(n12761) );
  NAND2_X1 U14730 ( .A1(n12261), .A2(n12393), .ZN(n12263) );
  AOI22_X1 U14731 ( .A1(n12855), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n12294), 
        .B2(n14887), .ZN(n12262) );
  INV_X1 U14732 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n12269) );
  INV_X1 U14733 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n12264) );
  NAND2_X1 U14734 ( .A1(n12265), .A2(n12264), .ZN(n12266) );
  NAND2_X1 U14735 ( .A1(n12276), .A2(n12266), .ZN(n15144) );
  OR2_X1 U14736 ( .A1(n15144), .A2(n11447), .ZN(n12268) );
  AOI22_X1 U14737 ( .A1(n12410), .A2(P1_REG0_REG_16__SCAN_IN), .B1(n11451), 
        .B2(P1_REG1_REG_16__SCAN_IN), .ZN(n12267) );
  OAI211_X1 U14738 ( .C1(n12161), .C2(n12269), .A(n12268), .B(n12267), .ZN(
        n14778) );
  INV_X1 U14739 ( .A(n14778), .ZN(n15129) );
  XNOR2_X1 U14740 ( .A(n15302), .B(n15129), .ZN(n15149) );
  NAND2_X1 U14741 ( .A1(n15302), .A2(n15129), .ZN(n12271) );
  NAND2_X1 U14742 ( .A1(n12272), .A2(n12393), .ZN(n12274) );
  AOI22_X1 U14743 ( .A1(n12855), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n12294), 
        .B2(n14902), .ZN(n12273) );
  NAND2_X2 U14744 ( .A1(n12274), .A2(n12273), .ZN(n15298) );
  NAND2_X1 U14745 ( .A1(n12276), .A2(n12275), .ZN(n12277) );
  AND2_X1 U14746 ( .A1(n12286), .A2(n12277), .ZN(n15135) );
  NAND2_X1 U14747 ( .A1(n15135), .A2(n12158), .ZN(n12280) );
  AOI22_X1 U14748 ( .A1(n12448), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n11451), 
        .B2(P1_REG1_REG_17__SCAN_IN), .ZN(n12279) );
  NAND2_X1 U14749 ( .A1(n12410), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n12278) );
  XNOR2_X1 U14750 ( .A(n15298), .B(n14680), .ZN(n15126) );
  OR2_X1 U14751 ( .A1(n15298), .A2(n14680), .ZN(n12767) );
  NAND2_X1 U14752 ( .A1(n12282), .A2(n12393), .ZN(n12284) );
  AOI22_X1 U14753 ( .A1(n12855), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n12294), 
        .B2(n15808), .ZN(n12283) );
  INV_X1 U14754 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n12285) );
  NAND2_X1 U14755 ( .A1(n12286), .A2(n12285), .ZN(n12287) );
  NAND2_X1 U14756 ( .A1(n12304), .A2(n12287), .ZN(n15116) );
  OR2_X1 U14757 ( .A1(n15116), .A2(n11447), .ZN(n12292) );
  INV_X1 U14758 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n16098) );
  NAND2_X1 U14759 ( .A1(n12448), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n12289) );
  NAND2_X1 U14760 ( .A1(n11451), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n12288) );
  OAI211_X1 U14761 ( .C1(n16098), .C2(n10700), .A(n12289), .B(n12288), .ZN(
        n12290) );
  INV_X1 U14762 ( .A(n12290), .ZN(n12291) );
  NAND2_X1 U14763 ( .A1(n15294), .A2(n15131), .ZN(n12780) );
  NAND2_X1 U14764 ( .A1(n12779), .A2(n12780), .ZN(n15105) );
  INV_X1 U14765 ( .A(n15105), .ZN(n15109) );
  NAND2_X1 U14766 ( .A1(n12293), .A2(n12393), .ZN(n12296) );
  AOI22_X1 U14767 ( .A1(n12855), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n12672), 
        .B2(n12294), .ZN(n12295) );
  XNOR2_X1 U14768 ( .A(n12304), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n15091) );
  INV_X1 U14769 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n15807) );
  NAND2_X1 U14770 ( .A1(n12410), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n12298) );
  NAND2_X1 U14771 ( .A1(n12448), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n12297) );
  OAI211_X1 U14772 ( .C1(n12413), .C2(n15807), .A(n12298), .B(n12297), .ZN(
        n12299) );
  AOI21_X1 U14773 ( .B1(n15091), .B2(n12158), .A(n12299), .ZN(n15070) );
  INV_X1 U14774 ( .A(n15070), .ZN(n14776) );
  NAND2_X1 U14775 ( .A1(n6576), .A2(n12785), .ZN(n15100) );
  INV_X1 U14776 ( .A(n12785), .ZN(n12300) );
  NAND2_X1 U14777 ( .A1(n12855), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12302) );
  INV_X1 U14778 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n12303) );
  OAI21_X1 U14779 ( .B1(n12304), .B2(n12303), .A(n14705), .ZN(n12305) );
  AND2_X1 U14780 ( .A1(n12305), .A2(n12316), .ZN(n15079) );
  NAND2_X1 U14781 ( .A1(n15079), .A2(n12158), .ZN(n12310) );
  INV_X1 U14782 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n16014) );
  NAND2_X1 U14783 ( .A1(n12448), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n12307) );
  NAND2_X1 U14784 ( .A1(n12410), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n12306) );
  OAI211_X1 U14785 ( .C1(n12413), .C2(n16014), .A(n12307), .B(n12306), .ZN(
        n12308) );
  INV_X1 U14786 ( .A(n12308), .ZN(n12309) );
  OR2_X1 U14787 ( .A1(n15278), .A2(n15090), .ZN(n12311) );
  NAND2_X1 U14788 ( .A1(n12312), .A2(n12393), .ZN(n12314) );
  NAND2_X1 U14789 ( .A1(n12855), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12313) );
  INV_X1 U14790 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n15949) );
  NAND2_X1 U14791 ( .A1(n12316), .A2(n15949), .ZN(n12317) );
  AND2_X1 U14792 ( .A1(n12330), .A2(n12317), .ZN(n15057) );
  NAND2_X1 U14793 ( .A1(n15057), .A2(n12158), .ZN(n12323) );
  INV_X1 U14794 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n12320) );
  NAND2_X1 U14795 ( .A1(n11451), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n12319) );
  NAND2_X1 U14796 ( .A1(n12448), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n12318) );
  OAI211_X1 U14797 ( .C1(n12320), .C2(n10700), .A(n12319), .B(n12318), .ZN(
        n12321) );
  INV_X1 U14798 ( .A(n12321), .ZN(n12322) );
  XNOR2_X1 U14799 ( .A(n15271), .B(n14775), .ZN(n15062) );
  NAND2_X1 U14800 ( .A1(n15059), .A2(n14775), .ZN(n12324) );
  OR2_X1 U14801 ( .A1(n12326), .A2(n12325), .ZN(n12327) );
  XNOR2_X1 U14802 ( .A(n12327), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15382) );
  INV_X1 U14803 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n16040) );
  NAND2_X1 U14804 ( .A1(n12330), .A2(n16040), .ZN(n12331) );
  NAND2_X1 U14805 ( .A1(n12343), .A2(n12331), .ZN(n15040) );
  INV_X1 U14806 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n12334) );
  NAND2_X1 U14807 ( .A1(n12448), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n12333) );
  NAND2_X1 U14808 ( .A1(n11031), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n12332) );
  OAI211_X1 U14809 ( .C1(n12334), .C2(n10700), .A(n12333), .B(n12332), .ZN(
        n12335) );
  INV_X1 U14810 ( .A(n12335), .ZN(n12336) );
  NAND2_X1 U14811 ( .A1(n15044), .A2(n15051), .ZN(n12338) );
  NAND2_X1 U14812 ( .A1(n12340), .A2(n12393), .ZN(n12342) );
  NAND2_X1 U14813 ( .A1(n12855), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12341) );
  INV_X1 U14814 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14614) );
  NAND2_X1 U14815 ( .A1(n12343), .A2(n14614), .ZN(n12344) );
  AND2_X1 U14816 ( .A1(n12363), .A2(n12344), .ZN(n15021) );
  NAND2_X1 U14817 ( .A1(n15021), .A2(n12158), .ZN(n12349) );
  INV_X1 U14818 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n16071) );
  NAND2_X1 U14819 ( .A1(n12410), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n12346) );
  NAND2_X1 U14820 ( .A1(n12448), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n12345) );
  OAI211_X1 U14821 ( .C1(n12413), .C2(n16071), .A(n12346), .B(n12345), .ZN(
        n12347) );
  INV_X1 U14822 ( .A(n12347), .ZN(n12348) );
  NAND2_X1 U14823 ( .A1(n12350), .A2(n11018), .ZN(n12352) );
  NAND2_X1 U14824 ( .A1(n12855), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12351) );
  INV_X1 U14825 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n12353) );
  NAND2_X1 U14826 ( .A1(n12365), .A2(n12353), .ZN(n12354) );
  NAND2_X1 U14827 ( .A1(n14995), .A2(n12158), .ZN(n12359) );
  INV_X1 U14828 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n15919) );
  NAND2_X1 U14829 ( .A1(n12448), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n12356) );
  NAND2_X1 U14830 ( .A1(n12410), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n12355) );
  OAI211_X1 U14831 ( .C1(n12413), .C2(n15919), .A(n12356), .B(n12355), .ZN(
        n12357) );
  INV_X1 U14832 ( .A(n12357), .ZN(n12358) );
  NAND2_X1 U14833 ( .A1(n12678), .A2(n14748), .ZN(n14968) );
  NAND2_X1 U14834 ( .A1(n12360), .A2(n11018), .ZN(n12362) );
  NAND2_X1 U14835 ( .A1(n12855), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12361) );
  INV_X1 U14836 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14699) );
  NAND2_X1 U14837 ( .A1(n12363), .A2(n14699), .ZN(n12364) );
  NAND2_X1 U14838 ( .A1(n12365), .A2(n12364), .ZN(n15012) );
  INV_X1 U14839 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n12368) );
  NAND2_X1 U14840 ( .A1(n12448), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n12367) );
  NAND2_X1 U14841 ( .A1(n11031), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n12366) );
  OAI211_X1 U14842 ( .C1(n12368), .C2(n10700), .A(n12367), .B(n12366), .ZN(
        n12369) );
  INV_X1 U14843 ( .A(n12369), .ZN(n12370) );
  NAND2_X2 U14844 ( .A1(n12371), .A2(n12370), .ZN(n14773) );
  NAND2_X1 U14845 ( .A1(n15253), .A2(n14989), .ZN(n12434) );
  INV_X1 U14846 ( .A(n14967), .ZN(n12384) );
  AOI21_X1 U14847 ( .B1(n14748), .B2(n14967), .A(n12678), .ZN(n12383) );
  NAND2_X1 U14848 ( .A1(n12372), .A2(n12393), .ZN(n12374) );
  NAND2_X1 U14849 ( .A1(n12855), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12373) );
  INV_X1 U14850 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14749) );
  NAND2_X1 U14851 ( .A1(n12375), .A2(n14749), .ZN(n12376) );
  NAND2_X1 U14852 ( .A1(n12400), .A2(n12376), .ZN(n14976) );
  INV_X1 U14853 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n12379) );
  NAND2_X1 U14854 ( .A1(n12448), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n12378) );
  NAND2_X1 U14855 ( .A1(n11451), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n12377) );
  OAI211_X1 U14856 ( .C1(n12379), .C2(n10700), .A(n12378), .B(n12377), .ZN(
        n12380) );
  INV_X1 U14857 ( .A(n12380), .ZN(n12381) );
  AOI211_X1 U14858 ( .C1(n12384), .C2(n14772), .A(n12383), .B(n14969), .ZN(
        n12385) );
  XNOR2_X1 U14859 ( .A(n12400), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n14958) );
  NAND2_X1 U14860 ( .A1(n14958), .A2(n12158), .ZN(n12392) );
  INV_X1 U14861 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n12389) );
  NAND2_X1 U14862 ( .A1(n12448), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n12388) );
  NAND2_X1 U14863 ( .A1(n12410), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n12387) );
  OAI211_X1 U14864 ( .C1(n12413), .C2(n12389), .A(n12388), .B(n12387), .ZN(
        n12390) );
  INV_X1 U14865 ( .A(n12390), .ZN(n12391) );
  NAND2_X1 U14866 ( .A1(n12394), .A2(n12393), .ZN(n12396) );
  NAND2_X1 U14867 ( .A1(n12855), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12395) );
  NAND2_X1 U14868 ( .A1(n12461), .A2(n11018), .ZN(n12398) );
  NAND2_X1 U14869 ( .A1(n12855), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12397) );
  INV_X1 U14870 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n12580) );
  INV_X1 U14871 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n14642) );
  OAI21_X1 U14872 ( .B1(n12400), .B2(n12580), .A(n14642), .ZN(n12402) );
  NAND2_X1 U14873 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n12399) );
  INV_X1 U14874 ( .A(n12456), .ZN(n12401) );
  NAND2_X1 U14875 ( .A1(n12402), .A2(n12401), .ZN(n14944) );
  INV_X1 U14876 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n15876) );
  NAND2_X1 U14877 ( .A1(n12448), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n12404) );
  NAND2_X1 U14878 ( .A1(n11031), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n12403) );
  OAI211_X1 U14879 ( .C1(n15876), .C2(n10700), .A(n12404), .B(n12403), .ZN(
        n12405) );
  INV_X1 U14880 ( .A(n12405), .ZN(n12406) );
  NAND2_X1 U14881 ( .A1(n14586), .A2(n12393), .ZN(n12409) );
  NAND2_X1 U14882 ( .A1(n12855), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12408) );
  INV_X1 U14883 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n12414) );
  NAND2_X1 U14884 ( .A1(n12448), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n12412) );
  NAND2_X1 U14885 ( .A1(n12410), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n12411) );
  OAI211_X1 U14886 ( .C1(n12414), .C2(n12413), .A(n12412), .B(n12411), .ZN(
        n12415) );
  AOI21_X1 U14887 ( .B1(n12456), .B2(n12158), .A(n12415), .ZN(n14940) );
  INV_X1 U14888 ( .A(n14940), .ZN(n14768) );
  INV_X1 U14889 ( .A(n14758), .ZN(n14779) );
  NAND2_X1 U14890 ( .A1(n15314), .A2(n14779), .ZN(n12417) );
  OR2_X1 U14891 ( .A1(n15308), .A2(n15179), .ZN(n12418) );
  OR2_X1 U14892 ( .A1(n15302), .A2(n14778), .ZN(n12419) );
  NOR2_X1 U14893 ( .A1(n15298), .A2(n15151), .ZN(n12422) );
  NAND2_X1 U14894 ( .A1(n15298), .A2(n15151), .ZN(n12421) );
  AND2_X1 U14895 ( .A1(n15294), .A2(n14777), .ZN(n12423) );
  NAND2_X1 U14896 ( .A1(n15099), .A2(n15100), .ZN(n12425) );
  OR2_X1 U14897 ( .A1(n15287), .A2(n14776), .ZN(n12424) );
  NAND2_X1 U14898 ( .A1(n12425), .A2(n12424), .ZN(n15060) );
  NAND2_X1 U14899 ( .A1(n15278), .A2(n15050), .ZN(n15061) );
  OAI21_X1 U14900 ( .B1(n15059), .B2(n15071), .A(n15061), .ZN(n12426) );
  INV_X1 U14901 ( .A(n12426), .ZN(n12427) );
  NAND2_X1 U14902 ( .A1(n15060), .A2(n12427), .ZN(n12431) );
  OAI21_X1 U14903 ( .B1(n15278), .B2(n15050), .A(n14775), .ZN(n12429) );
  INV_X1 U14904 ( .A(n15278), .ZN(n12782) );
  AND2_X1 U14905 ( .A1(n15071), .A2(n15090), .ZN(n12428) );
  AOI22_X1 U14906 ( .A1(n15059), .A2(n12429), .B1(n12782), .B2(n12428), .ZN(
        n12430) );
  OR2_X1 U14907 ( .A1(n15267), .A2(n15051), .ZN(n12432) );
  OR2_X1 U14908 ( .A1(n14619), .A2(n14729), .ZN(n12433) );
  INV_X1 U14909 ( .A(n14969), .ZN(n14972) );
  INV_X1 U14910 ( .A(n12895), .ZN(n12441) );
  INV_X1 U14911 ( .A(n12440), .ZN(n12436) );
  NAND2_X1 U14912 ( .A1(n12441), .A2(n12436), .ZN(n12437) );
  AND2_X1 U14913 ( .A1(n14962), .A2(n14939), .ZN(n14931) );
  NOR2_X1 U14914 ( .A1(n12438), .A2(n14931), .ZN(n12444) );
  OAI21_X1 U14915 ( .B1(n12440), .B2(n12444), .A(n12441), .ZN(n12439) );
  OAI21_X1 U14916 ( .B1(n12441), .B2(n12440), .A(n12439), .ZN(n12442) );
  NAND3_X1 U14917 ( .A1(n14954), .A2(n12444), .A3(n12895), .ZN(n12445) );
  INV_X1 U14918 ( .A(n15302), .ZN(n15148) );
  AND2_X2 U14919 ( .A1(n15169), .A2(n15148), .ZN(n15142) );
  INV_X1 U14920 ( .A(n15298), .ZN(n15137) );
  NOR2_X1 U14921 ( .A1(n15207), .A2(n15056), .ZN(n12459) );
  INV_X1 U14922 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n12453) );
  INV_X1 U14923 ( .A(P1_B_REG_SCAN_IN), .ZN(n12446) );
  NOR2_X1 U14924 ( .A1(n6762), .A2(n12446), .ZN(n12447) );
  NOR2_X1 U14925 ( .A1(n15130), .A2(n12447), .ZN(n14919) );
  INV_X1 U14926 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n12451) );
  NAND2_X1 U14927 ( .A1(n12448), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n12450) );
  NAND2_X1 U14928 ( .A1(n11451), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n12449) );
  OAI211_X1 U14929 ( .C1(n10700), .C2(n12451), .A(n12450), .B(n12449), .ZN(
        n14767) );
  NAND2_X1 U14930 ( .A1(n14919), .A2(n14767), .ZN(n15208) );
  OAI22_X1 U14931 ( .A1(n15097), .A2(n12453), .B1(n15208), .B2(n12452), .ZN(
        n12455) );
  NAND2_X1 U14932 ( .A1(n14769), .A2(n15180), .ZN(n15209) );
  NOR2_X1 U14933 ( .A1(n15209), .A2(n15512), .ZN(n12454) );
  AOI211_X1 U14934 ( .C1(n15513), .C2(n12456), .A(n12455), .B(n12454), .ZN(
        n12457) );
  OAI21_X1 U14935 ( .B1(n15210), .B2(n15147), .A(n12457), .ZN(n12458) );
  AOI211_X1 U14936 ( .C1(n15214), .C2(n15101), .A(n12459), .B(n12458), .ZN(
        n12460) );
  OAI21_X1 U14937 ( .B1(n15215), .B2(n15104), .A(n12460), .ZN(P1_U3356) );
  INV_X1 U14938 ( .A(n12461), .ZN(n14595) );
  OAI222_X1 U14939 ( .A1(n15370), .A2(n12462), .B1(n15379), .B2(n14595), .C1(
        P1_U3086), .C2(n10463), .ZN(P1_U3327) );
  OAI22_X1 U14940 ( .A1(n14962), .A2(n14638), .B1(n14939), .B2(n12463), .ZN(
        n12464) );
  XNOR2_X1 U14941 ( .A(n12464), .B(n11860), .ZN(n12468) );
  OR2_X1 U14942 ( .A1(n14962), .A2(n10379), .ZN(n12466) );
  OR2_X1 U14943 ( .A1(n14939), .A2(n14636), .ZN(n12465) );
  NAND2_X1 U14944 ( .A1(n12466), .A2(n12465), .ZN(n12467) );
  NOR2_X1 U14945 ( .A1(n12468), .A2(n12467), .ZN(n14649) );
  AOI21_X1 U14946 ( .B1(n12468), .B2(n12467), .A(n14649), .ZN(n12579) );
  INV_X1 U14947 ( .A(n12469), .ZN(n12472) );
  INV_X1 U14948 ( .A(n12470), .ZN(n12471) );
  NAND2_X1 U14949 ( .A1(n12472), .A2(n12471), .ZN(n12473) );
  OAI22_X1 U14950 ( .A1(n14723), .A2(n14638), .B1(n12754), .B2(n10699), .ZN(
        n12475) );
  XNOR2_X1 U14951 ( .A(n12475), .B(n11860), .ZN(n12477) );
  NOR2_X1 U14952 ( .A1(n14636), .A2(n12754), .ZN(n12476) );
  AOI21_X1 U14953 ( .B1(n15319), .B2(n12552), .A(n12476), .ZN(n12478) );
  XNOR2_X1 U14954 ( .A(n12477), .B(n12478), .ZN(n14713) );
  INV_X1 U14955 ( .A(n12477), .ZN(n12479) );
  OR2_X1 U14956 ( .A1(n12479), .A2(n12478), .ZN(n12480) );
  NAND2_X1 U14957 ( .A1(n14712), .A2(n12480), .ZN(n14600) );
  INV_X1 U14958 ( .A(n14600), .ZN(n12484) );
  INV_X1 U14959 ( .A(n15314), .ZN(n12482) );
  OAI22_X1 U14960 ( .A1(n12482), .A2(n14638), .B1(n14758), .B2(n10699), .ZN(
        n12481) );
  XNOR2_X1 U14961 ( .A(n12481), .B(n11860), .ZN(n12485) );
  OAI22_X1 U14962 ( .A1(n12482), .A2(n12463), .B1(n14758), .B2(n14636), .ZN(
        n12486) );
  XNOR2_X1 U14963 ( .A(n12485), .B(n12486), .ZN(n14601) );
  INV_X1 U14964 ( .A(n14601), .ZN(n12483) );
  NAND2_X2 U14965 ( .A1(n12484), .A2(n12483), .ZN(n14598) );
  INV_X1 U14966 ( .A(n12485), .ZN(n12488) );
  INV_X1 U14967 ( .A(n12486), .ZN(n12487) );
  NAND2_X1 U14968 ( .A1(n12488), .A2(n12487), .ZN(n12489) );
  NAND2_X1 U14969 ( .A1(n15308), .A2(n6553), .ZN(n12491) );
  NAND2_X1 U14970 ( .A1(n15179), .A2(n6554), .ZN(n12490) );
  NAND2_X1 U14971 ( .A1(n12491), .A2(n12490), .ZN(n12492) );
  XNOR2_X1 U14972 ( .A(n12492), .B(n11860), .ZN(n14674) );
  NAND2_X1 U14973 ( .A1(n15308), .A2(n12552), .ZN(n12494) );
  NAND2_X1 U14974 ( .A1(n12572), .A2(n15179), .ZN(n12493) );
  NAND2_X1 U14975 ( .A1(n12494), .A2(n12493), .ZN(n14755) );
  NAND2_X1 U14976 ( .A1(n15302), .A2(n6553), .ZN(n12496) );
  NAND2_X1 U14977 ( .A1(n14778), .A2(n12552), .ZN(n12495) );
  NAND2_X1 U14978 ( .A1(n12496), .A2(n12495), .ZN(n12497) );
  XNOR2_X1 U14979 ( .A(n12497), .B(n11860), .ZN(n14676) );
  NAND2_X1 U14980 ( .A1(n15302), .A2(n12552), .ZN(n12499) );
  NAND2_X1 U14981 ( .A1(n12572), .A2(n14778), .ZN(n12498) );
  NAND2_X1 U14982 ( .A1(n12499), .A2(n12498), .ZN(n14677) );
  AND2_X1 U14983 ( .A1(n14676), .A2(n14677), .ZN(n12500) );
  AOI21_X1 U14984 ( .B1(n14674), .B2(n14755), .A(n12500), .ZN(n12505) );
  INV_X1 U14985 ( .A(n12500), .ZN(n12502) );
  INV_X1 U14986 ( .A(n14755), .ZN(n12501) );
  NAND2_X1 U14987 ( .A1(n12502), .A2(n12501), .ZN(n12503) );
  OAI22_X1 U14988 ( .A1(n14674), .A2(n12503), .B1(n14677), .B2(n14676), .ZN(
        n12504) );
  AOI22_X1 U14989 ( .A1(n15298), .A2(n6553), .B1(n6554), .B2(n15151), .ZN(
        n12506) );
  XNOR2_X1 U14990 ( .A(n12506), .B(n11860), .ZN(n14687) );
  NOR2_X1 U14991 ( .A1(n14680), .A2(n14636), .ZN(n12507) );
  AOI21_X1 U14992 ( .B1(n15298), .B2(n6554), .A(n12507), .ZN(n14688) );
  NAND2_X1 U14993 ( .A1(n14687), .A2(n14688), .ZN(n12508) );
  INV_X1 U14994 ( .A(n15294), .ZN(n12510) );
  OAI22_X1 U14995 ( .A1(n12510), .A2(n14638), .B1(n15131), .B2(n12463), .ZN(
        n12509) );
  XNOR2_X1 U14996 ( .A(n12509), .B(n11860), .ZN(n12512) );
  OAI22_X1 U14997 ( .A1(n12510), .A2(n10699), .B1(n15131), .B2(n14636), .ZN(
        n12513) );
  XNOR2_X1 U14998 ( .A(n12512), .B(n12513), .ZN(n14736) );
  INV_X1 U14999 ( .A(n12512), .ZN(n12515) );
  INV_X1 U15000 ( .A(n12513), .ZN(n12514) );
  NAND2_X1 U15001 ( .A1(n12515), .A2(n12514), .ZN(n12516) );
  OAI22_X1 U15002 ( .A1(n15095), .A2(n14638), .B1(n15070), .B2(n10699), .ZN(
        n12517) );
  XNOR2_X1 U15003 ( .A(n12517), .B(n11860), .ZN(n12520) );
  OAI22_X1 U15004 ( .A1(n15095), .A2(n10379), .B1(n15070), .B2(n14636), .ZN(
        n12519) );
  XNOR2_X1 U15005 ( .A(n12520), .B(n12519), .ZN(n14632) );
  NAND2_X1 U15006 ( .A1(n12520), .A2(n12519), .ZN(n12521) );
  NAND2_X1 U15007 ( .A1(n15278), .A2(n6553), .ZN(n12523) );
  NAND2_X1 U15008 ( .A1(n15050), .A2(n12552), .ZN(n12522) );
  NAND2_X1 U15009 ( .A1(n12523), .A2(n12522), .ZN(n12524) );
  XNOR2_X1 U15010 ( .A(n12524), .B(n11860), .ZN(n12528) );
  NOR2_X1 U15011 ( .A1(n15090), .A2(n14636), .ZN(n12525) );
  AOI21_X1 U15012 ( .B1(n15278), .B2(n12552), .A(n12525), .ZN(n12526) );
  XNOR2_X1 U15013 ( .A(n12528), .B(n12526), .ZN(n14703) );
  INV_X1 U15014 ( .A(n12526), .ZN(n12527) );
  OAI22_X1 U15015 ( .A1(n15059), .A2(n14638), .B1(n15071), .B2(n10699), .ZN(
        n12529) );
  XNOR2_X1 U15016 ( .A(n12529), .B(n11860), .ZN(n12531) );
  OAI22_X1 U15017 ( .A1(n15059), .A2(n12463), .B1(n15071), .B2(n14636), .ZN(
        n12530) );
  NOR2_X1 U15018 ( .A1(n12531), .A2(n12530), .ZN(n14725) );
  AOI21_X1 U15019 ( .B1(n12531), .B2(n12530), .A(n14725), .ZN(n14656) );
  NAND2_X1 U15020 ( .A1(n15267), .A2(n6553), .ZN(n12533) );
  NAND2_X1 U15021 ( .A1(n15051), .A2(n12552), .ZN(n12532) );
  NAND2_X1 U15022 ( .A1(n12533), .A2(n12532), .ZN(n12535) );
  XNOR2_X1 U15023 ( .A(n12535), .B(n12534), .ZN(n12537) );
  AND2_X1 U15024 ( .A1(n15051), .A2(n12572), .ZN(n12536) );
  AOI21_X1 U15025 ( .B1(n15267), .B2(n6554), .A(n12536), .ZN(n12538) );
  NAND2_X1 U15026 ( .A1(n12537), .A2(n12538), .ZN(n14607) );
  INV_X1 U15027 ( .A(n12537), .ZN(n12540) );
  INV_X1 U15028 ( .A(n12538), .ZN(n12539) );
  NAND2_X1 U15029 ( .A1(n12540), .A2(n12539), .ZN(n12541) );
  NAND2_X1 U15030 ( .A1(n14606), .A2(n14607), .ZN(n12550) );
  OAI22_X1 U15031 ( .A1(n14619), .A2(n14638), .B1(n14729), .B2(n12463), .ZN(
        n12542) );
  XNOR2_X1 U15032 ( .A(n12542), .B(n12534), .ZN(n12545) );
  OR2_X1 U15033 ( .A1(n14619), .A2(n10699), .ZN(n12544) );
  NAND2_X1 U15034 ( .A1(n14774), .A2(n12572), .ZN(n12543) );
  NAND2_X1 U15035 ( .A1(n12545), .A2(n12546), .ZN(n14695) );
  INV_X1 U15036 ( .A(n12545), .ZN(n12548) );
  INV_X1 U15037 ( .A(n12546), .ZN(n12547) );
  NAND2_X1 U15038 ( .A1(n12548), .A2(n12547), .ZN(n12549) );
  NAND2_X1 U15039 ( .A1(n15253), .A2(n6553), .ZN(n12554) );
  NAND2_X1 U15040 ( .A1(n14773), .A2(n12552), .ZN(n12553) );
  NAND2_X1 U15041 ( .A1(n12554), .A2(n12553), .ZN(n12555) );
  XNOR2_X1 U15042 ( .A(n12555), .B(n12534), .ZN(n12557) );
  AND2_X1 U15043 ( .A1(n14773), .A2(n12572), .ZN(n12556) );
  AOI21_X1 U15044 ( .B1(n15253), .B2(n12552), .A(n12556), .ZN(n12558) );
  NAND2_X1 U15045 ( .A1(n12557), .A2(n12558), .ZN(n14664) );
  INV_X1 U15046 ( .A(n12557), .ZN(n12560) );
  INV_X1 U15047 ( .A(n12558), .ZN(n12559) );
  NAND2_X1 U15048 ( .A1(n12560), .A2(n12559), .ZN(n12561) );
  OAI22_X1 U15049 ( .A1(n15245), .A2(n14638), .B1(n14748), .B2(n10379), .ZN(
        n12562) );
  XNOR2_X1 U15050 ( .A(n12562), .B(n12534), .ZN(n12565) );
  OR2_X1 U15051 ( .A1(n15245), .A2(n10379), .ZN(n12564) );
  NAND2_X1 U15052 ( .A1(n14772), .A2(n12572), .ZN(n12563) );
  NAND2_X1 U15053 ( .A1(n12565), .A2(n12566), .ZN(n12570) );
  INV_X1 U15054 ( .A(n12565), .ZN(n12568) );
  INV_X1 U15055 ( .A(n12566), .ZN(n12567) );
  NAND2_X1 U15056 ( .A1(n12568), .A2(n12567), .ZN(n12569) );
  OAI22_X1 U15057 ( .A1(n14980), .A2(n14638), .B1(n14990), .B2(n10379), .ZN(
        n12571) );
  XNOR2_X1 U15058 ( .A(n12571), .B(n11860), .ZN(n12576) );
  OR2_X1 U15059 ( .A1(n14980), .A2(n10379), .ZN(n12574) );
  NAND2_X1 U15060 ( .A1(n14771), .A2(n12572), .ZN(n12573) );
  NAND2_X1 U15061 ( .A1(n12574), .A2(n12573), .ZN(n12575) );
  NOR2_X1 U15062 ( .A1(n12576), .A2(n12575), .ZN(n12577) );
  AOI21_X1 U15063 ( .B1(n12576), .B2(n12575), .A(n12577), .ZN(n14746) );
  NAND2_X1 U15064 ( .A1(n14745), .A2(n14746), .ZN(n14744) );
  INV_X1 U15065 ( .A(n12577), .ZN(n12578) );
  OAI22_X1 U15066 ( .A1(n14990), .A2(n14715), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12580), .ZN(n12581) );
  AOI21_X1 U15067 ( .B1(n14958), .B2(n14690), .A(n12581), .ZN(n12582) );
  OAI21_X1 U15068 ( .B1(n14959), .B2(n14706), .A(n12582), .ZN(n12583) );
  AOI21_X1 U15069 ( .B1(n15230), .B2(n14740), .A(n12583), .ZN(n12584) );
  NAND2_X1 U15070 ( .A1(n12585), .A2(n12584), .ZN(P1_U3214) );
  OAI222_X1 U15071 ( .A1(P1_U3086), .A2(n12588), .B1(n15379), .B2(n12587), 
        .C1(n12586), .C2(n15370), .ZN(P1_U3329) );
  NAND2_X1 U15072 ( .A1(n12589), .A2(n15750), .ZN(n12593) );
  OAI21_X1 U15073 ( .B1(n14111), .B2(n14514), .A(n12594), .ZN(P2_U3527) );
  INV_X1 U15074 ( .A(n12811), .ZN(n15373) );
  INV_X1 U15075 ( .A(n12596), .ZN(n12599) );
  INV_X1 U15076 ( .A(n12597), .ZN(n12598) );
  XNOR2_X1 U15077 ( .A(n14570), .B(n13789), .ZN(n12602) );
  NOR2_X1 U15078 ( .A1(n13812), .A2(n14293), .ZN(n12603) );
  XNOR2_X1 U15079 ( .A(n12602), .B(n12603), .ZN(n13881) );
  INV_X1 U15080 ( .A(n12602), .ZN(n12604) );
  NAND2_X1 U15081 ( .A1(n12604), .A2(n12603), .ZN(n12605) );
  NAND2_X1 U15082 ( .A1(n12606), .A2(n12605), .ZN(n13810) );
  XNOR2_X1 U15083 ( .A(n14357), .B(n12649), .ZN(n12607) );
  NAND2_X1 U15084 ( .A1(n13946), .A2(n6556), .ZN(n12608) );
  NAND2_X1 U15085 ( .A1(n12607), .A2(n12608), .ZN(n13809) );
  NAND2_X1 U15086 ( .A1(n13810), .A2(n13809), .ZN(n12611) );
  INV_X1 U15087 ( .A(n12607), .ZN(n12610) );
  INV_X1 U15088 ( .A(n12608), .ZN(n12609) );
  NAND2_X1 U15089 ( .A1(n12610), .A2(n12609), .ZN(n13808) );
  NAND2_X1 U15090 ( .A1(n12611), .A2(n13808), .ZN(n13863) );
  XNOR2_X1 U15091 ( .A(n14339), .B(n13789), .ZN(n12615) );
  NAND2_X1 U15092 ( .A1(n13945), .A2(n12612), .ZN(n12613) );
  XNOR2_X1 U15093 ( .A(n12615), .B(n12613), .ZN(n13862) );
  NAND2_X1 U15094 ( .A1(n13863), .A2(n13862), .ZN(n12617) );
  INV_X1 U15095 ( .A(n12613), .ZN(n12614) );
  NAND2_X1 U15096 ( .A1(n12615), .A2(n12614), .ZN(n12616) );
  XNOR2_X1 U15097 ( .A(n14481), .B(n12649), .ZN(n12618) );
  NAND2_X1 U15098 ( .A1(n13944), .A2(n12612), .ZN(n12619) );
  NAND2_X1 U15099 ( .A1(n12618), .A2(n12619), .ZN(n12624) );
  INV_X1 U15100 ( .A(n12618), .ZN(n12621) );
  INV_X1 U15101 ( .A(n12619), .ZN(n12620) );
  NAND2_X1 U15102 ( .A1(n12621), .A2(n12620), .ZN(n12622) );
  NAND2_X1 U15103 ( .A1(n12624), .A2(n12622), .ZN(n13758) );
  INV_X1 U15104 ( .A(n13758), .ZN(n12623) );
  XNOR2_X1 U15105 ( .A(n14306), .B(n12649), .ZN(n13821) );
  XNOR2_X1 U15106 ( .A(n14469), .B(n12649), .ZN(n12626) );
  NAND2_X1 U15107 ( .A1(n13942), .A2(n6556), .ZN(n12627) );
  NAND2_X1 U15108 ( .A1(n12626), .A2(n12627), .ZN(n13825) );
  INV_X1 U15109 ( .A(n13825), .ZN(n12625) );
  AND2_X1 U15110 ( .A1(n13943), .A2(n12612), .ZN(n13913) );
  NAND2_X1 U15111 ( .A1(n13825), .A2(n13913), .ZN(n12630) );
  OAI21_X1 U15112 ( .B1(n13821), .B2(n12625), .A(n12630), .ZN(n12632) );
  INV_X1 U15113 ( .A(n12626), .ZN(n12629) );
  INV_X1 U15114 ( .A(n12627), .ZN(n12628) );
  NAND2_X1 U15115 ( .A1(n12629), .A2(n12628), .ZN(n13824) );
  OAI21_X1 U15116 ( .B1(n13821), .B2(n12630), .A(n13824), .ZN(n12631) );
  XNOR2_X1 U15117 ( .A(n14274), .B(n12649), .ZN(n12633) );
  NAND2_X1 U15118 ( .A1(n13941), .A2(n12612), .ZN(n12634) );
  NAND2_X1 U15119 ( .A1(n12633), .A2(n12634), .ZN(n12638) );
  INV_X1 U15120 ( .A(n12633), .ZN(n12636) );
  INV_X1 U15121 ( .A(n12634), .ZN(n12635) );
  NAND2_X1 U15122 ( .A1(n12636), .A2(n12635), .ZN(n12637) );
  XNOR2_X1 U15123 ( .A(n14260), .B(n12649), .ZN(n12641) );
  NOR2_X1 U15124 ( .A1(n12639), .A2(n14293), .ZN(n12640) );
  XNOR2_X1 U15125 ( .A(n12641), .B(n12640), .ZN(n13890) );
  XNOR2_X1 U15126 ( .A(n14251), .B(n13789), .ZN(n12642) );
  NAND2_X1 U15127 ( .A1(n13939), .A2(n6556), .ZN(n12643) );
  NAND2_X1 U15128 ( .A1(n12642), .A2(n12643), .ZN(n12648) );
  INV_X1 U15129 ( .A(n12642), .ZN(n12645) );
  INV_X1 U15130 ( .A(n12643), .ZN(n12644) );
  NAND2_X1 U15131 ( .A1(n12645), .A2(n12644), .ZN(n12646) );
  NAND2_X1 U15132 ( .A1(n12648), .A2(n12646), .ZN(n13777) );
  INV_X1 U15133 ( .A(n13777), .ZN(n12647) );
  XNOR2_X1 U15134 ( .A(n14451), .B(n12649), .ZN(n12650) );
  NAND2_X1 U15135 ( .A1(n13938), .A2(n6556), .ZN(n12651) );
  NAND2_X1 U15136 ( .A1(n12650), .A2(n12651), .ZN(n13851) );
  INV_X1 U15137 ( .A(n12650), .ZN(n12653) );
  INV_X1 U15138 ( .A(n12651), .ZN(n12652) );
  NAND2_X1 U15139 ( .A1(n12653), .A2(n12652), .ZN(n13850) );
  XNOR2_X1 U15140 ( .A(n14548), .B(n13789), .ZN(n12657) );
  NOR2_X1 U15141 ( .A1(n12655), .A2(n14293), .ZN(n12660) );
  XNOR2_X1 U15142 ( .A(n12657), .B(n12660), .ZN(n13871) );
  XNOR2_X1 U15143 ( .A(n14545), .B(n13789), .ZN(n13873) );
  OR2_X1 U15144 ( .A1(n13801), .A2(n14293), .ZN(n13872) );
  NAND2_X1 U15145 ( .A1(n13873), .A2(n13872), .ZN(n12656) );
  INV_X1 U15146 ( .A(n12657), .ZN(n12661) );
  NAND2_X1 U15147 ( .A1(n12661), .A2(n12660), .ZN(n13869) );
  NAND2_X1 U15148 ( .A1(n13869), .A2(n13872), .ZN(n12659) );
  INV_X1 U15149 ( .A(n13873), .ZN(n12658) );
  NAND2_X1 U15150 ( .A1(n12659), .A2(n12658), .ZN(n12663) );
  INV_X1 U15151 ( .A(n13801), .ZN(n13936) );
  NAND3_X1 U15152 ( .A1(n12661), .A2(n12660), .A3(n13936), .ZN(n12662) );
  XNOR2_X1 U15153 ( .A(n14541), .B(n13789), .ZN(n13733) );
  AND2_X1 U15154 ( .A1(n13729), .A2(n13733), .ZN(n12664) );
  XNOR2_X1 U15155 ( .A(n14167), .B(n13789), .ZN(n12665) );
  INV_X1 U15156 ( .A(n12665), .ZN(n13732) );
  NOR2_X1 U15157 ( .A1(n13768), .A2(n14293), .ZN(n13735) );
  XNOR2_X1 U15158 ( .A(n13732), .B(n13735), .ZN(n13843) );
  NAND2_X1 U15159 ( .A1(n13844), .A2(n13843), .ZN(n13842) );
  NAND2_X1 U15160 ( .A1(n12665), .A2(n13735), .ZN(n13728) );
  NAND2_X1 U15161 ( .A1(n13842), .A2(n13728), .ZN(n12667) );
  XNOR2_X1 U15162 ( .A(n14534), .B(n13789), .ZN(n13738) );
  NAND2_X1 U15163 ( .A1(n13933), .A2(n6556), .ZN(n13739) );
  XNOR2_X1 U15164 ( .A(n13738), .B(n13739), .ZN(n13737) );
  INV_X1 U15165 ( .A(n13737), .ZN(n12666) );
  XNOR2_X1 U15166 ( .A(n12667), .B(n12666), .ZN(n12671) );
  AOI22_X1 U15167 ( .A1(n13932), .A2(n13907), .B1(n13934), .B2(n13905), .ZN(
        n14144) );
  AOI22_X1 U15168 ( .A1(n14150), .A2(n13859), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12668) );
  OAI21_X1 U15169 ( .B1(n14144), .B2(n13855), .A(n12668), .ZN(n12669) );
  AOI21_X1 U15170 ( .B1(n14146), .B2(n13923), .A(n12669), .ZN(n12670) );
  OAI21_X1 U15171 ( .B1(n12671), .B2(n13925), .A(n12670), .ZN(P2_U3197) );
  XNOR2_X1 U15172 ( .A(n12673), .B(n12672), .ZN(n12676) );
  NAND2_X1 U15173 ( .A1(n12676), .A2(n12917), .ZN(n12816) );
  NAND2_X1 U15174 ( .A1(n12676), .A2(n12675), .ZN(n12677) );
  MUX2_X1 U15175 ( .A(n15245), .B(n14748), .S(n12799), .Z(n12824) );
  CLKBUF_X3 U15176 ( .A(n12681), .Z(n12821) );
  MUX2_X1 U15177 ( .A(n14772), .B(n12678), .S(n12681), .Z(n12823) );
  MUX2_X1 U15178 ( .A(n14619), .B(n14729), .S(n12821), .Z(n12801) );
  MUX2_X1 U15179 ( .A(n15071), .B(n15059), .S(n12862), .Z(n12792) );
  MUX2_X1 U15180 ( .A(n12681), .B(n12680), .S(n12679), .Z(n12686) );
  INV_X1 U15181 ( .A(n12688), .ZN(n12682) );
  NAND2_X1 U15182 ( .A1(n12686), .A2(n12685), .ZN(n12690) );
  MUX2_X1 U15183 ( .A(n12688), .B(n12687), .S(n12821), .Z(n12689) );
  MUX2_X1 U15184 ( .A(n14790), .B(n12691), .S(n12821), .Z(n12694) );
  INV_X1 U15185 ( .A(n12694), .ZN(n12693) );
  MUX2_X1 U15186 ( .A(n12691), .B(n14790), .S(n12821), .Z(n12692) );
  MUX2_X1 U15187 ( .A(n12697), .B(n12696), .S(n12821), .Z(n12698) );
  MUX2_X1 U15188 ( .A(n14788), .B(n12699), .S(n12821), .Z(n12703) );
  NAND2_X1 U15189 ( .A1(n12702), .A2(n12703), .ZN(n12701) );
  MUX2_X1 U15190 ( .A(n14788), .B(n12699), .S(n12862), .Z(n12700) );
  NAND2_X1 U15191 ( .A1(n12701), .A2(n12700), .ZN(n12707) );
  INV_X1 U15192 ( .A(n12702), .ZN(n12705) );
  INV_X1 U15193 ( .A(n12703), .ZN(n12704) );
  NAND2_X1 U15194 ( .A1(n12705), .A2(n12704), .ZN(n12706) );
  MUX2_X1 U15195 ( .A(n12708), .B(n14787), .S(n12821), .Z(n12710) );
  MUX2_X1 U15196 ( .A(n14787), .B(n12708), .S(n12821), .Z(n12709) );
  INV_X1 U15197 ( .A(n12710), .ZN(n12711) );
  MUX2_X1 U15198 ( .A(n14786), .B(n12712), .S(n12799), .Z(n12716) );
  NAND2_X1 U15199 ( .A1(n12715), .A2(n12716), .ZN(n12714) );
  MUX2_X1 U15200 ( .A(n14786), .B(n12712), .S(n12862), .Z(n12713) );
  NAND2_X1 U15201 ( .A1(n12714), .A2(n12713), .ZN(n12720) );
  INV_X1 U15202 ( .A(n12715), .ZN(n12718) );
  INV_X1 U15203 ( .A(n12716), .ZN(n12717) );
  NAND2_X1 U15204 ( .A1(n12718), .A2(n12717), .ZN(n12719) );
  MUX2_X1 U15205 ( .A(n14785), .B(n15516), .S(n12862), .Z(n12722) );
  MUX2_X1 U15206 ( .A(n14785), .B(n15516), .S(n12799), .Z(n12721) );
  INV_X1 U15207 ( .A(n12722), .ZN(n12723) );
  MUX2_X1 U15208 ( .A(n14784), .B(n12724), .S(n12799), .Z(n12728) );
  NAND2_X1 U15209 ( .A1(n12727), .A2(n12728), .ZN(n12726) );
  MUX2_X1 U15210 ( .A(n14784), .B(n12724), .S(n12862), .Z(n12725) );
  NAND2_X1 U15211 ( .A1(n12726), .A2(n12725), .ZN(n12732) );
  INV_X1 U15212 ( .A(n12727), .ZN(n12730) );
  INV_X1 U15213 ( .A(n12728), .ZN(n12729) );
  NAND2_X1 U15214 ( .A1(n12730), .A2(n12729), .ZN(n12731) );
  MUX2_X1 U15215 ( .A(n14783), .B(n15499), .S(n12862), .Z(n12734) );
  MUX2_X1 U15216 ( .A(n14783), .B(n15499), .S(n12799), .Z(n12733) );
  INV_X1 U15217 ( .A(n12734), .ZN(n12735) );
  MUX2_X1 U15218 ( .A(n14782), .B(n15336), .S(n12799), .Z(n12739) );
  MUX2_X1 U15219 ( .A(n14782), .B(n15336), .S(n12862), .Z(n12736) );
  AOI21_X1 U15220 ( .B1(n12740), .B2(n12739), .A(n12737), .ZN(n12738) );
  INV_X1 U15221 ( .A(n12738), .ZN(n12741) );
  MUX2_X1 U15222 ( .A(n14781), .B(n15331), .S(n12862), .Z(n12743) );
  MUX2_X1 U15223 ( .A(n14781), .B(n15331), .S(n12799), .Z(n12742) );
  INV_X1 U15224 ( .A(n12743), .ZN(n12744) );
  MUX2_X1 U15225 ( .A(n14780), .B(n12745), .S(n12799), .Z(n12749) );
  NAND2_X1 U15226 ( .A1(n12748), .A2(n12749), .ZN(n12747) );
  MUX2_X1 U15227 ( .A(n14780), .B(n12745), .S(n12862), .Z(n12746) );
  NAND2_X1 U15228 ( .A1(n12747), .A2(n12746), .ZN(n12753) );
  INV_X1 U15229 ( .A(n12748), .ZN(n12751) );
  INV_X1 U15230 ( .A(n12749), .ZN(n12750) );
  NAND2_X1 U15231 ( .A1(n12751), .A2(n12750), .ZN(n12752) );
  MUX2_X1 U15232 ( .A(n15181), .B(n15319), .S(n12862), .Z(n12756) );
  MUX2_X1 U15233 ( .A(n12754), .B(n14723), .S(n12799), .Z(n12755) );
  NAND2_X1 U15234 ( .A1(n12761), .A2(n12757), .ZN(n12759) );
  NAND2_X1 U15235 ( .A1(n12760), .A2(n15163), .ZN(n12758) );
  MUX2_X1 U15236 ( .A(n12759), .B(n12758), .S(n12799), .Z(n12763) );
  MUX2_X1 U15237 ( .A(n12761), .B(n12760), .S(n12862), .Z(n12762) );
  MUX2_X1 U15238 ( .A(n15129), .B(n15148), .S(n12799), .Z(n12773) );
  AND2_X1 U15239 ( .A1(n14778), .A2(n12821), .ZN(n12764) );
  AOI21_X1 U15240 ( .B1(n15302), .B2(n12862), .A(n12764), .ZN(n12766) );
  NAND2_X1 U15241 ( .A1(n15298), .A2(n14680), .ZN(n12765) );
  NAND3_X1 U15242 ( .A1(n12767), .A2(n12766), .A3(n12765), .ZN(n12774) );
  OAI21_X1 U15243 ( .B1(n15126), .B2(n12773), .A(n12774), .ZN(n12768) );
  NAND2_X1 U15244 ( .A1(n12769), .A2(n12768), .ZN(n12777) );
  AND2_X1 U15245 ( .A1(n15151), .A2(n12862), .ZN(n12771) );
  OAI21_X1 U15246 ( .B1(n12862), .B2(n15151), .A(n15298), .ZN(n12770) );
  OAI21_X1 U15247 ( .B1(n12771), .B2(n15298), .A(n12770), .ZN(n12772) );
  OAI21_X1 U15248 ( .B1(n12774), .B2(n12773), .A(n12772), .ZN(n12775) );
  NAND2_X1 U15249 ( .A1(n12777), .A2(n12776), .ZN(n12778) );
  NAND2_X1 U15250 ( .A1(n6576), .A2(n15090), .ZN(n12783) );
  NAND3_X1 U15251 ( .A1(n12783), .A2(n12782), .A3(n12821), .ZN(n12789) );
  NAND2_X1 U15252 ( .A1(n12785), .A2(n15050), .ZN(n12784) );
  NAND3_X1 U15253 ( .A1(n12784), .A2(n12862), .A3(n15278), .ZN(n12788) );
  OR3_X1 U15254 ( .A1(n6576), .A2(n15090), .A3(n12862), .ZN(n12787) );
  OR3_X1 U15255 ( .A1(n12785), .A2(n15050), .A3(n12821), .ZN(n12786) );
  NAND4_X1 U15256 ( .A1(n12789), .A2(n12788), .A3(n12787), .A4(n12786), .ZN(
        n12790) );
  MUX2_X1 U15257 ( .A(n14775), .B(n15271), .S(n12799), .Z(n12791) );
  INV_X1 U15258 ( .A(n12793), .ZN(n12798) );
  MUX2_X1 U15259 ( .A(n15051), .B(n15267), .S(n12799), .Z(n12795) );
  INV_X1 U15260 ( .A(n12795), .ZN(n12797) );
  INV_X1 U15261 ( .A(n15051), .ZN(n14659) );
  MUX2_X1 U15262 ( .A(n15044), .B(n14659), .S(n12821), .Z(n12794) );
  AOI21_X1 U15263 ( .B1(n12793), .B2(n12795), .A(n12794), .ZN(n12796) );
  MUX2_X1 U15264 ( .A(n14774), .B(n15259), .S(n12799), .Z(n12800) );
  MUX2_X1 U15265 ( .A(n14773), .B(n15253), .S(n12821), .Z(n12802) );
  MUX2_X1 U15266 ( .A(n15253), .B(n14773), .S(n12821), .Z(n12803) );
  AOI21_X1 U15267 ( .B1(n12824), .B2(n12823), .A(n12804), .ZN(n12854) );
  MUX2_X1 U15268 ( .A(n14939), .B(n14962), .S(n12862), .Z(n12833) );
  MUX2_X1 U15269 ( .A(n14770), .B(n15230), .S(n12821), .Z(n12832) );
  INV_X1 U15270 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n12807) );
  NAND2_X1 U15271 ( .A1(n12448), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n12806) );
  NAND2_X1 U15272 ( .A1(n11031), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n12805) );
  OAI211_X1 U15273 ( .C1(n10700), .C2(n12807), .A(n12806), .B(n12805), .ZN(
        n14918) );
  INV_X1 U15274 ( .A(n12808), .ZN(n12809) );
  OAI21_X1 U15275 ( .B1(n14918), .B2(n12809), .A(n14767), .ZN(n12810) );
  INV_X1 U15276 ( .A(n12810), .ZN(n12814) );
  NAND2_X1 U15277 ( .A1(n12811), .A2(n12393), .ZN(n12813) );
  NAND2_X1 U15278 ( .A1(n12855), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12812) );
  NAND2_X1 U15279 ( .A1(n12862), .A2(n14918), .ZN(n12817) );
  INV_X1 U15280 ( .A(n14767), .ZN(n12815) );
  AOI21_X1 U15281 ( .B1(n12817), .B2(n12816), .A(n12815), .ZN(n12818) );
  AOI21_X1 U15282 ( .B1(n14923), .B2(n12821), .A(n12818), .ZN(n12840) );
  MUX2_X1 U15283 ( .A(n14940), .B(n15210), .S(n12821), .Z(n12835) );
  MUX2_X1 U15284 ( .A(n14768), .B(n12819), .S(n12862), .Z(n12834) );
  NAND2_X1 U15285 ( .A1(n12835), .A2(n12834), .ZN(n12820) );
  MUX2_X1 U15286 ( .A(n14959), .B(n14947), .S(n12821), .Z(n12846) );
  MUX2_X1 U15287 ( .A(n14769), .B(n15220), .S(n12862), .Z(n12845) );
  AND2_X1 U15288 ( .A1(n12846), .A2(n12845), .ZN(n12822) );
  OAI21_X1 U15289 ( .B1(n12833), .B2(n12832), .A(n12831), .ZN(n12830) );
  MUX2_X1 U15290 ( .A(n14990), .B(n14980), .S(n12862), .Z(n12827) );
  MUX2_X1 U15291 ( .A(n14771), .B(n15236), .S(n12681), .Z(n12826) );
  OAI22_X1 U15292 ( .A1(n12827), .A2(n12826), .B1(n12824), .B2(n12823), .ZN(
        n12825) );
  INV_X1 U15293 ( .A(n12826), .ZN(n12829) );
  INV_X1 U15294 ( .A(n12827), .ZN(n12828) );
  NOR3_X1 U15295 ( .A1(n12830), .A2(n12829), .A3(n12828), .ZN(n12853) );
  INV_X1 U15296 ( .A(n12831), .ZN(n12851) );
  NAND2_X1 U15297 ( .A1(n12833), .A2(n12832), .ZN(n12850) );
  INV_X1 U15298 ( .A(n12834), .ZN(n12837) );
  INV_X1 U15299 ( .A(n12835), .ZN(n12836) );
  NAND2_X1 U15300 ( .A1(n12837), .A2(n12836), .ZN(n12839) );
  NAND2_X1 U15301 ( .A1(n12840), .A2(n12839), .ZN(n12844) );
  INV_X1 U15302 ( .A(n12838), .ZN(n12843) );
  INV_X1 U15303 ( .A(n12839), .ZN(n12842) );
  INV_X1 U15304 ( .A(n12840), .ZN(n12841) );
  AOI22_X1 U15305 ( .A1(n12844), .A2(n12843), .B1(n12842), .B2(n12841), .ZN(
        n12849) );
  OR3_X1 U15306 ( .A1(n12847), .A2(n12846), .A3(n12845), .ZN(n12848) );
  OAI211_X1 U15307 ( .C1(n12851), .C2(n12850), .A(n12849), .B(n12848), .ZN(
        n12852) );
  NAND2_X1 U15308 ( .A1(n14579), .A2(n12393), .ZN(n12857) );
  NAND2_X1 U15309 ( .A1(n12855), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n12856) );
  NOR2_X1 U15310 ( .A1(n14916), .A2(n12862), .ZN(n12902) );
  NAND2_X1 U15311 ( .A1(n12859), .A2(n12858), .ZN(n12860) );
  NAND2_X1 U15312 ( .A1(n12861), .A2(n12860), .ZN(n12903) );
  NAND2_X1 U15313 ( .A1(n12903), .A2(n12907), .ZN(n12898) );
  NAND2_X1 U15314 ( .A1(n14916), .A2(n12862), .ZN(n12900) );
  NOR2_X1 U15315 ( .A1(n12900), .A2(n14918), .ZN(n12863) );
  AOI211_X1 U15316 ( .C1(n12902), .C2(n14918), .A(n12898), .B(n12863), .ZN(
        n12864) );
  INV_X1 U15317 ( .A(n14918), .ZN(n12866) );
  XNOR2_X1 U15318 ( .A(n14916), .B(n12866), .ZN(n12868) );
  NOR2_X1 U15319 ( .A1(n12868), .A2(n12903), .ZN(n12867) );
  INV_X1 U15320 ( .A(n12868), .ZN(n12897) );
  NOR2_X1 U15321 ( .A1(n12870), .A2(n12869), .ZN(n12873) );
  NAND4_X1 U15322 ( .A1(n12874), .A2(n12873), .A3(n12872), .A4(n12871), .ZN(
        n12876) );
  NOR2_X1 U15323 ( .A1(n12876), .A2(n12875), .ZN(n12879) );
  NAND4_X1 U15324 ( .A1(n12880), .A2(n12879), .A3(n12878), .A4(n12877), .ZN(
        n12881) );
  NOR2_X1 U15325 ( .A1(n12882), .A2(n12881), .ZN(n12884) );
  NAND4_X1 U15326 ( .A1(n12886), .A2(n12885), .A3(n12884), .A4(n12883), .ZN(
        n12887) );
  OR4_X1 U15327 ( .A1(n15193), .A2(n15149), .A3(n12888), .A4(n12887), .ZN(
        n12889) );
  NOR2_X1 U15328 ( .A1(n15100), .A2(n12890), .ZN(n12891) );
  NAND4_X1 U15329 ( .A1(n14999), .A2(n12892), .A3(n15029), .A4(n15062), .ZN(
        n12893) );
  NOR4_X1 U15330 ( .A1(n14933), .A2(n14955), .A3(n14969), .A4(n12893), .ZN(
        n12896) );
  XNOR2_X1 U15331 ( .A(n14923), .B(n14767), .ZN(n12894) );
  NOR3_X1 U15332 ( .A1(n15201), .A2(n14918), .A3(n12898), .ZN(n12901) );
  NOR3_X1 U15333 ( .A1(n12900), .A2(n14918), .A3(n12903), .ZN(n12899) );
  AOI21_X1 U15334 ( .B1(n12901), .B2(n12900), .A(n12899), .ZN(n12906) );
  XOR2_X1 U15335 ( .A(n12903), .B(n12902), .Z(n12904) );
  NAND3_X1 U15336 ( .A1(n12904), .A2(n15201), .A3(n14918), .ZN(n12905) );
  OAI211_X1 U15337 ( .C1(n12908), .C2(n12907), .A(n12906), .B(n12905), .ZN(
        n12909) );
  NAND3_X1 U15338 ( .A1(n12913), .A2(n12912), .A3(n15180), .ZN(n12914) );
  OAI211_X1 U15339 ( .C1(n15381), .C2(n12915), .A(n12914), .B(P1_B_REG_SCAN_IN), .ZN(n12916) );
  OAI222_X1 U15340 ( .A1(n15370), .A2(n16016), .B1(n15379), .B2(n12918), .C1(
        P1_U3086), .C2(n12917), .ZN(P1_U3334) );
  XNOR2_X1 U15341 ( .A(n13566), .B(n12995), .ZN(n12991) );
  XNOR2_X1 U15342 ( .A(n12991), .B(n13089), .ZN(n12993) );
  XNOR2_X1 U15343 ( .A(n13649), .B(n12995), .ZN(n12973) );
  INV_X1 U15344 ( .A(n12919), .ZN(n12920) );
  NAND2_X1 U15345 ( .A1(n12920), .A2(n13059), .ZN(n12921) );
  XNOR2_X1 U15346 ( .A(n13555), .B(n12995), .ZN(n13056) );
  AND2_X1 U15347 ( .A1(n13056), .A2(n13534), .ZN(n12922) );
  XNOR2_X1 U15348 ( .A(n13689), .B(n7247), .ZN(n12923) );
  XNOR2_X1 U15349 ( .A(n12923), .B(n13100), .ZN(n12965) );
  NAND2_X1 U15350 ( .A1(n12923), .A2(n13548), .ZN(n12924) );
  NAND2_X1 U15351 ( .A1(n12925), .A2(n12924), .ZN(n13094) );
  XNOR2_X1 U15352 ( .A(n13685), .B(n7247), .ZN(n12926) );
  XNOR2_X1 U15353 ( .A(n12926), .B(n13111), .ZN(n13093) );
  NAND2_X1 U15354 ( .A1(n13094), .A2(n13093), .ZN(n12929) );
  INV_X1 U15355 ( .A(n12926), .ZN(n12927) );
  NAND2_X1 U15356 ( .A1(n12927), .A2(n13111), .ZN(n12928) );
  XNOR2_X1 U15357 ( .A(n13679), .B(n7247), .ZN(n12930) );
  XNOR2_X1 U15358 ( .A(n12930), .B(n13519), .ZN(n13019) );
  INV_X1 U15359 ( .A(n12930), .ZN(n12931) );
  NAND2_X1 U15360 ( .A1(n12931), .A2(n13519), .ZN(n12932) );
  XNOR2_X1 U15361 ( .A(n13672), .B(n7247), .ZN(n12934) );
  XNOR2_X1 U15362 ( .A(n12934), .B(n13504), .ZN(n13029) );
  NAND2_X1 U15363 ( .A1(n12934), .A2(n13504), .ZN(n12935) );
  XNOR2_X1 U15364 ( .A(n13597), .B(n7247), .ZN(n12936) );
  XNOR2_X1 U15365 ( .A(n12936), .B(n13490), .ZN(n13073) );
  INV_X1 U15366 ( .A(n12936), .ZN(n12937) );
  NAND2_X1 U15367 ( .A1(n12937), .A2(n13109), .ZN(n12938) );
  XNOR2_X1 U15368 ( .A(n13593), .B(n7247), .ZN(n12939) );
  XNOR2_X1 U15369 ( .A(n12939), .B(n13476), .ZN(n12983) );
  NAND2_X1 U15370 ( .A1(n12984), .A2(n12983), .ZN(n12941) );
  NAND2_X1 U15371 ( .A1(n12939), .A2(n13108), .ZN(n12940) );
  NAND2_X1 U15372 ( .A1(n12941), .A2(n12940), .ZN(n13048) );
  XNOR2_X1 U15373 ( .A(n13590), .B(n7247), .ZN(n12942) );
  NAND2_X1 U15374 ( .A1(n12942), .A2(n13460), .ZN(n13046) );
  NAND2_X1 U15375 ( .A1(n13048), .A2(n13046), .ZN(n12944) );
  INV_X1 U15376 ( .A(n12942), .ZN(n12943) );
  NAND2_X1 U15377 ( .A1(n12943), .A2(n13107), .ZN(n13047) );
  XNOR2_X1 U15378 ( .A(n13434), .B(n7247), .ZN(n12945) );
  XNOR2_X1 U15379 ( .A(n12945), .B(n13446), .ZN(n13006) );
  NAND2_X1 U15380 ( .A1(n12945), .A2(n13446), .ZN(n12946) );
  XNOR2_X1 U15381 ( .A(n13580), .B(n7247), .ZN(n12977) );
  INV_X1 U15382 ( .A(n12977), .ZN(n13036) );
  AOI22_X1 U15383 ( .A1(n13036), .A2(n13421), .B1(n12973), .B2(n13106), .ZN(
        n12949) );
  XNOR2_X1 U15384 ( .A(n13396), .B(n7247), .ZN(n13038) );
  INV_X1 U15385 ( .A(n13038), .ZN(n12952) );
  AOI21_X1 U15386 ( .B1(n12977), .B2(n13069), .A(n13406), .ZN(n12951) );
  NAND3_X1 U15387 ( .A1(n12977), .A2(n13069), .A3(n13406), .ZN(n12950) );
  XNOR2_X1 U15388 ( .A(n13636), .B(n12995), .ZN(n12956) );
  XNOR2_X1 U15389 ( .A(n12956), .B(n13085), .ZN(n13013) );
  INV_X1 U15390 ( .A(n12956), .ZN(n12957) );
  XNOR2_X1 U15391 ( .A(n13629), .B(n12995), .ZN(n12958) );
  XNOR2_X1 U15392 ( .A(n12958), .B(n13375), .ZN(n13084) );
  XOR2_X1 U15393 ( .A(n12993), .B(n12994), .Z(n12964) );
  NOR2_X1 U15394 ( .A1(n13353), .A2(n13099), .ZN(n12962) );
  AOI22_X1 U15395 ( .A1(n13357), .A2(n13095), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12960) );
  OAI21_X1 U15396 ( .B1(n13352), .B2(n13088), .A(n12960), .ZN(n12961) );
  AOI211_X1 U15397 ( .C1(n13566), .C2(n13102), .A(n12962), .B(n12961), .ZN(
        n12963) );
  OAI21_X1 U15398 ( .B1(n12964), .B2(n13104), .A(n12963), .ZN(P3_U3154) );
  XNOR2_X1 U15399 ( .A(n12966), .B(n12965), .ZN(n12972) );
  INV_X1 U15400 ( .A(n13689), .ZN(n13529) );
  NAND2_X1 U15401 ( .A1(n13095), .A2(n13528), .ZN(n12969) );
  NAND2_X1 U15402 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n13203)
         );
  OAI21_X1 U15403 ( .B1(n13088), .B2(n13536), .A(n13203), .ZN(n12967) );
  INV_X1 U15404 ( .A(n12967), .ZN(n12968) );
  OAI211_X1 U15405 ( .C1(n13534), .C2(n13099), .A(n12969), .B(n12968), .ZN(
        n12970) );
  AOI21_X1 U15406 ( .B1(n13529), .B2(n13102), .A(n12970), .ZN(n12971) );
  OAI21_X1 U15407 ( .B1(n12972), .B2(n13104), .A(n12971), .ZN(P3_U3155) );
  INV_X1 U15408 ( .A(n12973), .ZN(n12974) );
  AND2_X1 U15409 ( .A1(n12975), .A2(n12974), .ZN(n12976) );
  XNOR2_X1 U15410 ( .A(n13037), .B(n13069), .ZN(n12982) );
  NOR2_X1 U15411 ( .A1(n13406), .A2(n13088), .ZN(n12980) );
  AOI22_X1 U15412 ( .A1(n13411), .A2(n13095), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12978) );
  OAI21_X1 U15413 ( .B1(n13433), .B2(n13099), .A(n12978), .ZN(n12979) );
  AOI211_X1 U15414 ( .C1(n13580), .C2(n13102), .A(n12980), .B(n12979), .ZN(
        n12981) );
  OAI21_X1 U15415 ( .B1(n12982), .B2(n13104), .A(n12981), .ZN(P3_U3156) );
  XNOR2_X1 U15416 ( .A(n12984), .B(n12983), .ZN(n12990) );
  NAND2_X1 U15417 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13320)
         );
  OAI21_X1 U15418 ( .B1(n13490), .B2(n13099), .A(n13320), .ZN(n12985) );
  AOI21_X1 U15419 ( .B1(n13107), .B2(n13096), .A(n12985), .ZN(n12987) );
  NAND2_X1 U15420 ( .A1(n13466), .A2(n13095), .ZN(n12986) );
  OAI211_X1 U15421 ( .C1(n13593), .C2(n13081), .A(n12987), .B(n12986), .ZN(
        n12988) );
  INV_X1 U15422 ( .A(n12988), .ZN(n12989) );
  OAI21_X1 U15423 ( .B1(n12990), .B2(n13104), .A(n12989), .ZN(P3_U3159) );
  INV_X1 U15424 ( .A(n12991), .ZN(n12992) );
  XNOR2_X1 U15425 ( .A(n12996), .B(n12995), .ZN(n12997) );
  NOR2_X1 U15426 ( .A1(n13089), .A2(n13099), .ZN(n13001) );
  AOI22_X1 U15427 ( .A1(n13343), .A2(n13095), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12998) );
  OAI21_X1 U15428 ( .B1(n12999), .B2(n13088), .A(n12998), .ZN(n13000) );
  AOI211_X1 U15429 ( .C1(n13002), .C2(n13102), .A(n13001), .B(n13000), .ZN(
        n13003) );
  OAI21_X1 U15430 ( .B1(n13004), .B2(n13104), .A(n13003), .ZN(P3_U3160) );
  XOR2_X1 U15431 ( .A(n13005), .B(n13006), .Z(n13011) );
  AOI22_X1 U15432 ( .A1(n13107), .A2(n13066), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13008) );
  NAND2_X1 U15433 ( .A1(n13435), .A2(n13095), .ZN(n13007) );
  OAI211_X1 U15434 ( .C1(n13433), .C2(n13088), .A(n13008), .B(n13007), .ZN(
        n13009) );
  AOI21_X1 U15435 ( .B1(n13434), .B2(n13102), .A(n13009), .ZN(n13010) );
  OAI21_X1 U15436 ( .B1(n13011), .B2(n13104), .A(n13010), .ZN(P3_U3163) );
  XOR2_X1 U15437 ( .A(n13013), .B(n13012), .Z(n13018) );
  AOI22_X1 U15438 ( .A1(n13379), .A2(n13095), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13015) );
  NAND2_X1 U15439 ( .A1(n13374), .A2(n13066), .ZN(n13014) );
  OAI211_X1 U15440 ( .C1(n13353), .C2(n13088), .A(n13015), .B(n13014), .ZN(
        n13016) );
  AOI21_X1 U15441 ( .B1(n13636), .B2(n13102), .A(n13016), .ZN(n13017) );
  OAI21_X1 U15442 ( .B1(n13018), .B2(n13104), .A(n13017), .ZN(P3_U3165) );
  XNOR2_X1 U15443 ( .A(n6774), .B(n13019), .ZN(n13025) );
  NAND2_X1 U15444 ( .A1(n13066), .A2(n13111), .ZN(n13021) );
  NAND2_X1 U15445 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13247)
         );
  OAI211_X1 U15446 ( .C1(n13504), .C2(n13088), .A(n13021), .B(n13247), .ZN(
        n13022) );
  AOI21_X1 U15447 ( .B1(n13508), .B2(n13095), .A(n13022), .ZN(n13024) );
  NAND2_X1 U15448 ( .A1(n13679), .A2(n13102), .ZN(n13023) );
  OAI211_X1 U15449 ( .C1(n13025), .C2(n13104), .A(n13024), .B(n13023), .ZN(
        P3_U3166) );
  INV_X1 U15450 ( .A(n13026), .ZN(n13027) );
  AOI21_X1 U15451 ( .B1(n13029), .B2(n13028), .A(n13027), .ZN(n13034) );
  AND2_X1 U15452 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13276) );
  AOI21_X1 U15453 ( .B1(n13109), .B2(n13096), .A(n13276), .ZN(n13031) );
  NAND2_X1 U15454 ( .A1(n13095), .A2(n13495), .ZN(n13030) );
  OAI211_X1 U15455 ( .C1(n13489), .C2(n13099), .A(n13031), .B(n13030), .ZN(
        n13032) );
  AOI21_X1 U15456 ( .B1(n13672), .B2(n13102), .A(n13032), .ZN(n13033) );
  OAI21_X1 U15457 ( .B1(n13034), .B2(n13104), .A(n13033), .ZN(P3_U3168) );
  XNOR2_X1 U15458 ( .A(n13038), .B(n13406), .ZN(n13039) );
  XNOR2_X1 U15459 ( .A(n13040), .B(n13039), .ZN(n13045) );
  NOR2_X1 U15460 ( .A1(n13085), .A2(n13088), .ZN(n13043) );
  AOI22_X1 U15461 ( .A1(n13397), .A2(n13095), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13041) );
  OAI21_X1 U15462 ( .B1(n13069), .B2(n13099), .A(n13041), .ZN(n13042) );
  AOI211_X1 U15463 ( .C1(n13396), .C2(n13102), .A(n13043), .B(n13042), .ZN(
        n13044) );
  OAI21_X1 U15464 ( .B1(n13045), .B2(n13104), .A(n13044), .ZN(P3_U3169) );
  NAND2_X1 U15465 ( .A1(n13047), .A2(n13046), .ZN(n13049) );
  XOR2_X1 U15466 ( .A(n13049), .B(n13048), .Z(n13054) );
  AOI22_X1 U15467 ( .A1(n13108), .A2(n13066), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13051) );
  NAND2_X1 U15468 ( .A1(n13451), .A2(n13095), .ZN(n13050) );
  OAI211_X1 U15469 ( .C1(n13446), .C2(n13088), .A(n13051), .B(n13050), .ZN(
        n13052) );
  AOI21_X1 U15470 ( .B1(n13590), .B2(n13102), .A(n13052), .ZN(n13053) );
  OAI21_X1 U15471 ( .B1(n13054), .B2(n13104), .A(n13053), .ZN(P3_U3173) );
  XNOR2_X1 U15472 ( .A(n13055), .B(n13534), .ZN(n13057) );
  XNOR2_X1 U15473 ( .A(n13057), .B(n13056), .ZN(n13063) );
  NAND2_X1 U15474 ( .A1(n13096), .A2(n13548), .ZN(n13058) );
  NAND2_X1 U15475 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n13177)
         );
  OAI211_X1 U15476 ( .C1(n13059), .C2(n13099), .A(n13058), .B(n13177), .ZN(
        n13061) );
  NOR2_X1 U15477 ( .A1(n13555), .A2(n13081), .ZN(n13060) );
  AOI211_X1 U15478 ( .C1(n13556), .C2(n13095), .A(n13061), .B(n13060), .ZN(
        n13062) );
  OAI21_X1 U15479 ( .B1(n13063), .B2(n13104), .A(n13062), .ZN(P3_U3174) );
  XNOR2_X1 U15480 ( .A(n13064), .B(n13106), .ZN(n13072) );
  AOI22_X1 U15481 ( .A1(n13420), .A2(n13066), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13068) );
  NAND2_X1 U15482 ( .A1(n13424), .A2(n13095), .ZN(n13067) );
  OAI211_X1 U15483 ( .C1(n13069), .C2(n13088), .A(n13068), .B(n13067), .ZN(
        n13070) );
  AOI21_X1 U15484 ( .B1(n13649), .B2(n13102), .A(n13070), .ZN(n13071) );
  OAI21_X1 U15485 ( .B1(n13072), .B2(n13104), .A(n13071), .ZN(P3_U3175) );
  INV_X1 U15486 ( .A(n13597), .ZN(n13082) );
  AOI21_X1 U15487 ( .B1(n13074), .B2(n13073), .A(n13104), .ZN(n13076) );
  NAND2_X1 U15488 ( .A1(n13076), .A2(n13075), .ZN(n13080) );
  AND2_X1 U15489 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13297) );
  AOI21_X1 U15490 ( .B1(n13108), .B2(n13096), .A(n13297), .ZN(n13077) );
  OAI21_X1 U15491 ( .B1(n13504), .B2(n13099), .A(n13077), .ZN(n13078) );
  AOI21_X1 U15492 ( .B1(n13477), .B2(n13095), .A(n13078), .ZN(n13079) );
  OAI211_X1 U15493 ( .C1(n13082), .C2(n13081), .A(n13080), .B(n13079), .ZN(
        P3_U3178) );
  XOR2_X1 U15494 ( .A(n13084), .B(n13083), .Z(n13092) );
  OAI22_X1 U15495 ( .A1(n13085), .A2(n13099), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n16003), .ZN(n13086) );
  AOI21_X1 U15496 ( .B1(n13366), .B2(n13095), .A(n13086), .ZN(n13087) );
  OAI21_X1 U15497 ( .B1(n13089), .B2(n13088), .A(n13087), .ZN(n13090) );
  AOI21_X1 U15498 ( .B1(n13629), .B2(n13102), .A(n13090), .ZN(n13091) );
  OAI21_X1 U15499 ( .B1(n13092), .B2(n13104), .A(n13091), .ZN(P3_U3180) );
  XNOR2_X1 U15500 ( .A(n13094), .B(n13093), .ZN(n13105) );
  NAND2_X1 U15501 ( .A1(n13095), .A2(n13513), .ZN(n13098) );
  AND2_X1 U15502 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13232) );
  AOI21_X1 U15503 ( .B1(n13096), .B2(n13519), .A(n13232), .ZN(n13097) );
  OAI211_X1 U15504 ( .C1(n13100), .C2(n13099), .A(n13098), .B(n13097), .ZN(
        n13101) );
  AOI21_X1 U15505 ( .B1(n13685), .B2(n13102), .A(n13101), .ZN(n13103) );
  OAI21_X1 U15506 ( .B1(n13105), .B2(n13104), .A(n13103), .ZN(P3_U3181) );
  MUX2_X1 U15507 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n13375), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U15508 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n13374), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15509 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n13421), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U15510 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n13106), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15511 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13420), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U15512 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13107), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15513 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n13108), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U15514 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13109), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15515 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13110), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U15516 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13519), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U15517 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n13111), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U15518 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13550), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15519 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n13112), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15520 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n13113), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15521 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n13114), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15522 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n13116), .S(n13115), .Z(
        P3_U3498) );
  MUX2_X1 U15523 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13117), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15524 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13118), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15525 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n13119), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U15526 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13120), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15527 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n13121), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15528 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n13122), .S(P3_U3897), .Z(
        P3_U3491) );
  AOI21_X1 U15529 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n13124), .A(n13123), 
        .ZN(n13125) );
  INV_X1 U15530 ( .A(n13153), .ZN(n13128) );
  NOR2_X1 U15531 ( .A1(n13125), .A2(n13128), .ZN(n13161) );
  AND2_X1 U15532 ( .A1(n13125), .A2(n13128), .ZN(n13126) );
  NAND2_X1 U15533 ( .A1(n13127), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n13165) );
  OAI21_X1 U15534 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n13127), .A(n13165), 
        .ZN(n13145) );
  NAND2_X1 U15535 ( .A1(n13323), .A2(n13128), .ZN(n13130) );
  OAI211_X1 U15536 ( .C1(n13131), .C2(n13321), .A(n13130), .B(n13129), .ZN(
        n13144) );
  AOI21_X1 U15537 ( .B1(n13136), .B2(n13135), .A(n6641), .ZN(n13142) );
  MUX2_X1 U15538 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13724), .Z(n13154) );
  XNOR2_X1 U15539 ( .A(n13153), .B(n13154), .ZN(n13155) );
  INV_X1 U15540 ( .A(n13137), .ZN(n13139) );
  AOI21_X1 U15541 ( .B1(n13140), .B2(n13139), .A(n13138), .ZN(n13156) );
  XOR2_X1 U15542 ( .A(n13155), .B(n13156), .Z(n13141) );
  OAI22_X1 U15543 ( .A1(n13142), .A2(n13190), .B1(n13141), .B2(n13210), .ZN(
        n13143) );
  AOI211_X1 U15544 ( .C1(n13318), .C2(n13145), .A(n13144), .B(n13143), .ZN(
        n13146) );
  INV_X1 U15545 ( .A(n13146), .ZN(P3_U3193) );
  INV_X1 U15546 ( .A(n13147), .ZN(n13149) );
  XNOR2_X1 U15547 ( .A(n13171), .B(P3_REG1_REG_12__SCAN_IN), .ZN(n13148) );
  NOR3_X1 U15548 ( .A1(n6641), .A2(n13149), .A3(n13148), .ZN(n13150) );
  OAI21_X1 U15549 ( .B1(n13170), .B2(n13150), .A(n13313), .ZN(n13169) );
  OAI21_X1 U15550 ( .B1(n13321), .B2(n13152), .A(n13151), .ZN(n13160) );
  MUX2_X1 U15551 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13724), .Z(n13175) );
  XOR2_X1 U15552 ( .A(n13171), .B(n13175), .Z(n13158) );
  OAI22_X1 U15553 ( .A1(n13156), .A2(n13155), .B1(n13154), .B2(n13153), .ZN(
        n13157) );
  NOR2_X1 U15554 ( .A1(n13157), .A2(n13158), .ZN(n13174) );
  AOI211_X1 U15555 ( .C1(n13158), .C2(n13157), .A(n13210), .B(n13174), .ZN(
        n13159) );
  AOI211_X1 U15556 ( .C1(n13323), .C2(n13171), .A(n13160), .B(n13159), .ZN(
        n13168) );
  INV_X1 U15557 ( .A(n13161), .ZN(n13163) );
  XNOR2_X1 U15558 ( .A(n13171), .B(n13162), .ZN(n13164) );
  AND3_X1 U15559 ( .A1(n13165), .A2(n13164), .A3(n13163), .ZN(n13166) );
  OAI21_X1 U15560 ( .B1(n13182), .B2(n13166), .A(n13318), .ZN(n13167) );
  NAND3_X1 U15561 ( .A1(n13169), .A2(n13168), .A3(n13167), .ZN(P3_U3194) );
  NAND2_X1 U15562 ( .A1(n13172), .A2(n13207), .ZN(n13196) );
  AOI21_X1 U15563 ( .B1(n13613), .B2(n13173), .A(n13199), .ZN(n13191) );
  MUX2_X1 U15564 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13724), .Z(n13208) );
  XOR2_X1 U15565 ( .A(n13207), .B(n13208), .Z(n13176) );
  OAI21_X1 U15566 ( .B1(n6743), .B2(n13176), .A(n13206), .ZN(n13181) );
  INV_X1 U15567 ( .A(n13207), .ZN(n13184) );
  NAND2_X1 U15568 ( .A1(n13323), .A2(n13184), .ZN(n13178) );
  OAI211_X1 U15569 ( .C1(n13179), .C2(n13321), .A(n13178), .B(n13177), .ZN(
        n13180) );
  AOI21_X1 U15570 ( .B1(n13181), .B2(n13332), .A(n13180), .ZN(n13189) );
  OAI21_X1 U15571 ( .B1(P3_REG2_REG_13__SCAN_IN), .B2(n13186), .A(n13194), 
        .ZN(n13187) );
  NAND2_X1 U15572 ( .A1(n13187), .A2(n13318), .ZN(n13188) );
  OAI211_X1 U15573 ( .C1(n13191), .C2(n13190), .A(n13189), .B(n13188), .ZN(
        P3_U3195) );
  NAND2_X1 U15574 ( .A1(n13202), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n13226) );
  OAI21_X1 U15575 ( .B1(n13202), .B2(P3_REG2_REG_14__SCAN_IN), .A(n13226), 
        .ZN(n13204) );
  INV_X1 U15576 ( .A(n13204), .ZN(n13192) );
  NOR2_X1 U15577 ( .A1(n13193), .A2(n13192), .ZN(n13195) );
  AOI21_X1 U15578 ( .B1(n13195), .B2(n13194), .A(n13220), .ZN(n13218) );
  INV_X1 U15579 ( .A(n13196), .ZN(n13197) );
  NAND2_X1 U15580 ( .A1(n13202), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13227) );
  OAI21_X1 U15581 ( .B1(n13202), .B2(P3_REG1_REG_14__SCAN_IN), .A(n13227), 
        .ZN(n13205) );
  INV_X1 U15582 ( .A(n13205), .ZN(n13198) );
  INV_X1 U15583 ( .A(n13222), .ZN(n13201) );
  NOR3_X1 U15584 ( .A1(n13199), .A2(n13198), .A3(n13197), .ZN(n13200) );
  OAI21_X1 U15585 ( .B1(n13201), .B2(n13200), .A(n13313), .ZN(n13217) );
  INV_X1 U15586 ( .A(n13202), .ZN(n13215) );
  INV_X1 U15587 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n16031) );
  OAI21_X1 U15588 ( .B1(n13321), .B2(n16031), .A(n13203), .ZN(n13214) );
  MUX2_X1 U15589 ( .A(n13205), .B(n13204), .S(n13328), .Z(n13212) );
  INV_X1 U15590 ( .A(n13229), .ZN(n13209) );
  AOI211_X1 U15591 ( .C1(n13212), .C2(n13211), .A(n13210), .B(n13209), .ZN(
        n13213) );
  AOI211_X1 U15592 ( .C1(n13323), .C2(n13215), .A(n13214), .B(n13213), .ZN(
        n13216) );
  OAI211_X1 U15593 ( .C1(n13218), .C2(n13283), .A(n13217), .B(n13216), .ZN(
        P3_U3196) );
  INV_X1 U15594 ( .A(n13226), .ZN(n13219) );
  AOI21_X1 U15595 ( .B1(n7675), .B2(n7676), .A(n13251), .ZN(n13239) );
  NAND2_X1 U15596 ( .A1(n13223), .A2(n13235), .ZN(n13242) );
  OAI21_X1 U15597 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n13225), .A(n13243), 
        .ZN(n13237) );
  MUX2_X1 U15598 ( .A(n13227), .B(n13226), .S(n13328), .Z(n13228) );
  XNOR2_X1 U15599 ( .A(n13254), .B(n13256), .ZN(n13231) );
  MUX2_X1 U15600 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n13724), .Z(n13230) );
  NAND2_X1 U15601 ( .A1(n13231), .A2(n13230), .ZN(n13255) );
  OAI211_X1 U15602 ( .C1(n13231), .C2(n13230), .A(n13255), .B(n13332), .ZN(
        n13234) );
  AOI21_X1 U15603 ( .B1(n15751), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n13232), 
        .ZN(n13233) );
  OAI211_X1 U15604 ( .C1(n13295), .C2(n13235), .A(n13234), .B(n13233), .ZN(
        n13236) );
  AOI21_X1 U15605 ( .B1(n13237), .B2(n13313), .A(n13236), .ZN(n13238) );
  OAI21_X1 U15606 ( .B1(n13239), .B2(n13283), .A(n13238), .ZN(P3_U3197) );
  INV_X1 U15607 ( .A(n13243), .ZN(n13241) );
  INV_X1 U15608 ( .A(n13242), .ZN(n13240) );
  INV_X1 U15609 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13605) );
  XNOR2_X1 U15610 ( .A(n13257), .B(n13605), .ZN(n13244) );
  NOR3_X1 U15611 ( .A1(n13241), .A2(n13240), .A3(n13244), .ZN(n13246) );
  INV_X1 U15612 ( .A(n13268), .ZN(n13245) );
  OAI21_X1 U15613 ( .B1(n13246), .B2(n13245), .A(n13313), .ZN(n13263) );
  INV_X1 U15614 ( .A(n13257), .ZN(n13273) );
  INV_X1 U15615 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15436) );
  OAI21_X1 U15616 ( .B1(n13321), .B2(n15436), .A(n13247), .ZN(n13248) );
  AOI21_X1 U15617 ( .B1(n13273), .B2(n13323), .A(n13248), .ZN(n13262) );
  INV_X1 U15618 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13507) );
  XNOR2_X1 U15619 ( .A(n13257), .B(n13507), .ZN(n13249) );
  INV_X1 U15620 ( .A(n13264), .ZN(n13253) );
  NOR3_X1 U15621 ( .A1(n13251), .A2(n13250), .A3(n13249), .ZN(n13252) );
  OAI21_X1 U15622 ( .B1(n13253), .B2(n13252), .A(n13318), .ZN(n13261) );
  MUX2_X1 U15623 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n13724), .Z(n13270) );
  XOR2_X1 U15624 ( .A(n13270), .B(n13257), .Z(n13258) );
  OAI211_X1 U15625 ( .C1(n13259), .C2(n13258), .A(n13271), .B(n13332), .ZN(
        n13260) );
  NAND4_X1 U15626 ( .A1(n13263), .A2(n13262), .A3(n13261), .A4(n13260), .ZN(
        P3_U3198) );
  INV_X1 U15627 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13494) );
  OAI21_X1 U15628 ( .B1(n13273), .B2(n13507), .A(n13264), .ZN(n13265) );
  NAND2_X1 U15629 ( .A1(n13265), .A2(n13279), .ZN(n13287) );
  INV_X1 U15630 ( .A(n13288), .ZN(n13266) );
  AOI21_X1 U15631 ( .B1(n13494), .B2(n13267), .A(n13266), .ZN(n13284) );
  OAI21_X1 U15632 ( .B1(n13273), .B2(n13605), .A(n13268), .ZN(n13269) );
  INV_X1 U15633 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13601) );
  OAI21_X1 U15634 ( .B1(n6593), .B2(P3_REG1_REG_17__SCAN_IN), .A(n13293), .ZN(
        n13281) );
  INV_X1 U15635 ( .A(n13270), .ZN(n13272) );
  MUX2_X1 U15636 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13724), .Z(n13298) );
  XNOR2_X1 U15637 ( .A(n13301), .B(n13298), .ZN(n13274) );
  OAI211_X1 U15638 ( .C1(n13275), .C2(n13274), .A(n13299), .B(n13332), .ZN(
        n13278) );
  AOI21_X1 U15639 ( .B1(n15751), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n13276), 
        .ZN(n13277) );
  OAI211_X1 U15640 ( .C1(n13295), .C2(n13279), .A(n13278), .B(n13277), .ZN(
        n13280) );
  AOI21_X1 U15641 ( .B1(n13281), .B2(n13313), .A(n13280), .ZN(n13282) );
  OAI21_X1 U15642 ( .B1(n13284), .B2(n13283), .A(n13282), .ZN(P3_U3199) );
  INV_X1 U15643 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13478) );
  OR2_X1 U15644 ( .A1(n13302), .A2(n13478), .ZN(n13315) );
  NAND2_X1 U15645 ( .A1(n13302), .A2(n13478), .ZN(n13285) );
  NAND2_X1 U15646 ( .A1(n13315), .A2(n13285), .ZN(n13286) );
  OAI21_X1 U15647 ( .B1(n13316), .B2(n13289), .A(n13318), .ZN(n13309) );
  INV_X1 U15648 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13599) );
  OR2_X1 U15649 ( .A1(n13302), .A2(n13599), .ZN(n13310) );
  NAND2_X1 U15650 ( .A1(n13302), .A2(n13599), .ZN(n13290) );
  NAND2_X1 U15651 ( .A1(n13310), .A2(n13290), .ZN(n13291) );
  AND3_X1 U15652 ( .A1(n13293), .A2(n13292), .A3(n13291), .ZN(n13294) );
  OAI21_X1 U15653 ( .B1(n13311), .B2(n13294), .A(n13313), .ZN(n13308) );
  NOR2_X1 U15654 ( .A1(n13295), .A2(n13326), .ZN(n13296) );
  AOI211_X1 U15655 ( .C1(n15751), .C2(P3_ADDR_REG_18__SCAN_IN), .A(n13297), 
        .B(n13296), .ZN(n13307) );
  INV_X1 U15656 ( .A(n13298), .ZN(n13300) );
  MUX2_X1 U15657 ( .A(n13478), .B(n13599), .S(n13724), .Z(n13303) );
  NAND2_X1 U15658 ( .A1(n13304), .A2(n13303), .ZN(n13325) );
  OAI21_X1 U15659 ( .B1(n13304), .B2(n13303), .A(n13325), .ZN(n13305) );
  NAND2_X1 U15660 ( .A1(n13305), .A2(n13332), .ZN(n13306) );
  XNOR2_X1 U15661 ( .A(n13324), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13330) );
  XNOR2_X1 U15662 ( .A(n13312), .B(n13330), .ZN(n13314) );
  XNOR2_X1 U15663 ( .A(n13324), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13329) );
  XNOR2_X1 U15664 ( .A(n13317), .B(n13329), .ZN(n13319) );
  NAND2_X1 U15665 ( .A1(n13319), .A2(n13318), .ZN(n13334) );
  OAI21_X1 U15666 ( .B1(n13321), .B2(n7792), .A(n13320), .ZN(n13322) );
  AOI21_X1 U15667 ( .B1(n13324), .B2(n13323), .A(n13322), .ZN(n13333) );
  MUX2_X1 U15668 ( .A(n13330), .B(n13329), .S(n13328), .Z(n13331) );
  AOI21_X1 U15669 ( .B1(n13619), .B2(n13553), .A(n13337), .ZN(n13341) );
  NAND2_X1 U15670 ( .A1(n13540), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13338) );
  OAI211_X1 U15671 ( .C1(n13339), .C2(n13456), .A(n13341), .B(n13338), .ZN(
        P3_U3202) );
  NAND2_X1 U15672 ( .A1(n13540), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13340) );
  OAI211_X1 U15673 ( .C1(n13565), .C2(n13456), .A(n13341), .B(n13340), .ZN(
        P3_U3203) );
  INV_X1 U15674 ( .A(n13342), .ZN(n13349) );
  AOI22_X1 U15675 ( .A1(n13343), .A2(n13557), .B1(P3_REG2_REG_28__SCAN_IN), 
        .B2(n13540), .ZN(n13344) );
  OAI21_X1 U15676 ( .B1(n13345), .B2(n13456), .A(n13344), .ZN(n13346) );
  AOI21_X1 U15677 ( .B1(n13347), .B2(n13553), .A(n13346), .ZN(n13348) );
  OAI21_X1 U15678 ( .B1(n13561), .B2(n13349), .A(n13348), .ZN(P3_U3205) );
  OAI21_X1 U15679 ( .B1(n13356), .B2(n13355), .A(n13354), .ZN(n13567) );
  AOI22_X1 U15680 ( .A1(n13357), .A2(n13557), .B1(P3_REG2_REG_27__SCAN_IN), 
        .B2(n13540), .ZN(n13358) );
  OAI21_X1 U15681 ( .B1(n9690), .B2(n13456), .A(n13358), .ZN(n13359) );
  AOI21_X1 U15682 ( .B1(n13567), .B2(n13360), .A(n13359), .ZN(n13361) );
  OAI21_X1 U15683 ( .B1(n6616), .B2(n13540), .A(n13361), .ZN(P3_U3206) );
  XNOR2_X1 U15684 ( .A(n13362), .B(n13363), .ZN(n13632) );
  INV_X1 U15685 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n13365) );
  XNOR2_X1 U15686 ( .A(n6637), .B(n13363), .ZN(n13364) );
  AOI222_X1 U15687 ( .A1(n13552), .A2(n13364), .B1(n9803), .B2(n13547), .C1(
        n13386), .C2(n13549), .ZN(n13627) );
  MUX2_X1 U15688 ( .A(n13365), .B(n13627), .S(n13553), .Z(n13368) );
  AOI22_X1 U15689 ( .A1(n13629), .A2(n13558), .B1(n13557), .B2(n13366), .ZN(
        n13367) );
  OAI211_X1 U15690 ( .C1(n13632), .C2(n13561), .A(n13368), .B(n13367), .ZN(
        P3_U3207) );
  XNOR2_X1 U15691 ( .A(n13369), .B(n13370), .ZN(n13637) );
  INV_X1 U15692 ( .A(n13637), .ZN(n13382) );
  NAND2_X1 U15693 ( .A1(n13371), .A2(n13370), .ZN(n13372) );
  NAND2_X1 U15694 ( .A1(n13372), .A2(n13552), .ZN(n13373) );
  OR2_X1 U15695 ( .A1(n6707), .A2(n13373), .ZN(n13377) );
  AOI22_X1 U15696 ( .A1(n13375), .A2(n13547), .B1(n13549), .B2(n13374), .ZN(
        n13376) );
  NAND2_X1 U15697 ( .A1(n13377), .A2(n13376), .ZN(n13633) );
  MUX2_X1 U15698 ( .A(n13633), .B(P3_REG2_REG_25__SCAN_IN), .S(n13540), .Z(
        n13378) );
  INV_X1 U15699 ( .A(n13378), .ZN(n13381) );
  AOI22_X1 U15700 ( .A1(n13636), .A2(n13558), .B1(n13557), .B2(n13379), .ZN(
        n13380) );
  OAI211_X1 U15701 ( .C1(n13561), .C2(n13382), .A(n13381), .B(n13380), .ZN(
        P3_U3208) );
  INV_X1 U15702 ( .A(n13383), .ZN(n13384) );
  AOI21_X1 U15703 ( .B1(n13390), .B2(n13385), .A(n13384), .ZN(n13395) );
  AOI22_X1 U15704 ( .A1(n13386), .A2(n13547), .B1(n13549), .B2(n13421), .ZN(
        n13393) );
  NAND2_X1 U15705 ( .A1(n13388), .A2(n13387), .ZN(n13389) );
  XOR2_X1 U15706 ( .A(n13390), .B(n13389), .Z(n13391) );
  NAND2_X1 U15707 ( .A1(n13391), .A2(n13552), .ZN(n13392) );
  OAI211_X1 U15708 ( .C1(n13395), .C2(n13394), .A(n13393), .B(n13392), .ZN(
        n13575) );
  INV_X1 U15709 ( .A(n13575), .ZN(n13402) );
  INV_X1 U15710 ( .A(n13395), .ZN(n13576) );
  INV_X1 U15711 ( .A(n13396), .ZN(n13643) );
  AOI22_X1 U15712 ( .A1(n13397), .A2(n13557), .B1(n13540), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n13398) );
  OAI21_X1 U15713 ( .B1(n13643), .B2(n13456), .A(n13398), .ZN(n13399) );
  AOI21_X1 U15714 ( .B1(n13576), .B2(n13400), .A(n13399), .ZN(n13401) );
  OAI21_X1 U15715 ( .B1(n13402), .B2(n13540), .A(n13401), .ZN(P3_U3209) );
  XNOR2_X1 U15716 ( .A(n13403), .B(n13404), .ZN(n13405) );
  OAI222_X1 U15717 ( .A1(n13533), .A2(n13433), .B1(n13535), .B2(n13406), .C1(
        n13405), .C2(n13502), .ZN(n13579) );
  OR2_X1 U15718 ( .A1(n13408), .A2(n13407), .ZN(n13409) );
  NAND2_X1 U15719 ( .A1(n13410), .A2(n13409), .ZN(n13646) );
  AOI22_X1 U15720 ( .A1(n13411), .A2(n13557), .B1(n13540), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n13413) );
  NAND2_X1 U15721 ( .A1(n13580), .A2(n13558), .ZN(n13412) );
  OAI211_X1 U15722 ( .C1(n13646), .C2(n13561), .A(n13413), .B(n13412), .ZN(
        n13414) );
  AOI21_X1 U15723 ( .B1(n13579), .B2(n13553), .A(n13414), .ZN(n13415) );
  INV_X1 U15724 ( .A(n13415), .ZN(P3_U3210) );
  XNOR2_X1 U15725 ( .A(n13416), .B(n13417), .ZN(n13652) );
  INV_X1 U15726 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13423) );
  XNOR2_X1 U15727 ( .A(n13419), .B(n13418), .ZN(n13422) );
  AOI222_X1 U15728 ( .A1(n13552), .A2(n13422), .B1(n13421), .B2(n13547), .C1(
        n13420), .C2(n13549), .ZN(n13647) );
  MUX2_X1 U15729 ( .A(n13423), .B(n13647), .S(n13553), .Z(n13426) );
  AOI22_X1 U15730 ( .A1(n13649), .A2(n13558), .B1(n13557), .B2(n13424), .ZN(
        n13425) );
  OAI211_X1 U15731 ( .C1(n13652), .C2(n13561), .A(n13426), .B(n13425), .ZN(
        P3_U3211) );
  XOR2_X1 U15732 ( .A(n13427), .B(n13431), .Z(n13587) );
  INV_X1 U15733 ( .A(n13587), .ZN(n13439) );
  INV_X1 U15734 ( .A(n13428), .ZN(n13429) );
  AOI21_X1 U15735 ( .B1(n13431), .B2(n13430), .A(n13429), .ZN(n13432) );
  OAI222_X1 U15736 ( .A1(n13535), .A2(n13433), .B1(n13533), .B2(n13460), .C1(
        n13502), .C2(n13432), .ZN(n13586) );
  INV_X1 U15737 ( .A(n13434), .ZN(n13656) );
  AOI22_X1 U15738 ( .A1(n13435), .A2(n13557), .B1(n13540), .B2(
        P3_REG2_REG_21__SCAN_IN), .ZN(n13436) );
  OAI21_X1 U15739 ( .B1(n13656), .B2(n13456), .A(n13436), .ZN(n13437) );
  AOI21_X1 U15740 ( .B1(n13586), .B2(n13553), .A(n13437), .ZN(n13438) );
  OAI21_X1 U15741 ( .B1(n13439), .B2(n13561), .A(n13438), .ZN(P3_U3212) );
  OAI21_X1 U15742 ( .B1(n13442), .B2(n13441), .A(n13440), .ZN(n13658) );
  OAI211_X1 U15743 ( .C1(n13445), .C2(n13444), .A(n13443), .B(n13552), .ZN(
        n13449) );
  OAI22_X1 U15744 ( .A1(n13446), .A2(n13535), .B1(n13476), .B2(n13533), .ZN(
        n13447) );
  INV_X1 U15745 ( .A(n13447), .ZN(n13448) );
  NAND2_X1 U15746 ( .A1(n13449), .A2(n13448), .ZN(n13659) );
  MUX2_X1 U15747 ( .A(n13659), .B(P3_REG2_REG_20__SCAN_IN), .S(n13540), .Z(
        n13450) );
  INV_X1 U15748 ( .A(n13450), .ZN(n13453) );
  AOI22_X1 U15749 ( .A1(n13590), .A2(n13558), .B1(n13557), .B2(n13451), .ZN(
        n13452) );
  OAI211_X1 U15750 ( .C1(n13658), .C2(n13561), .A(n13453), .B(n13452), .ZN(
        P3_U3213) );
  NAND2_X1 U15751 ( .A1(n13470), .A2(n13454), .ZN(n13455) );
  XOR2_X1 U15752 ( .A(n13458), .B(n13455), .Z(n13666) );
  NOR2_X1 U15753 ( .A1(n13593), .A2(n13456), .ZN(n13465) );
  OAI211_X1 U15754 ( .C1(n13459), .C2(n13458), .A(n13457), .B(n13552), .ZN(
        n13463) );
  OAI22_X1 U15755 ( .A1(n13460), .A2(n13535), .B1(n13490), .B2(n13533), .ZN(
        n13461) );
  INV_X1 U15756 ( .A(n13461), .ZN(n13462) );
  NAND2_X1 U15757 ( .A1(n13463), .A2(n13462), .ZN(n13662) );
  MUX2_X1 U15758 ( .A(n13662), .B(P3_REG2_REG_19__SCAN_IN), .S(n13540), .Z(
        n13464) );
  AOI211_X1 U15759 ( .C1(n13557), .C2(n13466), .A(n13465), .B(n13464), .ZN(
        n13467) );
  OAI21_X1 U15760 ( .B1(n13666), .B2(n13561), .A(n13467), .ZN(P3_U3214) );
  NAND2_X1 U15761 ( .A1(n13468), .A2(n13473), .ZN(n13469) );
  NAND2_X1 U15762 ( .A1(n13470), .A2(n13469), .ZN(n13669) );
  OAI21_X1 U15763 ( .B1(n6620), .B2(n13472), .A(n13471), .ZN(n13474) );
  XNOR2_X1 U15764 ( .A(n13474), .B(n13473), .ZN(n13475) );
  OAI222_X1 U15765 ( .A1(n13533), .A2(n13504), .B1(n13535), .B2(n13476), .C1(
        n13475), .C2(n13502), .ZN(n13596) );
  NAND2_X1 U15766 ( .A1(n13596), .A2(n13553), .ZN(n13483) );
  INV_X1 U15767 ( .A(n13477), .ZN(n13480) );
  OAI22_X1 U15768 ( .A1(n13480), .A2(n13479), .B1(n13553), .B2(n13478), .ZN(
        n13481) );
  AOI21_X1 U15769 ( .B1(n13597), .B2(n13558), .A(n13481), .ZN(n13482) );
  OAI211_X1 U15770 ( .C1(n13669), .C2(n13561), .A(n13483), .B(n13482), .ZN(
        P3_U3215) );
  XNOR2_X1 U15771 ( .A(n13484), .B(n13485), .ZN(n13674) );
  INV_X1 U15772 ( .A(n13674), .ZN(n13498) );
  NOR3_X1 U15773 ( .A1(n13501), .A2(n13488), .A3(n13487), .ZN(n13486) );
  NOR2_X1 U15774 ( .A1(n13486), .A2(n13502), .ZN(n13493) );
  OAI21_X1 U15775 ( .B1(n13501), .B2(n13488), .A(n13487), .ZN(n13492) );
  OAI22_X1 U15776 ( .A1(n13490), .A2(n13535), .B1(n13489), .B2(n13533), .ZN(
        n13491) );
  AOI21_X1 U15777 ( .B1(n13493), .B2(n13492), .A(n13491), .ZN(n13670) );
  MUX2_X1 U15778 ( .A(n13494), .B(n13670), .S(n13553), .Z(n13497) );
  AOI22_X1 U15779 ( .A1(n13672), .A2(n13558), .B1(n13557), .B2(n13495), .ZN(
        n13496) );
  OAI211_X1 U15780 ( .C1(n13498), .C2(n13561), .A(n13497), .B(n13496), .ZN(
        P3_U3216) );
  XNOR2_X1 U15781 ( .A(n13500), .B(n13499), .ZN(n13682) );
  AOI211_X1 U15782 ( .C1(n13503), .C2(n6620), .A(n13502), .B(n13501), .ZN(
        n13506) );
  OAI22_X1 U15783 ( .A1(n13504), .A2(n13535), .B1(n13536), .B2(n13533), .ZN(
        n13505) );
  NOR2_X1 U15784 ( .A1(n13506), .A2(n13505), .ZN(n13677) );
  MUX2_X1 U15785 ( .A(n13507), .B(n13677), .S(n13553), .Z(n13510) );
  AOI22_X1 U15786 ( .A1(n13679), .A2(n13558), .B1(n13557), .B2(n13508), .ZN(
        n13509) );
  OAI211_X1 U15787 ( .C1(n13682), .C2(n13561), .A(n13510), .B(n13509), .ZN(
        P3_U3217) );
  NOR2_X1 U15788 ( .A1(n13526), .A2(n13527), .ZN(n13525) );
  NOR2_X1 U15789 ( .A1(n13525), .A2(n13511), .ZN(n13512) );
  XOR2_X1 U15790 ( .A(n13515), .B(n13512), .Z(n13687) );
  AOI22_X1 U15791 ( .A1(n13685), .A2(n13558), .B1(n13557), .B2(n13513), .ZN(
        n13524) );
  NAND3_X1 U15792 ( .A1(n13514), .A2(n6888), .A3(n13516), .ZN(n13517) );
  NAND3_X1 U15793 ( .A1(n13518), .A2(n13552), .A3(n13517), .ZN(n13521) );
  AOI22_X1 U15794 ( .A1(n13519), .A2(n13547), .B1(n13549), .B2(n13548), .ZN(
        n13520) );
  NAND2_X1 U15795 ( .A1(n13521), .A2(n13520), .ZN(n13683) );
  INV_X1 U15796 ( .A(n13683), .ZN(n13522) );
  MUX2_X1 U15797 ( .A(n13522), .B(n7675), .S(n13540), .Z(n13523) );
  OAI211_X1 U15798 ( .C1(n13687), .C2(n13561), .A(n13524), .B(n13523), .ZN(
        P3_U3218) );
  AOI21_X1 U15799 ( .B1(n13527), .B2(n13526), .A(n13525), .ZN(n13690) );
  AOI22_X1 U15800 ( .A1(n13529), .A2(n13558), .B1(n13557), .B2(n13528), .ZN(
        n13543) );
  NAND2_X1 U15801 ( .A1(n13531), .A2(n13530), .ZN(n13532) );
  NAND3_X1 U15802 ( .A1(n13514), .A2(n13552), .A3(n13532), .ZN(n13539) );
  OAI22_X1 U15803 ( .A1(n13536), .A2(n13535), .B1(n13534), .B2(n13533), .ZN(
        n13537) );
  INV_X1 U15804 ( .A(n13537), .ZN(n13538) );
  NAND2_X1 U15805 ( .A1(n13539), .A2(n13538), .ZN(n13691) );
  MUX2_X1 U15806 ( .A(n13691), .B(P3_REG2_REG_14__SCAN_IN), .S(n13540), .Z(
        n13541) );
  INV_X1 U15807 ( .A(n13541), .ZN(n13542) );
  OAI211_X1 U15808 ( .C1(n13690), .C2(n13561), .A(n13543), .B(n13542), .ZN(
        P3_U3219) );
  XNOR2_X1 U15809 ( .A(n13545), .B(n13544), .ZN(n13700) );
  XNOR2_X1 U15810 ( .A(n13546), .B(n7443), .ZN(n13551) );
  AOI222_X1 U15811 ( .A1(n13552), .A2(n13551), .B1(n13550), .B2(n13549), .C1(
        n13548), .C2(n13547), .ZN(n13694) );
  MUX2_X1 U15812 ( .A(n13554), .B(n13694), .S(n13553), .Z(n13560) );
  INV_X1 U15813 ( .A(n13555), .ZN(n13696) );
  AOI22_X1 U15814 ( .A1(n13696), .A2(n13558), .B1(n13557), .B2(n13556), .ZN(
        n13559) );
  OAI211_X1 U15815 ( .C1(n13700), .C2(n13561), .A(n13560), .B(n13559), .ZN(
        P3_U3220) );
  NAND2_X1 U15816 ( .A1(n13618), .A2(n13614), .ZN(n13562) );
  NAND2_X1 U15817 ( .A1(n13619), .A2(n15804), .ZN(n13563) );
  OAI211_X1 U15818 ( .C1(n15804), .C2(n16010), .A(n13562), .B(n13563), .ZN(
        P3_U3490) );
  NAND2_X1 U15819 ( .A1(n15801), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n13564) );
  OAI211_X1 U15820 ( .C1(n13565), .C2(n13610), .A(n13564), .B(n13563), .ZN(
        P3_U3489) );
  AOI22_X1 U15821 ( .A1(n13567), .A2(n15755), .B1(n13598), .B2(n13566), .ZN(
        n13568) );
  NAND2_X1 U15822 ( .A1(n6616), .A2(n13568), .ZN(n13626) );
  MUX2_X1 U15823 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n13626), .S(n15804), .Z(
        P3_U3486) );
  INV_X1 U15824 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13569) );
  MUX2_X1 U15825 ( .A(n13569), .B(n13627), .S(n15804), .Z(n13571) );
  NAND2_X1 U15826 ( .A1(n13629), .A2(n13614), .ZN(n13570) );
  OAI211_X1 U15827 ( .C1(n13617), .C2(n13632), .A(n13571), .B(n13570), .ZN(
        P3_U3485) );
  MUX2_X1 U15828 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13633), .S(n15804), .Z(
        n13572) );
  INV_X1 U15829 ( .A(n13572), .ZN(n13574) );
  AOI22_X1 U15830 ( .A1(n13637), .A2(n13602), .B1(n13614), .B2(n13636), .ZN(
        n13573) );
  NAND2_X1 U15831 ( .A1(n13574), .A2(n13573), .ZN(P3_U3484) );
  INV_X1 U15832 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13577) );
  AOI21_X1 U15833 ( .B1(n15784), .B2(n13576), .A(n13575), .ZN(n13640) );
  MUX2_X1 U15834 ( .A(n13577), .B(n13640), .S(n15804), .Z(n13578) );
  OAI21_X1 U15835 ( .B1(n13643), .B2(n13610), .A(n13578), .ZN(P3_U3483) );
  INV_X1 U15836 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13581) );
  AOI21_X1 U15837 ( .B1(n13598), .B2(n13580), .A(n13579), .ZN(n13644) );
  MUX2_X1 U15838 ( .A(n13581), .B(n13644), .S(n15804), .Z(n13582) );
  OAI21_X1 U15839 ( .B1(n13617), .B2(n13646), .A(n13582), .ZN(P3_U3482) );
  INV_X1 U15840 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13583) );
  MUX2_X1 U15841 ( .A(n13583), .B(n13647), .S(n15804), .Z(n13585) );
  NAND2_X1 U15842 ( .A1(n13649), .A2(n13614), .ZN(n13584) );
  OAI211_X1 U15843 ( .C1(n13652), .C2(n13617), .A(n13585), .B(n13584), .ZN(
        P3_U3481) );
  INV_X1 U15844 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13588) );
  AOI21_X1 U15845 ( .B1(n15755), .B2(n13587), .A(n13586), .ZN(n13653) );
  MUX2_X1 U15846 ( .A(n13588), .B(n13653), .S(n15804), .Z(n13589) );
  OAI21_X1 U15847 ( .B1(n13656), .B2(n13610), .A(n13589), .ZN(P3_U3480) );
  INV_X1 U15848 ( .A(n13590), .ZN(n13657) );
  OAI22_X1 U15849 ( .A1(n13658), .A2(n13617), .B1(n13657), .B2(n13610), .ZN(
        n13592) );
  MUX2_X1 U15850 ( .A(n13659), .B(P3_REG1_REG_20__SCAN_IN), .S(n15801), .Z(
        n13591) );
  OR2_X1 U15851 ( .A1(n13592), .A2(n13591), .ZN(P3_U3479) );
  INV_X1 U15852 ( .A(n13593), .ZN(n13664) );
  MUX2_X1 U15853 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n13662), .S(n15804), .Z(
        n13594) );
  AOI21_X1 U15854 ( .B1(n13614), .B2(n13664), .A(n13594), .ZN(n13595) );
  OAI21_X1 U15855 ( .B1(n13666), .B2(n13617), .A(n13595), .ZN(P3_U3478) );
  AOI21_X1 U15856 ( .B1(n13598), .B2(n13597), .A(n13596), .ZN(n13667) );
  MUX2_X1 U15857 ( .A(n13599), .B(n13667), .S(n15804), .Z(n13600) );
  OAI21_X1 U15858 ( .B1(n13617), .B2(n13669), .A(n13600), .ZN(P3_U3477) );
  MUX2_X1 U15859 ( .A(n13601), .B(n13670), .S(n15804), .Z(n13604) );
  AOI22_X1 U15860 ( .A1(n13674), .A2(n13602), .B1(n13614), .B2(n13672), .ZN(
        n13603) );
  NAND2_X1 U15861 ( .A1(n13604), .A2(n13603), .ZN(P3_U3476) );
  MUX2_X1 U15862 ( .A(n13605), .B(n13677), .S(n15804), .Z(n13607) );
  NAND2_X1 U15863 ( .A1(n13679), .A2(n13614), .ZN(n13606) );
  OAI211_X1 U15864 ( .C1(n13617), .C2(n13682), .A(n13607), .B(n13606), .ZN(
        P3_U3475) );
  MUX2_X1 U15865 ( .A(n13683), .B(P3_REG1_REG_15__SCAN_IN), .S(n15801), .Z(
        n13608) );
  AOI21_X1 U15866 ( .B1(n13614), .B2(n13685), .A(n13608), .ZN(n13609) );
  OAI21_X1 U15867 ( .B1(n13687), .B2(n13617), .A(n13609), .ZN(P3_U3474) );
  OAI22_X1 U15868 ( .A1(n13690), .A2(n13617), .B1(n13689), .B2(n13610), .ZN(
        n13612) );
  MUX2_X1 U15869 ( .A(n13691), .B(P3_REG1_REG_14__SCAN_IN), .S(n15801), .Z(
        n13611) );
  OR2_X1 U15870 ( .A1(n13612), .A2(n13611), .ZN(P3_U3473) );
  MUX2_X1 U15871 ( .A(n13613), .B(n13694), .S(n15804), .Z(n13616) );
  NAND2_X1 U15872 ( .A1(n13696), .A2(n13614), .ZN(n13615) );
  OAI211_X1 U15873 ( .C1(n13617), .C2(n13700), .A(n13616), .B(n13615), .ZN(
        P3_U3472) );
  NAND2_X1 U15874 ( .A1(n13618), .A2(n13695), .ZN(n13620) );
  NAND2_X1 U15875 ( .A1(n13619), .A2(n15786), .ZN(n13623) );
  OAI211_X1 U15876 ( .C1(n15786), .C2(n13621), .A(n13620), .B(n13623), .ZN(
        P3_U3458) );
  NAND2_X1 U15877 ( .A1(n13622), .A2(n13695), .ZN(n13624) );
  OAI211_X1 U15878 ( .C1(n15786), .C2(n13625), .A(n13624), .B(n13623), .ZN(
        P3_U3457) );
  MUX2_X1 U15879 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n13626), .S(n15786), .Z(
        P3_U3454) );
  MUX2_X1 U15880 ( .A(n13628), .B(n13627), .S(n15786), .Z(n13631) );
  NAND2_X1 U15881 ( .A1(n13629), .A2(n13695), .ZN(n13630) );
  OAI211_X1 U15882 ( .C1(n13632), .C2(n13699), .A(n13631), .B(n13630), .ZN(
        P3_U3453) );
  INV_X1 U15883 ( .A(n13633), .ZN(n13635) );
  MUX2_X1 U15884 ( .A(n13635), .B(n13634), .S(n15788), .Z(n13639) );
  AOI22_X1 U15885 ( .A1(n13637), .A2(n13673), .B1(n13695), .B2(n13636), .ZN(
        n13638) );
  NAND2_X1 U15886 ( .A1(n13639), .A2(n13638), .ZN(P3_U3452) );
  MUX2_X1 U15887 ( .A(n13641), .B(n13640), .S(n15786), .Z(n13642) );
  OAI21_X1 U15888 ( .B1(n13643), .B2(n13688), .A(n13642), .ZN(P3_U3451) );
  MUX2_X1 U15889 ( .A(n15999), .B(n13644), .S(n15786), .Z(n13645) );
  OAI21_X1 U15890 ( .B1(n13646), .B2(n13699), .A(n13645), .ZN(P3_U3450) );
  MUX2_X1 U15891 ( .A(n13648), .B(n13647), .S(n15786), .Z(n13651) );
  NAND2_X1 U15892 ( .A1(n13649), .A2(n13695), .ZN(n13650) );
  OAI211_X1 U15893 ( .C1(n13652), .C2(n13699), .A(n13651), .B(n13650), .ZN(
        P3_U3449) );
  MUX2_X1 U15894 ( .A(n13654), .B(n13653), .S(n15786), .Z(n13655) );
  OAI21_X1 U15895 ( .B1(n13656), .B2(n13688), .A(n13655), .ZN(P3_U3448) );
  OAI22_X1 U15896 ( .A1(n13658), .A2(n13699), .B1(n13657), .B2(n13688), .ZN(
        n13661) );
  MUX2_X1 U15897 ( .A(n13659), .B(P3_REG0_REG_20__SCAN_IN), .S(n15788), .Z(
        n13660) );
  OR2_X1 U15898 ( .A1(n13661), .A2(n13660), .ZN(P3_U3447) );
  MUX2_X1 U15899 ( .A(n13662), .B(P3_REG0_REG_19__SCAN_IN), .S(n15788), .Z(
        n13663) );
  AOI21_X1 U15900 ( .B1(n13695), .B2(n13664), .A(n13663), .ZN(n13665) );
  OAI21_X1 U15901 ( .B1(n13666), .B2(n13699), .A(n13665), .ZN(P3_U3446) );
  MUX2_X1 U15902 ( .A(n16057), .B(n13667), .S(n15786), .Z(n13668) );
  OAI21_X1 U15903 ( .B1(n13669), .B2(n13699), .A(n13668), .ZN(P3_U3444) );
  MUX2_X1 U15904 ( .A(n13671), .B(n13670), .S(n15786), .Z(n13676) );
  AOI22_X1 U15905 ( .A1(n13674), .A2(n13673), .B1(n13695), .B2(n13672), .ZN(
        n13675) );
  NAND2_X1 U15906 ( .A1(n13676), .A2(n13675), .ZN(P3_U3441) );
  MUX2_X1 U15907 ( .A(n13678), .B(n13677), .S(n15786), .Z(n13681) );
  NAND2_X1 U15908 ( .A1(n13679), .A2(n13695), .ZN(n13680) );
  OAI211_X1 U15909 ( .C1(n13682), .C2(n13699), .A(n13681), .B(n13680), .ZN(
        P3_U3438) );
  MUX2_X1 U15910 ( .A(n13683), .B(P3_REG0_REG_15__SCAN_IN), .S(n15788), .Z(
        n13684) );
  AOI21_X1 U15911 ( .B1(n13695), .B2(n13685), .A(n13684), .ZN(n13686) );
  OAI21_X1 U15912 ( .B1(n13687), .B2(n13699), .A(n13686), .ZN(P3_U3435) );
  OAI22_X1 U15913 ( .A1(n13690), .A2(n13699), .B1(n13689), .B2(n13688), .ZN(
        n13693) );
  MUX2_X1 U15914 ( .A(n13691), .B(P3_REG0_REG_14__SCAN_IN), .S(n15788), .Z(
        n13692) );
  OR2_X1 U15915 ( .A1(n13693), .A2(n13692), .ZN(P3_U3432) );
  MUX2_X1 U15916 ( .A(n15873), .B(n13694), .S(n15786), .Z(n13698) );
  NAND2_X1 U15917 ( .A1(n13696), .A2(n13695), .ZN(n13697) );
  OAI211_X1 U15918 ( .C1(n13700), .C2(n13699), .A(n13698), .B(n13697), .ZN(
        P3_U3429) );
  MUX2_X1 U15919 ( .A(n13701), .B(P3_D_REG_1__SCAN_IN), .S(n13702), .Z(
        P3_U3377) );
  MUX2_X1 U15920 ( .A(n13703), .B(P3_D_REG_0__SCAN_IN), .S(n13702), .Z(
        P3_U3376) );
  INV_X1 U15921 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13704) );
  NAND3_X1 U15922 ( .A1(n13704), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n13706) );
  OAI22_X1 U15923 ( .A1(n13707), .A2(n13706), .B1(n13705), .B2(n13723), .ZN(
        n13708) );
  AOI21_X1 U15924 ( .B1(n13710), .B2(n13709), .A(n13708), .ZN(n13711) );
  INV_X1 U15925 ( .A(n13711), .ZN(P3_U3264) );
  INV_X1 U15926 ( .A(n13712), .ZN(n13713) );
  OAI222_X1 U15927 ( .A1(P3_U3151), .A2(n13714), .B1(n13723), .B2(n16017), 
        .C1(n13721), .C2(n13713), .ZN(P3_U3265) );
  INV_X1 U15928 ( .A(n13715), .ZN(n13717) );
  OAI222_X1 U15929 ( .A1(n13723), .A2(n13718), .B1(n13721), .B2(n13717), .C1(
        P3_U3151), .C2(n13716), .ZN(P3_U3267) );
  INV_X1 U15930 ( .A(n13719), .ZN(n13720) );
  OAI222_X1 U15931 ( .A1(P3_U3151), .A2(n13724), .B1(n13723), .B2(n13722), 
        .C1(n13721), .C2(n13720), .ZN(P3_U3268) );
  MUX2_X1 U15932 ( .A(n13725), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  NAND2_X1 U15933 ( .A1(n13726), .A2(n8018), .ZN(n13727) );
  NAND3_X1 U15934 ( .A1(n13729), .A2(n13728), .A3(n13727), .ZN(n13744) );
  OAI21_X1 U15935 ( .B1(n13934), .B2(n13935), .A(n6556), .ZN(n13730) );
  AOI21_X1 U15936 ( .B1(n13732), .B2(n13731), .A(n13730), .ZN(n13734) );
  OAI22_X1 U15937 ( .A1(n13843), .A2(n13735), .B1(n13734), .B2(n13726), .ZN(
        n13736) );
  NOR2_X1 U15938 ( .A1(n13737), .A2(n13736), .ZN(n13743) );
  INV_X1 U15939 ( .A(n13738), .ZN(n13741) );
  INV_X1 U15940 ( .A(n13739), .ZN(n13740) );
  AND2_X1 U15941 ( .A1(n13932), .A2(n6556), .ZN(n13746) );
  XNOR2_X1 U15942 ( .A(n14130), .B(n13789), .ZN(n13745) );
  NOR2_X1 U15943 ( .A1(n13745), .A2(n13746), .ZN(n13747) );
  AOI21_X1 U15944 ( .B1(n13746), .B2(n13745), .A(n13747), .ZN(n13901) );
  NAND2_X1 U15945 ( .A1(n13902), .A2(n13901), .ZN(n13900) );
  INV_X1 U15946 ( .A(n13747), .ZN(n13748) );
  NAND2_X1 U15947 ( .A1(n13931), .A2(n6556), .ZN(n13784) );
  XNOR2_X1 U15948 ( .A(n13752), .B(n13789), .ZN(n13783) );
  XOR2_X1 U15949 ( .A(n13784), .B(n13783), .Z(n13786) );
  XNOR2_X1 U15950 ( .A(n13787), .B(n13786), .ZN(n13754) );
  AOI22_X1 U15951 ( .A1(n14120), .A2(n13859), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13749) );
  OAI21_X1 U15952 ( .B1(n13750), .B2(n13855), .A(n13749), .ZN(n13751) );
  AOI21_X1 U15953 ( .B1(n13752), .B2(n13923), .A(n13751), .ZN(n13753) );
  OAI21_X1 U15954 ( .B1(n13754), .B2(n13925), .A(n13753), .ZN(P2_U3186) );
  INV_X1 U15955 ( .A(n13755), .ZN(n13756) );
  AOI21_X1 U15956 ( .B1(n13758), .B2(n13757), .A(n13756), .ZN(n13765) );
  NAND2_X1 U15957 ( .A1(n13943), .A2(n13907), .ZN(n13760) );
  NAND2_X1 U15958 ( .A1(n13945), .A2(n13905), .ZN(n13759) );
  NAND2_X1 U15959 ( .A1(n13760), .A2(n13759), .ZN(n14316) );
  AOI21_X1 U15960 ( .B1(n13919), .B2(n14316), .A(n13761), .ZN(n13762) );
  OAI21_X1 U15961 ( .B1(n14322), .B2(n13921), .A(n13762), .ZN(n13763) );
  AOI21_X1 U15962 ( .B1(n14481), .B2(n13923), .A(n13763), .ZN(n13764) );
  OAI21_X1 U15963 ( .B1(n13765), .B2(n13925), .A(n13764), .ZN(P2_U3187) );
  AOI21_X1 U15964 ( .B1(n8018), .B2(n13767), .A(n13766), .ZN(n13774) );
  OR2_X1 U15965 ( .A1(n13768), .A2(n13917), .ZN(n13770) );
  OR2_X1 U15966 ( .A1(n13801), .A2(n13915), .ZN(n13769) );
  NAND2_X1 U15967 ( .A1(n13770), .A2(n13769), .ZN(n14180) );
  OAI22_X1 U15968 ( .A1(n13921), .A2(n14181), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n16033), .ZN(n13772) );
  NOR2_X1 U15969 ( .A1(n14541), .A2(n13912), .ZN(n13771) );
  AOI211_X1 U15970 ( .C1(n13919), .C2(n14180), .A(n13772), .B(n13771), .ZN(
        n13773) );
  OAI21_X1 U15971 ( .B1(n13774), .B2(n13925), .A(n13773), .ZN(P2_U3188) );
  INV_X1 U15972 ( .A(n13775), .ZN(n13776) );
  AOI21_X1 U15973 ( .B1(n13778), .B2(n13777), .A(n13776), .ZN(n13782) );
  NOR2_X1 U15974 ( .A1(n13921), .A2(n14247), .ZN(n13780) );
  AOI22_X1 U15975 ( .A1(n13938), .A2(n13907), .B1(n13940), .B2(n13905), .ZN(
        n14242) );
  NAND2_X1 U15976 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14087)
         );
  OAI21_X1 U15977 ( .B1(n13855), .B2(n14242), .A(n14087), .ZN(n13779) );
  AOI211_X1 U15978 ( .C1(n14456), .C2(n13923), .A(n13780), .B(n13779), .ZN(
        n13781) );
  OAI21_X1 U15979 ( .B1(n13782), .B2(n13925), .A(n13781), .ZN(P2_U3191) );
  INV_X1 U15980 ( .A(n13783), .ZN(n13785) );
  OAI22_X1 U15981 ( .A1(n13787), .A2(n13786), .B1(n13785), .B2(n13784), .ZN(
        n13792) );
  NAND2_X1 U15982 ( .A1(n13930), .A2(n6556), .ZN(n13788) );
  XOR2_X1 U15983 ( .A(n13789), .B(n13788), .Z(n13790) );
  XNOR2_X1 U15984 ( .A(n14111), .B(n13790), .ZN(n13791) );
  XNOR2_X1 U15985 ( .A(n13792), .B(n13791), .ZN(n13799) );
  INV_X1 U15986 ( .A(n13793), .ZN(n14109) );
  AOI22_X1 U15987 ( .A1(n14109), .A2(n13859), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13794) );
  OAI21_X1 U15988 ( .B1(n13795), .B2(n13855), .A(n13794), .ZN(n13796) );
  AOI21_X1 U15989 ( .B1(n13797), .B2(n13923), .A(n13796), .ZN(n13798) );
  OAI21_X1 U15990 ( .B1(n13799), .B2(n13925), .A(n13798), .ZN(P2_U3192) );
  XNOR2_X1 U15991 ( .A(n13800), .B(n13871), .ZN(n13807) );
  OR2_X1 U15992 ( .A1(n13801), .A2(n13917), .ZN(n13803) );
  NAND2_X1 U15993 ( .A1(n13938), .A2(n13905), .ZN(n13802) );
  NAND2_X1 U15994 ( .A1(n13803), .A2(n13802), .ZN(n14206) );
  AOI22_X1 U15995 ( .A1(n14206), .A2(n13919), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13804) );
  OAI21_X1 U15996 ( .B1(n14209), .B2(n13921), .A(n13804), .ZN(n13805) );
  AOI21_X1 U15997 ( .B1(n14214), .B2(n13923), .A(n13805), .ZN(n13806) );
  OAI21_X1 U15998 ( .B1(n13807), .B2(n13925), .A(n13806), .ZN(P2_U3195) );
  NAND2_X1 U15999 ( .A1(n13809), .A2(n13808), .ZN(n13811) );
  XOR2_X1 U16000 ( .A(n13811), .B(n13810), .Z(n13820) );
  OR2_X1 U16001 ( .A1(n13812), .A2(n13915), .ZN(n13814) );
  NAND2_X1 U16002 ( .A1(n13945), .A2(n13907), .ZN(n13813) );
  AND2_X1 U16003 ( .A1(n13814), .A2(n13813), .ZN(n14349) );
  INV_X1 U16004 ( .A(n14351), .ZN(n13815) );
  NAND2_X1 U16005 ( .A1(n13859), .A2(n13815), .ZN(n13817) );
  OAI211_X1 U16006 ( .C1(n14349), .C2(n13855), .A(n13817), .B(n13816), .ZN(
        n13818) );
  AOI21_X1 U16007 ( .B1(n14357), .B2(n13923), .A(n13818), .ZN(n13819) );
  OAI21_X1 U16008 ( .B1(n13820), .B2(n13925), .A(n13819), .ZN(P2_U3196) );
  XNOR2_X1 U16009 ( .A(n13823), .B(n13821), .ZN(n13914) );
  INV_X1 U16010 ( .A(n13821), .ZN(n13822) );
  AOI22_X1 U16011 ( .A1(n13914), .A2(n13913), .B1(n13823), .B2(n13822), .ZN(
        n13827) );
  NAND2_X1 U16012 ( .A1(n13825), .A2(n13824), .ZN(n13826) );
  XNOR2_X1 U16013 ( .A(n13827), .B(n13826), .ZN(n13832) );
  AOI22_X1 U16014 ( .A1(n13941), .A2(n13907), .B1(n13943), .B2(n13905), .ZN(
        n14288) );
  NAND2_X1 U16015 ( .A1(n13859), .A2(n14292), .ZN(n13829) );
  OAI211_X1 U16016 ( .C1(n14288), .C2(n13855), .A(n13829), .B(n13828), .ZN(
        n13830) );
  AOI21_X1 U16017 ( .B1(n14469), .B2(n13923), .A(n13830), .ZN(n13831) );
  OAI21_X1 U16018 ( .B1(n13832), .B2(n13925), .A(n13831), .ZN(P2_U3198) );
  OAI21_X1 U16019 ( .B1(n13835), .B2(n13834), .A(n13833), .ZN(n13836) );
  NAND2_X1 U16020 ( .A1(n13836), .A2(n13903), .ZN(n13841) );
  INV_X1 U16021 ( .A(n13837), .ZN(n14275) );
  AOI22_X1 U16022 ( .A1(n13940), .A2(n13907), .B1(n13905), .B2(n13942), .ZN(
        n14269) );
  OAI21_X1 U16023 ( .B1(n13855), .B2(n14269), .A(n13838), .ZN(n13839) );
  AOI21_X1 U16024 ( .B1(n14275), .B2(n13859), .A(n13839), .ZN(n13840) );
  OAI211_X1 U16025 ( .C1(n14555), .C2(n13912), .A(n13841), .B(n13840), .ZN(
        P2_U3200) );
  OAI211_X1 U16026 ( .C1(n13844), .C2(n13843), .A(n13842), .B(n13903), .ZN(
        n13849) );
  AND2_X1 U16027 ( .A1(n13935), .A2(n13905), .ZN(n13845) );
  AOI21_X1 U16028 ( .B1(n13933), .B2(n13907), .A(n13845), .ZN(n14161) );
  OAI22_X1 U16029 ( .A1(n14161), .A2(n13855), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13846), .ZN(n13847) );
  AOI21_X1 U16030 ( .B1(n14168), .B2(n13859), .A(n13847), .ZN(n13848) );
  OAI211_X1 U16031 ( .C1(n14537), .C2(n13912), .A(n13849), .B(n13848), .ZN(
        P2_U3201) );
  NAND2_X1 U16032 ( .A1(n13851), .A2(n13850), .ZN(n13853) );
  XOR2_X1 U16033 ( .A(n13853), .B(n13852), .Z(n13861) );
  AOI22_X1 U16034 ( .A1(n13937), .A2(n13907), .B1(n13905), .B2(n13939), .ZN(
        n14227) );
  OAI22_X1 U16035 ( .A1(n14227), .A2(n13855), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13854), .ZN(n13858) );
  NOR2_X1 U16036 ( .A1(n13856), .A2(n13912), .ZN(n13857) );
  AOI211_X1 U16037 ( .C1(n13859), .C2(n14232), .A(n13858), .B(n13857), .ZN(
        n13860) );
  OAI21_X1 U16038 ( .B1(n13861), .B2(n13925), .A(n13860), .ZN(P2_U3205) );
  XNOR2_X1 U16039 ( .A(n13863), .B(n13862), .ZN(n13868) );
  OAI22_X1 U16040 ( .A1(n13864), .A2(n13915), .B1(n13916), .B2(n13917), .ZN(
        n14334) );
  AOI22_X1 U16041 ( .A1(n13919), .A2(n14334), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13865) );
  OAI21_X1 U16042 ( .B1(n14340), .B2(n13921), .A(n13865), .ZN(n13866) );
  AOI21_X1 U16043 ( .B1(n14339), .B2(n13923), .A(n13866), .ZN(n13867) );
  OAI21_X1 U16044 ( .B1(n13868), .B2(n13925), .A(n13867), .ZN(P2_U3206) );
  INV_X1 U16045 ( .A(n13869), .ZN(n13870) );
  AOI21_X1 U16046 ( .B1(n13800), .B2(n13871), .A(n13870), .ZN(n13875) );
  XNOR2_X1 U16047 ( .A(n13873), .B(n13872), .ZN(n13874) );
  XNOR2_X1 U16048 ( .A(n13875), .B(n13874), .ZN(n13880) );
  AOI22_X1 U16049 ( .A1(n13935), .A2(n13907), .B1(n13937), .B2(n13905), .ZN(
        n14192) );
  INV_X1 U16050 ( .A(n14192), .ZN(n13876) );
  AOI22_X1 U16051 ( .A1(n13876), .A2(n13919), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13877) );
  OAI21_X1 U16052 ( .B1(n14198), .B2(n13921), .A(n13877), .ZN(n13878) );
  AOI21_X1 U16053 ( .B1(n14194), .B2(n13923), .A(n13878), .ZN(n13879) );
  OAI21_X1 U16054 ( .B1(n13880), .B2(n13925), .A(n13879), .ZN(P2_U3207) );
  XNOR2_X1 U16055 ( .A(n13882), .B(n13881), .ZN(n13889) );
  AND2_X1 U16056 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n14051) );
  AOI21_X1 U16057 ( .B1(n13919), .B2(n13883), .A(n14051), .ZN(n13884) );
  OAI21_X1 U16058 ( .B1(n13885), .B2(n13921), .A(n13884), .ZN(n13886) );
  AOI21_X1 U16059 ( .B1(n13887), .B2(n13923), .A(n13886), .ZN(n13888) );
  OAI21_X1 U16060 ( .B1(n13889), .B2(n13925), .A(n13888), .ZN(P2_U3208) );
  XNOR2_X1 U16061 ( .A(n13891), .B(n13890), .ZN(n13899) );
  INV_X1 U16062 ( .A(n14258), .ZN(n13896) );
  OAI22_X1 U16063 ( .A1(n13893), .A2(n13917), .B1(n13892), .B2(n13915), .ZN(
        n14255) );
  NOR2_X1 U16064 ( .A1(n13894), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14064) );
  AOI21_X1 U16065 ( .B1(n13919), .B2(n14255), .A(n14064), .ZN(n13895) );
  OAI21_X1 U16066 ( .B1(n13896), .B2(n13921), .A(n13895), .ZN(n13897) );
  AOI21_X1 U16067 ( .B1(n14460), .B2(n13923), .A(n13897), .ZN(n13898) );
  OAI21_X1 U16068 ( .B1(n13899), .B2(n13925), .A(n13898), .ZN(P2_U3210) );
  OAI21_X1 U16069 ( .B1(n13902), .B2(n13901), .A(n13900), .ZN(n13904) );
  NAND2_X1 U16070 ( .A1(n13904), .A2(n13903), .ZN(n13911) );
  AND2_X1 U16071 ( .A1(n13933), .A2(n13905), .ZN(n13906) );
  AOI21_X1 U16072 ( .B1(n13931), .B2(n13907), .A(n13906), .ZN(n14137) );
  INV_X1 U16073 ( .A(n14137), .ZN(n13909) );
  OAI22_X1 U16074 ( .A1(n14132), .A2(n13921), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15965), .ZN(n13908) );
  AOI21_X1 U16075 ( .B1(n13909), .B2(n13919), .A(n13908), .ZN(n13910) );
  OAI211_X1 U16076 ( .C1(n14530), .C2(n13912), .A(n13911), .B(n13910), .ZN(
        P2_U3212) );
  XNOR2_X1 U16077 ( .A(n13914), .B(n13913), .ZN(n13926) );
  OAI22_X1 U16078 ( .A1(n13918), .A2(n13917), .B1(n13916), .B2(n13915), .ZN(
        n14300) );
  AOI22_X1 U16079 ( .A1(n13919), .A2(n14300), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13920) );
  OAI21_X1 U16080 ( .B1(n14307), .B2(n13921), .A(n13920), .ZN(n13922) );
  AOI21_X1 U16081 ( .B1(n14306), .B2(n13923), .A(n13922), .ZN(n13924) );
  OAI21_X1 U16082 ( .B1(n13926), .B2(n13925), .A(n13924), .ZN(P2_U3213) );
  MUX2_X1 U16083 ( .A(n13927), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13957), .Z(
        P2_U3562) );
  MUX2_X1 U16084 ( .A(n13928), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13957), .Z(
        P2_U3561) );
  MUX2_X1 U16085 ( .A(n13929), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13957), .Z(
        P2_U3560) );
  MUX2_X1 U16086 ( .A(n13930), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13957), .Z(
        P2_U3559) );
  MUX2_X1 U16087 ( .A(n13931), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13957), .Z(
        P2_U3558) );
  MUX2_X1 U16088 ( .A(n13932), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13957), .Z(
        P2_U3557) );
  MUX2_X1 U16089 ( .A(n13933), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13957), .Z(
        P2_U3556) );
  MUX2_X1 U16090 ( .A(n13934), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13957), .Z(
        P2_U3555) );
  MUX2_X1 U16091 ( .A(n13935), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13957), .Z(
        P2_U3554) );
  MUX2_X1 U16092 ( .A(n13936), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13957), .Z(
        P2_U3553) );
  MUX2_X1 U16093 ( .A(n13937), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13957), .Z(
        P2_U3552) );
  MUX2_X1 U16094 ( .A(n13938), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13957), .Z(
        P2_U3551) );
  MUX2_X1 U16095 ( .A(n13939), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13957), .Z(
        P2_U3550) );
  MUX2_X1 U16096 ( .A(n13940), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13957), .Z(
        P2_U3549) );
  INV_X2 U16097 ( .A(P2_U3947), .ZN(n13957) );
  MUX2_X1 U16098 ( .A(n13941), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13957), .Z(
        P2_U3548) );
  MUX2_X1 U16099 ( .A(n13942), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13957), .Z(
        P2_U3547) );
  MUX2_X1 U16100 ( .A(n13943), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13957), .Z(
        P2_U3546) );
  MUX2_X1 U16101 ( .A(n13944), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13957), .Z(
        P2_U3545) );
  MUX2_X1 U16102 ( .A(n13945), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13957), .Z(
        P2_U3544) );
  MUX2_X1 U16103 ( .A(n13946), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13957), .Z(
        P2_U3543) );
  MUX2_X1 U16104 ( .A(n13947), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13957), .Z(
        P2_U3542) );
  MUX2_X1 U16105 ( .A(n13948), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13957), .Z(
        P2_U3541) );
  MUX2_X1 U16106 ( .A(n13949), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13957), .Z(
        P2_U3540) );
  MUX2_X1 U16107 ( .A(n13950), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13957), .Z(
        P2_U3539) );
  MUX2_X1 U16108 ( .A(n13951), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13957), .Z(
        P2_U3538) );
  MUX2_X1 U16109 ( .A(n13952), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13957), .Z(
        P2_U3537) );
  MUX2_X1 U16110 ( .A(n13953), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13957), .Z(
        P2_U3536) );
  MUX2_X1 U16111 ( .A(n13954), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13957), .Z(
        P2_U3535) );
  MUX2_X1 U16112 ( .A(n13955), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13957), .Z(
        P2_U3534) );
  MUX2_X1 U16113 ( .A(n13956), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13957), .Z(
        P2_U3533) );
  MUX2_X1 U16114 ( .A(n8781), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13957), .Z(
        P2_U3532) );
  MUX2_X1 U16115 ( .A(n8788), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13957), .Z(
        P2_U3531) );
  OAI22_X1 U16116 ( .A1(n15658), .A2(n15469), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13958), .ZN(n13959) );
  AOI21_X1 U16117 ( .B1(n13960), .B2(n15651), .A(n13959), .ZN(n13971) );
  OAI211_X1 U16118 ( .C1(n13963), .C2(n13962), .A(n15644), .B(n13961), .ZN(
        n13970) );
  MUX2_X1 U16119 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10435), .S(n13964), .Z(
        n13966) );
  NAND3_X1 U16120 ( .A1(n15636), .A2(n13966), .A3(n13965), .ZN(n13967) );
  NAND3_X1 U16121 ( .A1(n15653), .A2(n13968), .A3(n13967), .ZN(n13969) );
  NAND3_X1 U16122 ( .A1(n13971), .A2(n13970), .A3(n13969), .ZN(P2_U3216) );
  AND2_X1 U16123 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n13973) );
  NOR2_X1 U16124 ( .A1(n14082), .A2(n13977), .ZN(n13972) );
  AOI211_X1 U16125 ( .C1(n15629), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n13973), .B(
        n13972), .ZN(n13983) );
  OAI211_X1 U16126 ( .C1(n13976), .C2(n13975), .A(n15644), .B(n13974), .ZN(
        n13982) );
  MUX2_X1 U16127 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11629), .S(n13977), .Z(
        n13979) );
  NAND3_X1 U16128 ( .A1(n13979), .A2(n15652), .A3(n13978), .ZN(n13980) );
  NAND3_X1 U16129 ( .A1(n15653), .A2(n13993), .A3(n13980), .ZN(n13981) );
  NAND3_X1 U16130 ( .A1(n13983), .A2(n13982), .A3(n13981), .ZN(P2_U3218) );
  AND2_X1 U16131 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n13986) );
  NOR2_X1 U16132 ( .A1(n15658), .A2(n13984), .ZN(n13985) );
  AOI211_X1 U16133 ( .C1(n15651), .C2(n13990), .A(n13986), .B(n13985), .ZN(
        n13997) );
  OAI211_X1 U16134 ( .C1(n13989), .C2(n13988), .A(n15644), .B(n13987), .ZN(
        n13996) );
  MUX2_X1 U16135 ( .A(n11965), .B(P2_REG2_REG_5__SCAN_IN), .S(n13990), .Z(
        n13991) );
  NAND3_X1 U16136 ( .A1(n13993), .A2(n13992), .A3(n13991), .ZN(n13994) );
  NAND3_X1 U16137 ( .A1(n15653), .A2(n14007), .A3(n13994), .ZN(n13995) );
  NAND3_X1 U16138 ( .A1(n13997), .A2(n13996), .A3(n13995), .ZN(P2_U3219) );
  INV_X1 U16139 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n13999) );
  OAI21_X1 U16140 ( .B1(n15658), .B2(n13999), .A(n13998), .ZN(n14000) );
  AOI21_X1 U16141 ( .B1(n14004), .B2(n15651), .A(n14000), .ZN(n14011) );
  OAI211_X1 U16142 ( .C1(n14003), .C2(n14002), .A(n15644), .B(n14001), .ZN(
        n14010) );
  MUX2_X1 U16143 ( .A(n10444), .B(P2_REG2_REG_6__SCAN_IN), .S(n14004), .Z(
        n14005) );
  NAND3_X1 U16144 ( .A1(n14007), .A2(n14006), .A3(n14005), .ZN(n14008) );
  NAND3_X1 U16145 ( .A1(n15653), .A2(n14017), .A3(n14008), .ZN(n14009) );
  NAND3_X1 U16146 ( .A1(n14011), .A2(n14010), .A3(n14009), .ZN(P2_U3220) );
  OAI211_X1 U16147 ( .C1(n14014), .C2(n14013), .A(n15644), .B(n14012), .ZN(
        n14024) );
  MUX2_X1 U16148 ( .A(n11996), .B(P2_REG2_REG_7__SCAN_IN), .S(n14020), .Z(
        n14015) );
  NAND3_X1 U16149 ( .A1(n14017), .A2(n14016), .A3(n14015), .ZN(n14018) );
  NAND3_X1 U16150 ( .A1(n15653), .A2(n14036), .A3(n14018), .ZN(n14023) );
  AOI21_X1 U16151 ( .B1(n15629), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n14019), .ZN(
        n14022) );
  NAND2_X1 U16152 ( .A1(n15651), .A2(n14020), .ZN(n14021) );
  NAND4_X1 U16153 ( .A1(n14024), .A2(n14023), .A3(n14022), .A4(n14021), .ZN(
        P2_U3221) );
  INV_X1 U16154 ( .A(n14025), .ZN(n14028) );
  NOR2_X1 U16155 ( .A1(n15658), .A2(n14026), .ZN(n14027) );
  AOI211_X1 U16156 ( .C1(n15651), .C2(n14029), .A(n14028), .B(n14027), .ZN(
        n14041) );
  OAI211_X1 U16157 ( .C1(n14032), .C2(n14031), .A(n14030), .B(n15644), .ZN(
        n14040) );
  MUX2_X1 U16158 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11693), .S(n14033), .Z(
        n14034) );
  NAND3_X1 U16159 ( .A1(n14036), .A2(n14035), .A3(n14034), .ZN(n14037) );
  NAND3_X1 U16160 ( .A1(n15653), .A2(n14038), .A3(n14037), .ZN(n14039) );
  NAND3_X1 U16161 ( .A1(n14041), .A2(n14040), .A3(n14039), .ZN(P2_U3222) );
  OAI211_X1 U16162 ( .C1(n14044), .C2(n14043), .A(n14042), .B(n15644), .ZN(
        n14055) );
  OAI21_X1 U16163 ( .B1(n14047), .B2(n14046), .A(n14045), .ZN(n14048) );
  NAND2_X1 U16164 ( .A1(n14048), .A2(n15653), .ZN(n14054) );
  NOR2_X1 U16165 ( .A1(n15658), .A2(n14049), .ZN(n14050) );
  AOI211_X1 U16166 ( .C1(n15651), .C2(n14052), .A(n14051), .B(n14050), .ZN(
        n14053) );
  NAND3_X1 U16167 ( .A1(n14055), .A2(n14054), .A3(n14053), .ZN(P2_U3225) );
  NAND2_X1 U16168 ( .A1(n14065), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n14056) );
  NAND2_X1 U16169 ( .A1(n14057), .A2(n14056), .ZN(n14058) );
  OR2_X1 U16170 ( .A1(n14058), .A2(n14067), .ZN(n14076) );
  NAND2_X1 U16171 ( .A1(n14058), .A2(n14067), .ZN(n14059) );
  NAND2_X1 U16172 ( .A1(n14076), .A2(n14059), .ZN(n14061) );
  INV_X1 U16173 ( .A(n14077), .ZN(n14060) );
  AOI21_X1 U16174 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n14061), .A(n14060), 
        .ZN(n14075) );
  NOR2_X1 U16175 ( .A1(n14082), .A2(n14062), .ZN(n14063) );
  AOI211_X1 U16176 ( .C1(n15629), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n14064), 
        .B(n14063), .ZN(n14074) );
  NAND2_X1 U16177 ( .A1(n14068), .A2(n14067), .ZN(n14079) );
  OR2_X1 U16178 ( .A1(n14068), .A2(n14067), .ZN(n14069) );
  NAND2_X1 U16179 ( .A1(n14079), .A2(n14069), .ZN(n14071) );
  INV_X1 U16180 ( .A(n14071), .ZN(n14072) );
  INV_X1 U16181 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14070) );
  OAI211_X1 U16182 ( .C1(n14072), .C2(P2_REG1_REG_18__SCAN_IN), .A(n15644), 
        .B(n14080), .ZN(n14073) );
  OAI211_X1 U16183 ( .C1(n14075), .C2(n15623), .A(n14074), .B(n14073), .ZN(
        P2_U3232) );
  NAND2_X1 U16184 ( .A1(n14077), .A2(n14076), .ZN(n14078) );
  XNOR2_X1 U16185 ( .A(n14078), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n14085) );
  NAND2_X1 U16186 ( .A1(n14080), .A2(n14079), .ZN(n14081) );
  XNOR2_X1 U16187 ( .A(n14081), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n14083) );
  INV_X1 U16188 ( .A(n14083), .ZN(n14084) );
  NAND2_X1 U16189 ( .A1(n14088), .A2(n14401), .ZN(n14091) );
  INV_X1 U16190 ( .A(n14089), .ZN(n14409) );
  NOR2_X1 U16191 ( .A1(n6557), .A2(n14409), .ZN(n14096) );
  AOI21_X1 U16192 ( .B1(P2_REG2_REG_31__SCAN_IN), .B2(n6557), .A(n14096), .ZN(
        n14090) );
  OAI211_X1 U16193 ( .C1(n14408), .C2(n14399), .A(n14091), .B(n14090), .ZN(
        P2_U3234) );
  OAI211_X1 U16194 ( .C1(n14093), .C2(n14526), .A(n14470), .B(n14092), .ZN(
        n14410) );
  NOR2_X1 U16195 ( .A1(n14285), .A2(n14094), .ZN(n14095) );
  AOI211_X1 U16196 ( .C1(n14097), .C2(n14368), .A(n14096), .B(n14095), .ZN(
        n14098) );
  OAI21_X1 U16197 ( .B1(n14410), .B2(n14370), .A(n14098), .ZN(P2_U3235) );
  INV_X1 U16198 ( .A(n14099), .ZN(n14107) );
  NAND2_X1 U16199 ( .A1(n14100), .A2(n14401), .ZN(n14103) );
  AOI22_X1 U16200 ( .A1(n14101), .A2(n15666), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n6557), .ZN(n14102) );
  OAI211_X1 U16201 ( .C1(n7520), .C2(n14399), .A(n14103), .B(n14102), .ZN(
        n14104) );
  AOI21_X1 U16202 ( .B1(n14105), .B2(n14285), .A(n14104), .ZN(n14106) );
  OAI21_X1 U16203 ( .B1(n14107), .B2(n14361), .A(n14106), .ZN(P2_U3236) );
  AOI21_X1 U16204 ( .B1(n14109), .B2(n15666), .A(n14108), .ZN(n14117) );
  INV_X1 U16205 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n14110) );
  OAI22_X1 U16206 ( .A1(n14111), .A2(n14399), .B1(n14110), .B2(n14285), .ZN(
        n14112) );
  AOI21_X1 U16207 ( .B1(n14113), .B2(n14401), .A(n14112), .ZN(n14116) );
  NAND2_X1 U16208 ( .A1(n14114), .A2(n14312), .ZN(n14115) );
  OAI211_X1 U16209 ( .C1(n14117), .C2(n6557), .A(n14116), .B(n14115), .ZN(
        P2_U3237) );
  INV_X1 U16210 ( .A(n14118), .ZN(n14126) );
  NAND2_X1 U16211 ( .A1(n14119), .A2(n14401), .ZN(n14122) );
  AOI22_X1 U16212 ( .A1(n14120), .A2(n15666), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n6557), .ZN(n14121) );
  OAI211_X1 U16213 ( .C1(n14414), .C2(n14399), .A(n14122), .B(n14121), .ZN(
        n14123) );
  AOI21_X1 U16214 ( .B1(n14124), .B2(n14285), .A(n14123), .ZN(n14125) );
  OAI21_X1 U16215 ( .B1(n14126), .B2(n14361), .A(n14125), .ZN(P2_U3238) );
  XOR2_X1 U16216 ( .A(n14127), .B(n14136), .Z(n14417) );
  INV_X1 U16217 ( .A(n14417), .ZN(n14140) );
  INV_X1 U16218 ( .A(n14149), .ZN(n14129) );
  AOI211_X1 U16219 ( .C1(n14130), .C2(n14129), .A(n14338), .B(n14128), .ZN(
        n14416) );
  NOR2_X1 U16220 ( .A1(n14530), .A2(n14399), .ZN(n14134) );
  OAI22_X1 U16221 ( .A1(n14132), .A2(n14398), .B1(n14131), .B2(n14285), .ZN(
        n14133) );
  AOI211_X1 U16222 ( .C1(n14416), .C2(n14401), .A(n14134), .B(n14133), .ZN(
        n14139) );
  NAND2_X1 U16223 ( .A1(n14415), .A2(n14285), .ZN(n14138) );
  OAI211_X1 U16224 ( .C1(n14140), .C2(n14361), .A(n14139), .B(n14138), .ZN(
        P2_U3239) );
  XNOR2_X1 U16225 ( .A(n14141), .B(n14142), .ZN(n14422) );
  INV_X1 U16226 ( .A(n14422), .ZN(n14155) );
  XNOR2_X1 U16227 ( .A(n14143), .B(n14142), .ZN(n14145) );
  OAI21_X1 U16228 ( .B1(n14145), .B2(n14375), .A(n14144), .ZN(n14420) );
  NAND2_X1 U16229 ( .A1(n14166), .A2(n14146), .ZN(n14147) );
  NAND2_X1 U16230 ( .A1(n14147), .A2(n14470), .ZN(n14148) );
  NOR2_X1 U16231 ( .A1(n14149), .A2(n14148), .ZN(n14421) );
  NAND2_X1 U16232 ( .A1(n14421), .A2(n14401), .ZN(n14152) );
  AOI22_X1 U16233 ( .A1(n14150), .A2(n15666), .B1(n6557), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n14151) );
  OAI211_X1 U16234 ( .C1(n14534), .C2(n14399), .A(n14152), .B(n14151), .ZN(
        n14153) );
  AOI21_X1 U16235 ( .B1(n14420), .B2(n14285), .A(n14153), .ZN(n14154) );
  OAI21_X1 U16236 ( .B1(n14155), .B2(n14361), .A(n14154), .ZN(P2_U3240) );
  NAND2_X1 U16237 ( .A1(n14190), .A2(n14157), .ZN(n14176) );
  NAND2_X1 U16238 ( .A1(n14178), .A2(n14158), .ZN(n14160) );
  XNOR2_X1 U16239 ( .A(n14160), .B(n14159), .ZN(n14162) );
  INV_X1 U16240 ( .A(n14425), .ZN(n14173) );
  AOI211_X1 U16241 ( .C1(n14167), .C2(n6587), .A(n14338), .B(n6829), .ZN(
        n14426) );
  NAND2_X1 U16242 ( .A1(n14426), .A2(n14401), .ZN(n14170) );
  AOI22_X1 U16243 ( .A1(n6557), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n14168), 
        .B2(n15666), .ZN(n14169) );
  OAI211_X1 U16244 ( .C1(n14537), .C2(n14399), .A(n14170), .B(n14169), .ZN(
        n14171) );
  AOI21_X1 U16245 ( .B1(n14427), .B2(n14312), .A(n14171), .ZN(n14172) );
  OAI21_X1 U16246 ( .B1(n14173), .B2(n6557), .A(n14172), .ZN(P2_U3241) );
  XNOR2_X1 U16247 ( .A(n14174), .B(n14175), .ZN(n14434) );
  NAND2_X1 U16248 ( .A1(n14176), .A2(n14175), .ZN(n14177) );
  NAND2_X1 U16249 ( .A1(n14178), .A2(n14177), .ZN(n14179) );
  NAND2_X1 U16250 ( .A1(n14179), .A2(n15662), .ZN(n14433) );
  INV_X1 U16251 ( .A(n14180), .ZN(n14430) );
  OAI211_X1 U16252 ( .C1(n14398), .C2(n14181), .A(n14433), .B(n14430), .ZN(
        n14185) );
  OAI211_X1 U16253 ( .C1(n14197), .C2(n14541), .A(n14470), .B(n6587), .ZN(
        n14431) );
  AOI22_X1 U16254 ( .A1(n14182), .A2(n14368), .B1(n6557), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n14183) );
  OAI21_X1 U16255 ( .B1(n14431), .B2(n14370), .A(n14183), .ZN(n14184) );
  AOI21_X1 U16256 ( .B1(n14185), .B2(n14285), .A(n14184), .ZN(n14186) );
  OAI21_X1 U16257 ( .B1(n14434), .B2(n14361), .A(n14186), .ZN(P2_U3242) );
  NAND2_X1 U16258 ( .A1(n14187), .A2(n14191), .ZN(n14188) );
  NAND2_X1 U16259 ( .A1(n14189), .A2(n14188), .ZN(n14437) );
  OAI211_X1 U16260 ( .C1(n14156), .C2(n14191), .A(n14190), .B(n15662), .ZN(
        n14193) );
  NAND2_X1 U16261 ( .A1(n14193), .A2(n14192), .ZN(n14440) );
  NAND2_X1 U16262 ( .A1(n14440), .A2(n14285), .ZN(n14203) );
  NAND2_X1 U16263 ( .A1(n14216), .A2(n14194), .ZN(n14195) );
  NAND2_X1 U16264 ( .A1(n14195), .A2(n14470), .ZN(n14196) );
  NOR2_X1 U16265 ( .A1(n14197), .A2(n14196), .ZN(n14438) );
  INV_X1 U16266 ( .A(n14198), .ZN(n14199) );
  AOI22_X1 U16267 ( .A1(n6557), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n14199), 
        .B2(n15666), .ZN(n14200) );
  OAI21_X1 U16268 ( .B1(n14545), .B2(n14399), .A(n14200), .ZN(n14201) );
  AOI21_X1 U16269 ( .B1(n14438), .B2(n14401), .A(n14201), .ZN(n14202) );
  OAI211_X1 U16270 ( .C1(n14437), .C2(n14361), .A(n14203), .B(n14202), .ZN(
        P2_U3243) );
  XNOR2_X1 U16271 ( .A(n14204), .B(n14213), .ZN(n14205) );
  NAND2_X1 U16272 ( .A1(n14205), .A2(n15662), .ZN(n14208) );
  INV_X1 U16273 ( .A(n14206), .ZN(n14207) );
  NAND2_X1 U16274 ( .A1(n14208), .A2(n14207), .ZN(n14444) );
  NAND2_X1 U16275 ( .A1(n14444), .A2(n14285), .ZN(n14220) );
  INV_X1 U16276 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n14210) );
  OAI22_X1 U16277 ( .A1(n14285), .A2(n14210), .B1(n14209), .B2(n14398), .ZN(
        n14211) );
  AOI21_X1 U16278 ( .B1(n14214), .B2(n14368), .A(n14211), .ZN(n14219) );
  XNOR2_X1 U16279 ( .A(n14212), .B(n14213), .ZN(n14443) );
  NAND2_X1 U16280 ( .A1(n14443), .A2(n14312), .ZN(n14218) );
  AOI21_X1 U16281 ( .B1(n14230), .B2(n14214), .A(n14338), .ZN(n14215) );
  AND2_X1 U16282 ( .A1(n14216), .A2(n14215), .ZN(n14445) );
  NAND2_X1 U16283 ( .A1(n14445), .A2(n14401), .ZN(n14217) );
  NAND4_X1 U16284 ( .A1(n14220), .A2(n14219), .A3(n14218), .A4(n14217), .ZN(
        P2_U3244) );
  XNOR2_X1 U16285 ( .A(n14221), .B(n14222), .ZN(n14453) );
  INV_X1 U16286 ( .A(n14223), .ZN(n14224) );
  AOI21_X1 U16287 ( .B1(n14226), .B2(n14225), .A(n14224), .ZN(n14228) );
  OAI21_X1 U16288 ( .B1(n14228), .B2(n14375), .A(n14227), .ZN(n14449) );
  NAND2_X1 U16289 ( .A1(n14449), .A2(n14285), .ZN(n14238) );
  AOI21_X1 U16290 ( .B1(n14229), .B2(n14451), .A(n14338), .ZN(n14231) );
  AND2_X1 U16291 ( .A1(n14231), .A2(n14230), .ZN(n14450) );
  INV_X1 U16292 ( .A(n14232), .ZN(n14235) );
  NAND2_X1 U16293 ( .A1(n14451), .A2(n14368), .ZN(n14234) );
  NAND2_X1 U16294 ( .A1(n6557), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n14233) );
  OAI211_X1 U16295 ( .C1(n14398), .C2(n14235), .A(n14234), .B(n14233), .ZN(
        n14236) );
  AOI21_X1 U16296 ( .B1(n14450), .B2(n14401), .A(n14236), .ZN(n14237) );
  OAI211_X1 U16297 ( .C1(n14453), .C2(n14361), .A(n14238), .B(n14237), .ZN(
        P2_U3245) );
  XNOR2_X1 U16298 ( .A(n14239), .B(n14240), .ZN(n14458) );
  XOR2_X1 U16299 ( .A(n14241), .B(n14240), .Z(n14243) );
  OAI21_X1 U16300 ( .B1(n14243), .B2(n14375), .A(n14242), .ZN(n14454) );
  INV_X1 U16301 ( .A(n14244), .ZN(n14246) );
  INV_X1 U16302 ( .A(n14229), .ZN(n14245) );
  AOI211_X1 U16303 ( .C1(n14456), .C2(n14246), .A(n14338), .B(n14245), .ZN(
        n14455) );
  NAND2_X1 U16304 ( .A1(n14455), .A2(n14401), .ZN(n14250) );
  INV_X1 U16305 ( .A(n14247), .ZN(n14248) );
  AOI22_X1 U16306 ( .A1(n6557), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14248), 
        .B2(n15666), .ZN(n14249) );
  OAI211_X1 U16307 ( .C1(n14251), .C2(n14399), .A(n14250), .B(n14249), .ZN(
        n14252) );
  AOI21_X1 U16308 ( .B1(n14454), .B2(n14285), .A(n14252), .ZN(n14253) );
  OAI21_X1 U16309 ( .B1(n14361), .B2(n14458), .A(n14253), .ZN(P2_U3246) );
  XOR2_X1 U16310 ( .A(n14254), .B(n14264), .Z(n14256) );
  AOI21_X1 U16311 ( .B1(n14256), .B2(n15662), .A(n14255), .ZN(n14462) );
  INV_X1 U16312 ( .A(n14273), .ZN(n14257) );
  AOI211_X1 U16313 ( .C1(n14460), .C2(n14257), .A(n14338), .B(n14244), .ZN(
        n14459) );
  AOI22_X1 U16314 ( .A1(n6557), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14258), 
        .B2(n15666), .ZN(n14259) );
  OAI21_X1 U16315 ( .B1(n14260), .B2(n14399), .A(n14259), .ZN(n14266) );
  INV_X1 U16316 ( .A(n14261), .ZN(n14262) );
  AOI21_X1 U16317 ( .B1(n14264), .B2(n14263), .A(n14262), .ZN(n14463) );
  NOR2_X1 U16318 ( .A1(n14463), .A2(n14361), .ZN(n14265) );
  AOI211_X1 U16319 ( .C1(n14459), .C2(n14401), .A(n14266), .B(n14265), .ZN(
        n14267) );
  OAI21_X1 U16320 ( .B1(n6557), .B2(n14462), .A(n14267), .ZN(P2_U3247) );
  XNOR2_X1 U16321 ( .A(n14268), .B(n14272), .ZN(n14270) );
  OAI21_X1 U16322 ( .B1(n14270), .B2(n14375), .A(n14269), .ZN(n14464) );
  INV_X1 U16323 ( .A(n14464), .ZN(n14280) );
  XOR2_X1 U16324 ( .A(n14271), .B(n14272), .Z(n14466) );
  AOI211_X1 U16325 ( .C1(n14274), .C2(n7515), .A(n14338), .B(n14273), .ZN(
        n14465) );
  NAND2_X1 U16326 ( .A1(n14465), .A2(n14401), .ZN(n14277) );
  AOI22_X1 U16327 ( .A1(n6557), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n14275), 
        .B2(n15666), .ZN(n14276) );
  OAI211_X1 U16328 ( .C1(n14555), .C2(n14399), .A(n14277), .B(n14276), .ZN(
        n14278) );
  AOI21_X1 U16329 ( .B1(n14466), .B2(n14312), .A(n14278), .ZN(n14279) );
  OAI21_X1 U16330 ( .B1(n14280), .B2(n6557), .A(n14279), .ZN(P2_U3248) );
  OAI21_X1 U16331 ( .B1(n14303), .B2(n7154), .A(n14282), .ZN(n14283) );
  XNOR2_X1 U16332 ( .A(n14283), .B(n14287), .ZN(n14474) );
  NOR2_X1 U16333 ( .A1(n14285), .A2(n14284), .ZN(n14296) );
  XOR2_X1 U16334 ( .A(n14287), .B(n14286), .Z(n14290) );
  INV_X1 U16335 ( .A(n14288), .ZN(n14289) );
  AOI21_X1 U16336 ( .B1(n14290), .B2(n15662), .A(n14289), .ZN(n14473) );
  AOI21_X1 U16337 ( .B1(n14469), .B2(n14304), .A(n14291), .ZN(n14471) );
  AOI22_X1 U16338 ( .A1(n14471), .A2(n14293), .B1(n14292), .B2(n15666), .ZN(
        n14294) );
  AOI21_X1 U16339 ( .B1(n14473), .B2(n14294), .A(n6557), .ZN(n14295) );
  AOI211_X1 U16340 ( .C1(n14368), .C2(n14469), .A(n14296), .B(n14295), .ZN(
        n14297) );
  OAI21_X1 U16341 ( .B1(n14361), .B2(n14474), .A(n14297), .ZN(P2_U3249) );
  XNOR2_X1 U16342 ( .A(n14299), .B(n14298), .ZN(n14302) );
  INV_X1 U16343 ( .A(n14300), .ZN(n14301) );
  OAI21_X1 U16344 ( .B1(n14302), .B2(n14375), .A(n14301), .ZN(n14475) );
  INV_X1 U16345 ( .A(n14475), .ZN(n14314) );
  XNOR2_X1 U16346 ( .A(n14303), .B(n7154), .ZN(n14477) );
  INV_X1 U16347 ( .A(n14306), .ZN(n14560) );
  INV_X1 U16348 ( .A(n14304), .ZN(n14305) );
  AOI211_X1 U16349 ( .C1(n14306), .C2(n14319), .A(n14338), .B(n14305), .ZN(
        n14476) );
  NAND2_X1 U16350 ( .A1(n14476), .A2(n14401), .ZN(n14310) );
  INV_X1 U16351 ( .A(n14307), .ZN(n14308) );
  AOI22_X1 U16352 ( .A1(n6557), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n14308), 
        .B2(n15666), .ZN(n14309) );
  OAI211_X1 U16353 ( .C1(n14560), .C2(n14399), .A(n14310), .B(n14309), .ZN(
        n14311) );
  AOI21_X1 U16354 ( .B1(n14312), .B2(n14477), .A(n14311), .ZN(n14313) );
  OAI21_X1 U16355 ( .B1(n14314), .B2(n6557), .A(n14313), .ZN(P2_U3250) );
  XNOR2_X1 U16356 ( .A(n14315), .B(n14326), .ZN(n14317) );
  AOI21_X1 U16357 ( .B1(n14317), .B2(n15662), .A(n14316), .ZN(n14483) );
  INV_X1 U16358 ( .A(n14318), .ZN(n14321) );
  INV_X1 U16359 ( .A(n14319), .ZN(n14320) );
  AOI211_X1 U16360 ( .C1(n14481), .C2(n14321), .A(n14338), .B(n14320), .ZN(
        n14480) );
  INV_X1 U16361 ( .A(n14322), .ZN(n14323) );
  AOI22_X1 U16362 ( .A1(n6557), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n14323), 
        .B2(n15666), .ZN(n14324) );
  OAI21_X1 U16363 ( .B1(n14325), .B2(n14399), .A(n14324), .ZN(n14329) );
  XOR2_X1 U16364 ( .A(n14327), .B(n14326), .Z(n14485) );
  NOR2_X1 U16365 ( .A1(n14485), .A2(n14361), .ZN(n14328) );
  AOI211_X1 U16366 ( .C1(n14480), .C2(n14401), .A(n14329), .B(n14328), .ZN(
        n14330) );
  OAI21_X1 U16367 ( .B1(n6557), .B2(n14483), .A(n14330), .ZN(P2_U3251) );
  XNOR2_X1 U16368 ( .A(n14331), .B(n14332), .ZN(n14488) );
  INV_X1 U16369 ( .A(n14488), .ZN(n14345) );
  XOR2_X1 U16370 ( .A(n14333), .B(n14332), .Z(n14336) );
  INV_X1 U16371 ( .A(n14334), .ZN(n14335) );
  OAI21_X1 U16372 ( .B1(n14336), .B2(n14375), .A(n14335), .ZN(n14486) );
  NAND2_X1 U16373 ( .A1(n14486), .A2(n14285), .ZN(n14344) );
  INV_X1 U16374 ( .A(n14337), .ZN(n14353) );
  AOI211_X1 U16375 ( .C1(n14339), .C2(n14353), .A(n14338), .B(n14318), .ZN(
        n14487) );
  NOR2_X1 U16376 ( .A1(n14564), .A2(n14399), .ZN(n14342) );
  OAI22_X1 U16377 ( .A1(n14285), .A2(n10835), .B1(n14340), .B2(n14398), .ZN(
        n14341) );
  AOI211_X1 U16378 ( .C1(n14487), .C2(n14401), .A(n14342), .B(n14341), .ZN(
        n14343) );
  OAI211_X1 U16379 ( .C1(n14345), .C2(n14361), .A(n14344), .B(n14343), .ZN(
        P2_U3252) );
  XOR2_X1 U16380 ( .A(n14346), .B(n14348), .Z(n14495) );
  INV_X1 U16381 ( .A(n14495), .ZN(n14360) );
  XOR2_X1 U16382 ( .A(n14347), .B(n14348), .Z(n14350) );
  OAI21_X1 U16383 ( .B1(n14350), .B2(n14375), .A(n14349), .ZN(n14493) );
  NAND2_X1 U16384 ( .A1(n14493), .A2(n14285), .ZN(n14359) );
  OAI22_X1 U16385 ( .A1(n14285), .A2(n14352), .B1(n14351), .B2(n14398), .ZN(
        n14356) );
  INV_X1 U16386 ( .A(n14357), .ZN(n14492) );
  OAI211_X1 U16387 ( .C1(n14492), .C2(n14354), .A(n14353), .B(n14470), .ZN(
        n14491) );
  NOR2_X1 U16388 ( .A1(n14491), .A2(n14370), .ZN(n14355) );
  AOI211_X1 U16389 ( .C1(n14368), .C2(n14357), .A(n14356), .B(n14355), .ZN(
        n14358) );
  OAI211_X1 U16390 ( .C1(n14361), .C2(n14360), .A(n14359), .B(n14358), .ZN(
        P2_U3253) );
  XNOR2_X1 U16391 ( .A(n14362), .B(n14363), .ZN(n14507) );
  OAI211_X1 U16392 ( .C1(n14364), .C2(n14504), .A(n14470), .B(n11735), .ZN(
        n14503) );
  INV_X1 U16393 ( .A(n14365), .ZN(n14366) );
  AOI22_X1 U16394 ( .A1(n14368), .A2(n14367), .B1(n14366), .B2(n15666), .ZN(
        n14369) );
  OAI21_X1 U16395 ( .B1(n14503), .B2(n14370), .A(n14369), .ZN(n14381) );
  NAND2_X1 U16396 ( .A1(n14372), .A2(n14371), .ZN(n14390) );
  NAND2_X1 U16397 ( .A1(n14390), .A2(n14391), .ZN(n14389) );
  NAND3_X1 U16398 ( .A1(n14389), .A2(n14374), .A3(n14373), .ZN(n14376) );
  AOI21_X1 U16399 ( .B1(n14376), .B2(n11729), .A(n14375), .ZN(n14379) );
  AND2_X1 U16400 ( .A1(n14507), .A2(n15713), .ZN(n14378) );
  OR3_X1 U16401 ( .A1(n14379), .A2(n14378), .A3(n14377), .ZN(n14505) );
  MUX2_X1 U16402 ( .A(n14505), .B(P2_REG2_REG_10__SCAN_IN), .S(n6557), .Z(
        n14380) );
  AOI211_X1 U16403 ( .C1(n14507), .C2(n15667), .A(n14381), .B(n14380), .ZN(
        n14382) );
  INV_X1 U16404 ( .A(n14382), .ZN(P2_U3255) );
  INV_X1 U16405 ( .A(n14383), .ZN(n14386) );
  OAI21_X1 U16406 ( .B1(n14386), .B2(n14385), .A(n14384), .ZN(n14388) );
  XNOR2_X1 U16407 ( .A(n14387), .B(n14388), .ZN(n14511) );
  OAI21_X1 U16408 ( .B1(n14391), .B2(n14390), .A(n14389), .ZN(n14394) );
  NOR2_X1 U16409 ( .A1(n14511), .A2(n15715), .ZN(n14392) );
  AOI211_X1 U16410 ( .C1(n15662), .C2(n14394), .A(n14393), .B(n14392), .ZN(
        n14510) );
  MUX2_X1 U16411 ( .A(n10483), .B(n14510), .S(n14285), .Z(n14404) );
  INV_X1 U16412 ( .A(n14364), .ZN(n14395) );
  OAI211_X1 U16413 ( .C1(n14513), .C2(n14396), .A(n14395), .B(n14470), .ZN(
        n14509) );
  INV_X1 U16414 ( .A(n14509), .ZN(n14402) );
  OAI22_X1 U16415 ( .A1(n14399), .A2(n14513), .B1(n14398), .B2(n14397), .ZN(
        n14400) );
  AOI21_X1 U16416 ( .B1(n14402), .B2(n14401), .A(n14400), .ZN(n14403) );
  OAI211_X1 U16417 ( .C1(n14511), .C2(n14405), .A(n14404), .B(n14403), .ZN(
        P2_U3256) );
  OAI21_X1 U16418 ( .B1(n14408), .B2(n14514), .A(n14407), .ZN(P2_U3530) );
  AND2_X1 U16419 ( .A1(n14410), .A2(n14409), .ZN(n14523) );
  MUX2_X1 U16420 ( .A(n14411), .B(n14523), .S(n15750), .Z(n14412) );
  OAI21_X1 U16421 ( .B1(n14526), .B2(n14514), .A(n14412), .ZN(P2_U3529) );
  INV_X1 U16422 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n14418) );
  MUX2_X1 U16423 ( .A(n14418), .B(n14527), .S(n15750), .Z(n14419) );
  OAI21_X1 U16424 ( .B1(n14530), .B2(n14514), .A(n14419), .ZN(P2_U3525) );
  AOI211_X1 U16425 ( .C1(n15740), .C2(n14422), .A(n14421), .B(n14420), .ZN(
        n14531) );
  MUX2_X1 U16426 ( .A(n14423), .B(n14531), .S(n15750), .Z(n14424) );
  OAI21_X1 U16427 ( .B1(n14534), .B2(n14514), .A(n14424), .ZN(P2_U3524) );
  INV_X1 U16428 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n14428) );
  OAI21_X1 U16429 ( .B1(n14537), .B2(n14514), .A(n14429), .ZN(P2_U3523) );
  AND2_X1 U16430 ( .A1(n14431), .A2(n14430), .ZN(n14432) );
  OAI211_X1 U16431 ( .C1(n14484), .C2(n14434), .A(n14433), .B(n14432), .ZN(
        n14538) );
  MUX2_X1 U16432 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14538), .S(n15750), .Z(
        n14435) );
  INV_X1 U16433 ( .A(n14435), .ZN(n14436) );
  OAI21_X1 U16434 ( .B1(n14541), .B2(n14514), .A(n14436), .ZN(P2_U3522) );
  NOR2_X1 U16435 ( .A1(n14437), .A2(n14484), .ZN(n14439) );
  NOR3_X1 U16436 ( .A1(n14440), .A2(n14439), .A3(n14438), .ZN(n14542) );
  MUX2_X1 U16437 ( .A(n14542), .B(n14441), .S(n12591), .Z(n14442) );
  OAI21_X1 U16438 ( .B1(n14545), .B2(n14514), .A(n14442), .ZN(P2_U3521) );
  AND2_X1 U16439 ( .A1(n14443), .A2(n15740), .ZN(n14446) );
  MUX2_X1 U16440 ( .A(n14447), .B(n8033), .S(n15750), .Z(n14448) );
  OAI21_X1 U16441 ( .B1(n14548), .B2(n14514), .A(n14448), .ZN(P2_U3520) );
  AOI211_X1 U16442 ( .C1(n14451), .C2(n14518), .A(n14450), .B(n14449), .ZN(
        n14452) );
  OAI21_X1 U16443 ( .B1(n14484), .B2(n14453), .A(n14452), .ZN(n14549) );
  MUX2_X1 U16444 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14549), .S(n15750), .Z(
        P2_U3519) );
  AOI211_X1 U16445 ( .C1(n14456), .C2(n14518), .A(n14455), .B(n14454), .ZN(
        n14457) );
  OAI21_X1 U16446 ( .B1(n14484), .B2(n14458), .A(n14457), .ZN(n14550) );
  MUX2_X1 U16447 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14550), .S(n15750), .Z(
        P2_U3518) );
  AOI21_X1 U16448 ( .B1(n14460), .B2(n14518), .A(n14459), .ZN(n14461) );
  OAI211_X1 U16449 ( .C1(n14484), .C2(n14463), .A(n14462), .B(n14461), .ZN(
        n14551) );
  MUX2_X1 U16450 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14551), .S(n15750), .Z(
        P2_U3517) );
  AOI211_X1 U16451 ( .C1(n15740), .C2(n14466), .A(n14465), .B(n14464), .ZN(
        n14552) );
  MUX2_X1 U16452 ( .A(n14467), .B(n14552), .S(n15750), .Z(n14468) );
  OAI21_X1 U16453 ( .B1(n14555), .B2(n14514), .A(n14468), .ZN(P2_U3516) );
  AOI22_X1 U16454 ( .A1(n14471), .A2(n14470), .B1(n14469), .B2(n14518), .ZN(
        n14472) );
  OAI211_X1 U16455 ( .C1(n14484), .C2(n14474), .A(n14473), .B(n14472), .ZN(
        n14556) );
  MUX2_X1 U16456 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14556), .S(n15750), .Z(
        P2_U3515) );
  AOI211_X1 U16457 ( .C1(n15740), .C2(n14477), .A(n14476), .B(n14475), .ZN(
        n14557) );
  MUX2_X1 U16458 ( .A(n14478), .B(n14557), .S(n15750), .Z(n14479) );
  OAI21_X1 U16459 ( .B1(n14560), .B2(n14514), .A(n14479), .ZN(P2_U3514) );
  AOI21_X1 U16460 ( .B1(n14481), .B2(n14518), .A(n14480), .ZN(n14482) );
  OAI211_X1 U16461 ( .C1(n14485), .C2(n14484), .A(n14483), .B(n14482), .ZN(
        n14561) );
  MUX2_X1 U16462 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14561), .S(n15750), .Z(
        P2_U3513) );
  AOI211_X1 U16463 ( .C1(n15740), .C2(n14488), .A(n14487), .B(n14486), .ZN(
        n14562) );
  MUX2_X1 U16464 ( .A(n14489), .B(n14562), .S(n15750), .Z(n14490) );
  OAI21_X1 U16465 ( .B1(n14564), .B2(n14514), .A(n14490), .ZN(P2_U3512) );
  INV_X1 U16466 ( .A(n14518), .ZN(n15737) );
  OAI21_X1 U16467 ( .B1(n14492), .B2(n15737), .A(n14491), .ZN(n14494) );
  AOI211_X1 U16468 ( .C1(n14495), .C2(n15740), .A(n14494), .B(n14493), .ZN(
        n14566) );
  NAND2_X1 U16469 ( .A1(n12591), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n14496) );
  OAI21_X1 U16470 ( .B1(n14566), .B2(n12591), .A(n14496), .ZN(P2_U3511) );
  INV_X1 U16471 ( .A(n15716), .ZN(n15733) );
  INV_X1 U16472 ( .A(n14497), .ZN(n14498) );
  AOI211_X1 U16473 ( .C1(n15733), .C2(n14500), .A(n14499), .B(n14498), .ZN(
        n14567) );
  MUX2_X1 U16474 ( .A(n14501), .B(n14567), .S(n15750), .Z(n14502) );
  OAI21_X1 U16475 ( .B1(n14570), .B2(n14514), .A(n14502), .ZN(P2_U3510) );
  OAI21_X1 U16476 ( .B1(n14504), .B2(n15737), .A(n14503), .ZN(n14506) );
  AOI211_X1 U16477 ( .C1(n15733), .C2(n14507), .A(n14506), .B(n14505), .ZN(
        n14572) );
  NAND2_X1 U16478 ( .A1(n12591), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n14508) );
  OAI21_X1 U16479 ( .B1(n14572), .B2(n12591), .A(n14508), .ZN(P2_U3509) );
  OAI211_X1 U16480 ( .C1(n14511), .C2(n15716), .A(n14510), .B(n14509), .ZN(
        n14573) );
  OAI22_X1 U16481 ( .A1(n14514), .A2(n14513), .B1(n15750), .B2(n14512), .ZN(
        n14515) );
  AOI21_X1 U16482 ( .B1(n14573), .B2(n15750), .A(n14515), .ZN(n14516) );
  INV_X1 U16483 ( .A(n14516), .ZN(P2_U3508) );
  AOI21_X1 U16484 ( .B1(n14519), .B2(n14518), .A(n14517), .ZN(n14520) );
  OAI211_X1 U16485 ( .C1(n15716), .C2(n14522), .A(n14521), .B(n14520), .ZN(
        n14578) );
  MUX2_X1 U16486 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n14578), .S(n15750), .Z(
        P2_U3507) );
  MUX2_X1 U16487 ( .A(n14524), .B(n14523), .S(n15743), .Z(n14525) );
  OAI21_X1 U16488 ( .B1(n14526), .B2(n14574), .A(n14525), .ZN(P2_U3497) );
  INV_X1 U16489 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n14528) );
  OAI21_X1 U16490 ( .B1(n14530), .B2(n14574), .A(n14529), .ZN(P2_U3493) );
  INV_X1 U16491 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14532) );
  MUX2_X1 U16492 ( .A(n14532), .B(n14531), .S(n15743), .Z(n14533) );
  OAI21_X1 U16493 ( .B1(n14534), .B2(n14574), .A(n14533), .ZN(P2_U3492) );
  INV_X1 U16494 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n14536) );
  MUX2_X1 U16495 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14538), .S(n15743), .Z(
        n14539) );
  INV_X1 U16496 ( .A(n14539), .ZN(n14540) );
  OAI21_X1 U16497 ( .B1(n14541), .B2(n14574), .A(n14540), .ZN(P2_U3490) );
  INV_X1 U16498 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n14543) );
  MUX2_X1 U16499 ( .A(n14543), .B(n14542), .S(n15743), .Z(n14544) );
  OAI21_X1 U16500 ( .B1(n14545), .B2(n14574), .A(n14544), .ZN(P2_U3489) );
  INV_X1 U16501 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n14546) );
  MUX2_X1 U16502 ( .A(n14546), .B(n8033), .S(n15743), .Z(n14547) );
  OAI21_X1 U16503 ( .B1(n14548), .B2(n14574), .A(n14547), .ZN(P2_U3488) );
  MUX2_X1 U16504 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14549), .S(n15743), .Z(
        P2_U3487) );
  MUX2_X1 U16505 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14550), .S(n15743), .Z(
        P2_U3486) );
  MUX2_X1 U16506 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14551), .S(n15743), .Z(
        P2_U3484) );
  INV_X1 U16507 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14553) );
  MUX2_X1 U16508 ( .A(n14553), .B(n14552), .S(n15743), .Z(n14554) );
  OAI21_X1 U16509 ( .B1(n14555), .B2(n14574), .A(n14554), .ZN(P2_U3481) );
  MUX2_X1 U16510 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14556), .S(n15743), .Z(
        P2_U3478) );
  MUX2_X1 U16511 ( .A(n14558), .B(n14557), .S(n15743), .Z(n14559) );
  OAI21_X1 U16512 ( .B1(n14560), .B2(n14574), .A(n14559), .ZN(P2_U3475) );
  MUX2_X1 U16513 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n14561), .S(n15743), .Z(
        P2_U3472) );
  MUX2_X1 U16514 ( .A(n15879), .B(n14562), .S(n15743), .Z(n14563) );
  OAI21_X1 U16515 ( .B1(n14564), .B2(n14574), .A(n14563), .ZN(P2_U3469) );
  NAND2_X1 U16516 ( .A1(n15741), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n14565) );
  OAI21_X1 U16517 ( .B1(n14566), .B2(n15741), .A(n14565), .ZN(P2_U3466) );
  MUX2_X1 U16518 ( .A(n14568), .B(n14567), .S(n15743), .Z(n14569) );
  OAI21_X1 U16519 ( .B1(n14570), .B2(n14574), .A(n14569), .ZN(P2_U3463) );
  NAND2_X1 U16520 ( .A1(n15741), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n14571) );
  OAI21_X1 U16521 ( .B1(n14572), .B2(n15741), .A(n14571), .ZN(P2_U3460) );
  INV_X1 U16522 ( .A(n14573), .ZN(n14577) );
  AOI22_X1 U16523 ( .A1(n8433), .A2(n14575), .B1(P2_REG0_REG_9__SCAN_IN), .B2(
        n15741), .ZN(n14576) );
  OAI21_X1 U16524 ( .B1(n14577), .B2(n15741), .A(n14576), .ZN(P2_U3457) );
  MUX2_X1 U16525 ( .A(P2_REG0_REG_8__SCAN_IN), .B(n14578), .S(n15743), .Z(
        P2_U3454) );
  INV_X1 U16526 ( .A(n14579), .ZN(n15369) );
  NAND3_X1 U16527 ( .A1(n14581), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n14583) );
  OAI22_X1 U16528 ( .A1(n14580), .A2(n14583), .B1(n14582), .B2(n14590), .ZN(
        n14584) );
  INV_X1 U16529 ( .A(n14584), .ZN(n14585) );
  OAI21_X1 U16530 ( .B1(n15369), .B2(n14594), .A(n14585), .ZN(P2_U3296) );
  INV_X1 U16531 ( .A(n14586), .ZN(n15375) );
  OAI222_X1 U16532 ( .A1(n14590), .A2(n14589), .B1(P2_U3088), .B2(n14587), 
        .C1(n14594), .C2(n15375), .ZN(P2_U3298) );
  AOI21_X1 U16533 ( .B1(n14592), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n14591), 
        .ZN(n14593) );
  OAI21_X1 U16534 ( .B1(n14595), .B2(n14594), .A(n14593), .ZN(P2_U3299) );
  INV_X1 U16535 ( .A(n14596), .ZN(n14597) );
  MUX2_X1 U16536 ( .A(n14597), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  INV_X1 U16537 ( .A(n14598), .ZN(n14599) );
  AOI21_X1 U16538 ( .B1(n14601), .B2(n14600), .A(n14599), .ZN(n14605) );
  AOI22_X1 U16539 ( .A1(n14627), .A2(n15181), .B1(n14690), .B2(n15188), .ZN(
        n14602) );
  NAND2_X1 U16540 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n14857)
         );
  OAI211_X1 U16541 ( .C1(n14681), .C2(n14706), .A(n14602), .B(n14857), .ZN(
        n14603) );
  AOI21_X1 U16542 ( .B1(n15314), .B2(n14740), .A(n14603), .ZN(n14604) );
  OAI21_X1 U16543 ( .B1(n14605), .B2(n14742), .A(n14604), .ZN(P1_U3215) );
  INV_X1 U16544 ( .A(n14606), .ZN(n14727) );
  INV_X1 U16545 ( .A(n14607), .ZN(n14609) );
  NOR3_X1 U16546 ( .A1(n14727), .A2(n14609), .A3(n14608), .ZN(n14611) );
  INV_X1 U16547 ( .A(n14610), .ZN(n14697) );
  OAI21_X1 U16548 ( .B1(n14611), .B2(n14697), .A(n14753), .ZN(n14618) );
  NAND2_X1 U16549 ( .A1(n14773), .A2(n15178), .ZN(n14613) );
  NAND2_X1 U16550 ( .A1(n15051), .A2(n15180), .ZN(n14612) );
  NAND2_X1 U16551 ( .A1(n14613), .A2(n14612), .ZN(n15258) );
  INV_X1 U16552 ( .A(n15021), .ZN(n14615) );
  OAI22_X1 U16553 ( .A1(n14615), .A2(n14759), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14614), .ZN(n14616) );
  AOI21_X1 U16554 ( .B1(n15258), .B2(n14762), .A(n14616), .ZN(n14617) );
  OAI211_X1 U16555 ( .C1(n14619), .C2(n14765), .A(n14618), .B(n14617), .ZN(
        P1_U3216) );
  OAI211_X1 U16556 ( .C1(n14622), .C2(n14621), .A(n14620), .B(n14753), .ZN(
        n14626) );
  AOI22_X1 U16557 ( .A1(n14740), .A2(n14623), .B1(n14762), .B2(n15545), .ZN(
        n14625) );
  MUX2_X1 U16558 ( .A(n14759), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n14624) );
  NAND3_X1 U16559 ( .A1(n14626), .A2(n14625), .A3(n14624), .ZN(P1_U3218) );
  AOI22_X1 U16560 ( .A1(n14627), .A2(n14777), .B1(n14690), .B2(n15091), .ZN(
        n14628) );
  NAND2_X1 U16561 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n15820)
         );
  OAI211_X1 U16562 ( .C1(n15090), .C2(n14706), .A(n14628), .B(n15820), .ZN(
        n14634) );
  INV_X1 U16563 ( .A(n14629), .ZN(n14630) );
  AOI211_X1 U16564 ( .C1(n14632), .C2(n14631), .A(n14742), .B(n14630), .ZN(
        n14633) );
  AOI211_X1 U16565 ( .C1(n14740), .C2(n15287), .A(n14634), .B(n14633), .ZN(
        n14635) );
  INV_X1 U16566 ( .A(n14635), .ZN(P1_U3219) );
  INV_X1 U16567 ( .A(n14648), .ZN(n14641) );
  OAI22_X1 U16568 ( .A1(n14947), .A2(n10379), .B1(n14959), .B2(n14636), .ZN(
        n14637) );
  XNOR2_X1 U16569 ( .A(n14637), .B(n12534), .ZN(n14640) );
  OAI22_X1 U16570 ( .A1(n14947), .A2(n14638), .B1(n14959), .B2(n10379), .ZN(
        n14639) );
  XNOR2_X1 U16571 ( .A(n14640), .B(n14639), .ZN(n14650) );
  NAND3_X1 U16572 ( .A1(n14641), .A2(n14753), .A3(n14650), .ZN(n14654) );
  OAI22_X1 U16573 ( .A1(n14944), .A2(n14759), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14642), .ZN(n14643) );
  AOI21_X1 U16574 ( .B1(n14768), .B2(n14720), .A(n14643), .ZN(n14644) );
  OAI21_X1 U16575 ( .B1(n14939), .B2(n14715), .A(n14644), .ZN(n14645) );
  AOI21_X1 U16576 ( .B1(n15220), .B2(n14740), .A(n14645), .ZN(n14653) );
  INV_X1 U16577 ( .A(n14649), .ZN(n14647) );
  INV_X1 U16578 ( .A(n14650), .ZN(n14646) );
  NAND4_X1 U16579 ( .A1(n14648), .A2(n14753), .A3(n14647), .A4(n14646), .ZN(
        n14652) );
  NAND3_X1 U16580 ( .A1(n14650), .A2(n14753), .A3(n14649), .ZN(n14651) );
  NAND4_X1 U16581 ( .A1(n14654), .A2(n14653), .A3(n14652), .A4(n14651), .ZN(
        P1_U3220) );
  OAI21_X1 U16582 ( .B1(n14657), .B2(n14656), .A(n14655), .ZN(n14658) );
  NAND2_X1 U16583 ( .A1(n14658), .A2(n14753), .ZN(n14663) );
  NOR2_X1 U16584 ( .A1(n15090), .A2(n14715), .ZN(n14661) );
  OAI22_X1 U16585 ( .A1(n14659), .A2(n14706), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15949), .ZN(n14660) );
  AOI211_X1 U16586 ( .C1(n14690), .C2(n15057), .A(n14661), .B(n14660), .ZN(
        n14662) );
  OAI211_X1 U16587 ( .C1(n15059), .C2(n14765), .A(n14663), .B(n14662), .ZN(
        P1_U3223) );
  NOR3_X1 U16588 ( .A1(n6615), .A2(n7978), .A3(n14665), .ZN(n14668) );
  INV_X1 U16589 ( .A(n14666), .ZN(n14667) );
  OAI21_X1 U16590 ( .B1(n14668), .B2(n14667), .A(n14753), .ZN(n14672) );
  AOI22_X1 U16591 ( .A1(n14995), .A2(n14690), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14669) );
  OAI21_X1 U16592 ( .B1(n14989), .B2(n14715), .A(n14669), .ZN(n14670) );
  AOI21_X1 U16593 ( .B1(n14771), .B2(n14720), .A(n14670), .ZN(n14671) );
  OAI211_X1 U16594 ( .C1(n15245), .C2(n14765), .A(n14672), .B(n14671), .ZN(
        P1_U3225) );
  INV_X1 U16595 ( .A(n14674), .ZN(n14675) );
  XNOR2_X1 U16596 ( .A(n14673), .B(n14674), .ZN(n14756) );
  NAND2_X1 U16597 ( .A1(n14756), .A2(n14755), .ZN(n14754) );
  OAI21_X1 U16598 ( .B1(n14675), .B2(n14673), .A(n14754), .ZN(n14679) );
  XOR2_X1 U16599 ( .A(n14677), .B(n14676), .Z(n14678) );
  XNOR2_X1 U16600 ( .A(n14679), .B(n14678), .ZN(n14685) );
  NAND2_X1 U16601 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14880)
         );
  OAI21_X1 U16602 ( .B1(n14706), .B2(n14680), .A(n14880), .ZN(n14683) );
  OAI22_X1 U16603 ( .A1(n14759), .A2(n15144), .B1(n14681), .B2(n14715), .ZN(
        n14682) );
  AOI211_X1 U16604 ( .C1(n15302), .C2(n14740), .A(n14683), .B(n14682), .ZN(
        n14684) );
  OAI21_X1 U16605 ( .B1(n14685), .B2(n14742), .A(n14684), .ZN(P1_U3226) );
  XOR2_X1 U16606 ( .A(n14688), .B(n14687), .Z(n14689) );
  XNOR2_X1 U16607 ( .A(n14686), .B(n14689), .ZN(n14694) );
  AOI22_X1 U16608 ( .A1(n14720), .A2(n14777), .B1(n14690), .B2(n15135), .ZN(
        n14691) );
  NAND2_X1 U16609 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14895)
         );
  OAI211_X1 U16610 ( .C1(n15129), .C2(n14715), .A(n14691), .B(n14895), .ZN(
        n14692) );
  AOI21_X1 U16611 ( .B1(n15298), .B2(n14740), .A(n14692), .ZN(n14693) );
  OAI21_X1 U16612 ( .B1(n14694), .B2(n14742), .A(n14693), .ZN(P1_U3228) );
  NOR3_X1 U16613 ( .A1(n14697), .A2(n7979), .A3(n14696), .ZN(n14698) );
  OAI21_X1 U16614 ( .B1(n14698), .B2(n6615), .A(n14753), .ZN(n14702) );
  OAI22_X1 U16615 ( .A1(n14748), .A2(n15130), .B1(n14729), .B2(n15128), .ZN(
        n15252) );
  OAI22_X1 U16616 ( .A1(n15012), .A2(n14759), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14699), .ZN(n14700) );
  AOI21_X1 U16617 ( .B1(n15252), .B2(n14762), .A(n14700), .ZN(n14701) );
  OAI211_X1 U16618 ( .C1(n15016), .C2(n14765), .A(n14702), .B(n14701), .ZN(
        P1_U3229) );
  XNOR2_X1 U16619 ( .A(n14704), .B(n14703), .ZN(n14711) );
  OAI22_X1 U16620 ( .A1(n15071), .A2(n14706), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14705), .ZN(n14709) );
  INV_X1 U16621 ( .A(n15079), .ZN(n14707) );
  OAI22_X1 U16622 ( .A1(n14759), .A2(n14707), .B1(n15070), .B2(n14715), .ZN(
        n14708) );
  AOI211_X1 U16623 ( .C1(n15278), .C2(n14740), .A(n14709), .B(n14708), .ZN(
        n14710) );
  OAI21_X1 U16624 ( .B1(n14711), .B2(n14742), .A(n14710), .ZN(P1_U3233) );
  OAI211_X1 U16625 ( .C1(n14714), .C2(n14713), .A(n14712), .B(n14753), .ZN(
        n14722) );
  OAI22_X1 U16626 ( .A1(n14759), .A2(n14717), .B1(n14716), .B2(n14715), .ZN(
        n14718) );
  AOI211_X1 U16627 ( .C1(n14720), .C2(n14779), .A(n14719), .B(n14718), .ZN(
        n14721) );
  OAI211_X1 U16628 ( .C1(n14723), .C2(n14765), .A(n14722), .B(n14721), .ZN(
        P1_U3234) );
  INV_X1 U16629 ( .A(n14655), .ZN(n14726) );
  NOR3_X1 U16630 ( .A1(n14726), .A2(n14725), .A3(n14724), .ZN(n14728) );
  OAI21_X1 U16631 ( .B1(n14728), .B2(n14727), .A(n14753), .ZN(n14732) );
  OAI22_X1 U16632 ( .A1(n14729), .A2(n15130), .B1(n15071), .B2(n15128), .ZN(
        n15038) );
  OAI22_X1 U16633 ( .A1(n14759), .A2(n15040), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n16040), .ZN(n14730) );
  AOI21_X1 U16634 ( .B1(n15038), .B2(n14762), .A(n14730), .ZN(n14731) );
  OAI211_X1 U16635 ( .C1(n14765), .C2(n15044), .A(n14732), .B(n14731), .ZN(
        P1_U3235) );
  INV_X1 U16636 ( .A(n14734), .ZN(n14735) );
  AOI21_X1 U16637 ( .B1(n14736), .B2(n14733), .A(n14735), .ZN(n14743) );
  NOR2_X1 U16638 ( .A1(n14759), .A2(n15116), .ZN(n14739) );
  AOI22_X1 U16639 ( .A1(n14776), .A2(n15178), .B1(n15180), .B2(n15151), .ZN(
        n15110) );
  NAND2_X1 U16640 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14910)
         );
  OAI21_X1 U16641 ( .B1(n15110), .B2(n14737), .A(n14910), .ZN(n14738) );
  AOI211_X1 U16642 ( .C1(n15294), .C2(n14740), .A(n14739), .B(n14738), .ZN(
        n14741) );
  OAI21_X1 U16643 ( .B1(n14743), .B2(n14742), .A(n14741), .ZN(P1_U3238) );
  OAI21_X1 U16644 ( .B1(n14746), .B2(n14745), .A(n14744), .ZN(n14747) );
  NAND2_X1 U16645 ( .A1(n14747), .A2(n14753), .ZN(n14752) );
  OAI22_X1 U16646 ( .A1(n14939), .A2(n15130), .B1(n14748), .B2(n15128), .ZN(
        n15235) );
  OAI22_X1 U16647 ( .A1(n14976), .A2(n14759), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14749), .ZN(n14750) );
  AOI21_X1 U16648 ( .B1(n15235), .B2(n14762), .A(n14750), .ZN(n14751) );
  OAI211_X1 U16649 ( .C1(n14980), .C2(n14765), .A(n14752), .B(n14751), .ZN(
        P1_U3240) );
  INV_X1 U16650 ( .A(n15308), .ZN(n14766) );
  OAI211_X1 U16651 ( .C1(n14756), .C2(n14755), .A(n14754), .B(n14753), .ZN(
        n14764) );
  NAND2_X1 U16652 ( .A1(n14778), .A2(n15178), .ZN(n14757) );
  OAI21_X1 U16653 ( .B1(n14758), .B2(n15128), .A(n14757), .ZN(n15167) );
  NAND2_X1 U16654 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15488)
         );
  INV_X1 U16655 ( .A(n15488), .ZN(n14761) );
  NOR2_X1 U16656 ( .A1(n14759), .A2(n15171), .ZN(n14760) );
  AOI211_X1 U16657 ( .C1(n14762), .C2(n15167), .A(n14761), .B(n14760), .ZN(
        n14763) );
  OAI211_X1 U16658 ( .C1(n14766), .C2(n14765), .A(n14764), .B(n14763), .ZN(
        P1_U3241) );
  MUX2_X1 U16659 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14918), .S(n14791), .Z(
        P1_U3591) );
  MUX2_X1 U16660 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14767), .S(n14791), .Z(
        P1_U3590) );
  MUX2_X1 U16661 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14768), .S(n14791), .Z(
        P1_U3589) );
  MUX2_X1 U16662 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14769), .S(n14791), .Z(
        P1_U3588) );
  MUX2_X1 U16663 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14770), .S(n14791), .Z(
        P1_U3587) );
  MUX2_X1 U16664 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14771), .S(n14791), .Z(
        P1_U3586) );
  MUX2_X1 U16665 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14772), .S(n14791), .Z(
        P1_U3585) );
  MUX2_X1 U16666 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14773), .S(n14791), .Z(
        P1_U3584) );
  MUX2_X1 U16667 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14774), .S(n14791), .Z(
        P1_U3583) );
  MUX2_X1 U16668 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n15051), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16669 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14775), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16670 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n15050), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16671 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14776), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16672 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14777), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16673 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n15151), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16674 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14778), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16675 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n15179), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16676 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14779), .S(n14791), .Z(
        P1_U3574) );
  MUX2_X1 U16677 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n15181), .S(n14791), .Z(
        P1_U3573) );
  MUX2_X1 U16678 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14780), .S(n14791), .Z(
        P1_U3572) );
  MUX2_X1 U16679 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14781), .S(n14791), .Z(
        P1_U3571) );
  MUX2_X1 U16680 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14782), .S(n14791), .Z(
        P1_U3570) );
  MUX2_X1 U16681 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14783), .S(n14791), .Z(
        P1_U3569) );
  MUX2_X1 U16682 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14784), .S(n14791), .Z(
        P1_U3568) );
  MUX2_X1 U16683 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14785), .S(n14791), .Z(
        P1_U3567) );
  MUX2_X1 U16684 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14786), .S(n14791), .Z(
        P1_U3566) );
  MUX2_X1 U16685 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14787), .S(n14791), .Z(
        P1_U3565) );
  MUX2_X1 U16686 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14788), .S(n14791), .Z(
        P1_U3564) );
  MUX2_X1 U16687 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14789), .S(n14791), .Z(
        P1_U3563) );
  MUX2_X1 U16688 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14790), .S(n14791), .Z(
        P1_U3562) );
  MUX2_X1 U16689 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14792), .S(n14791), .Z(
        P1_U3561) );
  OAI22_X1 U16690 ( .A1(n15821), .A2(n14794), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14793), .ZN(n14795) );
  AOI21_X1 U16691 ( .B1(n14796), .B2(n15483), .A(n14795), .ZN(n14805) );
  OAI211_X1 U16692 ( .C1(n10236), .C2(n14799), .A(n15812), .B(n14798), .ZN(
        n14804) );
  OAI211_X1 U16693 ( .C1(n14802), .C2(n14801), .A(n15486), .B(n14800), .ZN(
        n14803) );
  NAND3_X1 U16694 ( .A1(n14805), .A2(n14804), .A3(n14803), .ZN(P1_U3244) );
  AOI22_X1 U16695 ( .A1(n15475), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n14817) );
  OAI21_X1 U16696 ( .B1(n14807), .B2(n14806), .A(n14825), .ZN(n14812) );
  OAI21_X1 U16697 ( .B1(n14810), .B2(n14809), .A(n14808), .ZN(n14811) );
  OAI22_X1 U16698 ( .A1(n15815), .A2(n14812), .B1(n15817), .B2(n14811), .ZN(
        n14813) );
  INV_X1 U16699 ( .A(n14813), .ZN(n14816) );
  NAND2_X1 U16700 ( .A1(n15483), .A2(n14814), .ZN(n14815) );
  NAND4_X1 U16701 ( .A1(n14818), .A2(n14817), .A3(n14816), .A4(n14815), .ZN(
        P1_U3245) );
  OAI211_X1 U16702 ( .C1(n14821), .C2(n14820), .A(n15486), .B(n14819), .ZN(
        n14834) );
  MUX2_X1 U16703 ( .A(n14822), .B(P1_REG2_REG_3__SCAN_IN), .S(n14828), .Z(
        n14823) );
  NAND3_X1 U16704 ( .A1(n14825), .A2(n14824), .A3(n14823), .ZN(n14826) );
  NAND3_X1 U16705 ( .A1(n15812), .A2(n14827), .A3(n14826), .ZN(n14833) );
  NAND2_X1 U16706 ( .A1(n15483), .A2(n14828), .ZN(n14832) );
  NOR2_X1 U16707 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14829), .ZN(n14830) );
  AOI21_X1 U16708 ( .B1(n15475), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n14830), .ZN(
        n14831) );
  NAND4_X1 U16709 ( .A1(n14834), .A2(n14833), .A3(n14832), .A4(n14831), .ZN(
        P1_U3246) );
  OAI21_X1 U16710 ( .B1(n14837), .B2(n14836), .A(n14835), .ZN(n14838) );
  NAND2_X1 U16711 ( .A1(n14838), .A2(n15486), .ZN(n14851) );
  OAI21_X1 U16712 ( .B1(n15821), .B2(n14840), .A(n14839), .ZN(n14841) );
  AOI21_X1 U16713 ( .B1(n14842), .B2(n15483), .A(n14841), .ZN(n14850) );
  MUX2_X1 U16714 ( .A(n10654), .B(P1_REG2_REG_9__SCAN_IN), .S(n14842), .Z(
        n14845) );
  INV_X1 U16715 ( .A(n14843), .ZN(n14844) );
  NAND2_X1 U16716 ( .A1(n14845), .A2(n14844), .ZN(n14847) );
  OAI211_X1 U16717 ( .C1(n14848), .C2(n14847), .A(n14846), .B(n15812), .ZN(
        n14849) );
  NAND3_X1 U16718 ( .A1(n14851), .A2(n14850), .A3(n14849), .ZN(P1_U3252) );
  XNOR2_X1 U16719 ( .A(n14868), .B(n14852), .ZN(n14855) );
  OAI21_X1 U16720 ( .B1(n14855), .B2(n14854), .A(n14867), .ZN(n14856) );
  NAND2_X1 U16721 ( .A1(n14856), .A2(n15486), .ZN(n14866) );
  INV_X1 U16722 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15906) );
  OAI21_X1 U16723 ( .B1(n15821), .B2(n15906), .A(n14857), .ZN(n14858) );
  AOI21_X1 U16724 ( .B1(n14868), .B2(n15483), .A(n14858), .ZN(n14865) );
  AND2_X1 U16725 ( .A1(n14859), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n14861) );
  MUX2_X1 U16726 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n15191), .S(n14868), .Z(
        n14860) );
  OAI21_X1 U16727 ( .B1(n14862), .B2(n14861), .A(n14860), .ZN(n14872) );
  OR3_X1 U16728 ( .A1(n14862), .A2(n14861), .A3(n14860), .ZN(n14863) );
  NAND3_X1 U16729 ( .A1(n14872), .A2(n15812), .A3(n14863), .ZN(n14864) );
  NAND3_X1 U16730 ( .A1(n14866), .A2(n14865), .A3(n14864), .ZN(P1_U3257) );
  XNOR2_X1 U16731 ( .A(n14887), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n14871) );
  AOI211_X1 U16732 ( .C1(n14871), .C2(n14870), .A(n15817), .B(n6736), .ZN(
        n14884) );
  OAI21_X1 U16733 ( .B1(n15191), .B2(n14873), .A(n14872), .ZN(n14874) );
  NOR2_X1 U16734 ( .A1(n14874), .A2(n15484), .ZN(n14875) );
  AOI21_X1 U16735 ( .B1(n15484), .B2(n14874), .A(n14875), .ZN(n15481) );
  INV_X1 U16736 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n15480) );
  INV_X1 U16737 ( .A(n14875), .ZN(n14876) );
  MUX2_X1 U16738 ( .A(n12269), .B(P1_REG2_REG_16__SCAN_IN), .S(n14887), .Z(
        n14877) );
  INV_X1 U16739 ( .A(n14890), .ZN(n14894) );
  AOI211_X1 U16740 ( .C1(n14878), .C2(n14877), .A(n15815), .B(n14894), .ZN(
        n14883) );
  NAND2_X1 U16741 ( .A1(n15475), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n14879) );
  OAI211_X1 U16742 ( .C1(n15814), .C2(n14881), .A(n14880), .B(n14879), .ZN(
        n14882) );
  OR3_X1 U16743 ( .A1(n14884), .A2(n14883), .A3(n14882), .ZN(P1_U3259) );
  XNOR2_X1 U16744 ( .A(n14902), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n14885) );
  AOI211_X1 U16745 ( .C1(n14886), .C2(n14885), .A(n15817), .B(n14901), .ZN(
        n14900) );
  NAND2_X1 U16746 ( .A1(n14887), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14889) );
  NAND2_X1 U16747 ( .A1(n14907), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14888) );
  OAI211_X1 U16748 ( .C1(P1_REG2_REG_17__SCAN_IN), .C2(n14907), .A(n14889), 
        .B(n14888), .ZN(n14893) );
  NAND2_X1 U16749 ( .A1(n14902), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14891) );
  OAI211_X1 U16750 ( .C1(n14902), .C2(P1_REG2_REG_17__SCAN_IN), .A(n14892), 
        .B(n14891), .ZN(n14906) );
  OAI211_X1 U16751 ( .C1(n14894), .C2(n14893), .A(n14906), .B(n15812), .ZN(
        n14898) );
  INV_X1 U16752 ( .A(n14895), .ZN(n14896) );
  AOI21_X1 U16753 ( .B1(n15475), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n14896), 
        .ZN(n14897) );
  OAI211_X1 U16754 ( .C1(n15814), .C2(n14907), .A(n14898), .B(n14897), .ZN(
        n14899) );
  OR2_X1 U16755 ( .A1(n14900), .A2(n14899), .ZN(P1_U3260) );
  NOR2_X1 U16756 ( .A1(n14904), .A2(n15808), .ZN(n14905) );
  OAI21_X1 U16757 ( .B1(n6735), .B2(P1_REG1_REG_18__SCAN_IN), .A(n15486), .ZN(
        n14915) );
  INV_X1 U16758 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14908) );
  OAI21_X1 U16759 ( .B1(n14908), .B2(n14907), .A(n14906), .ZN(n15809) );
  XNOR2_X1 U16760 ( .A(n15809), .B(n15808), .ZN(n15810) );
  XNOR2_X1 U16761 ( .A(n15810), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n14913) );
  NAND2_X1 U16762 ( .A1(n15475), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n14909) );
  OAI211_X1 U16763 ( .C1(n15814), .C2(n14911), .A(n14910), .B(n14909), .ZN(
        n14912) );
  AOI21_X1 U16764 ( .B1(n14913), .B2(n15812), .A(n14912), .ZN(n14914) );
  OAI21_X1 U16765 ( .B1(n14915), .B2(n15806), .A(n14914), .ZN(P1_U3261) );
  XNOR2_X1 U16766 ( .A(n14924), .B(n14916), .ZN(n14917) );
  NAND2_X1 U16767 ( .A1(n14917), .A2(n15517), .ZN(n15200) );
  NAND2_X1 U16768 ( .A1(n14919), .A2(n14918), .ZN(n15204) );
  NOR2_X1 U16769 ( .A1(n15512), .A2(n15204), .ZN(n14928) );
  NOR2_X1 U16770 ( .A1(n15201), .A2(n15147), .ZN(n14920) );
  AOI211_X1 U16771 ( .C1(n15525), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14928), 
        .B(n14920), .ZN(n14921) );
  OAI21_X1 U16772 ( .B1(n15082), .B2(n15200), .A(n14921), .ZN(P1_U3263) );
  INV_X1 U16773 ( .A(n14922), .ZN(n14926) );
  INV_X1 U16774 ( .A(n14924), .ZN(n14925) );
  OAI211_X1 U16775 ( .C1(n14926), .C2(n15206), .A(n14925), .B(n15517), .ZN(
        n15205) );
  NOR2_X1 U16776 ( .A1(n15206), .A2(n15147), .ZN(n14927) );
  AOI211_X1 U16777 ( .C1(n15525), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14928), 
        .B(n14927), .ZN(n14929) );
  OAI21_X1 U16778 ( .B1(n15082), .B2(n15205), .A(n14929), .ZN(P1_U3264) );
  INV_X1 U16779 ( .A(n15218), .ZN(n14952) );
  INV_X1 U16780 ( .A(n14931), .ZN(n14932) );
  NAND2_X1 U16781 ( .A1(n14954), .A2(n14932), .ZN(n14936) );
  INV_X1 U16782 ( .A(n14936), .ZN(n14934) );
  NAND2_X1 U16783 ( .A1(n14934), .A2(n14933), .ZN(n15216) );
  NAND2_X1 U16784 ( .A1(n14936), .A2(n14935), .ZN(n15217) );
  NAND3_X1 U16785 ( .A1(n15216), .A2(n15101), .A3(n15217), .ZN(n14951) );
  OAI21_X1 U16786 ( .B1(n14957), .B2(n14947), .A(n15517), .ZN(n14938) );
  INV_X1 U16787 ( .A(n15222), .ZN(n14949) );
  OR2_X1 U16788 ( .A1(n14939), .A2(n15128), .ZN(n14942) );
  OR2_X1 U16789 ( .A1(n14940), .A2(n15130), .ZN(n14941) );
  NAND2_X1 U16790 ( .A1(n14942), .A2(n14941), .ZN(n15219) );
  INV_X1 U16791 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n14943) );
  OAI22_X1 U16792 ( .A1(n14944), .A2(n15189), .B1(n14943), .B2(n15097), .ZN(
        n14945) );
  AOI21_X1 U16793 ( .B1(n15219), .B2(n15097), .A(n14945), .ZN(n14946) );
  OAI21_X1 U16794 ( .B1(n14947), .B2(n15147), .A(n14946), .ZN(n14948) );
  AOI21_X1 U16795 ( .B1(n14949), .B2(n15521), .A(n14948), .ZN(n14950) );
  OAI211_X1 U16796 ( .C1(n14952), .C2(n15104), .A(n14951), .B(n14950), .ZN(
        P1_U3265) );
  XOR2_X1 U16797 ( .A(n14955), .B(n14953), .Z(n15233) );
  OAI21_X1 U16798 ( .B1(n14956), .B2(n14955), .A(n14954), .ZN(n15227) );
  NAND2_X1 U16799 ( .A1(n15227), .A2(n15101), .ZN(n14965) );
  AOI211_X1 U16800 ( .C1(n15230), .C2(n14974), .A(n15538), .B(n14957), .ZN(
        n15228) );
  AOI22_X1 U16801 ( .A1(n14958), .A2(n15513), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n15512), .ZN(n14961) );
  OAI22_X1 U16802 ( .A1(n14959), .A2(n15130), .B1(n14990), .B2(n15128), .ZN(
        n15229) );
  NAND2_X1 U16803 ( .A1(n15229), .A2(n15097), .ZN(n14960) );
  OAI211_X1 U16804 ( .C1(n14962), .C2(n15147), .A(n14961), .B(n14960), .ZN(
        n14963) );
  AOI21_X1 U16805 ( .B1(n15228), .B2(n15521), .A(n14963), .ZN(n14964) );
  OAI211_X1 U16806 ( .C1(n15233), .C2(n15104), .A(n14965), .B(n14964), .ZN(
        P1_U3266) );
  NAND2_X1 U16807 ( .A1(n15249), .A2(n14967), .ZN(n14985) );
  INV_X1 U16808 ( .A(n14999), .ZN(n14984) );
  OR2_X2 U16809 ( .A1(n14985), .A2(n14984), .ZN(n14987) );
  NAND2_X1 U16810 ( .A1(n14987), .A2(n14968), .ZN(n14970) );
  XNOR2_X1 U16811 ( .A(n14970), .B(n14969), .ZN(n15240) );
  AOI21_X1 U16812 ( .B1(n14973), .B2(n14972), .A(n14971), .ZN(n15237) );
  NAND2_X1 U16813 ( .A1(n15237), .A2(n15101), .ZN(n14983) );
  INV_X1 U16814 ( .A(n14974), .ZN(n14975) );
  AOI211_X1 U16815 ( .C1(n15236), .C2(n14994), .A(n15538), .B(n14975), .ZN(
        n15234) );
  INV_X1 U16816 ( .A(n14976), .ZN(n14977) );
  AOI22_X1 U16817 ( .A1(n14977), .A2(n15513), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n15512), .ZN(n14979) );
  NAND2_X1 U16818 ( .A1(n15235), .A2(n15097), .ZN(n14978) );
  OAI211_X1 U16819 ( .C1(n14980), .C2(n15147), .A(n14979), .B(n14978), .ZN(
        n14981) );
  AOI21_X1 U16820 ( .B1(n15234), .B2(n15521), .A(n14981), .ZN(n14982) );
  OAI211_X1 U16821 ( .C1(n15240), .C2(n15104), .A(n14983), .B(n14982), .ZN(
        P1_U3267) );
  NAND2_X1 U16822 ( .A1(n14985), .A2(n14984), .ZN(n14986) );
  NAND2_X1 U16823 ( .A1(n14987), .A2(n14986), .ZN(n14988) );
  NAND2_X1 U16824 ( .A1(n14988), .A2(n15552), .ZN(n14993) );
  OAI22_X1 U16825 ( .A1(n14990), .A2(n15130), .B1(n14989), .B2(n15128), .ZN(
        n14991) );
  INV_X1 U16826 ( .A(n14991), .ZN(n14992) );
  NAND2_X1 U16827 ( .A1(n14993), .A2(n14992), .ZN(n15248) );
  INV_X1 U16828 ( .A(n15248), .ZN(n15004) );
  OAI211_X1 U16829 ( .C1(n15010), .C2(n15245), .A(n15517), .B(n14994), .ZN(
        n15244) );
  INV_X1 U16830 ( .A(n15244), .ZN(n14998) );
  AOI22_X1 U16831 ( .A1(n14995), .A2(n15513), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n15512), .ZN(n14996) );
  OAI21_X1 U16832 ( .B1(n15245), .B2(n15147), .A(n14996), .ZN(n14997) );
  AOI21_X1 U16833 ( .B1(n14998), .B2(n15521), .A(n14997), .ZN(n15003) );
  INV_X1 U16834 ( .A(n15243), .ZN(n15001) );
  NAND2_X1 U16835 ( .A1(n15000), .A2(n14999), .ZN(n15241) );
  NAND3_X1 U16836 ( .A1(n15001), .A2(n15101), .A3(n15241), .ZN(n15002) );
  OAI211_X1 U16837 ( .C1(n15004), .C2(n15512), .A(n15003), .B(n15002), .ZN(
        P1_U3268) );
  XNOR2_X1 U16838 ( .A(n15005), .B(n15007), .ZN(n15256) );
  INV_X1 U16839 ( .A(n15006), .ZN(n15008) );
  NAND2_X1 U16840 ( .A1(n15008), .A2(n15007), .ZN(n15250) );
  NAND3_X1 U16841 ( .A1(n15250), .A2(n15009), .A3(n15249), .ZN(n15019) );
  OAI21_X1 U16842 ( .B1(n15025), .B2(n15016), .A(n15517), .ZN(n15011) );
  NOR2_X1 U16843 ( .A1(n15011), .A2(n15010), .ZN(n15251) );
  INV_X1 U16844 ( .A(n15012), .ZN(n15013) );
  AOI22_X1 U16845 ( .A1(n15013), .A2(n15513), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n15525), .ZN(n15015) );
  NAND2_X1 U16846 ( .A1(n15252), .A2(n15097), .ZN(n15014) );
  OAI211_X1 U16847 ( .C1(n15016), .C2(n15147), .A(n15015), .B(n15014), .ZN(
        n15017) );
  AOI21_X1 U16848 ( .B1(n15251), .B2(n15521), .A(n15017), .ZN(n15018) );
  OAI211_X1 U16849 ( .C1(n15122), .C2(n15256), .A(n15019), .B(n15018), .ZN(
        P1_U3269) );
  XNOR2_X1 U16850 ( .A(n15020), .B(n15029), .ZN(n15257) );
  INV_X1 U16851 ( .A(n15257), .ZN(n15033) );
  INV_X1 U16852 ( .A(n15258), .ZN(n15023) );
  AOI22_X1 U16853 ( .A1(n15021), .A2(n15513), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n15512), .ZN(n15022) );
  OAI21_X1 U16854 ( .B1(n15023), .B2(n15512), .A(n15022), .ZN(n15028) );
  NAND2_X1 U16855 ( .A1(n6630), .A2(n15259), .ZN(n15024) );
  NAND2_X1 U16856 ( .A1(n15024), .A2(n15517), .ZN(n15026) );
  OR2_X1 U16857 ( .A1(n15026), .A2(n15025), .ZN(n15262) );
  NOR2_X1 U16858 ( .A1(n15262), .A2(n15082), .ZN(n15027) );
  AOI211_X1 U16859 ( .C1(n15515), .C2(n15259), .A(n15028), .B(n15027), .ZN(
        n15032) );
  NAND2_X1 U16860 ( .A1(n15030), .A2(n15029), .ZN(n15260) );
  NAND3_X1 U16861 ( .A1(n15261), .A2(n15260), .A3(n15101), .ZN(n15031) );
  OAI211_X1 U16862 ( .C1(n15033), .C2(n15104), .A(n15032), .B(n15031), .ZN(
        P1_U3270) );
  XNOR2_X1 U16863 ( .A(n15034), .B(n15037), .ZN(n15270) );
  OAI21_X1 U16864 ( .B1(n15037), .B2(n15036), .A(n15035), .ZN(n15039) );
  AOI21_X1 U16865 ( .B1(n15039), .B2(n15552), .A(n15038), .ZN(n15269) );
  OAI21_X1 U16866 ( .B1(n15040), .B2(n15189), .A(n15269), .ZN(n15041) );
  NAND2_X1 U16867 ( .A1(n15041), .A2(n15097), .ZN(n15047) );
  AOI21_X1 U16868 ( .B1(n15054), .B2(n15267), .A(n15538), .ZN(n15042) );
  AND2_X1 U16869 ( .A1(n15042), .A2(n6630), .ZN(n15266) );
  INV_X1 U16870 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n15043) );
  OAI22_X1 U16871 ( .A1(n15044), .A2(n15147), .B1(n15043), .B2(n15097), .ZN(
        n15045) );
  AOI21_X1 U16872 ( .B1(n15266), .B2(n15521), .A(n15045), .ZN(n15046) );
  OAI211_X1 U16873 ( .C1(n15270), .C2(n15195), .A(n15047), .B(n15046), .ZN(
        P1_U3271) );
  OAI211_X1 U16874 ( .C1(n15062), .C2(n15049), .A(n15048), .B(n15552), .ZN(
        n15053) );
  AOI22_X1 U16875 ( .A1(n15051), .A2(n15178), .B1(n15050), .B2(n15180), .ZN(
        n15052) );
  OR2_X1 U16876 ( .A1(n15076), .A2(n15059), .ZN(n15055) );
  AND2_X1 U16877 ( .A1(n15055), .A2(n15054), .ZN(n15272) );
  INV_X1 U16878 ( .A(n15056), .ZN(n15155) );
  AOI22_X1 U16879 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(n15512), .B1(n15057), 
        .B2(n15513), .ZN(n15058) );
  OAI21_X1 U16880 ( .B1(n15059), .B2(n15147), .A(n15058), .ZN(n15066) );
  NAND2_X1 U16881 ( .A1(n15277), .A2(n15061), .ZN(n15064) );
  INV_X1 U16882 ( .A(n15062), .ZN(n15063) );
  XNOR2_X1 U16883 ( .A(n15064), .B(n15063), .ZN(n15275) );
  NOR2_X1 U16884 ( .A1(n15275), .A2(n15195), .ZN(n15065) );
  AOI211_X1 U16885 ( .C1(n15272), .C2(n15155), .A(n15066), .B(n15065), .ZN(
        n15067) );
  OAI21_X1 U16886 ( .B1(n15525), .B2(n15274), .A(n15067), .ZN(P1_U3272) );
  OAI211_X1 U16887 ( .C1(n15069), .C2(n15075), .A(n15068), .B(n15552), .ZN(
        n15074) );
  OAI22_X1 U16888 ( .A1(n15071), .A2(n15130), .B1(n15070), .B2(n15128), .ZN(
        n15072) );
  INV_X1 U16889 ( .A(n15072), .ZN(n15073) );
  NAND2_X1 U16890 ( .A1(n15074), .A2(n15073), .ZN(n15283) );
  NAND2_X1 U16891 ( .A1(n15060), .A2(n15075), .ZN(n15276) );
  AND3_X1 U16892 ( .A1(n15277), .A2(n15101), .A3(n15276), .ZN(n15084) );
  INV_X1 U16893 ( .A(n15076), .ZN(n15078) );
  AOI21_X1 U16894 ( .B1(n15088), .B2(n15278), .A(n15538), .ZN(n15077) );
  NAND2_X1 U16895 ( .A1(n15078), .A2(n15077), .ZN(n15279) );
  AOI22_X1 U16896 ( .A1(n15525), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n15079), 
        .B2(n15513), .ZN(n15081) );
  NAND2_X1 U16897 ( .A1(n15278), .A2(n15515), .ZN(n15080) );
  OAI211_X1 U16898 ( .C1(n15279), .C2(n15082), .A(n15081), .B(n15080), .ZN(
        n15083) );
  AOI211_X1 U16899 ( .C1(n15283), .C2(n15097), .A(n15084), .B(n15083), .ZN(
        n15085) );
  INV_X1 U16900 ( .A(n15085), .ZN(P1_U3273) );
  AOI21_X1 U16901 ( .B1(n15100), .B2(n15087), .A(n15086), .ZN(n15291) );
  INV_X1 U16902 ( .A(n15088), .ZN(n15089) );
  AOI211_X1 U16903 ( .C1(n15287), .C2(n15113), .A(n15538), .B(n15089), .ZN(
        n15285) );
  INV_X1 U16904 ( .A(n15285), .ZN(n15093) );
  OAI22_X1 U16905 ( .A1(n15090), .A2(n15130), .B1(n15131), .B2(n15128), .ZN(
        n15286) );
  AOI21_X1 U16906 ( .B1(n15091), .B2(n15513), .A(n15286), .ZN(n15092) );
  OAI21_X1 U16907 ( .B1(n15093), .B2(n12672), .A(n15092), .ZN(n15098) );
  INV_X1 U16908 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n15094) );
  OAI22_X1 U16909 ( .A1(n15095), .A2(n15147), .B1(n15097), .B2(n15094), .ZN(
        n15096) );
  AOI21_X1 U16910 ( .B1(n15098), .B2(n15097), .A(n15096), .ZN(n15103) );
  XNOR2_X1 U16911 ( .A(n15099), .B(n15100), .ZN(n15288) );
  NAND2_X1 U16912 ( .A1(n15288), .A2(n15101), .ZN(n15102) );
  OAI211_X1 U16913 ( .C1(n15291), .C2(n15104), .A(n15103), .B(n15102), .ZN(
        P1_U3274) );
  XNOR2_X1 U16914 ( .A(n15106), .B(n15105), .ZN(n15296) );
  OAI211_X1 U16915 ( .C1(n15109), .C2(n15108), .A(n15107), .B(n15552), .ZN(
        n15111) );
  NAND2_X1 U16916 ( .A1(n15111), .A2(n15110), .ZN(n15292) );
  AOI21_X1 U16917 ( .B1(n15112), .B2(n15294), .A(n15538), .ZN(n15114) );
  AND2_X1 U16918 ( .A1(n15114), .A2(n15113), .ZN(n15293) );
  NAND2_X1 U16919 ( .A1(n15293), .A2(n15521), .ZN(n15119) );
  NAND2_X1 U16920 ( .A1(n15525), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n15115) );
  OAI21_X1 U16921 ( .B1(n15189), .B2(n15116), .A(n15115), .ZN(n15117) );
  AOI21_X1 U16922 ( .B1(n15294), .B2(n15515), .A(n15117), .ZN(n15118) );
  NAND2_X1 U16923 ( .A1(n15119), .A2(n15118), .ZN(n15120) );
  AOI21_X1 U16924 ( .B1(n15292), .B2(n15097), .A(n15120), .ZN(n15121) );
  OAI21_X1 U16925 ( .B1(n15122), .B2(n15296), .A(n15121), .ZN(P1_U3275) );
  XOR2_X1 U16926 ( .A(n15123), .B(n15126), .Z(n15301) );
  XNOR2_X1 U16927 ( .A(n15142), .B(n15137), .ZN(n15124) );
  NOR2_X1 U16928 ( .A1(n15124), .A2(n15538), .ZN(n15297) );
  INV_X1 U16929 ( .A(n15297), .ZN(n15134) );
  AOI21_X1 U16930 ( .B1(n15125), .B2(n15126), .A(n15558), .ZN(n15133) );
  OAI22_X1 U16931 ( .A1(n15131), .A2(n15130), .B1(n15129), .B2(n15128), .ZN(
        n15132) );
  AOI21_X1 U16932 ( .B1(n15133), .B2(n15127), .A(n15132), .ZN(n15300) );
  OAI21_X1 U16933 ( .B1(n12672), .B2(n15134), .A(n15300), .ZN(n15139) );
  AOI22_X1 U16934 ( .A1(n15525), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n15135), 
        .B2(n15513), .ZN(n15136) );
  OAI21_X1 U16935 ( .B1(n15137), .B2(n15147), .A(n15136), .ZN(n15138) );
  AOI21_X1 U16936 ( .B1(n15139), .B2(n15097), .A(n15138), .ZN(n15140) );
  OAI21_X1 U16937 ( .B1(n15195), .B2(n15301), .A(n15140), .ZN(P1_U3276) );
  XOR2_X1 U16938 ( .A(n15141), .B(n15149), .Z(n15306) );
  INV_X1 U16939 ( .A(n15169), .ZN(n15143) );
  AOI21_X1 U16940 ( .B1(n15302), .B2(n15143), .A(n15142), .ZN(n15303) );
  INV_X1 U16941 ( .A(n15144), .ZN(n15145) );
  AOI22_X1 U16942 ( .A1(n15525), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n15145), 
        .B2(n15513), .ZN(n15146) );
  OAI21_X1 U16943 ( .B1(n15148), .B2(n15147), .A(n15146), .ZN(n15154) );
  OAI21_X1 U16944 ( .B1(n6655), .B2(n12270), .A(n15150), .ZN(n15152) );
  AOI222_X1 U16945 ( .A1(n15152), .A2(n15552), .B1(n15151), .B2(n15178), .C1(
        n15179), .C2(n15180), .ZN(n15305) );
  NOR2_X1 U16946 ( .A1(n15305), .A2(n15512), .ZN(n15153) );
  AOI211_X1 U16947 ( .C1(n15303), .C2(n15155), .A(n15154), .B(n15153), .ZN(
        n15156) );
  OAI21_X1 U16948 ( .B1(n15195), .B2(n15306), .A(n15156), .ZN(P1_U3277) );
  INV_X1 U16949 ( .A(n15157), .ZN(n15158) );
  AOI21_X1 U16950 ( .B1(n7952), .B2(n15159), .A(n15158), .ZN(n15311) );
  INV_X1 U16951 ( .A(n15160), .ZN(n15161) );
  NAND2_X1 U16952 ( .A1(n15162), .A2(n15161), .ZN(n15186) );
  NAND2_X1 U16953 ( .A1(n15186), .A2(n15185), .ZN(n15184) );
  NAND3_X1 U16954 ( .A1(n15184), .A2(n15164), .A3(n15163), .ZN(n15165) );
  AND3_X1 U16955 ( .A1(n15166), .A2(n15165), .A3(n15552), .ZN(n15168) );
  NOR2_X1 U16956 ( .A1(n15168), .A2(n15167), .ZN(n15310) );
  AOI211_X1 U16957 ( .C1(n15308), .C2(n15176), .A(n15538), .B(n15169), .ZN(
        n15307) );
  NAND2_X1 U16958 ( .A1(n15307), .A2(n15819), .ZN(n15170) );
  OAI211_X1 U16959 ( .C1(n15189), .C2(n15171), .A(n15310), .B(n15170), .ZN(
        n15172) );
  NAND2_X1 U16960 ( .A1(n15172), .A2(n15097), .ZN(n15174) );
  AOI22_X1 U16961 ( .A1(n15308), .A2(n15515), .B1(P1_REG2_REG_15__SCAN_IN), 
        .B2(n15512), .ZN(n15173) );
  OAI211_X1 U16962 ( .C1(n15311), .C2(n15195), .A(n15174), .B(n15173), .ZN(
        P1_U3278) );
  AOI21_X1 U16963 ( .B1(n15175), .B2(n15314), .A(n15538), .ZN(n15177) );
  AND2_X1 U16964 ( .A1(n15177), .A2(n15176), .ZN(n15312) );
  NAND2_X1 U16965 ( .A1(n15179), .A2(n15178), .ZN(n15183) );
  NAND2_X1 U16966 ( .A1(n15181), .A2(n15180), .ZN(n15182) );
  NAND2_X1 U16967 ( .A1(n15183), .A2(n15182), .ZN(n15313) );
  OAI211_X1 U16968 ( .C1(n15186), .C2(n15185), .A(n15552), .B(n15184), .ZN(
        n15316) );
  INV_X1 U16969 ( .A(n15316), .ZN(n15187) );
  AOI211_X1 U16970 ( .C1(n15312), .C2(n15819), .A(n15313), .B(n15187), .ZN(
        n15199) );
  INV_X1 U16971 ( .A(n15188), .ZN(n15190) );
  OAI22_X1 U16972 ( .A1(n15097), .A2(n15191), .B1(n15190), .B2(n15189), .ZN(
        n15197) );
  OAI21_X1 U16973 ( .B1(n15194), .B2(n15193), .A(n15192), .ZN(n15317) );
  NOR2_X1 U16974 ( .A1(n15317), .A2(n15195), .ZN(n15196) );
  AOI211_X1 U16975 ( .C1(n15515), .C2(n15314), .A(n15197), .B(n15196), .ZN(
        n15198) );
  OAI21_X1 U16976 ( .B1(n15199), .B2(n15512), .A(n15198), .ZN(P1_U3279) );
  OAI211_X1 U16977 ( .C1(n15201), .C2(n15599), .A(n15200), .B(n15204), .ZN(
        n15342) );
  MUX2_X1 U16978 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15342), .S(n15622), .Z(
        P1_U3559) );
  OAI211_X1 U16979 ( .C1(n15206), .C2(n15599), .A(n15205), .B(n15204), .ZN(
        n15343) );
  MUX2_X1 U16980 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15343), .S(n15622), .Z(
        P1_U3558) );
  OAI211_X1 U16981 ( .C1(n15210), .C2(n15599), .A(n15209), .B(n15208), .ZN(
        n15211) );
  INV_X1 U16982 ( .A(n15211), .ZN(n15212) );
  NAND3_X1 U16983 ( .A1(n15217), .A2(n15216), .A3(n15561), .ZN(n15226) );
  NAND2_X1 U16984 ( .A1(n15218), .A2(n15552), .ZN(n15224) );
  AOI21_X1 U16985 ( .B1(n15220), .B2(n15530), .A(n15219), .ZN(n15221) );
  NAND2_X1 U16986 ( .A1(n15226), .A2(n15225), .ZN(n15344) );
  MUX2_X1 U16987 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15344), .S(n15622), .Z(
        P1_U3556) );
  NAND2_X1 U16988 ( .A1(n15227), .A2(n15561), .ZN(n15232) );
  OAI211_X1 U16989 ( .C1(n15558), .C2(n15233), .A(n15232), .B(n15231), .ZN(
        n15345) );
  MUX2_X1 U16990 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15345), .S(n15622), .Z(
        P1_U3555) );
  AOI211_X1 U16991 ( .C1(n15530), .C2(n15236), .A(n15235), .B(n15234), .ZN(
        n15239) );
  NAND2_X1 U16992 ( .A1(n15237), .A2(n15561), .ZN(n15238) );
  OAI211_X1 U16993 ( .C1(n15240), .C2(n15558), .A(n15239), .B(n15238), .ZN(
        n15346) );
  MUX2_X1 U16994 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15346), .S(n15622), .Z(
        P1_U3554) );
  NAND2_X1 U16995 ( .A1(n15241), .A2(n15561), .ZN(n15242) );
  NOR2_X1 U16996 ( .A1(n15243), .A2(n15242), .ZN(n15247) );
  OAI21_X1 U16997 ( .B1(n15245), .B2(n15599), .A(n15244), .ZN(n15246) );
  OR3_X2 U16998 ( .A1(n15248), .A2(n15247), .A3(n15246), .ZN(n15347) );
  MUX2_X1 U16999 ( .A(n15347), .B(P1_REG1_REG_25__SCAN_IN), .S(n15620), .Z(
        P1_U3553) );
  NAND3_X1 U17000 ( .A1(n15250), .A2(n15552), .A3(n15249), .ZN(n15255) );
  AOI211_X1 U17001 ( .C1(n15530), .C2(n15253), .A(n15252), .B(n15251), .ZN(
        n15254) );
  OAI211_X1 U17002 ( .C1(n15588), .C2(n15256), .A(n15255), .B(n15254), .ZN(
        n15348) );
  MUX2_X1 U17003 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15348), .S(n15622), .Z(
        P1_U3552) );
  NAND2_X1 U17004 ( .A1(n15257), .A2(n15552), .ZN(n15265) );
  AOI21_X1 U17005 ( .B1(n15259), .B2(n15530), .A(n15258), .ZN(n15264) );
  NAND3_X1 U17006 ( .A1(n15261), .A2(n15561), .A3(n15260), .ZN(n15263) );
  NAND4_X1 U17007 ( .A1(n15265), .A2(n15264), .A3(n15263), .A4(n15262), .ZN(
        n15349) );
  MUX2_X1 U17008 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15349), .S(n15622), .Z(
        P1_U3551) );
  AOI21_X1 U17009 ( .B1(n15530), .B2(n15267), .A(n15266), .ZN(n15268) );
  OAI211_X1 U17010 ( .C1(n15588), .C2(n15270), .A(n15269), .B(n15268), .ZN(
        n15350) );
  MUX2_X1 U17011 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15350), .S(n15622), .Z(
        P1_U3550) );
  AOI22_X1 U17012 ( .A1(n15272), .A2(n15517), .B1(n15530), .B2(n15271), .ZN(
        n15273) );
  OAI211_X1 U17013 ( .C1(n15588), .C2(n15275), .A(n15274), .B(n15273), .ZN(
        n15351) );
  MUX2_X1 U17014 ( .A(n15351), .B(P1_REG1_REG_21__SCAN_IN), .S(n15620), .Z(
        P1_U3549) );
  NAND3_X1 U17015 ( .A1(n15277), .A2(n15561), .A3(n15276), .ZN(n15281) );
  NAND2_X1 U17016 ( .A1(n15278), .A2(n15530), .ZN(n15280) );
  NAND3_X1 U17017 ( .A1(n15281), .A2(n15280), .A3(n15279), .ZN(n15282) );
  NOR2_X1 U17018 ( .A1(n15283), .A2(n15282), .ZN(n15352) );
  MUX2_X1 U17019 ( .A(n16014), .B(n15352), .S(n15622), .Z(n15284) );
  INV_X1 U17020 ( .A(n15284), .ZN(P1_U3548) );
  AOI211_X1 U17021 ( .C1(n15530), .C2(n15287), .A(n15286), .B(n15285), .ZN(
        n15290) );
  NAND2_X1 U17022 ( .A1(n15288), .A2(n15561), .ZN(n15289) );
  OAI211_X1 U17023 ( .C1(n15291), .C2(n15558), .A(n15290), .B(n15289), .ZN(
        n15355) );
  MUX2_X1 U17024 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15355), .S(n15622), .Z(
        P1_U3547) );
  AOI211_X1 U17025 ( .C1(n15530), .C2(n15294), .A(n15293), .B(n15292), .ZN(
        n15295) );
  OAI21_X1 U17026 ( .B1(n15588), .B2(n15296), .A(n15295), .ZN(n15356) );
  MUX2_X1 U17027 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15356), .S(n15622), .Z(
        P1_U3546) );
  AOI21_X1 U17028 ( .B1(n15530), .B2(n15298), .A(n15297), .ZN(n15299) );
  OAI211_X1 U17029 ( .C1(n15301), .C2(n15588), .A(n15300), .B(n15299), .ZN(
        n15357) );
  MUX2_X1 U17030 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15357), .S(n15622), .Z(
        P1_U3545) );
  AOI22_X1 U17031 ( .A1(n15303), .A2(n15517), .B1(n15530), .B2(n15302), .ZN(
        n15304) );
  OAI211_X1 U17032 ( .C1(n15588), .C2(n15306), .A(n15305), .B(n15304), .ZN(
        n15358) );
  MUX2_X1 U17033 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15358), .S(n15622), .Z(
        P1_U3544) );
  AOI21_X1 U17034 ( .B1(n15530), .B2(n15308), .A(n15307), .ZN(n15309) );
  OAI211_X1 U17035 ( .C1(n15588), .C2(n15311), .A(n15310), .B(n15309), .ZN(
        n15359) );
  MUX2_X1 U17036 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15359), .S(n15622), .Z(
        P1_U3543) );
  AOI211_X1 U17037 ( .C1(n15530), .C2(n15314), .A(n15313), .B(n15312), .ZN(
        n15315) );
  OAI211_X1 U17038 ( .C1(n15588), .C2(n15317), .A(n15316), .B(n15315), .ZN(
        n15360) );
  MUX2_X1 U17039 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15360), .S(n15622), .Z(
        P1_U3542) );
  AOI21_X1 U17040 ( .B1(n15530), .B2(n15319), .A(n15318), .ZN(n15320) );
  OAI211_X1 U17041 ( .C1(n15588), .C2(n15322), .A(n15321), .B(n15320), .ZN(
        n15361) );
  MUX2_X1 U17042 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15361), .S(n15622), .Z(
        P1_U3541) );
  AND2_X1 U17043 ( .A1(n15323), .A2(n15561), .ZN(n15327) );
  OAI21_X1 U17044 ( .B1(n15325), .B2(n15599), .A(n15324), .ZN(n15326) );
  MUX2_X1 U17045 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n15362), .S(n15622), .Z(
        P1_U3540) );
  AOI211_X1 U17046 ( .C1(n15530), .C2(n15331), .A(n15330), .B(n15329), .ZN(
        n15332) );
  OAI21_X1 U17047 ( .B1(n15588), .B2(n15333), .A(n15332), .ZN(n15363) );
  MUX2_X1 U17048 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n15363), .S(n15622), .Z(
        P1_U3539) );
  AOI211_X1 U17049 ( .C1(n15530), .C2(n15336), .A(n15335), .B(n15334), .ZN(
        n15339) );
  NAND3_X1 U17050 ( .A1(n12015), .A2(n15552), .A3(n15337), .ZN(n15338) );
  OAI211_X1 U17051 ( .C1(n15340), .C2(n15588), .A(n15339), .B(n15338), .ZN(
        n15364) );
  MUX2_X1 U17052 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n15364), .S(n15622), .Z(
        P1_U3538) );
  MUX2_X1 U17053 ( .A(n15341), .B(P1_REG1_REG_0__SCAN_IN), .S(n15620), .Z(
        P1_U3528) );
  MUX2_X1 U17054 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15342), .S(n15608), .Z(
        P1_U3527) );
  MUX2_X1 U17055 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15343), .S(n15608), .Z(
        P1_U3526) );
  MUX2_X1 U17056 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15344), .S(n15608), .Z(
        P1_U3524) );
  MUX2_X1 U17057 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15345), .S(n15608), .Z(
        P1_U3523) );
  MUX2_X1 U17058 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15346), .S(n15608), .Z(
        P1_U3522) );
  MUX2_X1 U17059 ( .A(n15347), .B(P1_REG0_REG_25__SCAN_IN), .S(n15606), .Z(
        P1_U3521) );
  MUX2_X1 U17060 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15348), .S(n15608), .Z(
        P1_U3520) );
  MUX2_X1 U17061 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15349), .S(n15608), .Z(
        P1_U3519) );
  MUX2_X1 U17062 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15350), .S(n15608), .Z(
        P1_U3518) );
  MUX2_X1 U17063 ( .A(n15351), .B(P1_REG0_REG_21__SCAN_IN), .S(n15606), .Z(
        P1_U3517) );
  INV_X1 U17064 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n15353) );
  MUX2_X1 U17065 ( .A(n15353), .B(n15352), .S(n15608), .Z(n15354) );
  INV_X1 U17066 ( .A(n15354), .ZN(P1_U3516) );
  MUX2_X1 U17067 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15355), .S(n15608), .Z(
        P1_U3515) );
  MUX2_X1 U17068 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15356), .S(n15608), .Z(
        P1_U3513) );
  MUX2_X1 U17069 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15357), .S(n15608), .Z(
        P1_U3510) );
  MUX2_X1 U17070 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15358), .S(n15608), .Z(
        P1_U3507) );
  MUX2_X1 U17071 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15359), .S(n15608), .Z(
        P1_U3504) );
  MUX2_X1 U17072 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15360), .S(n15608), .Z(
        P1_U3501) );
  MUX2_X1 U17073 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n15361), .S(n15608), .Z(
        P1_U3498) );
  MUX2_X1 U17074 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n15362), .S(n15608), .Z(
        P1_U3495) );
  MUX2_X1 U17075 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n15363), .S(n15608), .Z(
        P1_U3492) );
  MUX2_X1 U17076 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n15364), .S(n15608), .Z(
        P1_U3489) );
  NOR4_X1 U17077 ( .A1(n15365), .A2(P1_IR_REG_30__SCAN_IN), .A3(n10221), .A4(
        P1_U3086), .ZN(n15366) );
  AOI21_X1 U17078 ( .B1(n15367), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15366), 
        .ZN(n15368) );
  OAI21_X1 U17079 ( .B1(n15369), .B2(n15379), .A(n15368), .ZN(P1_U3324) );
  OAI222_X1 U17080 ( .A1(n15379), .A2(n15373), .B1(P1_U3086), .B2(n15372), 
        .C1(n15371), .C2(n15370), .ZN(P1_U3325) );
  OAI222_X1 U17081 ( .A1(n15370), .A2(n15376), .B1(n15379), .B2(n15375), .C1(
        n15374), .C2(P1_U3086), .ZN(P1_U3326) );
  OAI222_X1 U17082 ( .A1(n15370), .A2(n15380), .B1(n15379), .B2(n15378), .C1(
        n6762), .C2(P1_U3086), .ZN(P1_U3328) );
  MUX2_X1 U17083 ( .A(n15382), .B(n15381), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  XOR2_X1 U17084 ( .A(n15384), .B(n15383), .Z(SUB_1596_U59) );
  XOR2_X1 U17085 ( .A(n15385), .B(n15386), .Z(SUB_1596_U57) );
  XOR2_X1 U17086 ( .A(n15387), .B(n15388), .Z(SUB_1596_U56) );
  INV_X1 U17087 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15389) );
  NAND2_X1 U17088 ( .A1(n15390), .A2(n15389), .ZN(n15392) );
  INV_X1 U17089 ( .A(n15401), .ZN(n15399) );
  NAND2_X1 U17090 ( .A1(n15394), .A2(n15393), .ZN(n15396) );
  NAND2_X1 U17091 ( .A1(n15396), .A2(n15395), .ZN(n15410) );
  XNOR2_X1 U17092 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n15397) );
  XNOR2_X1 U17093 ( .A(n15410), .B(n15397), .ZN(n15400) );
  INV_X1 U17094 ( .A(n15400), .ZN(n15398) );
  INV_X1 U17095 ( .A(n15407), .ZN(n15406) );
  INV_X1 U17096 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15402) );
  INV_X1 U17097 ( .A(n15403), .ZN(n15404) );
  OAI21_X1 U17098 ( .B1(n15404), .B2(n15406), .A(P2_ADDR_REG_14__SCAN_IN), 
        .ZN(n15405) );
  OAI21_X1 U17099 ( .B1(n15406), .B2(n15408), .A(n15405), .ZN(SUB_1596_U66) );
  AND2_X1 U17100 ( .A1(P3_ADDR_REG_14__SCAN_IN), .A2(n15906), .ZN(n15409) );
  NAND2_X1 U17101 ( .A1(n16031), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n15411) );
  NAND2_X1 U17102 ( .A1(n15412), .A2(n15411), .ZN(n15423) );
  INV_X1 U17103 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15490) );
  NAND2_X1 U17104 ( .A1(n15490), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n15424) );
  INV_X1 U17105 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15413) );
  NAND2_X1 U17106 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n15413), .ZN(n15421) );
  AND2_X1 U17107 ( .A1(n15424), .A2(n15421), .ZN(n15414) );
  XNOR2_X1 U17108 ( .A(n15423), .B(n15414), .ZN(n15415) );
  NAND2_X1 U17109 ( .A1(n15416), .A2(n15415), .ZN(n15420) );
  NAND2_X1 U17110 ( .A1(n15419), .A2(n15420), .ZN(n15417) );
  XNOR2_X1 U17111 ( .A(n15417), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  INV_X1 U17112 ( .A(n15421), .ZN(n15422) );
  NAND2_X1 U17113 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n15436), .ZN(n15426) );
  OAI21_X1 U17114 ( .B1(n15436), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n15426), 
        .ZN(n15427) );
  XNOR2_X1 U17115 ( .A(n15439), .B(n15427), .ZN(n15428) );
  INV_X1 U17116 ( .A(n15428), .ZN(n15429) );
  NAND2_X1 U17117 ( .A1(n15433), .A2(n15434), .ZN(n15431) );
  XNOR2_X1 U17118 ( .A(n15431), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  OR2_X1 U17119 ( .A1(n15436), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n15438) );
  AND2_X1 U17120 ( .A1(n15436), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n15437) );
  AOI21_X1 U17121 ( .B1(n15439), .B2(n15438), .A(n15437), .ZN(n15447) );
  INV_X1 U17122 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15440) );
  XNOR2_X1 U17123 ( .A(n15447), .B(n15440), .ZN(n15445) );
  XNOR2_X1 U17124 ( .A(n15445), .B(P3_ADDR_REG_17__SCAN_IN), .ZN(n15441) );
  NAND2_X1 U17125 ( .A1(n15444), .A2(n15443), .ZN(n15442) );
  XNOR2_X1 U17126 ( .A(n15442), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  INV_X1 U17127 ( .A(n15445), .ZN(n15446) );
  NAND2_X1 U17128 ( .A1(n15446), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n15449) );
  NAND2_X1 U17129 ( .A1(n15447), .A2(n15440), .ZN(n15448) );
  NAND2_X1 U17130 ( .A1(n15449), .A2(n15448), .ZN(n15459) );
  INV_X1 U17131 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15450) );
  XNOR2_X1 U17132 ( .A(n15450), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(n15457) );
  XNOR2_X1 U17133 ( .A(n15459), .B(n15457), .ZN(n15451) );
  AOI21_X1 U17134 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n15452), .A(n15456), 
        .ZN(n15453) );
  INV_X1 U17135 ( .A(n15453), .ZN(SUB_1596_U62) );
  INV_X1 U17136 ( .A(n15454), .ZN(n15455) );
  INV_X1 U17137 ( .A(n15457), .ZN(n15458) );
  INV_X1 U17138 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15833) );
  AOI22_X1 U17139 ( .A1(n15459), .A2(n15458), .B1(P3_ADDR_REG_18__SCAN_IN), 
        .B2(n15833), .ZN(n15462) );
  XNOR2_X1 U17140 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n15460) );
  XNOR2_X1 U17141 ( .A(n15460), .B(n7792), .ZN(n15461) );
  XNOR2_X1 U17142 ( .A(n15462), .B(n15461), .ZN(n15463) );
  XNOR2_X1 U17143 ( .A(n15464), .B(n15463), .ZN(SUB_1596_U4) );
  AOI21_X1 U17144 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15465) );
  OAI21_X1 U17145 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15465), 
        .ZN(U28) );
  AOI21_X1 U17146 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15466) );
  OAI21_X1 U17147 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15466), 
        .ZN(U29) );
  AND2_X1 U17148 ( .A1(n15468), .A2(n15467), .ZN(n15470) );
  XNOR2_X1 U17149 ( .A(n15470), .B(n15469), .ZN(SUB_1596_U61) );
  INV_X1 U17150 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n15472) );
  AOI21_X1 U17151 ( .B1(n6762), .B2(n15472), .A(n15471), .ZN(n15474) );
  XNOR2_X1 U17152 ( .A(n15474), .B(P1_IR_REG_0__SCAN_IN), .ZN(n15477) );
  AOI22_X1 U17153 ( .A1(n15475), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15476) );
  OAI21_X1 U17154 ( .B1(n15478), .B2(n15477), .A(n15476), .ZN(P1_U3243) );
  OAI21_X1 U17155 ( .B1(n15481), .B2(n15480), .A(n15479), .ZN(n15487) );
  XNOR2_X1 U17156 ( .A(n15482), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n15485) );
  AOI222_X1 U17157 ( .A1(n15487), .A2(n15812), .B1(n15486), .B2(n15485), .C1(
        n15484), .C2(n15483), .ZN(n15489) );
  OAI211_X1 U17158 ( .C1(n15490), .C2(n15821), .A(n15489), .B(n15488), .ZN(
        P1_U3258) );
  XNOR2_X1 U17159 ( .A(n15491), .B(n15494), .ZN(n15604) );
  INV_X1 U17160 ( .A(n6740), .ZN(n15492) );
  AOI21_X1 U17161 ( .B1(n15494), .B2(n15493), .A(n15492), .ZN(n15496) );
  OAI21_X1 U17162 ( .B1(n15496), .B2(n15558), .A(n15495), .ZN(n15497) );
  AOI21_X1 U17163 ( .B1(n15576), .B2(n15604), .A(n15497), .ZN(n15601) );
  AOI222_X1 U17164 ( .A1(n15499), .A2(n15515), .B1(P1_REG2_REG_9__SCAN_IN), 
        .B2(n15512), .C1(n15513), .C2(n15498), .ZN(n15505) );
  INV_X1 U17165 ( .A(n15500), .ZN(n15522) );
  OAI211_X1 U17166 ( .C1(n15502), .C2(n15600), .A(n15517), .B(n15501), .ZN(
        n15598) );
  INV_X1 U17167 ( .A(n15598), .ZN(n15503) );
  AOI22_X1 U17168 ( .A1(n15604), .A2(n15522), .B1(n15521), .B2(n15503), .ZN(
        n15504) );
  OAI211_X1 U17169 ( .C1(n15525), .C2(n15601), .A(n15505), .B(n15504), .ZN(
        P1_U3284) );
  XNOR2_X1 U17170 ( .A(n15506), .B(n15508), .ZN(n15586) );
  XNOR2_X1 U17171 ( .A(n15507), .B(n15508), .ZN(n15510) );
  OAI21_X1 U17172 ( .B1(n15510), .B2(n15558), .A(n15509), .ZN(n15511) );
  AOI21_X1 U17173 ( .B1(n15576), .B2(n15586), .A(n15511), .ZN(n15583) );
  AOI222_X1 U17174 ( .A1(n15516), .A2(n15515), .B1(n15514), .B2(n15513), .C1(
        P1_REG2_REG_7__SCAN_IN), .C2(n15512), .ZN(n15524) );
  OAI211_X1 U17175 ( .C1(n15582), .C2(n15519), .A(n15518), .B(n15517), .ZN(
        n15581) );
  INV_X1 U17176 ( .A(n15581), .ZN(n15520) );
  AOI22_X1 U17177 ( .A1(n15586), .A2(n15522), .B1(n15521), .B2(n15520), .ZN(
        n15523) );
  OAI211_X1 U17178 ( .C1(n15525), .C2(n15583), .A(n15524), .B(n15523), .ZN(
        P1_U3286) );
  INV_X1 U17179 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15957) );
  NOR2_X1 U17180 ( .A1(n15526), .A2(n15957), .ZN(P1_U3294) );
  AND2_X1 U17181 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15527), .ZN(P1_U3295) );
  AND2_X1 U17182 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15527), .ZN(P1_U3296) );
  AND2_X1 U17183 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15527), .ZN(P1_U3297) );
  AND2_X1 U17184 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15527), .ZN(P1_U3298) );
  AND2_X1 U17185 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15527), .ZN(P1_U3299) );
  AND2_X1 U17186 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15527), .ZN(P1_U3300) );
  AND2_X1 U17187 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15527), .ZN(P1_U3301) );
  AND2_X1 U17188 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15527), .ZN(P1_U3302) );
  NOR2_X1 U17189 ( .A1(n15526), .A2(n16034), .ZN(P1_U3303) );
  NOR2_X1 U17190 ( .A1(n15526), .A2(n15894), .ZN(P1_U3304) );
  AND2_X1 U17191 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15527), .ZN(P1_U3305) );
  AND2_X1 U17192 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15527), .ZN(P1_U3306) );
  INV_X1 U17193 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15975) );
  NOR2_X1 U17194 ( .A1(n15526), .A2(n15975), .ZN(P1_U3307) );
  NOR2_X1 U17195 ( .A1(n15526), .A2(n16084), .ZN(P1_U3308) );
  AND2_X1 U17196 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15527), .ZN(P1_U3309) );
  NOR2_X1 U17197 ( .A1(n15526), .A2(n15980), .ZN(P1_U3310) );
  NOR2_X1 U17198 ( .A1(n15526), .A2(n15893), .ZN(P1_U3311) );
  AND2_X1 U17199 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15527), .ZN(P1_U3312) );
  AND2_X1 U17200 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15527), .ZN(P1_U3313) );
  AND2_X1 U17201 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15527), .ZN(P1_U3314) );
  AND2_X1 U17202 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15527), .ZN(P1_U3315) );
  NOR2_X1 U17203 ( .A1(n15526), .A2(n16039), .ZN(P1_U3316) );
  AND2_X1 U17204 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15527), .ZN(P1_U3317) );
  AND2_X1 U17205 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15527), .ZN(P1_U3318) );
  AND2_X1 U17206 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15527), .ZN(P1_U3319) );
  AND2_X1 U17207 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15527), .ZN(P1_U3320) );
  AND2_X1 U17208 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15527), .ZN(P1_U3321) );
  AND2_X1 U17209 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15527), .ZN(P1_U3322) );
  AND2_X1 U17210 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15527), .ZN(P1_U3323) );
  INV_X1 U17211 ( .A(n15565), .ZN(n15605) );
  INV_X1 U17212 ( .A(n15528), .ZN(n15536) );
  INV_X1 U17213 ( .A(n15529), .ZN(n15532) );
  NAND2_X1 U17214 ( .A1(n10668), .A2(n15530), .ZN(n15531) );
  OAI211_X1 U17215 ( .C1(n15538), .C2(n15533), .A(n15532), .B(n15531), .ZN(
        n15535) );
  AOI211_X1 U17216 ( .C1(n15605), .C2(n15536), .A(n15535), .B(n15534), .ZN(
        n15609) );
  AOI22_X1 U17217 ( .A1(n15608), .A2(n15609), .B1(n10359), .B2(n15606), .ZN(
        P1_U3462) );
  OAI22_X1 U17218 ( .A1(n15539), .A2(n15538), .B1(n15537), .B2(n15599), .ZN(
        n15541) );
  AOI211_X1 U17219 ( .C1(n15605), .C2(n15542), .A(n15541), .B(n15540), .ZN(
        n15611) );
  INV_X1 U17220 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15543) );
  AOI22_X1 U17221 ( .A1(n15608), .A2(n15611), .B1(n15543), .B2(n15606), .ZN(
        P1_U3465) );
  INV_X1 U17222 ( .A(n15544), .ZN(n15547) );
  INV_X1 U17223 ( .A(n15545), .ZN(n15546) );
  OAI211_X1 U17224 ( .C1(n15548), .C2(n15599), .A(n15547), .B(n15546), .ZN(
        n15551) );
  AOI21_X1 U17225 ( .B1(n15566), .B2(n15565), .A(n15549), .ZN(n15550) );
  AOI211_X1 U17226 ( .C1(n15553), .C2(n15552), .A(n15551), .B(n15550), .ZN(
        n15612) );
  AOI22_X1 U17227 ( .A1(n15608), .A2(n15612), .B1(n10701), .B2(n15606), .ZN(
        P1_U3468) );
  NOR2_X1 U17228 ( .A1(n15555), .A2(n15554), .ZN(n15557) );
  OAI211_X1 U17229 ( .C1(n15559), .C2(n15558), .A(n15557), .B(n15556), .ZN(
        n15560) );
  AOI21_X1 U17230 ( .B1(n15562), .B2(n15561), .A(n15560), .ZN(n15614) );
  INV_X1 U17231 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15563) );
  AOI22_X1 U17232 ( .A1(n15608), .A2(n15614), .B1(n15563), .B2(n15606), .ZN(
        P1_U3471) );
  AOI21_X1 U17233 ( .B1(n15566), .B2(n15565), .A(n15564), .ZN(n15570) );
  NOR4_X1 U17234 ( .A1(n15570), .A2(n15569), .A3(n15568), .A4(n15567), .ZN(
        n15615) );
  INV_X1 U17235 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15571) );
  AOI22_X1 U17236 ( .A1(n15608), .A2(n15615), .B1(n15571), .B2(n15606), .ZN(
        P1_U3474) );
  OAI21_X1 U17237 ( .B1(n15573), .B2(n15599), .A(n15572), .ZN(n15574) );
  INV_X1 U17238 ( .A(n15574), .ZN(n15578) );
  OAI21_X1 U17239 ( .B1(n15576), .B2(n15605), .A(n15575), .ZN(n15577) );
  INV_X1 U17240 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15580) );
  AOI22_X1 U17241 ( .A1(n15608), .A2(n15616), .B1(n15580), .B2(n15606), .ZN(
        P1_U3477) );
  OAI21_X1 U17242 ( .B1(n15582), .B2(n15599), .A(n15581), .ZN(n15585) );
  INV_X1 U17243 ( .A(n15583), .ZN(n15584) );
  AOI211_X1 U17244 ( .C1(n15605), .C2(n15586), .A(n15585), .B(n15584), .ZN(
        n15618) );
  INV_X1 U17245 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15587) );
  AOI22_X1 U17246 ( .A1(n15608), .A2(n15618), .B1(n15587), .B2(n15606), .ZN(
        P1_U3480) );
  NOR2_X1 U17247 ( .A1(n15589), .A2(n15588), .ZN(n15594) );
  INV_X1 U17248 ( .A(n15590), .ZN(n15591) );
  OAI21_X1 U17249 ( .B1(n15592), .B2(n15599), .A(n15591), .ZN(n15593) );
  NOR4_X1 U17250 ( .A1(n15596), .A2(n15595), .A3(n15594), .A4(n15593), .ZN(
        n15619) );
  INV_X1 U17251 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15597) );
  AOI22_X1 U17252 ( .A1(n15608), .A2(n15619), .B1(n15597), .B2(n15606), .ZN(
        P1_U3483) );
  OAI21_X1 U17253 ( .B1(n15600), .B2(n15599), .A(n15598), .ZN(n15603) );
  INV_X1 U17254 ( .A(n15601), .ZN(n15602) );
  AOI211_X1 U17255 ( .C1(n15605), .C2(n15604), .A(n15603), .B(n15602), .ZN(
        n15621) );
  INV_X1 U17256 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15607) );
  AOI22_X1 U17257 ( .A1(n15608), .A2(n15621), .B1(n15607), .B2(n15606), .ZN(
        P1_U3486) );
  AOI22_X1 U17258 ( .A1(n15622), .A2(n15609), .B1(n15996), .B2(n15620), .ZN(
        P1_U3529) );
  AOI22_X1 U17259 ( .A1(n15622), .A2(n15611), .B1(n15610), .B2(n15620), .ZN(
        P1_U3530) );
  AOI22_X1 U17260 ( .A1(n15622), .A2(n15612), .B1(n16062), .B2(n15620), .ZN(
        P1_U3531) );
  AOI22_X1 U17261 ( .A1(n15622), .A2(n15614), .B1(n15613), .B2(n15620), .ZN(
        P1_U3532) );
  AOI22_X1 U17262 ( .A1(n15622), .A2(n15615), .B1(n7499), .B2(n15620), .ZN(
        P1_U3533) );
  INV_X1 U17263 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n16024) );
  AOI22_X1 U17264 ( .A1(n15622), .A2(n15616), .B1(n16024), .B2(n15620), .ZN(
        P1_U3534) );
  INV_X1 U17265 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n15617) );
  AOI22_X1 U17266 ( .A1(n15622), .A2(n15618), .B1(n15617), .B2(n15620), .ZN(
        P1_U3535) );
  AOI22_X1 U17267 ( .A1(n15622), .A2(n15619), .B1(n15824), .B2(n15620), .ZN(
        P1_U3536) );
  AOI22_X1 U17268 ( .A1(n15622), .A2(n15621), .B1(n10650), .B2(n15620), .ZN(
        P1_U3537) );
  NOR2_X1 U17269 ( .A1(n15629), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U17270 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15653), .B1(n15644), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n15628) );
  AOI22_X1 U17271 ( .A1(n15629), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n15627) );
  OAI22_X1 U17272 ( .A1(n15624), .A2(P2_REG1_REG_0__SCAN_IN), .B1(
        P2_REG2_REG_0__SCAN_IN), .B2(n15623), .ZN(n15625) );
  OAI21_X1 U17273 ( .B1(n15651), .B2(n15625), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n15626) );
  OAI211_X1 U17274 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n15628), .A(n15627), .B(
        n15626), .ZN(P2_U3214) );
  AOI22_X1 U17275 ( .A1(n15629), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n15641) );
  XOR2_X1 U17276 ( .A(n15631), .B(n15630), .Z(n15635) );
  AND2_X1 U17277 ( .A1(n8398), .A2(n15632), .ZN(n15634) );
  AOI22_X1 U17278 ( .A1(n15644), .A2(n15635), .B1(n15634), .B2(n15633), .ZN(
        n15640) );
  OAI211_X1 U17279 ( .C1(n15638), .C2(n15637), .A(n15653), .B(n15636), .ZN(
        n15639) );
  NAND3_X1 U17280 ( .A1(n15641), .A2(n15640), .A3(n15639), .ZN(P2_U3215) );
  INV_X1 U17281 ( .A(n15642), .ZN(n15650) );
  AND2_X1 U17282 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n15649) );
  OAI211_X1 U17283 ( .C1(n15646), .C2(n15645), .A(n15644), .B(n15643), .ZN(
        n15647) );
  INV_X1 U17284 ( .A(n15647), .ZN(n15648) );
  AOI211_X1 U17285 ( .C1(n15651), .C2(n15650), .A(n15649), .B(n15648), .ZN(
        n15657) );
  OAI211_X1 U17286 ( .C1(n15655), .C2(n15654), .A(n15653), .B(n15652), .ZN(
        n15656) );
  OAI211_X1 U17287 ( .C1(n15658), .C2(n16124), .A(n15657), .B(n15656), .ZN(
        P2_U3217) );
  NOR2_X1 U17288 ( .A1(n15660), .A2(n15659), .ZN(n15704) );
  INV_X1 U17289 ( .A(n15661), .ZN(n15705) );
  OAI21_X1 U17290 ( .B1(n15713), .B2(n15662), .A(n15705), .ZN(n15664) );
  NAND2_X1 U17291 ( .A1(n15664), .A2(n15663), .ZN(n15703) );
  AOI21_X1 U17292 ( .B1(n15704), .B2(n15665), .A(n15703), .ZN(n15669) );
  AOI22_X1 U17293 ( .A1(n15667), .A2(n15705), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n15666), .ZN(n15668) );
  OAI221_X1 U17294 ( .B1(n6557), .B2(n15669), .C1(n14285), .C2(n8447), .A(
        n15668), .ZN(P2_U3265) );
  NOR2_X1 U17295 ( .A1(n15696), .A2(n16091), .ZN(P2_U3266) );
  INV_X1 U17296 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15671) );
  NOR2_X1 U17297 ( .A1(n15696), .A2(n15671), .ZN(P2_U3267) );
  INV_X1 U17298 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15672) );
  NOR2_X1 U17299 ( .A1(n15696), .A2(n15672), .ZN(P2_U3268) );
  INV_X1 U17300 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15673) );
  NOR2_X1 U17301 ( .A1(n15696), .A2(n15673), .ZN(P2_U3269) );
  NOR2_X1 U17302 ( .A1(n15696), .A2(n15674), .ZN(P2_U3270) );
  NOR2_X1 U17303 ( .A1(n15694), .A2(n16004), .ZN(P2_U3271) );
  INV_X1 U17304 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n15675) );
  NOR2_X1 U17305 ( .A1(n15694), .A2(n15675), .ZN(P2_U3272) );
  INV_X1 U17306 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15676) );
  NOR2_X1 U17307 ( .A1(n15694), .A2(n15676), .ZN(P2_U3273) );
  INV_X1 U17308 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15677) );
  NOR2_X1 U17309 ( .A1(n15694), .A2(n15677), .ZN(P2_U3274) );
  INV_X1 U17310 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n15891) );
  NOR2_X1 U17311 ( .A1(n15694), .A2(n15891), .ZN(P2_U3275) );
  INV_X1 U17312 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n15678) );
  NOR2_X1 U17313 ( .A1(n15694), .A2(n15678), .ZN(P2_U3276) );
  INV_X1 U17314 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15679) );
  NOR2_X1 U17315 ( .A1(n15694), .A2(n15679), .ZN(P2_U3277) );
  INV_X1 U17316 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15680) );
  NOR2_X1 U17317 ( .A1(n15696), .A2(n15680), .ZN(P2_U3278) );
  INV_X1 U17318 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n15681) );
  NOR2_X1 U17319 ( .A1(n15696), .A2(n15681), .ZN(P2_U3279) );
  INV_X1 U17320 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15682) );
  NOR2_X1 U17321 ( .A1(n15696), .A2(n15682), .ZN(P2_U3280) );
  INV_X1 U17322 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15683) );
  NOR2_X1 U17323 ( .A1(n15696), .A2(n15683), .ZN(P2_U3281) );
  INV_X1 U17324 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15684) );
  NOR2_X1 U17325 ( .A1(n15696), .A2(n15684), .ZN(P2_U3282) );
  INV_X1 U17326 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15685) );
  NOR2_X1 U17327 ( .A1(n15696), .A2(n15685), .ZN(P2_U3283) );
  INV_X1 U17328 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n15686) );
  NOR2_X1 U17329 ( .A1(n15696), .A2(n15686), .ZN(P2_U3284) );
  INV_X1 U17330 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n15889) );
  NOR2_X1 U17331 ( .A1(n15696), .A2(n15889), .ZN(P2_U3285) );
  INV_X1 U17332 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n15687) );
  NOR2_X1 U17333 ( .A1(n15696), .A2(n15687), .ZN(P2_U3286) );
  INV_X1 U17334 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n15688) );
  NOR2_X1 U17335 ( .A1(n15696), .A2(n15688), .ZN(P2_U3287) );
  INV_X1 U17336 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n15689) );
  NOR2_X1 U17337 ( .A1(n15696), .A2(n15689), .ZN(P2_U3288) );
  NOR2_X1 U17338 ( .A1(n15696), .A2(n15936), .ZN(P2_U3289) );
  INV_X1 U17339 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n15690) );
  NOR2_X1 U17340 ( .A1(n15694), .A2(n15690), .ZN(P2_U3290) );
  INV_X1 U17341 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15691) );
  NOR2_X1 U17342 ( .A1(n15694), .A2(n15691), .ZN(P2_U3291) );
  INV_X1 U17343 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n15692) );
  NOR2_X1 U17344 ( .A1(n15694), .A2(n15692), .ZN(P2_U3292) );
  INV_X1 U17345 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n15693) );
  NOR2_X1 U17346 ( .A1(n15694), .A2(n15693), .ZN(P2_U3293) );
  NOR2_X1 U17347 ( .A1(n15696), .A2(n15983), .ZN(P2_U3294) );
  INV_X1 U17348 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n15695) );
  NOR2_X1 U17349 ( .A1(n15696), .A2(n15695), .ZN(P2_U3295) );
  OAI21_X1 U17350 ( .B1(n15702), .B2(n15698), .A(n15697), .ZN(P2_U3416) );
  AOI22_X1 U17351 ( .A1(n15702), .A2(n15701), .B1(n15700), .B2(n15699), .ZN(
        P2_U3417) );
  AOI211_X1 U17352 ( .C1(n15705), .C2(n15733), .A(n15704), .B(n15703), .ZN(
        n15744) );
  AOI22_X1 U17353 ( .A1(n15743), .A2(n15744), .B1(n8444), .B2(n15741), .ZN(
        P2_U3430) );
  OAI21_X1 U17354 ( .B1(n15737), .B2(n15707), .A(n15706), .ZN(n15711) );
  INV_X1 U17355 ( .A(n15712), .ZN(n15709) );
  OAI21_X1 U17356 ( .B1(n15709), .B2(n15716), .A(n15708), .ZN(n15710) );
  AOI211_X1 U17357 ( .C1(n15713), .C2(n15712), .A(n15711), .B(n15710), .ZN(
        n15745) );
  AOI22_X1 U17358 ( .A1(n15743), .A2(n15745), .B1(n8439), .B2(n15741), .ZN(
        P2_U3433) );
  AOI21_X1 U17359 ( .B1(n15716), .B2(n15715), .A(n15714), .ZN(n15721) );
  NOR2_X1 U17360 ( .A1(n15737), .A2(n15717), .ZN(n15719) );
  NOR4_X1 U17361 ( .A1(n15721), .A2(n15720), .A3(n15719), .A4(n15718), .ZN(
        n15746) );
  INV_X1 U17362 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15722) );
  AOI22_X1 U17363 ( .A1(n15743), .A2(n15746), .B1(n15722), .B2(n15741), .ZN(
        P2_U3439) );
  OAI211_X1 U17364 ( .C1(n8148), .C2(n15737), .A(n15724), .B(n15723), .ZN(
        n15725) );
  AOI21_X1 U17365 ( .B1(n15726), .B2(n15740), .A(n15725), .ZN(n15747) );
  AOI22_X1 U17366 ( .A1(n15743), .A2(n15747), .B1(n8476), .B2(n15741), .ZN(
        P2_U3445) );
  INV_X1 U17367 ( .A(n15727), .ZN(n15732) );
  INV_X1 U17368 ( .A(n15728), .ZN(n15729) );
  OAI21_X1 U17369 ( .B1(n6823), .B2(n15737), .A(n15729), .ZN(n15731) );
  AOI211_X1 U17370 ( .C1(n15733), .C2(n15732), .A(n15731), .B(n15730), .ZN(
        n15748) );
  INV_X1 U17371 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15734) );
  AOI22_X1 U17372 ( .A1(n15743), .A2(n15748), .B1(n15734), .B2(n15741), .ZN(
        P2_U3448) );
  OAI211_X1 U17373 ( .C1(n7511), .C2(n15737), .A(n15736), .B(n15735), .ZN(
        n15738) );
  AOI21_X1 U17374 ( .B1(n15740), .B2(n15739), .A(n15738), .ZN(n15749) );
  INV_X1 U17375 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15742) );
  AOI22_X1 U17376 ( .A1(n15743), .A2(n15749), .B1(n15742), .B2(n15741), .ZN(
        P2_U3451) );
  AOI22_X1 U17377 ( .A1(n15750), .A2(n15744), .B1(n8445), .B2(n12591), .ZN(
        P2_U3499) );
  AOI22_X1 U17378 ( .A1(n15750), .A2(n15745), .B1(n10415), .B2(n12591), .ZN(
        P2_U3500) );
  AOI22_X1 U17379 ( .A1(n15750), .A2(n15746), .B1(n10417), .B2(n12591), .ZN(
        P2_U3502) );
  AOI22_X1 U17380 ( .A1(n15750), .A2(n15747), .B1(n8480), .B2(n12591), .ZN(
        P2_U3504) );
  AOI22_X1 U17381 ( .A1(n15750), .A2(n15748), .B1(n8491), .B2(n12591), .ZN(
        P2_U3505) );
  AOI22_X1 U17382 ( .A1(n15750), .A2(n15749), .B1(n8502), .B2(n12591), .ZN(
        P2_U3506) );
  NOR2_X1 U17383 ( .A1(P3_U3897), .A2(n15751), .ZN(P3_U3150) );
  AOI211_X1 U17384 ( .C1(n15755), .C2(n15754), .A(n15753), .B(n15752), .ZN(
        n15790) );
  AOI22_X1 U17385 ( .A1(n15788), .A2(n9168), .B1(n15790), .B2(n15786), .ZN(
        P3_U3393) );
  INV_X1 U17386 ( .A(n15756), .ZN(n15760) );
  INV_X1 U17387 ( .A(n15757), .ZN(n15759) );
  AOI211_X1 U17388 ( .C1(n15760), .C2(n15784), .A(n15759), .B(n15758), .ZN(
        n15792) );
  AOI22_X1 U17389 ( .A1(n15788), .A2(n9146), .B1(n15792), .B2(n15786), .ZN(
        P3_U3396) );
  INV_X1 U17390 ( .A(n15761), .ZN(n15762) );
  AOI211_X1 U17391 ( .C1(n15764), .C2(n15784), .A(n15763), .B(n15762), .ZN(
        n15794) );
  AOI22_X1 U17392 ( .A1(n15788), .A2(n9176), .B1(n15794), .B2(n15786), .ZN(
        P3_U3399) );
  INV_X1 U17393 ( .A(n15765), .ZN(n15767) );
  AOI211_X1 U17394 ( .C1(n15768), .C2(n15784), .A(n15767), .B(n15766), .ZN(
        n15796) );
  AOI22_X1 U17395 ( .A1(n15788), .A2(n9191), .B1(n15796), .B2(n15786), .ZN(
        P3_U3402) );
  INV_X1 U17396 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15775) );
  OAI22_X1 U17397 ( .A1(n15772), .A2(n15771), .B1(n15770), .B2(n15769), .ZN(
        n15773) );
  NOR2_X1 U17398 ( .A1(n15774), .A2(n15773), .ZN(n15798) );
  AOI22_X1 U17399 ( .A1(n15788), .A2(n15775), .B1(n15798), .B2(n15786), .ZN(
        P3_U3405) );
  INV_X1 U17400 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15780) );
  INV_X1 U17401 ( .A(n15776), .ZN(n15777) );
  AOI211_X1 U17402 ( .C1(n15779), .C2(n15784), .A(n15778), .B(n15777), .ZN(
        n15800) );
  AOI22_X1 U17403 ( .A1(n15788), .A2(n15780), .B1(n15800), .B2(n15786), .ZN(
        P3_U3408) );
  INV_X1 U17404 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15787) );
  INV_X1 U17405 ( .A(n15781), .ZN(n15782) );
  AOI211_X1 U17406 ( .C1(n15785), .C2(n15784), .A(n15783), .B(n15782), .ZN(
        n15803) );
  AOI22_X1 U17407 ( .A1(n15788), .A2(n15787), .B1(n15803), .B2(n15786), .ZN(
        P3_U3411) );
  AOI22_X1 U17408 ( .A1(n15804), .A2(n15790), .B1(n15789), .B2(n15801), .ZN(
        P3_U3460) );
  AOI22_X1 U17409 ( .A1(n15804), .A2(n15792), .B1(n15791), .B2(n15801), .ZN(
        P3_U3461) );
  AOI22_X1 U17410 ( .A1(n15804), .A2(n15794), .B1(n15793), .B2(n15801), .ZN(
        P3_U3462) );
  AOI22_X1 U17411 ( .A1(n15804), .A2(n15796), .B1(n15795), .B2(n15801), .ZN(
        P3_U3463) );
  AOI22_X1 U17412 ( .A1(n15804), .A2(n15798), .B1(n15797), .B2(n15801), .ZN(
        P3_U3464) );
  AOI22_X1 U17413 ( .A1(n15804), .A2(n15800), .B1(n15799), .B2(n15801), .ZN(
        P3_U3465) );
  AOI22_X1 U17414 ( .A1(n15804), .A2(n15803), .B1(n15802), .B2(n15801), .ZN(
        P3_U3466) );
  INV_X1 U17415 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n16058) );
  NAND2_X1 U17416 ( .A1(n15809), .A2(n15808), .ZN(n15811) );
  NAND2_X1 U17417 ( .A1(n15816), .A2(n15812), .ZN(n15813) );
  NAND4_X1 U17418 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(P1_REG1_REG_6__SCAN_IN), 
        .A3(P1_REG1_REG_0__SCAN_IN), .A4(P1_REG1_REG_1__SCAN_IN), .ZN(n15822)
         );
  OR3_X1 U17419 ( .A1(n15822), .A2(P2_REG2_REG_24__SCAN_IN), .A3(
        P3_REG1_REG_27__SCAN_IN), .ZN(n15831) );
  NAND4_X1 U17420 ( .A1(n7645), .A2(n16060), .A3(P3_REG0_REG_18__SCAN_IN), 
        .A4(P3_IR_REG_22__SCAN_IN), .ZN(n15829) );
  NAND4_X1 U17421 ( .A1(n15824), .A2(n15823), .A3(P1_IR_REG_17__SCAN_IN), .A4(
        P1_IR_REG_26__SCAN_IN), .ZN(n15828) );
  NOR4_X1 U17422 ( .A1(P3_REG2_REG_23__SCAN_IN), .A2(n16077), .A3(n16075), 
        .A4(n16071), .ZN(n15825) );
  NAND4_X1 U17423 ( .A1(n15826), .A2(n15825), .A3(P1_ADDR_REG_7__SCAN_IN), 
        .A4(P1_REG2_REG_14__SCAN_IN), .ZN(n15827) );
  OR4_X1 U17424 ( .A1(n15829), .A2(n15828), .A3(n15827), .A4(
        P3_DATAO_REG_31__SCAN_IN), .ZN(n15830) );
  NOR4_X1 U17425 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P1_REG1_REG_18__SCAN_IN), 
        .A3(n15831), .A4(n15830), .ZN(n15870) );
  NOR4_X1 U17426 ( .A1(SI_27_), .A2(P3_REG2_REG_5__SCAN_IN), .A3(
        P2_REG0_REG_1__SCAN_IN), .A4(n15926), .ZN(n15832) );
  NAND3_X1 U17427 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P1_REG3_REG_2__SCAN_IN), 
        .A3(n15832), .ZN(n15844) );
  NAND4_X1 U17428 ( .A1(n15964), .A2(SI_0_), .A3(P2_REG3_REG_26__SCAN_IN), 
        .A4(P2_REG0_REG_18__SCAN_IN), .ZN(n15834) );
  NOR3_X1 U17429 ( .A1(n15834), .A2(P3_DATAO_REG_30__SCAN_IN), .A3(n15833), 
        .ZN(n15842) );
  NAND4_X1 U17430 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(
        P3_DATAO_REG_14__SCAN_IN), .A3(n15955), .A4(n15954), .ZN(n15840) );
  NAND4_X1 U17431 ( .A1(P1_REG3_REG_21__SCAN_IN), .A2(P3_DATAO_REG_28__SCAN_IN), .A3(n8035), .A4(n15835), .ZN(n15839) );
  NAND4_X1 U17432 ( .A1(n15837), .A2(P1_D_REG_15__SCAN_IN), .A3(n15836), .A4(
        n15981), .ZN(n15838) );
  NOR4_X1 U17433 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(n15840), .A3(n15839), .A4(
        n15838), .ZN(n15841) );
  NAND4_X1 U17434 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(P2_REG3_REG_0__SCAN_IN), 
        .A3(n15842), .A4(n15841), .ZN(n15843) );
  NOR4_X1 U17435 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n15938), .A3(n15844), 
        .A4(n15843), .ZN(n15869) );
  NAND4_X1 U17436 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(P3_REG2_REG_28__SCAN_IN), .A3(SI_8_), .A4(P2_REG2_REG_26__SCAN_IN), .ZN(n15867) );
  NAND4_X1 U17437 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(P2_REG1_REG_5__SCAN_IN), 
        .A3(P1_D_REG_17__SCAN_IN), .A4(n15845), .ZN(n15866) );
  NAND4_X1 U17438 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(P1_REG3_REG_11__SCAN_IN), 
        .A3(P1_REG0_REG_18__SCAN_IN), .A4(n16097), .ZN(n15846) );
  NOR3_X1 U17439 ( .A1(SI_10_), .A2(P1_ADDR_REG_8__SCAN_IN), .A3(n15846), .ZN(
        n15852) );
  NAND4_X1 U17440 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(P1_REG1_REG_20__SCAN_IN), .A3(n7390), .A4(n16017), .ZN(n15850) );
  NAND4_X1 U17441 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P1_REG3_REG_0__SCAN_IN), 
        .A3(n16010), .A4(n16012), .ZN(n15849) );
  NAND4_X1 U17442 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P2_DATAO_REG_17__SCAN_IN), 
        .A3(P2_DATAO_REG_15__SCAN_IN), .A4(P1_REG0_REG_3__SCAN_IN), .ZN(n15848) );
  NAND4_X1 U17443 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(n15999), .A3(n16000), 
        .A4(n15997), .ZN(n15847) );
  NOR4_X1 U17444 ( .A1(n15850), .A2(n15849), .A3(n15848), .A4(n15847), .ZN(
        n15851) );
  NAND4_X1 U17445 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(P2_REG1_REG_27__SCAN_IN), 
        .A3(n15852), .A4(n15851), .ZN(n15865) );
  INV_X1 U17446 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n15874) );
  NOR4_X1 U17447 ( .A1(P3_REG0_REG_13__SCAN_IN), .A2(P1_DATAO_REG_16__SCAN_IN), 
        .A3(n15874), .A4(n15876), .ZN(n15856) );
  NOR4_X1 U17448 ( .A1(n16023), .A2(n15877), .A3(n15879), .A4(n15880), .ZN(
        n15855) );
  NOR4_X1 U17449 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P3_DATAO_REG_25__SCAN_IN), 
        .A3(n15918), .A4(n15924), .ZN(n15854) );
  NOR4_X1 U17450 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P1_REG1_REG_27__SCAN_IN), 
        .A3(P1_REG1_REG_25__SCAN_IN), .A4(P1_ADDR_REG_14__SCAN_IN), .ZN(n15853) );
  NAND4_X1 U17451 ( .A1(n15856), .A2(n15855), .A3(n15854), .A4(n15853), .ZN(
        n15860) );
  NOR4_X1 U17452 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .A3(P3_ADDR_REG_14__SCAN_IN), .A4(P3_DATAO_REG_29__SCAN_IN), .ZN(
        n15857) );
  NAND3_X1 U17453 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P2_REG2_REG_1__SCAN_IN), 
        .A3(n15857), .ZN(n15859) );
  NAND4_X1 U17454 ( .A1(n16040), .A2(P2_DATAO_REG_4__SCAN_IN), .A3(
        P3_REG1_REG_12__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n15858) );
  NOR3_X1 U17455 ( .A1(n15860), .A2(n15859), .A3(n15858), .ZN(n15863) );
  INV_X1 U17456 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n15897) );
  NAND4_X1 U17457 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), 
        .A3(P3_DATAO_REG_9__SCAN_IN), .A4(n15897), .ZN(n15861) );
  NOR3_X1 U17458 ( .A1(P3_DATAO_REG_3__SCAN_IN), .A2(n15910), .A3(n15861), 
        .ZN(n15862) );
  NAND2_X1 U17459 ( .A1(n15863), .A2(n15862), .ZN(n15864) );
  NOR4_X1 U17460 ( .A1(n15867), .A2(n15866), .A3(n15865), .A4(n15864), .ZN(
        n15868) );
  NAND4_X1 U17461 ( .A1(n15871), .A2(n15870), .A3(n15869), .A4(n15868), .ZN(
        n16118) );
  AOI22_X1 U17462 ( .A1(n15874), .A2(keyinput17), .B1(keyinput44), .B2(n15873), 
        .ZN(n15872) );
  OAI221_X1 U17463 ( .B1(n15874), .B2(keyinput17), .C1(n15873), .C2(keyinput44), .A(n15872), .ZN(n15886) );
  AOI22_X1 U17464 ( .A1(n15877), .A2(keyinput95), .B1(keyinput52), .B2(n15876), 
        .ZN(n15875) );
  OAI221_X1 U17465 ( .B1(n15877), .B2(keyinput95), .C1(n15876), .C2(keyinput52), .A(n15875), .ZN(n15885) );
  AOI22_X1 U17466 ( .A1(n15880), .A2(keyinput84), .B1(n15879), .B2(keyinput18), 
        .ZN(n15878) );
  OAI221_X1 U17467 ( .B1(n15880), .B2(keyinput84), .C1(n15879), .C2(keyinput18), .A(n15878), .ZN(n15884) );
  XNOR2_X1 U17468 ( .A(P1_REG1_REG_18__SCAN_IN), .B(keyinput59), .ZN(n15882)
         );
  XNOR2_X1 U17469 ( .A(P1_REG1_REG_0__SCAN_IN), .B(keyinput8), .ZN(n15881) );
  NAND2_X1 U17470 ( .A1(n15882), .A2(n15881), .ZN(n15883) );
  NOR4_X1 U17471 ( .A1(n15886), .A2(n15885), .A3(n15884), .A4(n15883), .ZN(
        n15934) );
  AOI22_X1 U17472 ( .A1(n15889), .A2(keyinput116), .B1(n15888), .B2(keyinput35), .ZN(n15887) );
  OAI221_X1 U17473 ( .B1(n15889), .B2(keyinput116), .C1(n15888), .C2(
        keyinput35), .A(n15887), .ZN(n15901) );
  AOI22_X1 U17474 ( .A1(n15824), .A2(keyinput120), .B1(n15891), .B2(keyinput77), .ZN(n15890) );
  OAI221_X1 U17475 ( .B1(n15824), .B2(keyinput120), .C1(n15891), .C2(
        keyinput77), .A(n15890), .ZN(n15900) );
  AOI22_X1 U17476 ( .A1(n15894), .A2(keyinput122), .B1(keyinput104), .B2(
        n15893), .ZN(n15892) );
  OAI221_X1 U17477 ( .B1(n15894), .B2(keyinput122), .C1(n15893), .C2(
        keyinput104), .A(n15892), .ZN(n15899) );
  AOI22_X1 U17478 ( .A1(n15897), .A2(keyinput91), .B1(keyinput108), .B2(n15896), .ZN(n15895) );
  OAI221_X1 U17479 ( .B1(n15897), .B2(keyinput91), .C1(n15896), .C2(
        keyinput108), .A(n15895), .ZN(n15898) );
  NOR4_X1 U17480 ( .A1(n15901), .A2(n15900), .A3(n15899), .A4(n15898), .ZN(
        n15933) );
  AOI22_X1 U17481 ( .A1(n15904), .A2(keyinput88), .B1(keyinput79), .B2(n15903), 
        .ZN(n15902) );
  OAI221_X1 U17482 ( .B1(n15904), .B2(keyinput88), .C1(n15903), .C2(keyinput79), .A(n15902), .ZN(n15916) );
  AOI22_X1 U17483 ( .A1(n15907), .A2(keyinput13), .B1(keyinput92), .B2(n15906), 
        .ZN(n15905) );
  OAI221_X1 U17484 ( .B1(n15907), .B2(keyinput13), .C1(n15906), .C2(keyinput92), .A(n15905), .ZN(n15915) );
  AOI22_X1 U17485 ( .A1(n15910), .A2(keyinput89), .B1(keyinput1), .B2(n15909), 
        .ZN(n15908) );
  OAI221_X1 U17486 ( .B1(n15910), .B2(keyinput89), .C1(n15909), .C2(keyinput1), 
        .A(n15908), .ZN(n15914) );
  XNOR2_X1 U17487 ( .A(P3_IR_REG_15__SCAN_IN), .B(keyinput110), .ZN(n15912) );
  XNOR2_X1 U17488 ( .A(P1_REG1_REG_27__SCAN_IN), .B(keyinput68), .ZN(n15911)
         );
  NAND2_X1 U17489 ( .A1(n15912), .A2(n15911), .ZN(n15913) );
  NOR4_X1 U17490 ( .A1(n15916), .A2(n15915), .A3(n15914), .A4(n15913), .ZN(
        n15932) );
  AOI22_X1 U17491 ( .A1(n15919), .A2(keyinput61), .B1(n15918), .B2(keyinput4), 
        .ZN(n15917) );
  OAI221_X1 U17492 ( .B1(n15919), .B2(keyinput61), .C1(n15918), .C2(keyinput4), 
        .A(n15917), .ZN(n15930) );
  AOI22_X1 U17493 ( .A1(n15922), .A2(keyinput42), .B1(keyinput90), .B2(n15921), 
        .ZN(n15920) );
  OAI221_X1 U17494 ( .B1(n15922), .B2(keyinput42), .C1(n15921), .C2(keyinput90), .A(n15920), .ZN(n15929) );
  AOI22_X1 U17495 ( .A1(n15924), .A2(keyinput53), .B1(keyinput87), .B2(n8439), 
        .ZN(n15923) );
  OAI221_X1 U17496 ( .B1(n15924), .B2(keyinput53), .C1(n8439), .C2(keyinput87), 
        .A(n15923), .ZN(n15928) );
  AOI22_X1 U17497 ( .A1(n15926), .A2(keyinput72), .B1(n13722), .B2(keyinput118), .ZN(n15925) );
  OAI221_X1 U17498 ( .B1(n15926), .B2(keyinput72), .C1(n13722), .C2(
        keyinput118), .A(n15925), .ZN(n15927) );
  NOR4_X1 U17499 ( .A1(n15930), .A2(n15929), .A3(n15928), .A4(n15927), .ZN(
        n15931) );
  NAND4_X1 U17500 ( .A1(n15934), .A2(n15933), .A3(n15932), .A4(n15931), .ZN(
        n16116) );
  AOI22_X1 U17501 ( .A1(n15191), .A2(keyinput98), .B1(n15936), .B2(keyinput119), .ZN(n15935) );
  OAI221_X1 U17502 ( .B1(n15191), .B2(keyinput98), .C1(n15936), .C2(
        keyinput119), .A(n15935), .ZN(n15947) );
  AOI22_X1 U17503 ( .A1(n15939), .A2(keyinput37), .B1(keyinput11), .B2(n15938), 
        .ZN(n15937) );
  OAI221_X1 U17504 ( .B1(n15939), .B2(keyinput37), .C1(n15938), .C2(keyinput11), .A(n15937), .ZN(n15946) );
  XOR2_X1 U17505 ( .A(n15940), .B(keyinput5), .Z(n15944) );
  XNOR2_X1 U17506 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput56), .ZN(n15943)
         );
  XNOR2_X1 U17507 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(keyinput22), .ZN(n15942)
         );
  XNOR2_X1 U17508 ( .A(P3_IR_REG_26__SCAN_IN), .B(keyinput10), .ZN(n15941) );
  NAND4_X1 U17509 ( .A1(n15944), .A2(n15943), .A3(n15942), .A4(n15941), .ZN(
        n15945) );
  NOR3_X1 U17510 ( .A1(n15947), .A2(n15946), .A3(n15945), .ZN(n15994) );
  AOI22_X1 U17511 ( .A1(n15950), .A2(keyinput33), .B1(n15949), .B2(keyinput50), 
        .ZN(n15948) );
  OAI221_X1 U17512 ( .B1(n15950), .B2(keyinput33), .C1(n15949), .C2(keyinput50), .A(n15948), .ZN(n15962) );
  AOI22_X1 U17513 ( .A1(n8035), .A2(keyinput66), .B1(keyinput30), .B2(n15952), 
        .ZN(n15951) );
  OAI221_X1 U17514 ( .B1(n8035), .B2(keyinput66), .C1(n15952), .C2(keyinput30), 
        .A(n15951), .ZN(n15961) );
  AOI22_X1 U17515 ( .A1(n15955), .A2(keyinput64), .B1(keyinput83), .B2(n15954), 
        .ZN(n15953) );
  OAI221_X1 U17516 ( .B1(n15955), .B2(keyinput64), .C1(n15954), .C2(keyinput83), .A(n15953), .ZN(n15960) );
  AOI22_X1 U17517 ( .A1(n15958), .A2(keyinput15), .B1(keyinput96), .B2(n15957), 
        .ZN(n15956) );
  OAI221_X1 U17518 ( .B1(n15958), .B2(keyinput15), .C1(n15957), .C2(keyinput96), .A(n15956), .ZN(n15959) );
  NOR4_X1 U17519 ( .A1(n15962), .A2(n15961), .A3(n15960), .A4(n15959), .ZN(
        n15993) );
  XNOR2_X1 U17520 ( .A(n15963), .B(keyinput58), .ZN(n15968) );
  XNOR2_X1 U17521 ( .A(n15964), .B(keyinput34), .ZN(n15967) );
  XNOR2_X1 U17522 ( .A(n15965), .B(keyinput117), .ZN(n15966) );
  NOR3_X1 U17523 ( .A1(n15968), .A2(n15967), .A3(n15966), .ZN(n15971) );
  XNOR2_X1 U17524 ( .A(SI_0_), .B(keyinput60), .ZN(n15970) );
  XNOR2_X1 U17525 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(keyinput126), .ZN(n15969)
         );
  NAND3_X1 U17526 ( .A1(n15971), .A2(n15970), .A3(n15969), .ZN(n15978) );
  INV_X1 U17527 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n15974) );
  AOI22_X1 U17528 ( .A1(n15974), .A2(keyinput49), .B1(keyinput29), .B2(n15973), 
        .ZN(n15972) );
  OAI221_X1 U17529 ( .B1(n15974), .B2(keyinput49), .C1(n15973), .C2(keyinput29), .A(n15972), .ZN(n15977) );
  XNOR2_X1 U17530 ( .A(n15975), .B(keyinput57), .ZN(n15976) );
  NOR3_X1 U17531 ( .A1(n15978), .A2(n15977), .A3(n15976), .ZN(n15992) );
  AOI22_X1 U17532 ( .A1(n15981), .A2(keyinput106), .B1(n15980), .B2(keyinput86), .ZN(n15979) );
  OAI221_X1 U17533 ( .B1(n15981), .B2(keyinput106), .C1(n15980), .C2(
        keyinput86), .A(n15979), .ZN(n15990) );
  AOI22_X1 U17534 ( .A1(n15983), .A2(keyinput62), .B1(keyinput69), .B2(n8391), 
        .ZN(n15982) );
  OAI221_X1 U17535 ( .B1(n15983), .B2(keyinput62), .C1(n8391), .C2(keyinput69), 
        .A(n15982), .ZN(n15989) );
  XNOR2_X1 U17536 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput9), .ZN(n15987) );
  XNOR2_X1 U17537 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput113), .ZN(n15986)
         );
  XNOR2_X1 U17538 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput94), .ZN(n15985) );
  XNOR2_X1 U17539 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(keyinput47), .ZN(n15984)
         );
  NAND4_X1 U17540 ( .A1(n15987), .A2(n15986), .A3(n15985), .A4(n15984), .ZN(
        n15988) );
  NOR3_X1 U17541 ( .A1(n15990), .A2(n15989), .A3(n15988), .ZN(n15991) );
  NAND4_X1 U17542 ( .A1(n15994), .A2(n15993), .A3(n15992), .A4(n15991), .ZN(
        n16115) );
  AOI22_X1 U17543 ( .A1(n15997), .A2(keyinput6), .B1(n15996), .B2(keyinput70), 
        .ZN(n15995) );
  OAI221_X1 U17544 ( .B1(n15997), .B2(keyinput6), .C1(n15996), .C2(keyinput70), 
        .A(n15995), .ZN(n16008) );
  AOI22_X1 U17545 ( .A1(n16000), .A2(keyinput100), .B1(keyinput3), .B2(n15999), 
        .ZN(n15998) );
  OAI221_X1 U17546 ( .B1(n16000), .B2(keyinput100), .C1(n15999), .C2(keyinput3), .A(n15998), .ZN(n16007) );
  AOI22_X1 U17547 ( .A1(n10701), .A2(keyinput46), .B1(keyinput28), .B2(n7645), 
        .ZN(n16001) );
  OAI221_X1 U17548 ( .B1(n10701), .B2(keyinput46), .C1(n7645), .C2(keyinput28), 
        .A(n16001), .ZN(n16006) );
  AOI22_X1 U17549 ( .A1(n16004), .A2(keyinput20), .B1(n16003), .B2(keyinput36), 
        .ZN(n16002) );
  OAI221_X1 U17550 ( .B1(n16004), .B2(keyinput20), .C1(n16003), .C2(keyinput36), .A(n16002), .ZN(n16005) );
  NOR4_X1 U17551 ( .A1(n16008), .A2(n16007), .A3(n16006), .A4(n16005), .ZN(
        n16055) );
  AOI22_X1 U17552 ( .A1(n16010), .A2(keyinput43), .B1(n7662), .B2(keyinput54), 
        .ZN(n16009) );
  OAI221_X1 U17553 ( .B1(n16010), .B2(keyinput43), .C1(n7662), .C2(keyinput54), 
        .A(n16009), .ZN(n16021) );
  AOI22_X1 U17554 ( .A1(n16012), .A2(keyinput80), .B1(n11315), .B2(keyinput31), 
        .ZN(n16011) );
  OAI221_X1 U17555 ( .B1(n16012), .B2(keyinput80), .C1(n11315), .C2(keyinput31), .A(n16011), .ZN(n16020) );
  AOI22_X1 U17556 ( .A1(n7390), .A2(keyinput124), .B1(keyinput2), .B2(n16014), 
        .ZN(n16013) );
  OAI221_X1 U17557 ( .B1(n7390), .B2(keyinput124), .C1(n16014), .C2(keyinput2), 
        .A(n16013), .ZN(n16019) );
  AOI22_X1 U17558 ( .A1(n16017), .A2(keyinput23), .B1(n16016), .B2(keyinput45), 
        .ZN(n16015) );
  OAI221_X1 U17559 ( .B1(n16017), .B2(keyinput23), .C1(n16016), .C2(keyinput45), .A(n16015), .ZN(n16018) );
  NOR4_X1 U17560 ( .A1(n16021), .A2(n16020), .A3(n16019), .A4(n16018), .ZN(
        n16054) );
  AOI22_X1 U17561 ( .A1(n16024), .A2(keyinput65), .B1(n16023), .B2(keyinput41), 
        .ZN(n16022) );
  OAI221_X1 U17562 ( .B1(n16024), .B2(keyinput65), .C1(n16023), .C2(keyinput41), .A(n16022), .ZN(n16029) );
  XNOR2_X1 U17563 ( .A(n16025), .B(keyinput21), .ZN(n16028) );
  XNOR2_X1 U17564 ( .A(n16026), .B(keyinput0), .ZN(n16027) );
  OR3_X1 U17565 ( .A1(n16029), .A2(n16028), .A3(n16027), .ZN(n16037) );
  AOI22_X1 U17566 ( .A1(n16031), .A2(keyinput16), .B1(n15440), .B2(keyinput26), 
        .ZN(n16030) );
  OAI221_X1 U17567 ( .B1(n16031), .B2(keyinput16), .C1(n15440), .C2(keyinput26), .A(n16030), .ZN(n16036) );
  AOI22_X1 U17568 ( .A1(n16034), .A2(keyinput127), .B1(n16033), .B2(keyinput32), .ZN(n16032) );
  OAI221_X1 U17569 ( .B1(n16034), .B2(keyinput127), .C1(n16033), .C2(
        keyinput32), .A(n16032), .ZN(n16035) );
  NOR3_X1 U17570 ( .A1(n16037), .A2(n16036), .A3(n16035), .ZN(n16053) );
  AOI22_X1 U17571 ( .A1(n16040), .A2(keyinput12), .B1(n16039), .B2(keyinput121), .ZN(n16038) );
  OAI221_X1 U17572 ( .B1(n16040), .B2(keyinput12), .C1(n16039), .C2(
        keyinput121), .A(n16038), .ZN(n16051) );
  AOI22_X1 U17573 ( .A1(n16043), .A2(keyinput74), .B1(keyinput111), .B2(n16042), .ZN(n16041) );
  OAI221_X1 U17574 ( .B1(n16043), .B2(keyinput74), .C1(n16042), .C2(
        keyinput111), .A(n16041), .ZN(n16050) );
  XNOR2_X1 U17575 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput81), .ZN(n16046)
         );
  XNOR2_X1 U17576 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput55), .ZN(n16045) );
  XNOR2_X1 U17577 ( .A(keyinput97), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n16044) );
  NAND3_X1 U17578 ( .A1(n16046), .A2(n16045), .A3(n16044), .ZN(n16049) );
  XNOR2_X1 U17579 ( .A(n16047), .B(keyinput24), .ZN(n16048) );
  NOR4_X1 U17580 ( .A1(n16051), .A2(n16050), .A3(n16049), .A4(n16048), .ZN(
        n16052) );
  NAND4_X1 U17581 ( .A1(n16055), .A2(n16054), .A3(n16053), .A4(n16052), .ZN(
        n16114) );
  AOI22_X1 U17582 ( .A1(n16058), .A2(keyinput93), .B1(keyinput112), .B2(n16057), .ZN(n16056) );
  OAI221_X1 U17583 ( .B1(n16058), .B2(keyinput93), .C1(n16057), .C2(
        keyinput112), .A(n16056), .ZN(n16069) );
  AOI22_X1 U17584 ( .A1(n16061), .A2(keyinput123), .B1(n16060), .B2(keyinput7), 
        .ZN(n16059) );
  OAI221_X1 U17585 ( .B1(n16061), .B2(keyinput123), .C1(n16060), .C2(keyinput7), .A(n16059), .ZN(n16068) );
  XOR2_X1 U17586 ( .A(n16062), .B(keyinput107), .Z(n16066) );
  XNOR2_X1 U17587 ( .A(P3_IR_REG_22__SCAN_IN), .B(keyinput115), .ZN(n16065) );
  XNOR2_X1 U17588 ( .A(SI_10_), .B(keyinput99), .ZN(n16064) );
  XNOR2_X1 U17589 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(keyinput51), .ZN(n16063) );
  NAND4_X1 U17590 ( .A1(n16066), .A2(n16065), .A3(n16064), .A4(n16063), .ZN(
        n16067) );
  NOR3_X1 U17591 ( .A1(n16069), .A2(n16068), .A3(n16067), .ZN(n16112) );
  AOI22_X1 U17592 ( .A1(keyinput102), .A2(n16071), .B1(keyinput67), .B2(n16119), .ZN(n16070) );
  OAI21_X1 U17593 ( .B1(n16071), .B2(keyinput102), .A(n16070), .ZN(n16082) );
  AOI22_X1 U17594 ( .A1(n8658), .A2(keyinput101), .B1(n16073), .B2(keyinput78), 
        .ZN(n16072) );
  OAI221_X1 U17595 ( .B1(n8658), .B2(keyinput101), .C1(n16073), .C2(keyinput78), .A(n16072), .ZN(n16081) );
  AOI22_X1 U17596 ( .A1(n10616), .A2(keyinput25), .B1(n16075), .B2(keyinput14), 
        .ZN(n16074) );
  OAI221_X1 U17597 ( .B1(n10616), .B2(keyinput25), .C1(n16075), .C2(keyinput14), .A(n16074), .ZN(n16080) );
  INV_X1 U17598 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n16078) );
  AOI22_X1 U17599 ( .A1(n16078), .A2(keyinput105), .B1(n16077), .B2(keyinput82), .ZN(n16076) );
  OAI221_X1 U17600 ( .B1(n16078), .B2(keyinput105), .C1(n16077), .C2(
        keyinput82), .A(n16076), .ZN(n16079) );
  NOR4_X1 U17601 ( .A1(n16082), .A2(n16081), .A3(n16080), .A4(n16079), .ZN(
        n16111) );
  AOI22_X1 U17602 ( .A1(n8480), .A2(keyinput109), .B1(keyinput48), .B2(n16084), 
        .ZN(n16083) );
  OAI221_X1 U17603 ( .B1(n8480), .B2(keyinput109), .C1(n16084), .C2(keyinput48), .A(n16083), .ZN(n16095) );
  AOI22_X1 U17604 ( .A1(n16086), .A2(keyinput103), .B1(n14131), .B2(keyinput76), .ZN(n16085) );
  OAI221_X1 U17605 ( .B1(n16086), .B2(keyinput103), .C1(n14131), .C2(
        keyinput76), .A(n16085), .ZN(n16094) );
  INV_X1 U17606 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n16087) );
  XOR2_X1 U17607 ( .A(n16087), .B(keyinput125), .Z(n16090) );
  XNOR2_X1 U17608 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(keyinput73), .ZN(n16089)
         );
  XNOR2_X1 U17609 ( .A(SI_8_), .B(keyinput38), .ZN(n16088) );
  NAND3_X1 U17610 ( .A1(n16090), .A2(n16089), .A3(n16088), .ZN(n16093) );
  XNOR2_X1 U17611 ( .A(n16091), .B(keyinput63), .ZN(n16092) );
  NOR4_X1 U17612 ( .A1(n16095), .A2(n16094), .A3(n16093), .A4(n16092), .ZN(
        n16110) );
  AOI22_X1 U17613 ( .A1(n16098), .A2(keyinput27), .B1(n16097), .B2(keyinput39), 
        .ZN(n16096) );
  OAI221_X1 U17614 ( .B1(n16098), .B2(keyinput27), .C1(n16097), .C2(keyinput39), .A(n16096), .ZN(n16108) );
  AOI22_X1 U17615 ( .A1(n16101), .A2(keyinput75), .B1(n16100), .B2(keyinput40), 
        .ZN(n16099) );
  OAI221_X1 U17616 ( .B1(n16101), .B2(keyinput75), .C1(n16100), .C2(keyinput40), .A(n16099), .ZN(n16107) );
  XNOR2_X1 U17617 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput71), .ZN(n16105) );
  XNOR2_X1 U17618 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput114), .ZN(n16104)
         );
  XNOR2_X1 U17619 ( .A(P2_REG1_REG_13__SCAN_IN), .B(keyinput19), .ZN(n16103)
         );
  XNOR2_X1 U17620 ( .A(P1_REG3_REG_11__SCAN_IN), .B(keyinput85), .ZN(n16102)
         );
  NAND4_X1 U17621 ( .A1(n16105), .A2(n16104), .A3(n16103), .A4(n16102), .ZN(
        n16106) );
  NOR3_X1 U17622 ( .A1(n16108), .A2(n16107), .A3(n16106), .ZN(n16109) );
  NAND4_X1 U17623 ( .A1(n16112), .A2(n16111), .A3(n16110), .A4(n16109), .ZN(
        n16113) );
  NOR4_X1 U17624 ( .A1(n16116), .A2(n16115), .A3(n16114), .A4(n16113), .ZN(
        n16117) );
  OAI221_X1 U17625 ( .B1(n16119), .B2(keyinput67), .C1(n16119), .C2(n16118), 
        .A(n16117), .ZN(n16120) );
  XNOR2_X1 U17626 ( .A(n16121), .B(n16120), .ZN(P1_U3262) );
  AND2_X1 U17627 ( .A1(n16122), .A2(n16123), .ZN(n16125) );
  XNOR2_X1 U17628 ( .A(n16125), .B(n16124), .ZN(SUB_1596_U60) );
  XOR2_X1 U17629 ( .A(n16127), .B(n16126), .Z(SUB_1596_U5) );
  CLKBUF_X1 U7309 ( .A(n10022), .Z(n6556) );
  CLKBUF_X2 U7311 ( .A(n8455), .Z(n8944) );
  CLKBUF_X1 U7321 ( .A(n8921), .Z(n8961) );
  INV_X1 U7329 ( .A(n8395), .ZN(n8437) );
  OAI22_X1 U7371 ( .A1(n14254), .A2(n8719), .B1(n14260), .B2(n13940), .ZN(
        n14241) );
  CLKBUF_X1 U7382 ( .A(n10910), .Z(n12572) );
  AND2_X2 U7417 ( .A1(n12328), .A2(n10052), .ZN(n11018) );
  OR2_X1 U7616 ( .A1(n10223), .A2(n10221), .ZN(n10222) );
  INV_X1 U9154 ( .A(n9131), .ZN(n13714) );
  AND3_X1 U10090 ( .A1(n9170), .A2(n9169), .A3(n9171), .ZN(n16132) );
  CLKBUF_X1 U10128 ( .A(n15694), .Z(n15696) );
endmodule

