

module b21_C_gen_AntiSAT_k_128_4 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, 
        keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, 
        keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, 
        keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, 
        keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, 
        keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, 
        keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, 
        keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, 
        keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, 
        keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, 
        keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, 
        keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, 
        keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128;

  INV_X4 U4817 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  CLKBUF_X1 U4818 ( .A(n5058), .Z(n7604) );
  OR2_X1 U4819 ( .A1(n5095), .A2(n5096), .ZN(n5097) );
  CLKBUF_X1 U4820 ( .A(n5743), .Z(n4317) );
  BUF_X2 U4821 ( .A(n5356), .Z(n5132) );
  CLKBUF_X1 U4822 ( .A(n5743), .Z(n4316) );
  CLKBUF_X2 U4823 ( .A(n4710), .Z(n7589) );
  INV_X4 U4824 ( .A(n9968), .ZN(n9944) );
  INV_X1 U4825 ( .A(n9266), .ZN(n4313) );
  INV_X1 U4827 ( .A(n7797), .ZN(n7791) );
  XNOR2_X1 U4828 ( .A(n8183), .B(n5132), .ZN(n5096) );
  INV_X1 U4830 ( .A(n5806), .ZN(n5962) );
  INV_X1 U4831 ( .A(n7584), .ZN(n6326) );
  AND2_X1 U4832 ( .A1(n8154), .A2(n8694), .ZN(n5416) );
  NAND2_X1 U4833 ( .A1(n8113), .A2(n7284), .ZN(n9982) );
  AND2_X1 U4834 ( .A1(n5646), .A2(n5648), .ZN(n6035) );
  NAND2_X1 U4835 ( .A1(n9268), .A2(n5645), .ZN(n5746) );
  NAND2_X1 U4836 ( .A1(n7368), .A2(n7367), .ZN(n9626) );
  INV_X1 U4837 ( .A(n5733), .ZN(n5718) );
  INV_X1 U4838 ( .A(n7027), .ZN(n9835) );
  INV_X1 U4839 ( .A(n5416), .ZN(n7584) );
  INV_X1 U4840 ( .A(n5575), .ZN(n9962) );
  OR2_X1 U4841 ( .A1(n4936), .A2(n4933), .ZN(n4935) );
  NAND2_X2 U4842 ( .A1(n6256), .A2(n6355), .ZN(n6275) );
  AND2_X1 U4843 ( .A1(n5161), .A2(n5160), .ZN(n10011) );
  AND2_X2 U4844 ( .A1(n9612), .A2(n9611), .ZN(n9614) );
  OR2_X2 U4845 ( .A1(n4963), .A2(n9982), .ZN(n5058) );
  CLKBUF_X2 U4846 ( .A(n4337), .Z(n4315) );
  AND2_X2 U4847 ( .A1(n7130), .A2(n10005), .ZN(n7169) );
  NAND4_X2 U4848 ( .A1(n5652), .A2(n5651), .A3(n5650), .A4(n5649), .ZN(n8827)
         );
  OAI211_X2 U4849 ( .C1(n4465), .C2(n4466), .A(n4463), .B(n5188), .ZN(n4998)
         );
  OAI22_X2 U4850 ( .A1(n9138), .A2(n4835), .B1(n4343), .B2(n4837), .ZN(n9093)
         );
  OAI21_X2 U4851 ( .B1(n7354), .B2(n4818), .A(n4816), .ZN(n7458) );
  OR2_X1 U4852 ( .A1(n6292), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9266) );
  AOI21_X2 U4853 ( .B1(n9003), .B2(n4349), .A(n4847), .ZN(n8965) );
  NAND2_X1 U4854 ( .A1(n5648), .A2(n5645), .ZN(n5743) );
  INV_X1 U4855 ( .A(n5678), .ZN(n4318) );
  AND2_X1 U4856 ( .A1(n5696), .A2(n5660), .ZN(n5678) );
  XNOR2_X2 U4857 ( .A(n5422), .B(n5413), .ZN(n8130) );
  NAND2_X2 U4858 ( .A1(n4722), .A2(n4724), .ZN(n5422) );
  AND2_X1 U4859 ( .A1(n5696), .A2(n5660), .ZN(n4319) );
  NAND2_X1 U4861 ( .A1(n7533), .A2(n4723), .ZN(n4730) );
  NAND2_X1 U4862 ( .A1(n6181), .A2(n6180), .ZN(n9172) );
  NAND2_X1 U4863 ( .A1(n6160), .A2(n6159), .ZN(n9175) );
  INV_X1 U4864 ( .A(n4502), .ZN(n4321) );
  INV_X1 U4865 ( .A(n9015), .ZN(n8982) );
  NAND2_X1 U4866 ( .A1(n4777), .A2(n4778), .ZN(n8119) );
  INV_X1 U4867 ( .A(n9957), .ZN(n9912) );
  INV_X1 U4868 ( .A(n8750), .ZN(n9842) );
  INV_X1 U4869 ( .A(n6842), .ZN(n6633) );
  NAND2_X2 U4870 ( .A1(n6466), .A2(n7589), .ZN(n7594) );
  NAND2_X1 U4871 ( .A1(n8240), .A2(n8241), .ZN(n8158) );
  NAND2_X1 U4872 ( .A1(n6099), .A2(n6098), .ZN(n8782) );
  XNOR2_X1 U4873 ( .A(n7571), .B(n7570), .ZN(n8692) );
  XNOR2_X1 U4874 ( .A(n7562), .B(n7561), .ZN(n9271) );
  AOI21_X1 U4875 ( .B1(n4481), .B2(n4480), .A(n4479), .ZN(n8454) );
  NAND2_X1 U4876 ( .A1(n5523), .A2(n5522), .ZN(n7562) );
  NAND2_X1 U4877 ( .A1(n4747), .A2(n4749), .ZN(n7450) );
  NAND2_X1 U4878 ( .A1(n5521), .A2(n5520), .ZN(n5523) );
  NAND2_X1 U4879 ( .A1(n4904), .A2(n4902), .ZN(n8515) );
  OR2_X1 U4880 ( .A1(n5939), .A2(n5938), .ZN(n7540) );
  NAND2_X1 U4881 ( .A1(n4498), .A2(n4495), .ZN(n5939) );
  NAND2_X1 U4882 ( .A1(n7350), .A2(n7349), .ZN(n7397) );
  NAND2_X1 U4883 ( .A1(n7311), .A2(n7618), .ZN(n7350) );
  NAND2_X1 U4884 ( .A1(n4772), .A2(n4506), .ZN(n4502) );
  NAND2_X1 U4885 ( .A1(n5376), .A2(n5375), .ZN(n8638) );
  AND2_X1 U4886 ( .A1(n5903), .A2(n5879), .ZN(n4772) );
  NAND2_X1 U4887 ( .A1(n7069), .A2(n5204), .ZN(n7065) );
  NAND2_X1 U4888 ( .A1(n5332), .A2(n5331), .ZN(n8656) );
  NAND2_X1 U4889 ( .A1(n5926), .A2(n5925), .ZN(n9232) );
  NAND2_X1 U4890 ( .A1(n6804), .A2(n5151), .ZN(n6807) );
  NAND2_X1 U4891 ( .A1(n5283), .A2(n5282), .ZN(n9536) );
  NAND2_X1 U4892 ( .A1(n5887), .A2(n5886), .ZN(n9237) );
  NAND2_X1 U4893 ( .A1(n5846), .A2(n5845), .ZN(n9522) );
  OR2_X1 U4894 ( .A1(n7035), .A2(n7034), .ZN(n7898) );
  NAND2_X1 U4895 ( .A1(n5178), .A2(n5177), .ZN(n10017) );
  AND2_X1 U4896 ( .A1(n6661), .A2(n5666), .ZN(n5680) );
  NAND2_X1 U4897 ( .A1(n5079), .A2(n5083), .ZN(n4400) );
  AND2_X1 U4898 ( .A1(n7668), .A2(n7650), .ZN(n7664) );
  NAND2_X1 U4899 ( .A1(n4784), .A2(n4981), .ZN(n5142) );
  AND2_X1 U4900 ( .A1(n5662), .A2(n5661), .ZN(n6663) );
  AND4_X1 U4901 ( .A1(n5103), .A2(n5102), .A3(n5101), .A4(n5100), .ZN(n9917)
         );
  AND4_X1 U4902 ( .A1(n5088), .A2(n5087), .A3(n5086), .A4(n5085), .ZN(n6796)
         );
  AND4_X1 U4903 ( .A1(n5053), .A2(n5052), .A3(n5051), .A4(n5050), .ZN(n4913)
         );
  NAND2_X1 U4904 ( .A1(n4534), .A2(n5674), .ZN(n7835) );
  CLKBUF_X3 U4905 ( .A(n4325), .Z(n7580) );
  INV_X1 U4906 ( .A(n7594), .ZN(n5353) );
  NAND2_X1 U4907 ( .A1(n4912), .A2(n4712), .ZN(n8187) );
  NAND2_X1 U4908 ( .A1(n6223), .A2(n5624), .ZN(n6354) );
  AND2_X1 U4909 ( .A1(n5646), .A2(n9268), .ZN(n6085) );
  NAND2_X2 U4910 ( .A1(n4941), .A2(n4940), .ZN(n5098) );
  INV_X1 U4911 ( .A(n8113), .ZN(n7815) );
  INV_X1 U4912 ( .A(n7284), .ZN(n7643) );
  XNOR2_X1 U4913 ( .A(n4761), .B(n4760), .ZN(n7284) );
  NAND2_X1 U4914 ( .A1(n6275), .A2(n7589), .ZN(n5806) );
  NAND2_X1 U4915 ( .A1(n4956), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4955) );
  CLKBUF_X1 U4916 ( .A(n6256), .Z(n9711) );
  NAND2_X1 U4917 ( .A1(n8688), .A2(n4939), .ZN(n8694) );
  NAND2_X1 U4918 ( .A1(n5623), .A2(n5622), .ZN(n7528) );
  XNOR2_X1 U4919 ( .A(n4935), .B(n4934), .ZN(n8154) );
  XNOR2_X1 U4920 ( .A(n5643), .B(n5642), .ZN(n9268) );
  AND2_X1 U4921 ( .A1(n5543), .A2(n4883), .ZN(n5038) );
  XNOR2_X1 U4922 ( .A(n5042), .B(n5041), .ZN(n8701) );
  OAI21_X1 U4923 ( .B1(n6292), .B2(n4422), .A(n4421), .ZN(n4420) );
  OAI21_X1 U4924 ( .B1(n5628), .B2(n5630), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4533) );
  AND2_X1 U4925 ( .A1(n5618), .A2(n4822), .ZN(n5639) );
  INV_X1 U4926 ( .A(n5725), .ZN(n5597) );
  NOR2_X1 U4927 ( .A1(n4930), .A2(n4929), .ZN(n4931) );
  AND2_X1 U4928 ( .A1(n5596), .A2(n4860), .ZN(n4859) );
  AND4_X1 U4929 ( .A1(n5600), .A2(n5599), .A3(n5790), .A4(n5598), .ZN(n5601)
         );
  AND2_X1 U4930 ( .A1(n5612), .A2(n5615), .ZN(n4531) );
  NAND2_X1 U4931 ( .A1(n4783), .A2(n5615), .ZN(n4782) );
  NOR2_X1 U4932 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n4927) );
  NOR2_X1 U4933 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5599) );
  INV_X1 U4934 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5541) );
  NOR2_X1 U4935 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5595) );
  INV_X2 U4936 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4937 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4954) );
  INV_X1 U4938 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5225) );
  INV_X1 U4939 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5654) );
  INV_X1 U4940 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5941) );
  INV_X1 U4941 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4919) );
  INV_X1 U4942 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4957) );
  INV_X1 U4943 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5158) );
  INV_X1 U4944 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5279) );
  NOR2_X1 U4945 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4920) );
  INV_X1 U4946 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5315) );
  INV_X1 U4947 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5538) );
  AND2_X1 U4948 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9500) );
  INV_X1 U4949 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5210) );
  INV_X1 U4950 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4760) );
  NOR2_X2 U4951 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9501) );
  AND2_X2 U4952 ( .A1(n4402), .A2(n4401), .ZN(n8240) );
  OR2_X2 U4953 ( .A1(n8142), .A2(n5534), .ZN(n5082) );
  NAND2_X1 U4954 ( .A1(n4962), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4761) );
  XNOR2_X1 U4955 ( .A(n5082), .B(n5080), .ZN(n8188) );
  NAND2_X2 U4956 ( .A1(n7065), .A2(n7066), .ZN(n6985) );
  OAI21_X2 U4957 ( .B1(n9143), .B2(n9598), .A(n8911), .ZN(n9138) );
  INV_X4 U4958 ( .A(n5098), .ZN(n5084) );
  AND2_X1 U4959 ( .A1(n4941), .A2(n8694), .ZN(n4337) );
  NOR2_X2 U4960 ( .A1(n5329), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n5044) );
  NAND2_X1 U4962 ( .A1(n8188), .A2(n8189), .ZN(n8233) );
  NOR2_X4 U4963 ( .A1(n8577), .A2(n10027), .ZN(n9949) );
  OR2_X2 U4964 ( .A1(n8579), .A2(n10017), .ZN(n8577) );
  AOI21_X2 U4965 ( .B1(n7514), .B2(n5342), .A(n7513), .ZN(n7515) );
  NOR2_X1 U4966 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5613) );
  NOR2_X1 U4967 ( .A1(n4486), .A2(n8487), .ZN(n4485) );
  INV_X1 U4968 ( .A(n4488), .ZN(n4486) );
  NAND2_X1 U4969 ( .A1(n5370), .A2(n5369), .ZN(n5387) );
  NAND2_X1 U4970 ( .A1(n4648), .A2(n4647), .ZN(n5370) );
  AND2_X1 U4971 ( .A1(n5368), .A2(n5349), .ZN(n4647) );
  NOR2_X1 U4972 ( .A1(n4645), .A2(n4465), .ZN(n4464) );
  AND2_X1 U4973 ( .A1(n4642), .A2(n4467), .ZN(n4466) );
  INV_X1 U4974 ( .A(n5170), .ZN(n4467) );
  INV_X1 U4975 ( .A(n4645), .ZN(n4644) );
  OAI21_X1 U4976 ( .B1(n5141), .B2(n4646), .A(n5156), .ZN(n4645) );
  OR2_X1 U4977 ( .A1(n4341), .A2(n4903), .ZN(n4902) );
  INV_X1 U4978 ( .A(n4908), .ZN(n4903) );
  INV_X1 U4979 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U4980 ( .A1(n4988), .A2(n9364), .ZN(n4991) );
  NAND2_X1 U4981 ( .A1(n5460), .A2(n5459), .ZN(n5476) );
  NOR2_X1 U4982 ( .A1(n8367), .A2(n4579), .ZN(n4578) );
  INV_X1 U4983 ( .A(n7771), .ZN(n4579) );
  OR2_X1 U4984 ( .A1(n4809), .A2(n8389), .ZN(n4323) );
  INV_X1 U4985 ( .A(n4810), .ZN(n4809) );
  OR2_X1 U4986 ( .A1(n8617), .A2(n8392), .ZN(n7767) );
  OR2_X1 U4987 ( .A1(n8660), .A2(n8520), .ZN(n7731) );
  NOR2_X1 U4988 ( .A1(n7716), .A2(n4874), .ZN(n4873) );
  INV_X1 U4989 ( .A(n7396), .ZN(n4874) );
  NAND2_X1 U4990 ( .A1(n6633), .A2(n8231), .ZN(n7659) );
  NAND3_X1 U4991 ( .A1(n4497), .A2(n4500), .A3(n4496), .ZN(n4495) );
  NAND2_X1 U4992 ( .A1(n7335), .A2(n4499), .ZN(n4498) );
  NAND2_X1 U4993 ( .A1(n4501), .A2(n7438), .ZN(n4500) );
  OR3_X1 U4994 ( .A1(n9172), .A2(n9175), .A3(n9166), .ZN(n4583) );
  OR2_X1 U4995 ( .A1(n9172), .A2(n8927), .ZN(n8947) );
  NAND2_X1 U4996 ( .A1(n9175), .A2(n9015), .ZN(n4853) );
  NAND2_X1 U4997 ( .A1(n9180), .A2(n9025), .ZN(n8031) );
  OR2_X1 U4998 ( .A1(n9180), .A2(n9025), .ZN(n8943) );
  OR2_X1 U4999 ( .A1(n9237), .A2(n7370), .ZN(n7911) );
  AND2_X1 U5000 ( .A1(n5613), .A2(n4823), .ZN(n4530) );
  NAND2_X1 U5001 ( .A1(n5444), .A2(n5443), .ZN(n5461) );
  NAND2_X1 U5002 ( .A1(n4628), .A2(n4626), .ZN(n5444) );
  AOI21_X1 U5003 ( .B1(n4629), .B2(n4385), .A(n4627), .ZN(n4626) );
  AND2_X1 U5004 ( .A1(n5388), .A2(n5374), .ZN(n5386) );
  NAND2_X1 U5005 ( .A1(n5347), .A2(n5346), .ZN(n4648) );
  AND2_X1 U5006 ( .A1(n5032), .A2(n5031), .ZN(n5297) );
  AND2_X1 U5007 ( .A1(n5018), .A2(n5017), .ZN(n5261) );
  AND2_X1 U5008 ( .A1(n4637), .A2(n5007), .ZN(n4636) );
  AND2_X1 U5009 ( .A1(n5004), .A2(n5003), .ZN(n5208) );
  AND2_X1 U5010 ( .A1(n4997), .A2(n4996), .ZN(n5188) );
  INV_X1 U5011 ( .A(n4991), .ZN(n4465) );
  AOI21_X1 U5012 ( .B1(n4644), .B2(n4646), .A(n4372), .ZN(n4642) );
  NAND2_X1 U5013 ( .A1(n5057), .A2(n4614), .ZN(n4613) );
  INV_X1 U5014 ( .A(n5625), .ZN(n4615) );
  INV_X1 U5015 ( .A(n5488), .ZN(n5487) );
  NOR2_X1 U5016 ( .A1(n5250), .A2(n9374), .ZN(n5284) );
  AND2_X1 U5017 ( .A1(n7808), .A2(n7809), .ZN(n7810) );
  NAND2_X1 U5018 ( .A1(n8375), .A2(n8393), .ZN(n4901) );
  OR2_X1 U5019 ( .A1(n8403), .A2(n4458), .ZN(n4457) );
  NOR2_X1 U5020 ( .A1(n8617), .A2(n4459), .ZN(n4458) );
  NAND2_X1 U5021 ( .A1(n4377), .A2(n4493), .ZN(n4488) );
  AOI21_X1 U5022 ( .B1(n4909), .B2(n4910), .A(n4368), .ZN(n4907) );
  INV_X1 U5023 ( .A(n6466), .ZN(n6338) );
  AND2_X1 U5024 ( .A1(n6339), .A2(n5591), .ZN(n8478) );
  AND2_X1 U5025 ( .A1(n6080), .A2(n6094), .ZN(n4774) );
  XNOR2_X1 U5026 ( .A(n9162), .B(n8974), .ZN(n8950) );
  NOR3_X1 U5027 ( .A1(n9004), .A2(n9172), .A3(n9175), .ZN(n8983) );
  NAND2_X1 U5028 ( .A1(n8947), .A2(n7980), .ZN(n8978) );
  XNOR2_X1 U5029 ( .A(n9187), .B(n8923), .ZN(n9023) );
  NOR2_X1 U5030 ( .A1(n9192), .A2(n8919), .ZN(n8921) );
  OR2_X1 U5031 ( .A1(n9084), .A2(n9069), .ZN(n4914) );
  INV_X1 U5032 ( .A(n7877), .ZN(n6030) );
  INV_X1 U5033 ( .A(n6275), .ZN(n6029) );
  AND2_X1 U5034 ( .A1(n6685), .A2(n6684), .ZN(n9643) );
  INV_X1 U5035 ( .A(n9583), .ZN(n9638) );
  XNOR2_X1 U5036 ( .A(n4985), .B(SI_7_), .ZN(n5156) );
  NAND2_X1 U5037 ( .A1(n4428), .A2(n7881), .ZN(n4427) );
  NAND2_X1 U5038 ( .A1(n4407), .A2(n4406), .ZN(n4405) );
  INV_X1 U5039 ( .A(n7676), .ZN(n4406) );
  NAND2_X1 U5040 ( .A1(n7677), .A2(n7678), .ZN(n4407) );
  OAI211_X1 U5041 ( .C1(n7921), .C2(n7920), .A(n7919), .B(n7918), .ZN(n4444)
         );
  NAND2_X1 U5042 ( .A1(n7912), .A2(n7911), .ZN(n4442) );
  NOR2_X1 U5043 ( .A1(n7940), .A2(n7995), .ZN(n4453) );
  NAND2_X1 U5044 ( .A1(n7934), .A2(n4438), .ZN(n7932) );
  NOR2_X1 U5045 ( .A1(n4440), .A2(n4439), .ZN(n4438) );
  OAI21_X1 U5046 ( .B1(n7939), .B2(n7988), .A(n4842), .ZN(n4454) );
  MUX2_X1 U5047 ( .A(n7891), .B(n7890), .S(n7988), .Z(n7969) );
  NAND2_X1 U5048 ( .A1(n7969), .A2(n4434), .ZN(n4433) );
  INV_X1 U5049 ( .A(n8926), .ZN(n4434) );
  NAND2_X1 U5050 ( .A1(n4436), .A2(n7969), .ZN(n4435) );
  INV_X1 U5051 ( .A(n8978), .ZN(n4436) );
  INV_X1 U5052 ( .A(n4687), .ZN(n4680) );
  INV_X1 U5053 ( .A(n7919), .ZN(n4679) );
  NAND2_X1 U5054 ( .A1(n7799), .A2(n7788), .ZN(n7790) );
  NOR2_X1 U5055 ( .A1(n4321), .A2(n4501), .ZN(n4499) );
  AND2_X1 U5056 ( .A1(n7985), .A2(n7984), .ZN(n7993) );
  NOR2_X1 U5057 ( .A1(n4431), .A2(n4437), .ZN(n4430) );
  NAND2_X1 U5058 ( .A1(n8978), .A2(n4849), .ZN(n4848) );
  INV_X1 U5059 ( .A(n4850), .ZN(n4849) );
  OR2_X1 U5060 ( .A1(n9202), .A2(n9197), .ZN(n4590) );
  NOR2_X1 U5061 ( .A1(n5479), .A2(n4661), .ZN(n4660) );
  INV_X1 U5062 ( .A(n5464), .ZN(n4661) );
  INV_X1 U5063 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4823) );
  INV_X1 U5064 ( .A(n5297), .ZN(n4620) );
  AOI21_X1 U5065 ( .B1(n5243), .B2(n5013), .A(n4477), .ZN(n4476) );
  INV_X1 U5066 ( .A(n5261), .ZN(n4477) );
  INV_X1 U5067 ( .A(n4983), .ZN(n4646) );
  INV_X1 U5068 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4860) );
  NAND2_X1 U5069 ( .A1(n5384), .A2(n5385), .ZN(n4733) );
  OR2_X1 U5070 ( .A1(n9542), .A2(n8331), .ZN(n7798) );
  OR2_X1 U5071 ( .A1(n8597), .A2(n8368), .ZN(n7775) );
  AND2_X1 U5072 ( .A1(n7780), .A2(n7782), .ZN(n8343) );
  OR3_X1 U5073 ( .A1(n5526), .A2(n9469), .A3(n5588), .ZN(n5578) );
  NAND2_X1 U5074 ( .A1(n4580), .A2(n4578), .ZN(n4790) );
  AND2_X1 U5075 ( .A1(n7633), .A2(n7629), .ZN(n8100) );
  OR2_X1 U5076 ( .A1(n8614), .A2(n8415), .ZN(n7634) );
  OR2_X1 U5077 ( .A1(n8629), .A2(n8196), .ZN(n7754) );
  NAND2_X1 U5078 ( .A1(n8405), .A2(n4813), .ZN(n4812) );
  OR2_X1 U5079 ( .A1(n5414), .A2(n9392), .ZN(n5434) );
  NAND2_X1 U5080 ( .A1(n8649), .A2(n8253), .ZN(n4493) );
  OR2_X1 U5081 ( .A1(n8656), .A2(n8536), .ZN(n7641) );
  OR2_X1 U5082 ( .A1(n9536), .A2(n8092), .ZN(n7723) );
  AND2_X1 U5083 ( .A1(n7716), .A2(n7710), .ZN(n4819) );
  OR2_X1 U5084 ( .A1(n9901), .A2(n7402), .ZN(n7710) );
  OR2_X1 U5085 ( .A1(n9946), .A2(n7304), .ZN(n7696) );
  NAND2_X1 U5086 ( .A1(n4815), .A2(n4814), .ZN(n7687) );
  INV_X1 U5087 ( .A(n10017), .ZN(n4815) );
  AND2_X1 U5088 ( .A1(n7176), .A2(n7679), .ZN(n4565) );
  INV_X1 U5089 ( .A(n7680), .ZN(n7176) );
  NAND2_X1 U5090 ( .A1(n4376), .A2(n7123), .ZN(n4880) );
  NOR2_X1 U5091 ( .A1(n7167), .A2(n4881), .ZN(n4878) );
  INV_X1 U5092 ( .A(n7123), .ZN(n4881) );
  NAND2_X1 U5093 ( .A1(n7112), .A2(n8263), .ZN(n7668) );
  NAND2_X1 U5094 ( .A1(n8183), .A2(n6796), .ZN(n7650) );
  NAND2_X1 U5095 ( .A1(n6997), .A2(n9988), .ZN(n7648) );
  NAND2_X1 U5096 ( .A1(n4932), .A2(n5041), .ZN(n4885) );
  AND2_X1 U5097 ( .A1(n4396), .A2(n4532), .ZN(n5617) );
  INV_X1 U5098 ( .A(n8946), .ZN(n4692) );
  NAND2_X1 U5099 ( .A1(n9172), .A2(n8927), .ZN(n7980) );
  NOR2_X1 U5100 ( .A1(n9023), .A2(n7886), .ZN(n4698) );
  OR2_X1 U5101 ( .A1(n9197), .A2(n9070), .ZN(n8940) );
  NAND2_X1 U5102 ( .A1(n4672), .A2(n4669), .ZN(n4668) );
  OR2_X1 U5103 ( .A1(n9202), .A2(n9054), .ZN(n8033) );
  OAI21_X1 U5104 ( .B1(n4841), .B2(n4840), .A(n9113), .ZN(n4838) );
  NOR2_X1 U5105 ( .A1(n7841), .A2(n4688), .ZN(n4687) );
  NAND2_X1 U5106 ( .A1(n8123), .A2(n4445), .ZN(n8040) );
  INV_X1 U5107 ( .A(n8819), .ZN(n4445) );
  AND2_X1 U5108 ( .A1(n7913), .A2(n7916), .ZN(n8051) );
  INV_X1 U5109 ( .A(n7570), .ZN(n4654) );
  AOI21_X1 U5110 ( .B1(n7570), .B2(n4653), .A(n4395), .ZN(n4652) );
  INV_X1 U5111 ( .A(n7565), .ZN(n4653) );
  NAND2_X1 U5112 ( .A1(n7562), .A2(n7561), .ZN(n7566) );
  NAND2_X1 U5113 ( .A1(n5502), .A2(n5501), .ZN(n5521) );
  OAI21_X1 U5114 ( .B1(n5328), .B2(n5037), .A(n5036), .ZN(n5347) );
  INV_X1 U5115 ( .A(n4623), .ZN(n4622) );
  OAI21_X1 U5116 ( .B1(n4624), .B2(n4336), .A(n5026), .ZN(n4623) );
  AOI21_X1 U5117 ( .B1(n4476), .B2(n4474), .A(n4473), .ZN(n4472) );
  INV_X1 U5118 ( .A(n5013), .ZN(n4474) );
  INV_X1 U5119 ( .A(n4624), .ZN(n4473) );
  INV_X1 U5120 ( .A(n4476), .ZN(n4475) );
  NAND2_X1 U5121 ( .A1(n4471), .A2(n4476), .ZN(n5019) );
  NAND2_X1 U5122 ( .A1(n5244), .A2(n5013), .ZN(n4471) );
  INV_X1 U5123 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U5124 ( .A1(n4991), .A2(n4990), .ZN(n5170) );
  INV_X1 U5125 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n4984) );
  INV_X1 U5126 ( .A(SI_6_), .ZN(n9438) );
  XNOR2_X1 U5127 ( .A(n8231), .B(n4414), .ZN(n8178) );
  NAND2_X1 U5128 ( .A1(n5145), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5179) );
  OR2_X1 U5129 ( .A1(n5377), .A2(n9405), .ZN(n5394) );
  NOR2_X1 U5130 ( .A1(n4744), .A2(n4740), .ZN(n4739) );
  INV_X1 U5131 ( .A(n5222), .ZN(n4740) );
  INV_X1 U5132 ( .A(n5242), .ZN(n4744) );
  NAND2_X1 U5133 ( .A1(n7243), .A2(n5276), .ZN(n9533) );
  INV_X1 U5134 ( .A(n5325), .ZN(n4748) );
  NAND2_X1 U5135 ( .A1(n5326), .A2(n4751), .ZN(n4750) );
  NAND2_X1 U5136 ( .A1(n4328), .A2(n9532), .ZN(n4751) );
  AOI21_X1 U5137 ( .B1(n5431), .B2(n4755), .A(n5439), .ZN(n4754) );
  INV_X1 U5138 ( .A(n8167), .ZN(n4755) );
  NAND2_X1 U5139 ( .A1(n4726), .A2(n4725), .ZN(n4724) );
  INV_X1 U5140 ( .A(n5401), .ZN(n4725) );
  OR2_X1 U5141 ( .A1(n5232), .A2(n4943), .ZN(n5250) );
  NAND2_X1 U5142 ( .A1(n9542), .A2(n8331), .ZN(n7799) );
  OR2_X1 U5143 ( .A1(n7432), .A2(n7431), .ZN(n4537) );
  NAND2_X1 U5144 ( .A1(n7568), .A2(n7567), .ZN(n8327) );
  OR2_X1 U5145 ( .A1(n4790), .A2(n8340), .ZN(n4785) );
  INV_X1 U5146 ( .A(n4789), .ZN(n4788) );
  OAI21_X1 U5147 ( .B1(n8340), .B2(n7633), .A(n7775), .ZN(n4789) );
  NOR2_X1 U5148 ( .A1(n8100), .A2(n4581), .ZN(n4896) );
  INV_X1 U5149 ( .A(n4898), .ZN(n4897) );
  OAI21_X1 U5150 ( .B1(n8100), .B2(n4901), .A(n4899), .ZN(n4898) );
  NAND2_X1 U5151 ( .A1(n4900), .A2(n8242), .ZN(n4899) );
  AOI21_X1 U5152 ( .B1(n4322), .B2(n4323), .A(n4332), .ZN(n4576) );
  INV_X1 U5153 ( .A(n4790), .ZN(n8365) );
  INV_X1 U5154 ( .A(n8100), .ZN(n8367) );
  INV_X1 U5155 ( .A(n4807), .ZN(n4806) );
  OAI21_X1 U5156 ( .B1(n4808), .B2(n8389), .A(n7634), .ZN(n4807) );
  NAND2_X1 U5157 ( .A1(n4810), .A2(n4811), .ZN(n4808) );
  NAND2_X1 U5158 ( .A1(n4456), .A2(n4455), .ZN(n8374) );
  OR2_X1 U5159 ( .A1(n8614), .A2(n8251), .ZN(n4455) );
  NAND2_X1 U5160 ( .A1(n4457), .A2(n8389), .ZN(n4456) );
  NAND2_X1 U5161 ( .A1(n7767), .A2(n8425), .ZN(n4811) );
  NAND2_X1 U5162 ( .A1(n8624), .A2(n4460), .ZN(n8404) );
  NAND2_X1 U5163 ( .A1(n8622), .A2(n8252), .ZN(n4460) );
  NOR2_X1 U5164 ( .A1(n8404), .A2(n8405), .ZN(n8403) );
  NAND2_X1 U5165 ( .A1(n4560), .A2(n4558), .ZN(n8462) );
  AND2_X1 U5166 ( .A1(n8463), .A2(n4559), .ZN(n4558) );
  NAND2_X1 U5167 ( .A1(n4561), .A2(n4562), .ZN(n4559) );
  AOI21_X1 U5168 ( .B1(n4485), .B2(n4483), .A(n4373), .ZN(n4482) );
  INV_X1 U5169 ( .A(n4489), .ZN(n4483) );
  INV_X1 U5170 ( .A(n4485), .ZN(n4484) );
  NOR2_X1 U5171 ( .A1(n4490), .A2(n8514), .ZN(n4489) );
  INV_X1 U5172 ( .A(n4493), .ZN(n4490) );
  AND4_X1 U5173 ( .A1(n4952), .A2(n4951), .A3(n4950), .A4(n4949), .ZN(n8519)
         );
  NOR2_X1 U5174 ( .A1(n7558), .A2(n4799), .ZN(n4798) );
  INV_X1 U5175 ( .A(n8532), .ZN(n4905) );
  AND2_X1 U5176 ( .A1(n7731), .A2(n7732), .ZN(n8532) );
  NAND2_X1 U5177 ( .A1(n7556), .A2(n7723), .ZN(n8556) );
  NAND2_X1 U5178 ( .A1(n8556), .A2(n8557), .ZN(n8560) );
  NOR2_X1 U5179 ( .A1(n9536), .A2(n4911), .ZN(n4910) );
  INV_X1 U5180 ( .A(n8092), .ZN(n4911) );
  OR2_X1 U5181 ( .A1(n4706), .A2(n7459), .ZN(n4915) );
  NOR2_X1 U5182 ( .A1(n7456), .A2(n7721), .ZN(n8091) );
  AND2_X1 U5183 ( .A1(n7723), .A2(n7724), .ZN(n7721) );
  OAI21_X1 U5184 ( .B1(n7225), .B2(n4890), .A(n4886), .ZN(n9935) );
  AOI21_X1 U5185 ( .B1(n4889), .B2(n8575), .A(n4365), .ZN(n4886) );
  INV_X1 U5186 ( .A(n10022), .ZN(n4888) );
  NAND2_X1 U5187 ( .A1(n7174), .A2(n7173), .ZN(n4566) );
  AOI21_X1 U5188 ( .B1(n4870), .B2(n6755), .A(n4364), .ZN(n4869) );
  OR2_X1 U5189 ( .A1(n6448), .A2(n5591), .ZN(n8535) );
  INV_X1 U5190 ( .A(n8478), .ZN(n8537) );
  NOR2_X1 U5191 ( .A1(n6299), .A2(n6292), .ZN(n4709) );
  NAND2_X1 U5192 ( .A1(n7579), .A2(n7578), .ZN(n8587) );
  NAND2_X1 U5193 ( .A1(n5486), .A2(n5485), .ZN(n8608) );
  NAND2_X1 U5194 ( .A1(n7550), .A2(n5484), .ZN(n5486) );
  NAND2_X1 U5195 ( .A1(n5447), .A2(n5446), .ZN(n8617) );
  INV_X1 U5196 ( .A(n8511), .ZN(n8649) );
  NAND2_X1 U5197 ( .A1(n4478), .A2(n5321), .ZN(n8665) );
  NAND2_X1 U5198 ( .A1(n6721), .A2(n5484), .ZN(n4478) );
  OAI211_X2 U5199 ( .C1(n6466), .C2(n6303), .A(n5131), .B(n5130), .ZN(n9957)
         );
  INV_X1 U5200 ( .A(n10048), .ZN(n10018) );
  INV_X1 U5201 ( .A(n8187), .ZN(n9988) );
  OR2_X1 U5202 ( .A1(n7812), .A2(n9982), .ZN(n10048) );
  AND2_X1 U5203 ( .A1(n5551), .A2(n5549), .ZN(n9971) );
  OR2_X1 U5204 ( .A1(n5562), .A2(n5548), .ZN(n5549) );
  INV_X1 U5205 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4570) );
  NAND2_X1 U5206 ( .A1(n4919), .A2(n4868), .ZN(n4867) );
  INV_X1 U5207 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4868) );
  AND2_X1 U5208 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4966) );
  NAND2_X1 U5209 ( .A1(n4518), .A2(n4517), .ZN(n4516) );
  INV_X1 U5210 ( .A(n8116), .ZN(n4518) );
  INV_X1 U5211 ( .A(n8117), .ZN(n4517) );
  NAND2_X1 U5212 ( .A1(n4520), .A2(n4342), .ZN(n4519) );
  INV_X1 U5213 ( .A(n8119), .ZN(n4520) );
  NAND2_X1 U5214 ( .A1(n7335), .A2(n7334), .ZN(n5880) );
  INV_X1 U5215 ( .A(n5761), .ZN(n5763) );
  INV_X1 U5216 ( .A(n4777), .ZN(n4776) );
  NAND2_X1 U5217 ( .A1(n4357), .A2(n6028), .ZN(n8715) );
  INV_X1 U5218 ( .A(n5840), .ZN(n4765) );
  INV_X1 U5219 ( .A(n7157), .ZN(n4764) );
  INV_X1 U5220 ( .A(n5818), .ZN(n5821) );
  AND2_X1 U5221 ( .A1(n4525), .A2(n8731), .ZN(n4524) );
  OR2_X1 U5222 ( .A1(n8767), .A2(n4526), .ZN(n4525) );
  INV_X1 U5223 ( .A(n6139), .ZN(n4526) );
  NAND2_X1 U5224 ( .A1(n5940), .A2(n4767), .ZN(n9573) );
  NAND2_X1 U5225 ( .A1(n5940), .A2(n7539), .ZN(n4770) );
  INV_X1 U5226 ( .A(n6241), .ZN(n8087) );
  OAI21_X1 U5227 ( .B1(n4451), .B2(n4450), .A(n4446), .ZN(n4618) );
  INV_X1 U5228 ( .A(n8025), .ZN(n4450) );
  AOI21_X1 U5229 ( .B1(n4449), .B2(n4448), .A(n4447), .ZN(n4446) );
  INV_X1 U5230 ( .A(n7997), .ZN(n4451) );
  OR2_X1 U5231 ( .A1(n9753), .A2(n9754), .ZN(n4599) );
  OR2_X1 U5232 ( .A1(n6748), .A2(n6749), .ZN(n4602) );
  AND2_X1 U5233 ( .A1(n6835), .A2(n6836), .ZN(n7252) );
  OR2_X1 U5234 ( .A1(n8847), .A2(n8846), .ZN(n4596) );
  NAND2_X1 U5235 ( .A1(n7874), .A2(n7873), .ZN(n8901) );
  NAND2_X1 U5236 ( .A1(n7818), .A2(n7817), .ZN(n9162) );
  NOR2_X1 U5237 ( .A1(n9004), .A2(n4583), .ZN(n8966) );
  NAND2_X1 U5238 ( .A1(n4851), .A2(n4853), .ZN(n4850) );
  NAND2_X1 U5239 ( .A1(n8926), .A2(n4854), .ZN(n4851) );
  INV_X1 U5240 ( .A(n4697), .ZN(n4696) );
  OAI21_X1 U5241 ( .B1(n8944), .B2(n4698), .A(n8943), .ZN(n4697) );
  INV_X1 U5242 ( .A(n9034), .ZN(n4695) );
  NAND2_X1 U5243 ( .A1(n8943), .A2(n8031), .ZN(n9013) );
  INV_X1 U5244 ( .A(n8998), .ZN(n9025) );
  AND2_X1 U5245 ( .A1(n9034), .A2(n4698), .ZN(n9021) );
  OAI21_X1 U5246 ( .B1(n9065), .B2(n8941), .A(n8940), .ZN(n9036) );
  NAND2_X1 U5247 ( .A1(n9036), .A2(n9035), .ZN(n9034) );
  NAND2_X1 U5248 ( .A1(n4416), .A2(n4415), .ZN(n8922) );
  NAND2_X1 U5249 ( .A1(n9061), .A2(n9070), .ZN(n4415) );
  AOI21_X1 U5250 ( .B1(n9064), .B2(n9067), .A(n8917), .ZN(n9048) );
  AND2_X1 U5251 ( .A1(n9202), .A2(n9087), .ZN(n8917) );
  AOI21_X1 U5252 ( .B1(n4675), .B2(n4674), .A(n4673), .ZN(n4672) );
  INV_X1 U5253 ( .A(n8936), .ZN(n4674) );
  OR2_X1 U5254 ( .A1(n9094), .A2(n9205), .ZN(n9079) );
  AND2_X1 U5255 ( .A1(n4669), .A2(n8938), .ZN(n9085) );
  AOI21_X1 U5256 ( .B1(n9093), .B2(n8915), .A(n4844), .ZN(n9078) );
  NOR2_X1 U5257 ( .A1(n9210), .A2(n9088), .ZN(n4844) );
  NAND2_X1 U5258 ( .A1(n9132), .A2(n8936), .ZN(n4676) );
  AND2_X1 U5259 ( .A1(n8034), .A2(n8937), .ZN(n9101) );
  NOR2_X1 U5260 ( .A1(n8914), .A2(n4842), .ZN(n4841) );
  OR2_X1 U5261 ( .A1(n9595), .A2(n8909), .ZN(n8910) );
  NOR2_X1 U5262 ( .A1(n9605), .A2(n9622), .ZN(n9606) );
  NOR2_X1 U5263 ( .A1(n7500), .A2(n4830), .ZN(n4829) );
  INV_X1 U5264 ( .A(n7369), .ZN(n4830) );
  NAND2_X1 U5265 ( .A1(n4375), .A2(n4834), .ZN(n4831) );
  NAND2_X1 U5266 ( .A1(n4339), .A2(n7369), .ZN(n4832) );
  NAND2_X1 U5267 ( .A1(n7843), .A2(n7920), .ZN(n4677) );
  NAND2_X1 U5268 ( .A1(n7371), .A2(n4687), .ZN(n4683) );
  OAI22_X1 U5269 ( .A1(n7321), .A2(n7320), .B1(n8816), .B2(n7319), .ZN(n7366)
         );
  NAND3_X1 U5270 ( .A1(n7141), .A2(n4592), .A3(n4593), .ZN(n7327) );
  NOR2_X1 U5271 ( .A1(n7277), .A2(n7319), .ZN(n4592) );
  NAND2_X1 U5272 ( .A1(n7904), .A2(n8003), .ZN(n7095) );
  NAND2_X1 U5273 ( .A1(n7091), .A2(n7095), .ZN(n7104) );
  NAND2_X1 U5274 ( .A1(n6910), .A2(n8037), .ZN(n7040) );
  XNOR2_X1 U5275 ( .A(n8822), .B(n9835), .ZN(n7019) );
  NAND2_X1 U5276 ( .A1(n6868), .A2(n6867), .ZN(n6870) );
  OR2_X1 U5277 ( .A1(n6870), .A2(n8043), .ZN(n6908) );
  INV_X1 U5278 ( .A(n7835), .ZN(n6872) );
  NAND2_X1 U5279 ( .A1(n5969), .A2(n5968), .ZN(n9227) );
  INV_X1 U5280 ( .A(n8123), .ZN(n9846) );
  OR2_X1 U5281 ( .A1(n7995), .A2(n8078), .ZN(n9658) );
  INV_X1 U5282 ( .A(n6447), .ZN(n8084) );
  XNOR2_X1 U5283 ( .A(n7593), .B(n7592), .ZN(n8687) );
  NAND2_X1 U5284 ( .A1(n7588), .A2(n7587), .ZN(n7593) );
  AND2_X1 U5285 ( .A1(n5639), .A2(n5638), .ZN(n5641) );
  INV_X1 U5286 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5642) );
  XNOR2_X1 U5287 ( .A(n5521), .B(n5520), .ZN(n8700) );
  NAND2_X1 U5288 ( .A1(n4632), .A2(n5405), .ZN(n5425) );
  NAND2_X1 U5289 ( .A1(n5389), .A2(n4633), .ZN(n4632) );
  NAND2_X1 U5290 ( .A1(n5389), .A2(n5388), .ZN(n5407) );
  NAND2_X1 U5291 ( .A1(n4780), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5610) );
  NOR2_X1 U5292 ( .A1(n4782), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n4781) );
  NAND2_X1 U5293 ( .A1(n5881), .A2(n5604), .ZN(n5986) );
  OAI21_X1 U5294 ( .B1(n5244), .B2(n5243), .A(n5013), .ZN(n5262) );
  OAI21_X1 U5295 ( .B1(n4998), .B2(n4641), .A(n4638), .ZN(n5224) );
  OAI21_X1 U5296 ( .B1(n4462), .B2(n5142), .A(n4461), .ZN(n5189) );
  AOI21_X1 U5297 ( .B1(n4466), .B2(n4645), .A(n4465), .ZN(n4461) );
  INV_X1 U5298 ( .A(n4466), .ZN(n4462) );
  INV_X1 U5299 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5965) );
  XNOR2_X1 U5300 ( .A(n4982), .B(n9438), .ZN(n5141) );
  NAND2_X1 U5301 ( .A1(n4978), .A2(n4977), .ZN(n5129) );
  NAND2_X1 U5302 ( .A1(n4420), .A2(SI_2_), .ZN(n4969) );
  XNOR2_X1 U5303 ( .A(n4971), .B(SI_3_), .ZN(n5091) );
  NAND2_X1 U5304 ( .A1(n6807), .A2(n5155), .ZN(n6935) );
  CLKBUF_X1 U5305 ( .A(n6986), .Z(n7056) );
  INV_X1 U5306 ( .A(n8461), .ZN(n8093) );
  NAND2_X1 U5307 ( .A1(n5302), .A2(n5301), .ZN(n8660) );
  INV_X1 U5308 ( .A(n7810), .ZN(n4804) );
  INV_X1 U5309 ( .A(n7816), .ZN(n4802) );
  AOI21_X1 U5310 ( .B1(n7810), .B2(n4335), .A(n7814), .ZN(n4803) );
  AND2_X1 U5311 ( .A1(n5495), .A2(n5494), .ZN(n8393) );
  NAND4_X1 U5312 ( .A1(n5126), .A2(n5125), .A3(n5124), .A4(n5123), .ZN(n8261)
         );
  OAI21_X1 U5313 ( .B1(n8321), .B2(n9929), .A(n4356), .ZN(n4543) );
  OAI22_X1 U5314 ( .A1(n8323), .A2(n9929), .B1(n8322), .B2(n9928), .ZN(n4539)
         );
  OAI21_X1 U5315 ( .B1(n8325), .B2(n8326), .A(n8324), .ZN(n4541) );
  CLKBUF_X1 U5316 ( .A(n5575), .Z(n8383) );
  NOR2_X1 U5317 ( .A1(n8145), .A2(n8144), .ZN(n8143) );
  NAND2_X1 U5318 ( .A1(n6198), .A2(n6197), .ZN(n9166) );
  NOR2_X1 U5319 ( .A1(n4510), .A2(n4354), .ZN(n4509) );
  NAND2_X1 U5320 ( .A1(n6141), .A2(n6140), .ZN(n9180) );
  NAND2_X1 U5321 ( .A1(n8706), .A2(n8708), .ZN(n6119) );
  NAND2_X1 U5322 ( .A1(n4503), .A2(n4504), .ZN(n7441) );
  AND2_X1 U5323 ( .A1(n4502), .A2(n5904), .ZN(n4504) );
  OR2_X1 U5324 ( .A1(n7335), .A2(n4507), .ZN(n4503) );
  NAND2_X1 U5325 ( .A1(n7550), .A2(n5962), .ZN(n6160) );
  NAND2_X1 U5326 ( .A1(n4618), .A2(n4617), .ZN(n4616) );
  NAND2_X1 U5327 ( .A1(n6242), .A2(n8072), .ZN(n4617) );
  NAND4_X1 U5328 ( .A1(n5724), .A2(n5723), .A3(n5722), .A4(n5721), .ZN(n8821)
         );
  XNOR2_X1 U5329 ( .A(n6361), .B(n4603), .ZN(n6362) );
  OAI21_X1 U5330 ( .B1(n8891), .B2(n8890), .A(n8889), .ZN(n4608) );
  OAI21_X1 U5331 ( .B1(n8886), .B2(n9775), .A(n4612), .ZN(n4611) );
  OR2_X1 U5332 ( .A1(n8888), .A2(n9736), .ZN(n4612) );
  OAI21_X1 U5333 ( .B1(n4412), .B2(n9643), .A(n4409), .ZN(n9164) );
  AOI21_X1 U5334 ( .B1(n4411), .B2(n9641), .A(n4410), .ZN(n4409) );
  NOR2_X1 U5335 ( .A1(n8954), .A2(n8953), .ZN(n4410) );
  OR2_X1 U5336 ( .A1(n9169), .A2(n9156), .ZN(n4702) );
  AOI21_X1 U5337 ( .B1(n8975), .B2(n9613), .A(n4703), .ZN(n9168) );
  NAND2_X1 U5338 ( .A1(n4705), .A2(n4704), .ZN(n4703) );
  NAND2_X1 U5339 ( .A1(n8974), .A2(n9638), .ZN(n4704) );
  NAND2_X1 U5340 ( .A1(n6121), .A2(n6120), .ZN(n9187) );
  OAI211_X1 U5341 ( .C1(n6275), .C2(n6418), .A(n5793), .B(n5792), .ZN(n7102)
         );
  OR2_X1 U5342 ( .A1(n9149), .A2(n6929), .ZN(n9152) );
  INV_X1 U5343 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9260) );
  INV_X1 U5344 ( .A(n4782), .ZN(n4779) );
  OAI21_X1 U5345 ( .B1(n7672), .B2(n7671), .A(n7670), .ZN(n7675) );
  NAND2_X1 U5346 ( .A1(n4405), .A2(n4404), .ZN(n7685) );
  NOR2_X1 U5347 ( .A1(n7681), .A2(n7680), .ZN(n4404) );
  AND2_X1 U5348 ( .A1(n7721), .A2(n7720), .ZN(n4403) );
  NOR2_X1 U5349 ( .A1(n7925), .A2(n7926), .ZN(n4439) );
  NAND2_X1 U5350 ( .A1(n4443), .A2(n4441), .ZN(n7934) );
  AOI21_X1 U5351 ( .B1(n4442), .B2(n7988), .A(n7923), .ZN(n4441) );
  NAND2_X1 U5352 ( .A1(n4444), .A2(n7995), .ZN(n4443) );
  NAND2_X1 U5353 ( .A1(n4452), .A2(n7947), .ZN(n7952) );
  OAI21_X1 U5354 ( .B1(n4454), .B2(n4453), .A(n7945), .ZN(n4452) );
  NAND2_X1 U5355 ( .A1(n4656), .A2(n4655), .ZN(n7774) );
  NAND2_X1 U5356 ( .A1(n7637), .A2(n7791), .ZN(n4656) );
  OAI21_X1 U5357 ( .B1(n7636), .B2(n8376), .A(n7797), .ZN(n4655) );
  NOR2_X1 U5358 ( .A1(n7974), .A2(n7979), .ZN(n4431) );
  NAND2_X1 U5359 ( .A1(n7981), .A2(n8949), .ZN(n4437) );
  OAI22_X1 U5360 ( .A1(n4435), .A2(n4358), .B1(n7974), .B2(n4433), .ZN(n4432)
         );
  MUX2_X1 U5361 ( .A(n7793), .B(n7792), .S(n7791), .Z(n7794) );
  NOR2_X1 U5362 ( .A1(n8516), .A2(n4796), .ZN(n4795) );
  INV_X1 U5363 ( .A(n7732), .ZN(n4796) );
  INV_X1 U5364 ( .A(n4885), .ZN(n4883) );
  OR2_X1 U5365 ( .A1(n7437), .A2(n4505), .ZN(n4501) );
  NAND2_X1 U5366 ( .A1(n4772), .A2(n7438), .ZN(n4497) );
  OAI21_X1 U5367 ( .B1(n7371), .B2(n4681), .A(n4678), .ZN(n9612) );
  NOR2_X1 U5368 ( .A1(n4686), .A2(n7926), .ZN(n4682) );
  INV_X1 U5369 ( .A(n5441), .ZN(n4627) );
  NOR2_X1 U5370 ( .A1(n5022), .A2(n4625), .ZN(n4624) );
  INV_X1 U5371 ( .A(n5018), .ZN(n4625) );
  INV_X1 U5372 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4964) );
  NOR2_X1 U5373 ( .A1(n5431), .A2(n8167), .ZN(n4753) );
  INV_X1 U5374 ( .A(n8194), .ZN(n4727) );
  INV_X1 U5375 ( .A(n5402), .ZN(n4726) );
  NOR4_X1 U5376 ( .A1(n7625), .A2(n7790), .A3(n8346), .A4(n7624), .ZN(n7626)
         );
  NAND2_X1 U5377 ( .A1(n7286), .A2(n4549), .ZN(n7426) );
  OR2_X1 U5378 ( .A1(n7291), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4549) );
  NOR2_X1 U5379 ( .A1(n8649), .A2(n8656), .ZN(n4717) );
  NOR2_X1 U5380 ( .A1(n4794), .A2(n4909), .ZN(n4575) );
  INV_X1 U5381 ( .A(n4795), .ZN(n4794) );
  INV_X1 U5382 ( .A(n4791), .ZN(n4572) );
  AOI21_X1 U5383 ( .B1(n4795), .B2(n4793), .A(n4792), .ZN(n4791) );
  INV_X1 U5384 ( .A(n7641), .ZN(n4792) );
  INV_X1 U5385 ( .A(n4798), .ZN(n4793) );
  NAND2_X1 U5386 ( .A1(n8660), .A2(n8254), .ZN(n4908) );
  INV_X1 U5387 ( .A(n6635), .ZN(n4870) );
  NAND2_X1 U5388 ( .A1(n8406), .A2(n8400), .ZN(n8394) );
  OR2_X1 U5389 ( .A1(n6770), .A2(n6769), .ZN(n6945) );
  NAND2_X1 U5390 ( .A1(n6781), .A2(n7112), .ZN(n6770) );
  NAND2_X1 U5391 ( .A1(n4959), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4958) );
  INV_X1 U5392 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4953) );
  NAND2_X1 U5393 ( .A1(n8722), .A2(n8723), .ZN(n4775) );
  INV_X1 U5394 ( .A(n4514), .ZN(n4513) );
  OAI21_X1 U5395 ( .B1(n4516), .B2(n4515), .A(n6280), .ZN(n4514) );
  NAND2_X1 U5396 ( .A1(n4771), .A2(n6354), .ZN(n6217) );
  NAND2_X1 U5397 ( .A1(n7994), .A2(n8025), .ZN(n4449) );
  AND2_X1 U5398 ( .A1(n7996), .A2(n7988), .ZN(n4447) );
  NOR2_X1 U5399 ( .A1(n8070), .A2(n7988), .ZN(n4448) );
  OR2_X1 U5400 ( .A1(n8901), .A2(n8953), .ZN(n8068) );
  OR2_X1 U5401 ( .A1(n9166), .A2(n8981), .ZN(n7982) );
  OR2_X1 U5402 ( .A1(n9175), .A2(n9015), .ZN(n8926) );
  OR2_X1 U5403 ( .A1(n4590), .A2(n9192), .ZN(n4589) );
  NOR2_X1 U5404 ( .A1(n9595), .A2(n9227), .ZN(n4587) );
  NAND2_X1 U5405 ( .A1(n5971), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5990) );
  NOR2_X1 U5406 ( .A1(n8908), .A2(n8907), .ZN(n9587) );
  AND2_X1 U5407 ( .A1(n9232), .A2(n9616), .ZN(n4833) );
  INV_X1 U5408 ( .A(n4829), .ZN(n4825) );
  OR2_X1 U5409 ( .A1(n9522), .A2(n7322), .ZN(n7922) );
  OR2_X1 U5410 ( .A1(n5827), .A2(n5826), .ZN(n5848) );
  NAND2_X1 U5411 ( .A1(n7892), .A2(n7080), .ZN(n4663) );
  AND2_X1 U5412 ( .A1(n9855), .A2(n9846), .ZN(n4593) );
  OR2_X1 U5413 ( .A1(n8818), .A2(n9855), .ZN(n7904) );
  OR2_X1 U5414 ( .A1(n8820), .A2(n9842), .ZN(n7899) );
  NAND2_X1 U5415 ( .A1(n4848), .A2(n4367), .ZN(n4847) );
  NOR2_X1 U5416 ( .A1(n9079), .A2(n4589), .ZN(n9041) );
  NOR2_X1 U5417 ( .A1(n9079), .A2(n4590), .ZN(n9056) );
  NAND2_X1 U5418 ( .A1(n9599), .A2(n9598), .ZN(n9597) );
  OR2_X1 U5419 ( .A1(n9629), .A2(n9237), .ZN(n9605) );
  NAND2_X1 U5420 ( .A1(n4684), .A2(n7843), .ZN(n9637) );
  OR2_X1 U5421 ( .A1(n7371), .A2(n7920), .ZN(n4684) );
  NOR2_X1 U5422 ( .A1(n7327), .A2(n9522), .ZN(n9627) );
  INV_X1 U5423 ( .A(n6692), .ZN(n8039) );
  AOI21_X1 U5424 ( .B1(n4652), .B2(n4654), .A(n4651), .ZN(n4650) );
  INV_X1 U5425 ( .A(n7585), .ZN(n4651) );
  NAND2_X1 U5426 ( .A1(n4659), .A2(n4657), .ZN(n5500) );
  AOI21_X1 U5427 ( .B1(n4660), .B2(n4662), .A(n4658), .ZN(n4657) );
  INV_X1 U5428 ( .A(n5478), .ZN(n4658) );
  AND2_X1 U5429 ( .A1(n4823), .A2(n5631), .ZN(n4529) );
  AND2_X1 U5430 ( .A1(n4531), .A2(n5613), .ZN(n4528) );
  INV_X1 U5431 ( .A(n5462), .ZN(n4662) );
  NOR2_X1 U5432 ( .A1(n5406), .A2(n4634), .ZN(n4633) );
  INV_X1 U5433 ( .A(n5388), .ZN(n4634) );
  INV_X1 U5434 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U5435 ( .A1(n5033), .A2(n5032), .ZN(n5328) );
  NAND2_X1 U5436 ( .A1(n4621), .A2(n4619), .ZN(n5033) );
  AOI21_X1 U5437 ( .B1(n4622), .B2(n4336), .A(n4620), .ZN(n4619) );
  NAND2_X1 U5438 ( .A1(n5010), .A2(n5009), .ZN(n5013) );
  AOI21_X1 U5439 ( .B1(n5208), .B2(n4640), .A(n4639), .ZN(n4638) );
  INV_X1 U5440 ( .A(n5004), .ZN(n4639) );
  INV_X1 U5441 ( .A(n4997), .ZN(n4640) );
  INV_X1 U5442 ( .A(n5208), .ZN(n4641) );
  NAND2_X1 U5443 ( .A1(n4710), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4421) );
  INV_X1 U5444 ( .A(SI_2_), .ZN(n9427) );
  NAND2_X1 U5445 ( .A1(n4821), .A2(n4820), .ZN(n5043) );
  NAND2_X1 U5446 ( .A1(n9500), .A2(n4965), .ZN(n4820) );
  NAND2_X1 U5447 ( .A1(n9501), .A2(n4964), .ZN(n4821) );
  INV_X1 U5448 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4965) );
  INV_X1 U5449 ( .A(SI_8_), .ZN(n9364) );
  NOR2_X1 U5450 ( .A1(n5179), .A2(n4942), .ZN(n5193) );
  INV_X1 U5451 ( .A(n5394), .ZN(n5393) );
  OR2_X1 U5452 ( .A1(n4731), .A2(n4729), .ZN(n4728) );
  INV_X1 U5453 ( .A(n4733), .ZN(n4729) );
  AND2_X1 U5454 ( .A1(n8220), .A2(n4732), .ZN(n4731) );
  NAND2_X1 U5455 ( .A1(n7529), .A2(n7530), .ZN(n4732) );
  AND2_X1 U5456 ( .A1(n4733), .A2(n7530), .ZN(n4723) );
  AND2_X1 U5457 ( .A1(n5118), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5145) );
  NAND2_X1 U5458 ( .A1(n6807), .A2(n4758), .ZN(n6976) );
  NOR2_X1 U5459 ( .A1(n6934), .A2(n4759), .ZN(n4758) );
  INV_X1 U5460 ( .A(n5155), .ZN(n4759) );
  INV_X1 U5461 ( .A(n8232), .ZN(n4399) );
  AND2_X1 U5462 ( .A1(n9972), .A2(n6627), .ZN(n8137) );
  OR2_X1 U5463 ( .A1(n5333), .A2(n4946), .ZN(n5334) );
  INV_X1 U5464 ( .A(n5476), .ZN(n8205) );
  XNOR2_X1 U5465 ( .A(n8608), .B(n4414), .ZN(n8157) );
  NAND2_X1 U5466 ( .A1(n4387), .A2(n4328), .ZN(n7480) );
  AND2_X1 U5467 ( .A1(n7798), .A2(n7787), .ZN(n7792) );
  NAND2_X1 U5468 ( .A1(n4787), .A2(n4786), .ZN(n7569) );
  AOI21_X1 U5469 ( .B1(n4788), .B2(n8340), .A(n7778), .ZN(n4786) );
  OR2_X1 U5470 ( .A1(n8327), .A2(n8109), .ZN(n7780) );
  AND4_X1 U5471 ( .A1(n5237), .A2(n5236), .A3(n5235), .A4(n5234), .ZN(n7355)
         );
  AND4_X1 U5472 ( .A1(n5198), .A2(n5197), .A3(n5196), .A4(n5195), .ZN(n7305)
         );
  OR2_X1 U5473 ( .A1(n6557), .A2(n6556), .ZN(n4556) );
  OR2_X1 U5474 ( .A1(n6514), .A2(n6513), .ZN(n4547) );
  OR2_X1 U5475 ( .A1(n6569), .A2(n6568), .ZN(n4545) );
  NOR2_X1 U5476 ( .A1(n6674), .A2(n4551), .ZN(n6678) );
  AND2_X1 U5477 ( .A1(n6675), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4551) );
  NAND2_X1 U5478 ( .A1(n6678), .A2(n6677), .ZN(n6858) );
  NAND2_X1 U5479 ( .A1(n7004), .A2(n4550), .ZN(n7005) );
  OR2_X1 U5480 ( .A1(n7012), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4550) );
  NAND2_X1 U5481 ( .A1(n7005), .A2(n7006), .ZN(n7286) );
  XNOR2_X1 U5482 ( .A(n7426), .B(n4548), .ZN(n7288) );
  INV_X1 U5483 ( .A(n7427), .ZN(n4548) );
  OR2_X1 U5484 ( .A1(n8288), .A2(n8287), .ZN(n8294) );
  NAND2_X1 U5485 ( .A1(n8591), .A2(n8353), .ZN(n8352) );
  AND2_X1 U5486 ( .A1(n8340), .A2(n4896), .ZN(n4895) );
  NOR2_X1 U5487 ( .A1(n4897), .A2(n8107), .ZN(n4894) );
  AND2_X1 U5488 ( .A1(n5527), .A2(n5578), .ZN(n8103) );
  AND2_X1 U5489 ( .A1(n8105), .A2(n8362), .ZN(n8353) );
  OR2_X1 U5490 ( .A1(n8394), .A2(n8608), .ZN(n8380) );
  OR2_X1 U5491 ( .A1(n5449), .A2(n9346), .ZN(n5470) );
  NOR2_X1 U5492 ( .A1(n8423), .A2(n4812), .ZN(n8412) );
  AND2_X1 U5493 ( .A1(n8427), .A2(n8411), .ZN(n8406) );
  NOR2_X1 U5494 ( .A1(n8629), .A2(n8096), .ZN(n8097) );
  NOR2_X1 U5495 ( .A1(n8622), .A2(n8437), .ZN(n8427) );
  NOR2_X1 U5496 ( .A1(n8432), .A2(n8422), .ZN(n8423) );
  OR2_X1 U5497 ( .A1(n8455), .A2(n8629), .ZN(n8437) );
  INV_X1 U5498 ( .A(n8098), .ZN(n8443) );
  NAND2_X1 U5499 ( .A1(n8487), .A2(n7742), .ZN(n4562) );
  NAND2_X1 U5500 ( .A1(n4563), .A2(n7742), .ZN(n4561) );
  NAND2_X1 U5501 ( .A1(n4564), .A2(n7741), .ZN(n4563) );
  AND2_X1 U5502 ( .A1(n7759), .A2(n8444), .ZN(n8463) );
  NOR2_X1 U5503 ( .A1(n4484), .A2(n4564), .ZN(n4480) );
  OAI21_X1 U5504 ( .B1(n4482), .B2(n4564), .A(n4369), .ZN(n4479) );
  INV_X1 U5505 ( .A(n8515), .ZN(n4481) );
  AND2_X1 U5506 ( .A1(n8541), .A2(n4713), .ZN(n8471) );
  NOR2_X1 U5507 ( .A1(n8638), .A2(n4715), .ZN(n4713) );
  OR2_X1 U5508 ( .A1(n5358), .A2(n5357), .ZN(n5377) );
  AND4_X1 U5509 ( .A1(n5382), .A2(n5381), .A3(n5380), .A4(n5379), .ZN(n8493)
         );
  NOR2_X1 U5510 ( .A1(n8501), .A2(n7559), .ZN(n8491) );
  NOR2_X1 U5511 ( .A1(n8491), .A2(n8490), .ZN(n8489) );
  NAND2_X1 U5512 ( .A1(n8541), .A2(n4717), .ZN(n8506) );
  OAI21_X1 U5513 ( .B1(n7556), .B2(n4574), .A(n4571), .ZN(n8503) );
  AOI21_X1 U5514 ( .B1(n4575), .B2(n4573), .A(n4572), .ZN(n4571) );
  INV_X1 U5515 ( .A(n4575), .ZN(n4574) );
  INV_X1 U5516 ( .A(n7723), .ZN(n4573) );
  NAND2_X1 U5517 ( .A1(n8541), .A2(n8528), .ZN(n8521) );
  AND2_X1 U5518 ( .A1(n8550), .A2(n8546), .ZN(n8541) );
  AND2_X1 U5519 ( .A1(n8549), .A2(n8555), .ZN(n8550) );
  NAND2_X1 U5520 ( .A1(n7704), .A2(n7718), .ZN(n4818) );
  NAND2_X1 U5521 ( .A1(n4817), .A2(n7718), .ZN(n4816) );
  INV_X1 U5522 ( .A(n4819), .ZN(n4817) );
  NAND2_X1 U5523 ( .A1(n7401), .A2(n4819), .ZN(n7457) );
  NAND2_X1 U5524 ( .A1(n7397), .A2(n7396), .ZN(n7399) );
  NOR2_X1 U5525 ( .A1(n7347), .A2(n9946), .ZN(n4708) );
  NAND2_X1 U5526 ( .A1(n9949), .A2(n4324), .ZN(n7408) );
  OR2_X1 U5527 ( .A1(n7354), .A2(n7694), .ZN(n7401) );
  AND2_X1 U5528 ( .A1(n9949), .A2(n10034), .ZN(n9947) );
  NAND2_X1 U5529 ( .A1(n7220), .A2(n7219), .ZN(n8569) );
  INV_X1 U5530 ( .A(n4876), .ZN(n4875) );
  NOR2_X1 U5531 ( .A1(n6945), .A2(n9957), .ZN(n7130) );
  AOI21_X1 U5532 ( .B1(n6763), .B2(n7664), .A(n6762), .ZN(n6765) );
  NAND2_X1 U5533 ( .A1(n7653), .A2(n7124), .ZN(n7608) );
  NAND2_X1 U5534 ( .A1(n4913), .A2(n8139), .ZN(n6996) );
  OR2_X1 U5535 ( .A1(n10049), .A2(n8383), .ZN(n6759) );
  NAND2_X1 U5536 ( .A1(n5525), .A2(n5524), .ZN(n8597) );
  NAND2_X1 U5537 ( .A1(n9271), .A2(n5484), .ZN(n5525) );
  NAND2_X1 U5538 ( .A1(n8700), .A2(n5484), .ZN(n5507) );
  NAND2_X1 U5539 ( .A1(n5469), .A2(n5468), .ZN(n8614) );
  OR2_X1 U5540 ( .A1(n9982), .A2(n7627), .ZN(n10049) );
  INV_X1 U5541 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4882) );
  NOR2_X1 U5542 ( .A1(n4885), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4884) );
  CLKBUF_X1 U5543 ( .A(n5586), .Z(n5587) );
  INV_X1 U5544 ( .A(n5543), .ZN(n5544) );
  NAND2_X1 U5545 ( .A1(n5299), .A2(n4953), .ZN(n5329) );
  OR3_X1 U5546 ( .A1(n5245), .A2(P2_IR_REG_10__SCAN_IN), .A3(
        P2_IR_REG_11__SCAN_IN), .ZN(n5263) );
  OR2_X1 U5547 ( .A1(n5172), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5173) );
  NOR2_X1 U5548 ( .A1(n5173), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5211) );
  INV_X1 U5549 ( .A(n5104), .ZN(n4866) );
  NAND2_X1 U5550 ( .A1(n5768), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5784) );
  INV_X1 U5551 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5783) );
  OR2_X1 U5552 ( .A1(n6662), .A2(n5733), .ZN(n5666) );
  AND2_X1 U5553 ( .A1(n8774), .A2(n8716), .ZN(n4512) );
  AND2_X1 U5554 ( .A1(n8774), .A2(n4511), .ZN(n4510) );
  INV_X1 U5555 ( .A(n7334), .ZN(n4506) );
  AND2_X1 U5556 ( .A1(n6178), .A2(n6177), .ZN(n8802) );
  NAND2_X1 U5557 ( .A1(n5964), .A2(n5617), .ZN(n6236) );
  AND2_X1 U5558 ( .A1(n6249), .A2(n6447), .ZN(n6703) );
  INV_X1 U5559 ( .A(n4618), .ZN(n7998) );
  OR2_X1 U5560 ( .A1(n5992), .A2(n8991), .ZN(n6168) );
  NOR2_X1 U5561 ( .A1(n9763), .A2(n4606), .ZN(n9778) );
  AND2_X1 U5562 ( .A1(n9769), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4606) );
  NOR2_X1 U5563 ( .A1(n9778), .A2(n9777), .ZN(n9776) );
  NOR2_X1 U5564 ( .A1(n7252), .A2(n4600), .ZN(n8829) );
  NOR2_X1 U5565 ( .A1(n4601), .A2(n9610), .ZN(n4600) );
  INV_X1 U5566 ( .A(n7256), .ZN(n4601) );
  INV_X1 U5567 ( .A(n8981), .ZN(n4411) );
  NAND2_X1 U5568 ( .A1(n7982), .A2(n7983), .ZN(n8972) );
  NAND2_X1 U5569 ( .A1(n8997), .A2(n9641), .ZN(n4705) );
  AOI21_X1 U5570 ( .B1(n4691), .B2(n8944), .A(n7819), .ZN(n4690) );
  AND2_X1 U5571 ( .A1(n4696), .A2(n4692), .ZN(n4691) );
  NOR3_X1 U5572 ( .A1(n9079), .A2(n9187), .A3(n4589), .ZN(n9026) );
  NAND2_X1 U5573 ( .A1(n9026), .A2(n9010), .ZN(n9004) );
  NAND2_X1 U5574 ( .A1(n6123), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6145) );
  INV_X1 U5575 ( .A(n6104), .ZN(n6105) );
  NAND2_X1 U5576 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n6105), .ZN(n6125) );
  NOR2_X1 U5577 ( .A1(n6069), .A2(n8724), .ZN(n6083) );
  INV_X1 U5578 ( .A(n4665), .ZN(n4664) );
  OAI21_X1 U5579 ( .B1(n4668), .B2(n4675), .A(n8938), .ZN(n4665) );
  NOR2_X1 U5580 ( .A1(n9066), .A2(n9067), .ZN(n9065) );
  NAND2_X1 U5581 ( .A1(n8033), .A2(n9049), .ZN(n9067) );
  AND2_X1 U5582 ( .A1(n9599), .A2(n4586), .ZN(n9117) );
  AND2_X1 U5583 ( .A1(n4329), .A2(n9121), .ZN(n4586) );
  OR2_X1 U5584 ( .A1(n4840), .A2(n4343), .ZN(n4835) );
  INV_X1 U5585 ( .A(n4838), .ZN(n4837) );
  OR2_X1 U5586 ( .A1(n5990), .A2(n8760), .ZN(n6011) );
  NAND2_X1 U5587 ( .A1(n9599), .A2(n4587), .ZN(n9145) );
  NOR2_X1 U5588 ( .A1(n5927), .A2(n7261), .ZN(n5950) );
  AND2_X1 U5589 ( .A1(n7935), .A2(n8932), .ZN(n9588) );
  AND2_X1 U5590 ( .A1(n9606), .A2(n8906), .ZN(n9599) );
  OAI21_X1 U5591 ( .B1(n9626), .B2(n4826), .A(n4824), .ZN(n8905) );
  INV_X1 U5592 ( .A(n4827), .ZN(n4826) );
  AOI21_X1 U5593 ( .B1(n4827), .B2(n4825), .A(n4360), .ZN(n4824) );
  AND2_X1 U5594 ( .A1(n4831), .A2(n4379), .ZN(n4827) );
  OR2_X1 U5595 ( .A1(n5910), .A2(n5909), .ZN(n5927) );
  OR2_X1 U5596 ( .A1(n5848), .A2(n7209), .ZN(n5866) );
  NOR2_X1 U5597 ( .A1(n5866), .A2(n5865), .ZN(n5888) );
  AND2_X1 U5598 ( .A1(n7098), .A2(n7103), .ZN(n4857) );
  NAND2_X1 U5599 ( .A1(n4663), .A2(n7829), .ZN(n7837) );
  NAND2_X1 U5600 ( .A1(n7141), .A2(n4593), .ZN(n7105) );
  AND2_X1 U5601 ( .A1(n7150), .A2(n7041), .ZN(n7043) );
  NAND2_X1 U5602 ( .A1(n7902), .A2(n8040), .ZN(n7042) );
  AND2_X1 U5603 ( .A1(n7141), .A2(n9846), .ZN(n7085) );
  NOR2_X1 U5604 ( .A1(n7047), .A2(n8750), .ZN(n7141) );
  NOR2_X1 U5605 ( .A1(n6878), .A2(n6716), .ZN(n7024) );
  NAND2_X1 U5606 ( .A1(n6691), .A2(n6692), .ZN(n6868) );
  INV_X1 U5607 ( .A(n6243), .ZN(n8072) );
  NAND2_X1 U5608 ( .A1(n6872), .A2(n6666), .ZN(n6878) );
  NAND2_X1 U5609 ( .A1(n7104), .A2(n7103), .ZN(n7276) );
  OR2_X1 U5610 ( .A1(n5806), .A2(n6299), .ZN(n5674) );
  OAI21_X1 U5611 ( .B1(n7877), .B2(n6296), .A(n4351), .ZN(n4535) );
  INV_X1 U5612 ( .A(n9854), .ZN(n9563) );
  XNOR2_X1 U5613 ( .A(n7586), .B(n7585), .ZN(n8152) );
  NAND2_X1 U5614 ( .A1(n7566), .A2(n7565), .ZN(n7571) );
  XNOR2_X1 U5615 ( .A(n5500), .B(n5499), .ZN(n7550) );
  INV_X1 U5616 ( .A(n5405), .ZN(n4631) );
  INV_X1 U5617 ( .A(n4630), .ZN(n4629) );
  OAI21_X1 U5618 ( .B1(n4633), .B2(n4385), .A(n5423), .ZN(n4630) );
  NAND2_X1 U5619 ( .A1(n4648), .A2(n5349), .ZN(n5366) );
  OAI21_X1 U5620 ( .B1(n5019), .B2(n4336), .A(n4622), .ZN(n5298) );
  AOI21_X1 U5621 ( .B1(n4472), .B2(n4475), .A(n4362), .ZN(n4470) );
  CLKBUF_X1 U5622 ( .A(n5883), .Z(n5884) );
  INV_X1 U5623 ( .A(n5601), .ZN(n4858) );
  NAND2_X1 U5624 ( .A1(n4998), .A2(n4997), .ZN(n5209) );
  OR2_X1 U5625 ( .A1(n5807), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5809) );
  OR2_X1 U5626 ( .A1(n5809), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5841) );
  NAND2_X1 U5627 ( .A1(n4468), .A2(n4642), .ZN(n5171) );
  NAND2_X1 U5628 ( .A1(n5142), .A2(n4644), .ZN(n4468) );
  XNOR2_X1 U5629 ( .A(n4980), .B(n4979), .ZN(n5128) );
  INV_X1 U5630 ( .A(SI_5_), .ZN(n4979) );
  NAND2_X1 U5631 ( .A1(n4972), .A2(SI_3_), .ZN(n4973) );
  XNOR2_X1 U5632 ( .A(n4975), .B(SI_4_), .ZN(n5108) );
  NAND2_X1 U5633 ( .A1(n5597), .A2(n5596), .ZN(n5727) );
  NAND2_X1 U5634 ( .A1(n4613), .A2(SI_1_), .ZN(n4967) );
  XNOR2_X1 U5635 ( .A(n5440), .B(n5431), .ZN(n8168) );
  NAND2_X1 U5636 ( .A1(n5094), .A2(n4418), .ZN(n8183) );
  BUF_X1 U5637 ( .A(n7533), .Z(n4398) );
  NAND2_X1 U5638 ( .A1(n8160), .A2(n5519), .ZN(n4757) );
  NAND2_X1 U5639 ( .A1(n4730), .A2(n4728), .ZN(n8195) );
  NAND2_X1 U5640 ( .A1(n4738), .A2(n4741), .ZN(n9903) );
  AND2_X1 U5641 ( .A1(n4742), .A2(n9894), .ZN(n4741) );
  NAND2_X1 U5642 ( .A1(n4743), .A2(n5242), .ZN(n4742) );
  NAND2_X1 U5643 ( .A1(n4750), .A2(n4352), .ZN(n4749) );
  NAND2_X1 U5644 ( .A1(n5192), .A2(n5191), .ZN(n10027) );
  AND4_X1 U5645 ( .A1(n5363), .A2(n5362), .A3(n5361), .A4(n5360), .ZN(n8505)
         );
  AND4_X1 U5646 ( .A1(n5255), .A2(n5254), .A3(n5253), .A4(n5252), .ZN(n7402)
         );
  OR3_X1 U5647 ( .A1(n5570), .A2(n5583), .A3(n5569), .ZN(n9909) );
  AND4_X1 U5648 ( .A1(n5217), .A2(n5216), .A3(n5215), .A4(n5214), .ZN(n7304)
         );
  NAND2_X1 U5649 ( .A1(n7056), .A2(n5222), .ZN(n4745) );
  INV_X1 U5650 ( .A(n4400), .ZN(n8235) );
  OR2_X1 U5651 ( .A1(n7594), .A2(n4422), .ZN(n5074) );
  INV_X1 U5652 ( .A(n9923), .ZN(n8222) );
  NAND2_X1 U5653 ( .A1(n5568), .A2(n5567), .ZN(n9913) );
  AND2_X1 U5654 ( .A1(n5585), .A2(n5584), .ZN(n9892) );
  AND4_X1 U5655 ( .A1(n5292), .A2(n5291), .A3(n5290), .A4(n5289), .ZN(n8092)
         );
  AND4_X1 U5656 ( .A1(n5269), .A2(n5268), .A3(n5267), .A4(n5266), .ZN(n7459)
         );
  NAND2_X1 U5657 ( .A1(n5416), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n4863) );
  NAND2_X1 U5658 ( .A1(n4325), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4862) );
  OR3_X1 U5659 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n5089) );
  NOR2_X1 U5660 ( .A1(n6539), .A2(n4557), .ZN(n6557) );
  AND2_X1 U5661 ( .A1(n6544), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4557) );
  INV_X1 U5662 ( .A(n4556), .ZN(n6555) );
  NOR2_X1 U5663 ( .A1(n6527), .A2(n6526), .ZN(n6525) );
  AND2_X1 U5664 ( .A1(n4556), .A2(n4555), .ZN(n6527) );
  NAND2_X1 U5665 ( .A1(n6560), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4555) );
  INV_X1 U5666 ( .A(n4547), .ZN(n6512) );
  AND2_X1 U5667 ( .A1(n4547), .A2(n4546), .ZN(n6569) );
  NAND2_X1 U5668 ( .A1(n6517), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4546) );
  INV_X1 U5669 ( .A(n4545), .ZN(n6567) );
  AND2_X1 U5670 ( .A1(n4545), .A2(n4544), .ZN(n6491) );
  NAND2_X1 U5671 ( .A1(n6572), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4544) );
  NOR2_X1 U5672 ( .A1(n6611), .A2(n6610), .ZN(n6674) );
  NOR2_X1 U5673 ( .A1(n6607), .A2(n4552), .ZN(n6611) );
  NOR2_X1 U5674 ( .A1(n4554), .A2(n4553), .ZN(n4552) );
  INV_X1 U5675 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n4553) );
  INV_X1 U5676 ( .A(n6608), .ZN(n4554) );
  INV_X1 U5677 ( .A(n4537), .ZN(n8285) );
  AND2_X1 U5678 ( .A1(n4537), .A2(n4536), .ZN(n8288) );
  NAND2_X1 U5679 ( .A1(n8286), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4536) );
  INV_X1 U5680 ( .A(n8294), .ZN(n8293) );
  NAND2_X1 U5681 ( .A1(n7596), .A2(n7595), .ZN(n9542) );
  XNOR2_X1 U5682 ( .A(n8584), .B(n4721), .ZN(n9540) );
  INV_X1 U5683 ( .A(n9542), .ZN(n4721) );
  NAND2_X1 U5684 ( .A1(n4785), .A2(n4788), .ZN(n8345) );
  INV_X1 U5685 ( .A(n8597), .ZN(n8105) );
  NAND2_X1 U5686 ( .A1(n4893), .A2(n4897), .ZN(n8341) );
  NAND2_X1 U5687 ( .A1(n4577), .A2(n4576), .ZN(n8108) );
  NAND2_X1 U5688 ( .A1(n4580), .A2(n7771), .ZN(n8366) );
  INV_X1 U5689 ( .A(n4901), .ZN(n4892) );
  AOI21_X1 U5690 ( .B1(n8379), .B2(n8483), .A(n8378), .ZN(n8610) );
  NAND2_X1 U5691 ( .A1(n4582), .A2(n4806), .ZN(n8377) );
  INV_X1 U5692 ( .A(n8608), .ZN(n8375) );
  OAI21_X1 U5693 ( .B1(n8422), .B2(n4811), .A(n4810), .ZN(n8390) );
  INV_X1 U5694 ( .A(n4457), .ZN(n8388) );
  AND2_X1 U5695 ( .A1(n5392), .A2(n5391), .ZN(n8461) );
  INV_X1 U5696 ( .A(n8638), .ZN(n8474) );
  OAI21_X1 U5697 ( .B1(n8515), .B2(n4484), .A(n4482), .ZN(n8470) );
  NAND2_X1 U5698 ( .A1(n4487), .A2(n4488), .ZN(n8488) );
  NAND2_X1 U5699 ( .A1(n8515), .A2(n4489), .ZN(n4487) );
  AND2_X1 U5700 ( .A1(n5048), .A2(n5047), .ZN(n8511) );
  AND2_X1 U5701 ( .A1(n4491), .A2(n4494), .ZN(n8500) );
  NAND2_X1 U5702 ( .A1(n8515), .A2(n8516), .ZN(n4491) );
  NAND2_X1 U5703 ( .A1(n4797), .A2(n7732), .ZN(n8517) );
  NAND2_X1 U5704 ( .A1(n8560), .A2(n4798), .ZN(n4797) );
  NAND2_X1 U5705 ( .A1(n4906), .A2(n4907), .ZN(n8531) );
  NAND2_X1 U5706 ( .A1(n4320), .A2(n4909), .ZN(n4906) );
  INV_X1 U5707 ( .A(n7464), .ZN(n9960) );
  NOR2_X1 U5708 ( .A1(n4888), .A2(n4887), .ZN(n7227) );
  INV_X1 U5709 ( .A(n7226), .ZN(n4887) );
  NAND2_X1 U5710 ( .A1(n7225), .A2(n8566), .ZN(n10022) );
  NAND2_X1 U5711 ( .A1(n4566), .A2(n7679), .ZN(n7177) );
  NAND2_X1 U5712 ( .A1(n4879), .A2(n7123), .ZN(n7168) );
  OR2_X1 U5713 ( .A1(n7122), .A2(n4376), .ZN(n4879) );
  OR2_X1 U5714 ( .A1(n6768), .A2(n7604), .ZN(n8354) );
  NAND2_X1 U5715 ( .A1(n6637), .A2(n6778), .ZN(n4872) );
  NAND2_X1 U5716 ( .A1(n6768), .A2(n7464), .ZN(n9968) );
  OAI21_X1 U5717 ( .B1(n4709), .B2(n4711), .A(n6466), .ZN(n4712) );
  AND2_X1 U5718 ( .A1(n7589), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4711) );
  INV_X1 U5719 ( .A(n8554), .ZN(n9945) );
  INV_X1 U5720 ( .A(n8354), .ZN(n9951) );
  NOR3_X1 U5721 ( .A1(n4720), .A2(n9541), .A3(n4719), .ZN(n9558) );
  AND2_X1 U5722 ( .A1(n9542), .A2(n10018), .ZN(n4719) );
  NOR2_X1 U5723 ( .A1(n9540), .A2(n10049), .ZN(n4720) );
  OAI21_X1 U5724 ( .B1(n4569), .B2(n4568), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5042) );
  INV_X1 U5725 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U5726 ( .A1(n4519), .A2(n4516), .ZN(n6277) );
  NAND2_X1 U5727 ( .A1(n8700), .A2(n5962), .ZN(n6181) );
  NAND2_X1 U5728 ( .A1(n4766), .A2(n5840), .ZN(n7208) );
  NAND2_X1 U5729 ( .A1(n7156), .A2(n7157), .ZN(n4766) );
  OR2_X1 U5730 ( .A1(n7877), .A2(n6294), .ZN(n5715) );
  AND2_X1 U5731 ( .A1(n6028), .A2(n8791), .ZN(n4773) );
  AND2_X1 U5732 ( .A1(n6246), .A2(n9576), .ZN(n6247) );
  NAND2_X1 U5733 ( .A1(n5880), .A2(n5879), .ZN(n7387) );
  NAND2_X1 U5734 ( .A1(n8766), .A2(n8767), .ZN(n4523) );
  AND2_X1 U5735 ( .A1(n4769), .A2(n9572), .ZN(n8738) );
  AND2_X1 U5736 ( .A1(n4778), .A2(n5766), .ZN(n8746) );
  NAND2_X1 U5737 ( .A1(n6051), .A2(n6050), .ZN(n9205) );
  NAND2_X1 U5738 ( .A1(n6082), .A2(n6081), .ZN(n9197) );
  AOI21_X1 U5739 ( .B1(n4327), .B2(n4764), .A(n4371), .ZN(n4763) );
  NAND2_X1 U5740 ( .A1(n5776), .A2(n4361), .ZN(n8123) );
  AOI21_X1 U5741 ( .B1(n4524), .B2(n4526), .A(n4363), .ZN(n4522) );
  AND2_X1 U5742 ( .A1(n9570), .A2(n9563), .ZN(n8810) );
  OR2_X1 U5743 ( .A1(n6258), .A2(n9691), .ZN(n9568) );
  INV_X1 U5744 ( .A(n8812), .ZN(n9576) );
  INV_X1 U5745 ( .A(n4599), .ZN(n9752) );
  NAND2_X1 U5746 ( .A1(n6404), .A2(n6403), .ZN(n6425) );
  AND2_X1 U5747 ( .A1(n4599), .A2(n4598), .ZN(n6404) );
  NAND2_X1 U5748 ( .A1(n9749), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4598) );
  NAND2_X1 U5749 ( .A1(n6425), .A2(n4597), .ZN(n6427) );
  OR2_X1 U5750 ( .A1(n6429), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4597) );
  NOR2_X1 U5751 ( .A1(n9776), .A2(n4605), .ZN(n6583) );
  AND2_X1 U5752 ( .A1(n9782), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4605) );
  NAND2_X1 U5753 ( .A1(n6583), .A2(n6582), .ZN(n6746) );
  INV_X1 U5754 ( .A(n4602), .ZN(n6833) );
  NAND2_X1 U5755 ( .A1(n4602), .A2(n4392), .ZN(n6835) );
  NOR2_X1 U5756 ( .A1(n8843), .A2(n8844), .ZN(n8847) );
  INV_X1 U5757 ( .A(n4596), .ZN(n8860) );
  NOR2_X1 U5758 ( .A1(n8864), .A2(n8863), .ZN(n8878) );
  AND2_X1 U5759 ( .A1(n4596), .A2(n4595), .ZN(n8864) );
  NAND2_X1 U5760 ( .A1(n8866), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4595) );
  NAND2_X1 U5761 ( .A1(n7879), .A2(n7878), .ZN(n9157) );
  NAND2_X1 U5762 ( .A1(n4846), .A2(n4850), .ZN(n8977) );
  NAND2_X1 U5763 ( .A1(n9003), .A2(n4338), .ZN(n4846) );
  NAND2_X1 U5764 ( .A1(n4693), .A2(n4696), .ZN(n8996) );
  NAND2_X1 U5765 ( .A1(n4695), .A2(n4694), .ZN(n4693) );
  AOI21_X1 U5766 ( .B1(n9003), .B2(n9013), .A(n4852), .ZN(n8989) );
  NAND2_X1 U5767 ( .A1(n9034), .A2(n8942), .ZN(n9022) );
  INV_X1 U5768 ( .A(n8922), .ZN(n9033) );
  NAND2_X1 U5769 ( .A1(n6068), .A2(n6067), .ZN(n9202) );
  NAND2_X1 U5770 ( .A1(n4670), .A2(n4672), .ZN(n9086) );
  NAND2_X1 U5771 ( .A1(n4671), .A2(n4675), .ZN(n4670) );
  AND2_X1 U5772 ( .A1(n4676), .A2(n4348), .ZN(n9102) );
  NAND2_X1 U5773 ( .A1(n4676), .A2(n4675), .ZN(n9100) );
  NAND2_X1 U5774 ( .A1(n4836), .A2(n4839), .ZN(n9109) );
  NAND2_X1 U5775 ( .A1(n9138), .A2(n4841), .ZN(n4836) );
  AOI21_X1 U5776 ( .B1(n9138), .B2(n9137), .A(n4843), .ZN(n9124) );
  NAND2_X1 U5777 ( .A1(n4828), .A2(n4831), .ZN(n9604) );
  NAND2_X1 U5778 ( .A1(n9626), .A2(n4829), .ZN(n4828) );
  NAND2_X1 U5779 ( .A1(n5907), .A2(n5906), .ZN(n9622) );
  NAND2_X1 U5780 ( .A1(n4683), .A2(n4685), .ZN(n7506) );
  INV_X1 U5781 ( .A(n4686), .ZN(n4685) );
  OAI21_X1 U5782 ( .B1(n9626), .B2(n4339), .A(n7369), .ZN(n7501) );
  NAND2_X1 U5783 ( .A1(n5864), .A2(n5863), .ZN(n9650) );
  NAND2_X1 U5784 ( .A1(n5825), .A2(n5824), .ZN(n7319) );
  NAND2_X1 U5785 ( .A1(n7040), .A2(n7039), .ZN(n7152) );
  NAND2_X1 U5786 ( .A1(n6908), .A2(n6907), .ZN(n7020) );
  INV_X1 U5787 ( .A(n9152), .ZN(n9651) );
  INV_X1 U5788 ( .A(n8960), .ZN(n9631) );
  OR2_X1 U5789 ( .A1(n9161), .A2(n9873), .ZN(n4594) );
  NAND2_X1 U5790 ( .A1(n9160), .A2(n9875), .ZN(n4413) );
  NAND2_X1 U5791 ( .A1(n9262), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5640) );
  OR2_X1 U5792 ( .A1(n5641), .A2(n5965), .ZN(n5643) );
  XNOR2_X1 U5793 ( .A(n5442), .B(n5441), .ZN(n7384) );
  OAI21_X1 U5794 ( .B1(n5389), .B2(n4385), .A(n4629), .ZN(n5442) );
  CLKBUF_X1 U5795 ( .A(n6241), .Z(n6242) );
  INV_X1 U5796 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6314) );
  NAND2_X1 U5797 ( .A1(n4643), .A2(n4983), .ZN(n5157) );
  NAND2_X1 U5798 ( .A1(n5142), .A2(n5141), .ZN(n4643) );
  INV_X1 U5799 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6297) );
  INV_X1 U5800 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6294) );
  XNOR2_X1 U5801 ( .A(n5672), .B(n4604), .ZN(n6361) );
  NAND2_X1 U5802 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4604) );
  NOR2_X1 U5803 ( .A1(n9302), .A2(n10106), .ZN(n10105) );
  AOI21_X1 U5804 ( .B1(n4803), .B2(n4804), .A(n4802), .ZN(n4801) );
  INV_X1 U5805 ( .A(n4541), .ZN(n4540) );
  NAND2_X1 U5806 ( .A1(n4539), .A2(n8383), .ZN(n4538) );
  NAND2_X1 U5807 ( .A1(n4543), .A2(n9962), .ZN(n4542) );
  NAND2_X1 U5808 ( .A1(n4425), .A2(n4424), .ZN(P1_U3240) );
  AOI21_X1 U5809 ( .B1(n4428), .B2(n4330), .A(n4397), .ZN(n4424) );
  NAND2_X1 U5810 ( .A1(n4616), .A2(n4426), .ZN(n4425) );
  AOI21_X1 U5811 ( .B1(n9783), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n8892), .ZN(
        n4609) );
  NAND2_X1 U5812 ( .A1(n4611), .A2(n8000), .ZN(n4610) );
  NAND2_X1 U5813 ( .A1(n4608), .A2(n9073), .ZN(n4607) );
  OAI21_X1 U5814 ( .B1(n9168), .B2(n9647), .A(n4699), .ZN(P1_U3263) );
  NAND2_X1 U5815 ( .A1(n4702), .A2(n4701), .ZN(n4700) );
  INV_X1 U5816 ( .A(n8976), .ZN(n4701) );
  AND2_X1 U5817 ( .A1(n4344), .A2(n7633), .ZN(n4322) );
  AND2_X1 U5818 ( .A1(n4708), .A2(n4707), .ZN(n4324) );
  AND2_X1 U5819 ( .A1(n4940), .A2(n8154), .ZN(n4325) );
  OR2_X1 U5820 ( .A1(n8602), .A2(n8242), .ZN(n7633) );
  OR3_X1 U5821 ( .A1(n9004), .A2(n4583), .A3(n9162), .ZN(n4326) );
  AND2_X1 U5822 ( .A1(n4348), .A2(n9101), .ZN(n4675) );
  NOR2_X1 U5823 ( .A1(n5860), .A2(n4765), .ZN(n4327) );
  XNOR2_X1 U5824 ( .A(n5610), .B(n5609), .ZN(n5656) );
  NAND2_X1 U5825 ( .A1(n5296), .A2(n5295), .ZN(n4328) );
  OR2_X1 U5826 ( .A1(n8638), .A2(n8493), .ZN(n7742) );
  INV_X1 U5827 ( .A(n4840), .ZN(n4839) );
  OAI21_X1 U5828 ( .B1(n8914), .B2(n4845), .A(n4331), .ZN(n4840) );
  NAND2_X1 U5829 ( .A1(n7686), .A2(n7687), .ZN(n8566) );
  INV_X1 U5830 ( .A(n8566), .ZN(n8575) );
  AND2_X1 U5831 ( .A1(n4587), .A2(n9126), .ZN(n4329) );
  OR2_X1 U5832 ( .A1(n8076), .A2(n5656), .ZN(n4330) );
  INV_X1 U5833 ( .A(n8414), .ZN(n4813) );
  NAND2_X1 U5834 ( .A1(n7742), .A2(n7750), .ZN(n8476) );
  INV_X1 U5835 ( .A(n8476), .ZN(n4564) );
  OR2_X1 U5836 ( .A1(n9126), .A2(n9144), .ZN(n4331) );
  NOR2_X1 U5837 ( .A1(n4578), .A2(n7560), .ZN(n4332) );
  NAND2_X1 U5838 ( .A1(n6032), .A2(n6031), .ZN(n9210) );
  INV_X1 U5839 ( .A(n4890), .ZN(n4889) );
  NAND2_X1 U5840 ( .A1(n7300), .A2(n7226), .ZN(n4890) );
  AND2_X1 U5841 ( .A1(n8079), .A2(n5656), .ZN(n4333) );
  AND2_X1 U5842 ( .A1(n4324), .A2(n4706), .ZN(n4334) );
  AND2_X1 U5843 ( .A1(n7696), .A2(n7695), .ZN(n7614) );
  AND4_X1 U5844 ( .A1(n5658), .A2(n5616), .A3(n5941), .A4(n5654), .ZN(n4532)
         );
  NAND2_X1 U5845 ( .A1(n7302), .A2(n7690), .ZN(n9936) );
  AND3_X1 U5846 ( .A1(n5438), .A2(n5437), .A3(n5436), .ZN(n8448) );
  NAND2_X1 U5847 ( .A1(n5248), .A2(n5247), .ZN(n9901) );
  INV_X1 U5848 ( .A(n9901), .ZN(n4707) );
  AND2_X1 U5849 ( .A1(n7604), .A2(n7603), .ZN(n4335) );
  AND2_X2 U5850 ( .A1(n6687), .A2(n6354), .ZN(n5696) );
  OR2_X1 U5851 ( .A1(n5313), .A2(n4362), .ZN(n4336) );
  XNOR2_X1 U5852 ( .A(n8608), .B(n8393), .ZN(n8376) );
  INV_X1 U5853 ( .A(n8376), .ZN(n4581) );
  NAND2_X1 U5854 ( .A1(n4866), .A2(n4919), .ZN(n5106) );
  INV_X1 U5855 ( .A(n9172), .ZN(n4584) );
  AND2_X1 U5856 ( .A1(n4853), .A2(n9013), .ZN(n4338) );
  NAND2_X1 U5857 ( .A1(n5412), .A2(n5411), .ZN(n8629) );
  INV_X1 U5858 ( .A(n8340), .ZN(n8107) );
  XNOR2_X1 U5859 ( .A(n8622), .B(n8448), .ZN(n8432) );
  NOR2_X1 U5860 ( .A1(n9650), .A2(n8815), .ZN(n4339) );
  XOR2_X1 U5861 ( .A(n5757), .B(n5718), .Z(n4340) );
  INV_X1 U5862 ( .A(n8231), .ZN(n6634) );
  NAND2_X1 U5863 ( .A1(n4523), .A2(n6139), .ZN(n8730) );
  AND2_X1 U5864 ( .A1(n4907), .A2(n4905), .ZN(n4341) );
  NAND2_X1 U5865 ( .A1(n8117), .A2(n8116), .ZN(n4342) );
  XNOR2_X1 U5866 ( .A(n5006), .B(n5005), .ZN(n5223) );
  AND2_X1 U5867 ( .A1(n9217), .A2(n9104), .ZN(n4343) );
  NAND2_X1 U5868 ( .A1(n8715), .A2(n6049), .ZN(n8773) );
  INV_X1 U5869 ( .A(n9137), .ZN(n4842) );
  AND2_X1 U5870 ( .A1(n4806), .A2(n4581), .ZN(n4344) );
  INV_X1 U5871 ( .A(n7843), .ZN(n4688) );
  OR2_X1 U5872 ( .A1(n6275), .A2(n6410), .ZN(n4345) );
  NAND2_X1 U5873 ( .A1(n5355), .A2(n5354), .ZN(n8645) );
  INV_X1 U5874 ( .A(n8645), .ZN(n4716) );
  AND4_X1 U5875 ( .A1(n4528), .A2(n4532), .A3(n5614), .A4(n4529), .ZN(n4346)
         );
  NOR2_X1 U5876 ( .A1(n5093), .A2(n6293), .ZN(n4347) );
  NAND2_X1 U5877 ( .A1(n8934), .A2(n8935), .ZN(n4348) );
  AND2_X1 U5878 ( .A1(n8978), .A2(n4338), .ZN(n4349) );
  AND2_X1 U5879 ( .A1(n5343), .A2(n5344), .ZN(n4350) );
  INV_X1 U5880 ( .A(n8937), .ZN(n4673) );
  OR2_X1 U5881 ( .A1(n6275), .A2(n6361), .ZN(n4351) );
  AND4_X1 U5882 ( .A1(n5185), .A2(n5184), .A3(n5183), .A4(n5182), .ZN(n7218)
         );
  INV_X1 U5883 ( .A(n7218), .ZN(n4814) );
  INV_X1 U5884 ( .A(n8939), .ZN(n4669) );
  OR2_X1 U5885 ( .A1(n9192), .A2(n9055), .ZN(n8942) );
  INV_X1 U5886 ( .A(n8944), .ZN(n4694) );
  NAND2_X1 U5887 ( .A1(n8031), .A2(n9011), .ZN(n8944) );
  NOR2_X1 U5888 ( .A1(n5325), .A2(n5324), .ZN(n4352) );
  OR2_X1 U5889 ( .A1(n6466), .A2(n9516), .ZN(n4353) );
  AND2_X1 U5890 ( .A1(n6066), .A2(n6065), .ZN(n4354) );
  AND2_X1 U5891 ( .A1(n4757), .A2(n5573), .ZN(n4355) );
  INV_X1 U5892 ( .A(n9162), .ZN(n8955) );
  INV_X1 U5893 ( .A(n7924), .ZN(n4440) );
  NAND2_X1 U5894 ( .A1(n4812), .A2(n7767), .ZN(n4810) );
  AND2_X1 U5895 ( .A1(n8320), .A2(n9927), .ZN(n4356) );
  AND2_X1 U5896 ( .A1(n8791), .A2(n8716), .ZN(n4357) );
  AND2_X1 U5897 ( .A1(n7979), .A2(n4433), .ZN(n4358) );
  AND2_X1 U5898 ( .A1(n7634), .A2(n7635), .ZN(n8099) );
  AND2_X1 U5899 ( .A1(n8511), .A2(n8519), .ZN(n4359) );
  NOR2_X1 U5900 ( .A1(n9665), .A2(n7509), .ZN(n4360) );
  AND2_X1 U5901 ( .A1(n7719), .A2(n7718), .ZN(n7716) );
  AND2_X1 U5902 ( .A1(n5777), .A2(n4345), .ZN(n4361) );
  AND2_X1 U5903 ( .A1(n5021), .A2(SI_14_), .ZN(n4362) );
  AND2_X1 U5904 ( .A1(n6158), .A2(n6157), .ZN(n4363) );
  AND2_X1 U5905 ( .A1(n6796), .A2(n7112), .ZN(n4364) );
  NOR2_X1 U5906 ( .A1(n10027), .A2(n8258), .ZN(n4365) );
  NOR2_X1 U5907 ( .A1(n9004), .A2(n9175), .ZN(n4585) );
  INV_X1 U5908 ( .A(n7500), .ZN(n4834) );
  INV_X1 U5909 ( .A(n4854), .ZN(n4852) );
  NAND2_X1 U5910 ( .A1(n9010), .A2(n9025), .ZN(n4854) );
  NOR2_X1 U5911 ( .A1(n9164), .A2(n9163), .ZN(n4366) );
  NAND2_X1 U5912 ( .A1(n4584), .A2(n8927), .ZN(n4367) );
  NOR2_X1 U5913 ( .A1(n8665), .A2(n8255), .ZN(n4368) );
  NAND2_X1 U5914 ( .A1(n8638), .A2(n8465), .ZN(n4369) );
  INV_X1 U5915 ( .A(n4715), .ZN(n4714) );
  NAND2_X1 U5916 ( .A1(n4717), .A2(n4716), .ZN(n4715) );
  INV_X1 U5917 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5039) );
  NAND2_X1 U5918 ( .A1(n6278), .A2(n4342), .ZN(n4370) );
  INV_X1 U5919 ( .A(n4845), .ZN(n4843) );
  NAND2_X1 U5920 ( .A1(n9227), .A2(n8912), .ZN(n4845) );
  AND2_X1 U5921 ( .A1(n5859), .A2(n7205), .ZN(n4371) );
  OR2_X1 U5922 ( .A1(n9205), .A2(n9069), .ZN(n8938) );
  AND2_X1 U5923 ( .A1(n7767), .A2(n7765), .ZN(n8405) );
  AND2_X1 U5924 ( .A1(n4986), .A2(SI_7_), .ZN(n4372) );
  INV_X1 U5925 ( .A(n8487), .ZN(n8490) );
  AND2_X1 U5926 ( .A1(n7739), .A2(n7741), .ZN(n8487) );
  NOR2_X1 U5927 ( .A1(n4716), .A2(n8505), .ZN(n4373) );
  AND2_X1 U5928 ( .A1(n5073), .A2(n4353), .ZN(n4374) );
  INV_X1 U5929 ( .A(n4772), .ZN(n4507) );
  NAND2_X1 U5930 ( .A1(n8054), .A2(n4832), .ZN(n4375) );
  NOR2_X1 U5931 ( .A1(n8261), .A2(n9957), .ZN(n4376) );
  OR2_X1 U5932 ( .A1(n4492), .A2(n4359), .ZN(n4377) );
  AND2_X1 U5933 ( .A1(n4909), .A2(n4908), .ZN(n4378) );
  OR2_X1 U5934 ( .A1(n9622), .A2(n8814), .ZN(n4379) );
  AND2_X1 U5935 ( .A1(n4638), .A2(n5223), .ZN(n4380) );
  AND3_X1 U5936 ( .A1(n4748), .A2(n4328), .A3(n4746), .ZN(n4381) );
  INV_X1 U5937 ( .A(n9192), .ZN(n8920) );
  NAND2_X1 U5938 ( .A1(n6102), .A2(n6101), .ZN(n9192) );
  AND2_X1 U5939 ( .A1(n4884), .A2(n4882), .ZN(n4382) );
  NOR2_X1 U5940 ( .A1(n4894), .A2(n8342), .ZN(n4383) );
  INV_X1 U5941 ( .A(n7664), .ZN(n6755) );
  NAND2_X1 U5942 ( .A1(n6009), .A2(n6008), .ZN(n9217) );
  AND2_X1 U5943 ( .A1(n4728), .A2(n4727), .ZN(n4384) );
  INV_X1 U5944 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4932) );
  INV_X1 U5945 ( .A(n9128), .ZN(n9647) );
  NAND2_X1 U5946 ( .A1(n5265), .A2(n5264), .ZN(n7411) );
  INV_X1 U5947 ( .A(n7411), .ZN(n4706) );
  OR2_X1 U5948 ( .A1(n5424), .A2(n4631), .ZN(n4385) );
  NAND2_X1 U5949 ( .A1(n4745), .A2(n7055), .ZN(n7058) );
  INV_X1 U5950 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4422) );
  NAND2_X1 U5951 ( .A1(n5507), .A2(n5506), .ZN(n8602) );
  INV_X1 U5952 ( .A(n8602), .ZN(n4900) );
  NOR2_X1 U5953 ( .A1(n4320), .A2(n4910), .ZN(n4386) );
  NAND2_X1 U5954 ( .A1(n5988), .A2(n5987), .ZN(n9222) );
  OR2_X1 U5955 ( .A1(n9533), .A2(n9532), .ZN(n4387) );
  NAND2_X1 U5956 ( .A1(n5947), .A2(n5946), .ZN(n9595) );
  NAND2_X1 U5957 ( .A1(n4770), .A2(n5961), .ZN(n9572) );
  NAND2_X1 U5958 ( .A1(n7397), .A2(n4873), .ZN(n7455) );
  NAND2_X1 U5959 ( .A1(n9599), .A2(n4329), .ZN(n4588) );
  NAND2_X1 U5960 ( .A1(n8541), .A2(n4714), .ZN(n4718) );
  INV_X1 U5961 ( .A(n4591), .ZN(n9071) );
  NOR2_X1 U5962 ( .A1(n9079), .A2(n9202), .ZN(n4591) );
  AND2_X1 U5963 ( .A1(n4906), .A2(n4341), .ZN(n4388) );
  NAND2_X1 U5964 ( .A1(n5430), .A2(n5429), .ZN(n8622) );
  INV_X1 U5965 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n4603) );
  AND2_X1 U5966 ( .A1(n7401), .A2(n7710), .ZN(n4389) );
  AND2_X1 U5967 ( .A1(n5456), .A2(n5455), .ZN(n8392) );
  INV_X1 U5968 ( .A(n8392), .ZN(n4459) );
  AND3_X1 U5969 ( .A1(n7141), .A2(n4593), .A3(n7106), .ZN(n4390) );
  NAND2_X1 U5970 ( .A1(n5822), .A2(n7192), .ZN(n7156) );
  AND2_X1 U5971 ( .A1(n9949), .A2(n4708), .ZN(n4391) );
  INV_X1 U5972 ( .A(n4909), .ZN(n8557) );
  XNOR2_X1 U5973 ( .A(n8665), .B(n8538), .ZN(n4909) );
  NAND2_X1 U5974 ( .A1(n4776), .A2(n4778), .ZN(n8747) );
  NAND2_X1 U5975 ( .A1(n10022), .A2(n4889), .ZN(n7306) );
  OR2_X1 U5976 ( .A1(n6832), .A2(n6831), .ZN(n4392) );
  NAND2_X1 U5977 ( .A1(n4931), .A2(n5299), .ZN(n5546) );
  AND2_X1 U5978 ( .A1(n6277), .A2(n6278), .ZN(n4393) );
  INV_X1 U5979 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4783) );
  AND2_X1 U5980 ( .A1(n5880), .A2(n4772), .ZN(n4394) );
  AND2_X1 U5981 ( .A1(n7573), .A2(n9362), .ZN(n4395) );
  AND3_X1 U5982 ( .A1(n4531), .A2(n5614), .A3(n5613), .ZN(n4396) );
  INV_X1 U5983 ( .A(n5904), .ZN(n4505) );
  INV_X1 U5984 ( .A(n4494), .ZN(n4492) );
  NAND2_X1 U5985 ( .A1(n8528), .A2(n8536), .ZN(n4494) );
  INV_X1 U5986 ( .A(n9585), .ZN(n9641) );
  NAND2_X1 U5987 ( .A1(n6242), .A2(n9073), .ZN(n7995) );
  OR2_X1 U5988 ( .A1(n6243), .A2(n8078), .ZN(n6687) );
  OAI21_X1 U5989 ( .B1(n6779), .B2(n6637), .A(n7659), .ZN(n6763) );
  INV_X1 U5990 ( .A(n8142), .ZN(n6997) );
  NAND2_X1 U5991 ( .A1(n4872), .A2(n6635), .ZN(n6756) );
  NOR2_X1 U5992 ( .A1(n8089), .A2(n8088), .ZN(n4397) );
  INV_X1 U5993 ( .A(n5656), .ZN(n8078) );
  INV_X1 U5994 ( .A(n8000), .ZN(n9073) );
  NOR2_X1 U5995 ( .A1(n6337), .A2(P2_U3152), .ZN(n7811) );
  AOI21_X1 U5996 ( .B1(n9165), .B2(n9147), .A(n4700), .ZN(n4699) );
  NAND2_X1 U5997 ( .A1(n4615), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4614) );
  NAND2_X1 U5998 ( .A1(n5275), .A2(n7240), .ZN(n7243) );
  NAND2_X1 U5999 ( .A1(n5691), .A2(n5595), .ZN(n5725) );
  INV_X1 U6000 ( .A(n5883), .ZN(n5618) );
  NAND2_X1 U6001 ( .A1(n5639), .A2(n5636), .ZN(n5633) );
  NAND2_X1 U6002 ( .A1(n5633), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5634) );
  NOR2_X1 U6003 ( .A1(n9140), .A2(n8933), .ZN(n9132) );
  XNOR2_X2 U6004 ( .A(n8823), .B(n6716), .ZN(n8043) );
  XNOR2_X1 U6005 ( .A(n8952), .B(n8951), .ZN(n4412) );
  NOR2_X2 U6006 ( .A1(n4400), .A2(n4399), .ZN(n4737) );
  NAND2_X4 U6007 ( .A1(n5586), .A2(n8701), .ZN(n6466) );
  NAND2_X1 U6008 ( .A1(n6789), .A2(n5114), .ZN(n6794) );
  NAND2_X1 U6009 ( .A1(n5476), .A2(n8203), .ZN(n4417) );
  NAND2_X1 U6010 ( .A1(n4417), .A2(n8202), .ZN(n4401) );
  NAND2_X2 U6011 ( .A1(n7815), .A2(n9962), .ZN(n7806) );
  NOR2_X2 U6012 ( .A1(n7515), .A2(n4350), .ZN(n7533) );
  NAND2_X1 U6013 ( .A1(n8916), .A2(n4914), .ZN(n9064) );
  NAND2_X1 U6014 ( .A1(n9048), .A2(n8918), .ZN(n4416) );
  XNOR2_X1 U6015 ( .A(n5634), .B(n5637), .ZN(n6256) );
  NAND2_X1 U6016 ( .A1(n8205), .A2(n5477), .ZN(n4402) );
  NAND2_X1 U6017 ( .A1(n7722), .A2(n4403), .ZN(n7726) );
  NAND3_X1 U6018 ( .A1(n7776), .A2(n7777), .A3(n7775), .ZN(n7786) );
  NAND2_X1 U6019 ( .A1(n4408), .A2(n7763), .ZN(n7766) );
  NAND3_X1 U6020 ( .A1(n7761), .A2(n8425), .A3(n7762), .ZN(n4408) );
  OR2_X2 U6021 ( .A1(n7815), .A2(n7631), .ZN(n7797) );
  NAND2_X1 U6022 ( .A1(n4689), .A2(n4690), .ZN(n8979) );
  INV_X2 U6023 ( .A(n5673), .ZN(n6292) );
  INV_X1 U6024 ( .A(n5673), .ZN(n4710) );
  NOR2_X2 U6025 ( .A1(n9614), .A2(n7507), .ZN(n8931) );
  NAND3_X1 U6026 ( .A1(n4366), .A2(n4413), .A3(n4594), .ZN(n9244) );
  NAND2_X2 U6027 ( .A1(n7269), .A2(n7916), .ZN(n7371) );
  NAND2_X1 U6028 ( .A1(n6985), .A2(n6987), .ZN(n6986) );
  AND2_X2 U6029 ( .A1(n4567), .A2(n5299), .ZN(n5543) );
  INV_X2 U6030 ( .A(n5356), .ZN(n4414) );
  NAND2_X2 U6031 ( .A1(n4374), .A2(n5074), .ZN(n8231) );
  OAI22_X2 U6032 ( .A1(n9020), .A2(n8925), .B1(n9037), .B2(n9187), .ZN(n9003)
         );
  NAND3_X1 U6033 ( .A1(n7040), .A2(n7039), .A3(n7144), .ZN(n7150) );
  AND2_X2 U6034 ( .A1(n5112), .A2(n5097), .ZN(n8176) );
  NOR2_X1 U6035 ( .A1(n4347), .A2(n4419), .ZN(n4418) );
  NOR2_X1 U6036 ( .A1(n6466), .A2(n6290), .ZN(n4419) );
  NAND2_X1 U6037 ( .A1(n9533), .A2(n4381), .ZN(n4747) );
  NAND2_X1 U6038 ( .A1(n4931), .A2(n4570), .ZN(n4569) );
  XNOR2_X1 U6039 ( .A(n5040), .B(n5039), .ZN(n5586) );
  XNOR2_X1 U6040 ( .A(n4420), .B(n9427), .ZN(n5071) );
  INV_X1 U6041 ( .A(n8077), .ZN(n4423) );
  NOR2_X1 U6042 ( .A1(n4423), .A2(n4427), .ZN(n4426) );
  NOR2_X1 U6043 ( .A1(n8090), .A2(n4333), .ZN(n4428) );
  NAND2_X1 U6044 ( .A1(n7968), .A2(n4432), .ZN(n4429) );
  NAND2_X1 U6045 ( .A1(n4429), .A2(n4430), .ZN(n7985) );
  NAND2_X1 U6046 ( .A1(n5142), .A2(n4464), .ZN(n4463) );
  NAND2_X1 U6047 ( .A1(n5244), .A2(n4472), .ZN(n4469) );
  NAND2_X1 U6048 ( .A1(n4469), .A2(n4470), .ZN(n5314) );
  NAND2_X1 U6049 ( .A1(n4321), .A2(n7438), .ZN(n4496) );
  NAND3_X1 U6050 ( .A1(n6028), .A2(n8791), .A3(n4512), .ZN(n4508) );
  NAND2_X1 U6051 ( .A1(n4508), .A2(n4509), .ZN(n8722) );
  INV_X1 U6052 ( .A(n6049), .ZN(n4511) );
  INV_X1 U6053 ( .A(n6278), .ZN(n4515) );
  OAI21_X2 U6054 ( .B1(n8119), .B2(n4370), .A(n4513), .ZN(n5818) );
  NAND2_X1 U6055 ( .A1(n8766), .A2(n4524), .ZN(n4521) );
  NAND2_X1 U6056 ( .A1(n4521), .A2(n4522), .ZN(n8801) );
  AND2_X1 U6057 ( .A1(n4531), .A2(n5614), .ZN(n4527) );
  AND3_X1 U6058 ( .A1(n4530), .A2(n4532), .A3(n4527), .ZN(n4822) );
  NAND3_X1 U6059 ( .A1(n8782), .A2(n6100), .A3(n6115), .ZN(n8706) );
  XNOR2_X2 U6060 ( .A(n4533), .B(n5629), .ZN(n6355) );
  INV_X1 U6061 ( .A(n4535), .ZN(n4534) );
  NAND2_X1 U6062 ( .A1(n7835), .A2(n5696), .ZN(n5675) );
  NAND3_X1 U6063 ( .A1(n4542), .A2(n4540), .A3(n4538), .ZN(P2_U3264) );
  OAI21_X1 U6064 ( .B1(n8491), .B2(n4562), .A(n4561), .ZN(n8464) );
  NAND2_X1 U6065 ( .A1(n8491), .A2(n4561), .ZN(n4560) );
  NAND2_X1 U6066 ( .A1(n4566), .A2(n4565), .ZN(n7220) );
  INV_X1 U6067 ( .A(n4569), .ZN(n4567) );
  NAND2_X1 U6068 ( .A1(n5299), .A2(n4932), .ZN(n4568) );
  NOR2_X1 U6069 ( .A1(n8503), .A2(n8502), .ZN(n8501) );
  OR2_X1 U6070 ( .A1(n4805), .A2(n4323), .ZN(n4582) );
  NAND2_X1 U6071 ( .A1(n4805), .A2(n4322), .ZN(n4577) );
  NAND2_X1 U6072 ( .A1(n4582), .A2(n4344), .ZN(n4580) );
  INV_X1 U6073 ( .A(n4585), .ZN(n8990) );
  INV_X1 U6074 ( .A(n4588), .ZN(n9125) );
  NAND3_X1 U6075 ( .A1(n4610), .A2(n4609), .A3(n4607), .ZN(P1_U3260) );
  XNOR2_X1 U6076 ( .A(n4613), .B(n9437), .ZN(n5066) );
  NAND2_X1 U6077 ( .A1(n5019), .A2(n4622), .ZN(n4621) );
  NAND2_X1 U6078 ( .A1(n5019), .A2(n5018), .ZN(n5278) );
  NAND2_X1 U6079 ( .A1(n5389), .A2(n4629), .ZN(n4628) );
  NAND2_X1 U6080 ( .A1(n4998), .A2(n4380), .ZN(n4635) );
  NAND2_X1 U6081 ( .A1(n4635), .A2(n4636), .ZN(n5244) );
  NAND3_X1 U6082 ( .A1(n4638), .A2(n4641), .A3(n5223), .ZN(n4637) );
  NAND2_X1 U6083 ( .A1(n7566), .A2(n4652), .ZN(n4649) );
  OAI21_X1 U6084 ( .B1(n7566), .B2(n4654), .A(n4652), .ZN(n7586) );
  NAND2_X1 U6085 ( .A1(n4649), .A2(n4650), .ZN(n7588) );
  OAI21_X1 U6086 ( .B1(n5461), .B2(n4662), .A(n5464), .ZN(n5480) );
  NAND2_X1 U6087 ( .A1(n5461), .A2(n4660), .ZN(n4659) );
  XNOR2_X1 U6088 ( .A(n5480), .B(n5479), .ZN(n7523) );
  NAND3_X1 U6089 ( .A1(n4663), .A2(n7829), .A3(n7096), .ZN(n7097) );
  NAND2_X1 U6090 ( .A1(n9132), .A2(n4667), .ZN(n4666) );
  INV_X1 U6091 ( .A(n4668), .ZN(n4667) );
  INV_X1 U6092 ( .A(n9132), .ZN(n4671) );
  NAND2_X1 U6093 ( .A1(n4666), .A2(n4664), .ZN(n9066) );
  OAI21_X1 U6094 ( .B1(n7841), .B2(n4677), .A(n7851), .ZN(n4686) );
  AOI21_X1 U6095 ( .B1(n4682), .B2(n4680), .A(n4679), .ZN(n4678) );
  INV_X1 U6096 ( .A(n4682), .ZN(n4681) );
  NAND2_X1 U6097 ( .A1(n9034), .A2(n4691), .ZN(n4689) );
  NOR2_X2 U6098 ( .A1(n8380), .A2(n8602), .ZN(n8362) );
  NAND2_X1 U6099 ( .A1(n4334), .A2(n9949), .ZN(n8101) );
  NOR2_X2 U6100 ( .A1(n6846), .A2(n8231), .ZN(n6781) );
  NAND2_X2 U6101 ( .A1(n6466), .A2(n5673), .ZN(n5093) );
  INV_X1 U6102 ( .A(n4718), .ZN(n8494) );
  NOR2_X2 U6103 ( .A1(n8352), .A2(n8587), .ZN(n8584) );
  NAND2_X1 U6104 ( .A1(n4730), .A2(n4384), .ZN(n4722) );
  OAI21_X1 U6105 ( .B1(n4398), .B2(n7529), .A(n7530), .ZN(n8221) );
  NAND2_X1 U6106 ( .A1(n4737), .A2(n8233), .ZN(n8234) );
  AND2_X2 U6107 ( .A1(n4736), .A2(n4734), .ZN(n6789) );
  NAND2_X1 U6108 ( .A1(n8176), .A2(n4735), .ZN(n4734) );
  INV_X1 U6109 ( .A(n5083), .ZN(n4735) );
  NAND3_X1 U6110 ( .A1(n4737), .A2(n8176), .A3(n8233), .ZN(n4736) );
  INV_X1 U6111 ( .A(n7055), .ZN(n4743) );
  NAND2_X1 U6112 ( .A1(n6986), .A2(n4739), .ZN(n4738) );
  INV_X1 U6113 ( .A(n5324), .ZN(n4746) );
  NAND2_X2 U6114 ( .A1(n7450), .A2(n7449), .ZN(n7514) );
  NAND2_X1 U6115 ( .A1(n5440), .A2(n4753), .ZN(n4752) );
  OAI21_X2 U6116 ( .B1(n5440), .B2(n4754), .A(n4752), .ZN(n5458) );
  NAND2_X1 U6117 ( .A1(n8213), .A2(n8212), .ZN(n5460) );
  OAI21_X1 U6118 ( .B1(n4355), .B2(n4756), .A(n5594), .ZN(P2_U3222) );
  OAI21_X1 U6119 ( .B1(n4757), .B2(n5537), .A(n5574), .ZN(n4756) );
  XNOR2_X2 U6120 ( .A(n5539), .B(n5538), .ZN(n8113) );
  OAI21_X2 U6121 ( .B1(n4962), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5539) );
  AND2_X2 U6122 ( .A1(n4925), .A2(n5139), .ZN(n5299) );
  NAND2_X1 U6123 ( .A1(n6100), .A2(n8782), .ZN(n6118) );
  NAND3_X1 U6124 ( .A1(n5822), .A2(n4327), .A3(n7192), .ZN(n4762) );
  NAND2_X2 U6125 ( .A1(n4762), .A2(n4763), .ZN(n7335) );
  INV_X1 U6126 ( .A(n7539), .ZN(n4768) );
  NAND2_X1 U6127 ( .A1(n9573), .A2(n9574), .ZN(n4769) );
  NOR2_X1 U6128 ( .A1(n4768), .A2(n5961), .ZN(n4767) );
  NAND3_X1 U6129 ( .A1(n4769), .A2(n8739), .A3(n9572), .ZN(n8737) );
  INV_X1 U6130 ( .A(n6687), .ZN(n4771) );
  OAI21_X1 U6131 ( .B1(n8716), .B2(n4773), .A(n8715), .ZN(n8717) );
  NAND2_X1 U6132 ( .A1(n4775), .A2(n6080), .ZN(n6099) );
  NAND2_X1 U6133 ( .A1(n4775), .A2(n4774), .ZN(n8781) );
  NAND2_X2 U6134 ( .A1(n5759), .A2(n5758), .ZN(n4778) );
  NAND2_X1 U6135 ( .A1(n5766), .A2(n8748), .ZN(n4777) );
  NAND3_X1 U6136 ( .A1(n5881), .A2(n5604), .A3(n4779), .ZN(n5657) );
  NAND3_X1 U6137 ( .A1(n5881), .A2(n5604), .A3(n4781), .ZN(n4780) );
  NAND2_X1 U6138 ( .A1(n5129), .A2(n5128), .ZN(n4784) );
  NAND2_X1 U6139 ( .A1(n4790), .A2(n4788), .ZN(n4787) );
  NAND2_X1 U6140 ( .A1(n8560), .A2(n7557), .ZN(n8533) );
  INV_X1 U6141 ( .A(n7557), .ZN(n4799) );
  NAND2_X1 U6142 ( .A1(n4800), .A2(n4801), .ZN(P2_U3244) );
  NAND2_X1 U6143 ( .A1(n7605), .A2(n4803), .ZN(n4800) );
  INV_X1 U6144 ( .A(n8422), .ZN(n4805) );
  NAND3_X1 U6145 ( .A1(n7302), .A2(n7690), .A3(n7614), .ZN(n9937) );
  NAND2_X1 U6146 ( .A1(n9937), .A2(n7696), .ZN(n7352) );
  INV_X2 U6147 ( .A(n5043), .ZN(n5673) );
  NAND2_X1 U6148 ( .A1(n5043), .A2(SI_0_), .ZN(n5625) );
  NOR2_X2 U6149 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5691) );
  NAND2_X1 U6150 ( .A1(n5618), .A2(n4346), .ZN(n5628) );
  NOR2_X1 U6151 ( .A1(n8905), .A2(n4833), .ZN(n8908) );
  XNOR2_X2 U6152 ( .A(n8825), .B(n6872), .ZN(n6692) );
  NAND2_X1 U6153 ( .A1(n6870), .A2(n6907), .ZN(n4856) );
  NAND3_X1 U6154 ( .A1(n4856), .A2(n4855), .A3(n7019), .ZN(n7018) );
  NAND2_X1 U6155 ( .A1(n8043), .A2(n6907), .ZN(n4855) );
  NAND2_X1 U6156 ( .A1(n7104), .A2(n4857), .ZN(n7279) );
  NAND4_X1 U6157 ( .A1(n5601), .A2(n5597), .A3(n5611), .A4(n4859), .ZN(n5883)
         );
  NAND2_X1 U6158 ( .A1(n5597), .A2(n4859), .ZN(n4861) );
  NOR2_X2 U6159 ( .A1(n4858), .A2(n4861), .ZN(n5881) );
  INV_X1 U6160 ( .A(n4861), .ZN(n5774) );
  NAND4_X1 U6161 ( .A1(n4865), .A2(n4864), .A3(n4863), .A4(n4862), .ZN(n6842)
         );
  NAND2_X1 U6162 ( .A1(n4337), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4864) );
  NAND2_X1 U6163 ( .A1(n5084), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n4865) );
  NOR2_X2 U6164 ( .A1(n5104), .A2(n4867), .ZN(n5139) );
  NAND2_X1 U6165 ( .A1(n4871), .A2(n4869), .ZN(n6942) );
  NAND3_X1 U6166 ( .A1(n6637), .A2(n6778), .A3(n6755), .ZN(n4871) );
  NAND2_X1 U6167 ( .A1(n4877), .A2(n4875), .ZN(n7221) );
  OAI21_X1 U6168 ( .B1(n7167), .B2(n4880), .A(n7166), .ZN(n4876) );
  NAND2_X1 U6169 ( .A1(n7122), .A2(n4878), .ZN(n4877) );
  NAND2_X1 U6170 ( .A1(n5543), .A2(n4884), .ZN(n4937) );
  AND2_X2 U6171 ( .A1(n5543), .A2(n4382), .ZN(n4936) );
  NAND2_X1 U6172 ( .A1(n4891), .A2(n4383), .ZN(n8344) );
  NAND2_X1 U6173 ( .A1(n8374), .A2(n4895), .ZN(n4891) );
  NAND2_X1 U6174 ( .A1(n8374), .A2(n4896), .ZN(n4893) );
  AOI21_X1 U6175 ( .B1(n8374), .B2(n8376), .A(n4892), .ZN(n8361) );
  NAND2_X1 U6176 ( .A1(n4320), .A2(n4378), .ZN(n4904) );
  OR2_X1 U6177 ( .A1(n8143), .A2(n6245), .ZN(n6272) );
  NAND2_X1 U6178 ( .A1(n5680), .A2(n5681), .ZN(n6727) );
  NAND2_X1 U6179 ( .A1(n6027), .A2(n6026), .ZN(n8791) );
  INV_X1 U6180 ( .A(n6024), .ZN(n6027) );
  INV_X4 U6181 ( .A(n5746), .ZN(n6316) );
  INV_X1 U6182 ( .A(n9268), .ZN(n5648) );
  NAND4_X4 U6183 ( .A1(n5671), .A2(n5670), .A3(n5669), .A4(n5668), .ZN(n8825)
         );
  NOR2_X1 U6184 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4918) );
  OR2_X1 U6185 ( .A1(n5038), .A2(n4933), .ZN(n5040) );
  OAI222_X1 U6186 ( .A1(n8695), .A2(n8156), .B1(P2_U3152), .B2(n8154), .C1(
        n8153), .C2(n8704), .ZN(P2_U3328) );
  MUX2_X2 U6187 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8705), .S(n6466), .Z(n8139) );
  AOI21_X2 U6188 ( .B1(n8801), .B2(n8803), .A(n8802), .ZN(n8145) );
  INV_X1 U6189 ( .A(n7716), .ZN(n7398) );
  OR2_X1 U6190 ( .A1(n6466), .A2(n6477), .ZN(n4912) );
  INV_X1 U6191 ( .A(n8343), .ZN(n8346) );
  AND2_X1 U6192 ( .A1(n8443), .A2(n8444), .ZN(n4916) );
  AND3_X1 U6193 ( .A1(n5419), .A2(n5418), .A3(n5417), .ZN(n8196) );
  AND3_X1 U6194 ( .A1(n5400), .A2(n5399), .A3(n5398), .ZN(n8447) );
  OR2_X1 U6195 ( .A1(n5422), .A2(n5421), .ZN(n4917) );
  INV_X1 U6196 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5616) );
  INV_X1 U6197 ( .A(n6117), .ZN(n6115) );
  INV_X1 U6198 ( .A(n6098), .ZN(n6094) );
  AOI21_X1 U6199 ( .B1(n5763), .B2(n5762), .A(n4340), .ZN(n5764) );
  INV_X1 U6200 ( .A(n5434), .ZN(n5432) );
  INV_X1 U6201 ( .A(n8196), .ZN(n8096) );
  OR2_X1 U6202 ( .A1(n8665), .A2(n8538), .ZN(n7557) );
  INV_X1 U6203 ( .A(n7650), .ZN(n6762) );
  INV_X1 U6204 ( .A(n5819), .ZN(n5820) );
  INV_X1 U6205 ( .A(n6217), .ZN(n6199) );
  INV_X1 U6206 ( .A(n8972), .ZN(n8949) );
  INV_X1 U6207 ( .A(n6125), .ZN(n6123) );
  INV_X1 U6208 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5826) );
  AND2_X1 U6209 ( .A1(n9162), .A2(n9563), .ZN(n9163) );
  AND2_X1 U6210 ( .A1(n5603), .A2(n5611), .ZN(n5604) );
  INV_X1 U6211 ( .A(SI_9_), .ZN(n9440) );
  INV_X1 U6212 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5596) );
  INV_X1 U6213 ( .A(n8694), .ZN(n4940) );
  NAND2_X1 U6214 ( .A1(n4945), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6215 ( .A1(n8093), .A2(n8481), .ZN(n8094) );
  INV_X1 U6216 ( .A(n8405), .ZN(n8413) );
  NAND2_X1 U6217 ( .A1(n7642), .A2(n7648), .ZN(n6779) );
  NAND2_X1 U6218 ( .A1(n5821), .A2(n5820), .ZN(n7192) );
  AOI21_X1 U6219 ( .B1(n6199), .B2(n6930), .A(n5635), .ZN(n5662) );
  INV_X1 U6220 ( .A(n6025), .ZN(n6026) );
  NAND2_X1 U6221 ( .A1(n6162), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6204) );
  OR2_X1 U6222 ( .A1(n6052), .A2(n8775), .ZN(n6069) );
  INV_X1 U6223 ( .A(n9187), .ZN(n8924) );
  AOI21_X1 U6224 ( .B1(n9581), .B2(n8932), .A(n9137), .ZN(n9140) );
  AND2_X1 U6225 ( .A1(n7849), .A2(n7840), .ZN(n9611) );
  NAND2_X1 U6226 ( .A1(n6915), .A2(n6914), .ZN(n8005) );
  NAND2_X1 U6227 ( .A1(n5001), .A2(n9354), .ZN(n5004) );
  INV_X1 U6228 ( .A(n8159), .ZN(n5517) );
  INV_X1 U6229 ( .A(n5439), .ZN(n5431) );
  OR2_X1 U6230 ( .A1(n5470), .A2(n8207), .ZN(n5488) );
  NOR2_X1 U6231 ( .A1(n8157), .A2(n5496), .ZN(n5497) );
  INV_X1 U6232 ( .A(n8327), .ZN(n8591) );
  INV_X1 U6233 ( .A(n6769), .ZN(n9999) );
  AND2_X1 U6234 ( .A1(n7806), .A2(n7603), .ZN(n9939) );
  NOR2_X1 U6235 ( .A1(n5784), .A2(n5783), .ZN(n5800) );
  NOR2_X1 U6236 ( .A1(n6011), .A2(n6010), .ZN(n6033) );
  INV_X1 U6237 ( .A(n4317), .ZN(n6200) );
  INV_X1 U6238 ( .A(n9166), .ZN(n8971) );
  INV_X1 U6239 ( .A(n9180), .ZN(n9010) );
  INV_X1 U6240 ( .A(n8919), .ZN(n9055) );
  INV_X1 U6241 ( .A(n8814), .ZN(n7509) );
  AND3_X1 U6242 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5768) );
  OR2_X1 U6243 ( .A1(n7999), .A2(n9691), .ZN(n9583) );
  AND2_X1 U6244 ( .A1(n6690), .A2(n6689), .ZN(n9864) );
  OR2_X1 U6245 ( .A1(n6927), .A2(n6926), .ZN(n9854) );
  NOR2_X1 U6246 ( .A1(n8242), .A2(n9916), .ZN(n5592) );
  OR2_X1 U6247 ( .A1(n8196), .A2(n5534), .ZN(n5420) );
  INV_X1 U6248 ( .A(n9913), .ZN(n9902) );
  INV_X1 U6249 ( .A(n9909), .ZN(n9893) );
  AND2_X1 U6250 ( .A1(n5533), .A2(n5532), .ZN(n8368) );
  AND4_X1 U6251 ( .A1(n5306), .A2(n5305), .A3(n5304), .A4(n5303), .ZN(n8520)
         );
  AND2_X1 U6252 ( .A1(n6468), .A2(n6467), .ZN(n9924) );
  OAI21_X1 U6253 ( .B1(n8351), .B2(n9939), .A(n8350), .ZN(n8594) );
  INV_X1 U6254 ( .A(n8099), .ZN(n8389) );
  INV_X1 U6255 ( .A(n8535), .ZN(n8480) );
  NOR2_X1 U6256 ( .A1(n9974), .A2(n5550), .ZN(n6643) );
  INV_X1 U6257 ( .A(n10054), .ZN(n9983) );
  AND2_X1 U6258 ( .A1(n6449), .A2(n9979), .ZN(n9972) );
  AND2_X1 U6259 ( .A1(n5176), .A2(n5175), .ZN(n6572) );
  INV_X1 U6260 ( .A(n9568), .ZN(n8806) );
  INV_X1 U6261 ( .A(n9580), .ZN(n8798) );
  AND2_X1 U6262 ( .A1(n5950), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5971) );
  OR2_X1 U6263 ( .A1(n5992), .A2(n8146), .ZN(n6185) );
  OR2_X1 U6264 ( .A1(n5746), .A2(n5684), .ZN(n5690) );
  AND2_X1 U6265 ( .A1(n8942), .A2(n8032), .ZN(n9035) );
  INV_X1 U6266 ( .A(n9643), .ZN(n9613) );
  OR3_X1 U6267 ( .A1(n9658), .A2(n8072), .A3(n8084), .ZN(n9633) );
  INV_X1 U6268 ( .A(n9149), .ZN(n9128) );
  OR2_X1 U6269 ( .A1(n6927), .A2(n8078), .ZN(n9873) );
  INV_X1 U6270 ( .A(n9875), .ZN(n9240) );
  AND2_X1 U6271 ( .A1(n6222), .A2(n6223), .ZN(n6443) );
  INV_X1 U6272 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5790) );
  NOR2_X1 U6273 ( .A1(n9290), .A2(n9289), .ZN(n10122) );
  OR3_X1 U6274 ( .A1(n7496), .A2(n7552), .A3(n7524), .ZN(n6449) );
  NOR2_X1 U6275 ( .A1(n5593), .A2(n5592), .ZN(n5594) );
  INV_X1 U6276 ( .A(n8617), .ZN(n8411) );
  AND4_X1 U6277 ( .A1(n5339), .A2(n5338), .A3(n5337), .A4(n5336), .ZN(n8536)
         );
  AND2_X1 U6278 ( .A1(n6341), .A2(n6340), .ZN(n8325) );
  INV_X1 U6279 ( .A(n10077), .ZN(n10075) );
  INV_X1 U6280 ( .A(n10057), .ZN(n10055) );
  AND2_X1 U6281 ( .A1(n6337), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9979) );
  XNOR2_X1 U6282 ( .A(n5542), .B(n5541), .ZN(n7496) );
  INV_X1 U6283 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6301) );
  INV_X1 U6284 ( .A(n9210), .ZN(n9099) );
  AND2_X1 U6285 ( .A1(n6253), .A2(n6252), .ZN(n9580) );
  AND4_X1 U6286 ( .A1(n6212), .A2(n6211), .A3(n6210), .A4(n6209), .ZN(n8981)
         );
  OR3_X1 U6287 ( .A1(n6059), .A2(n6058), .A3(n6057), .ZN(n9103) );
  OR2_X1 U6288 ( .A1(P1_U3083), .A2(n9710), .ZN(n9802) );
  OR2_X1 U6289 ( .A1(n9149), .A2(n7092), .ZN(n9156) );
  AND2_X1 U6290 ( .A1(n6704), .A2(n9633), .ZN(n9149) );
  OR2_X1 U6291 ( .A1(n6866), .A2(n6865), .ZN(n9886) );
  AND2_X1 U6292 ( .A1(n9670), .A2(n9669), .ZN(n9682) );
  OR2_X1 U6293 ( .A1(n6866), .A2(n6375), .ZN(n9877) );
  CLKBUF_X1 U6294 ( .A(n9816), .Z(n9834) );
  AND2_X1 U6295 ( .A1(n6354), .A2(n6240), .ZN(n6447) );
  INV_X1 U6296 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6325) );
  NOR2_X1 U6297 ( .A1(n10105), .A2(n10104), .ZN(n10103) );
  NOR2_X2 U6298 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5069) );
  NAND2_X1 U6299 ( .A1(n5069), .A2(n4918), .ZN(n5104) );
  NOR2_X1 U6300 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4921) );
  NAND4_X1 U6301 ( .A1(n4921), .A2(n4920), .A3(n5210), .A4(n5279), .ZN(n4924)
         );
  INV_X1 U6302 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4922) );
  NAND4_X1 U6303 ( .A1(n4922), .A2(n5315), .A3(n5225), .A4(n5158), .ZN(n4923)
         );
  NOR2_X1 U6304 ( .A1(n4924), .A2(n4923), .ZN(n4925) );
  INV_X1 U6305 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4926) );
  NAND4_X1 U6306 ( .A1(n4927), .A2(n4954), .A3(n4926), .A4(n4953), .ZN(n4930)
         );
  INV_X1 U6307 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4928) );
  NAND4_X1 U6308 ( .A1(n4957), .A2(n4928), .A3(n5538), .A4(n5541), .ZN(n4929)
         );
  INV_X1 U6309 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4933) );
  INV_X1 U6310 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4934) );
  INV_X1 U6311 ( .A(n8154), .ZN(n4941) );
  INV_X1 U6312 ( .A(n4936), .ZN(n8688) );
  NAND2_X1 U6313 ( .A1(n4937), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4938) );
  MUX2_X1 U6314 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4938), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n4939) );
  NAND2_X1 U6315 ( .A1(n4315), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n4952) );
  NAND2_X1 U6316 ( .A1(n7580), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4951) );
  AND2_X1 U6317 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5118) );
  NAND2_X1 U6318 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .ZN(n4942) );
  NAND2_X1 U6319 ( .A1(n5193), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5232) );
  NAND2_X1 U6320 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n4943) );
  INV_X1 U6321 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9374) );
  AND2_X1 U6322 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_REG3_REG_13__SCAN_IN), 
        .ZN(n4944) );
  NAND2_X1 U6323 ( .A1(n5284), .A2(n4944), .ZN(n5307) );
  INV_X1 U6324 ( .A(n5307), .ZN(n4945) );
  NAND2_X1 U6325 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n4946) );
  INV_X1 U6326 ( .A(n5334), .ZN(n4947) );
  NAND2_X1 U6327 ( .A1(n4947), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5358) );
  INV_X1 U6328 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9473) );
  NAND2_X1 U6329 ( .A1(n5334), .A2(n9473), .ZN(n4948) );
  AND2_X1 U6330 ( .A1(n5358), .A2(n4948), .ZN(n8508) );
  NAND2_X1 U6331 ( .A1(n5084), .A2(n8508), .ZN(n4950) );
  NAND2_X1 U6332 ( .A1(n5416), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n4949) );
  NAND2_X1 U6333 ( .A1(n5044), .A2(n4928), .ZN(n4959) );
  NAND2_X1 U6334 ( .A1(n4958), .A2(n4957), .ZN(n4956) );
  XNOR2_X2 U6335 ( .A(n4955), .B(n4954), .ZN(n7802) );
  OAI21_X1 U6336 ( .B1(n4958), .B2(n4957), .A(n4956), .ZN(n5575) );
  AND2_X2 U6337 ( .A1(n7802), .A2(n5575), .ZN(n7812) );
  INV_X1 U6338 ( .A(n7812), .ZN(n4963) );
  INV_X1 U6339 ( .A(n4959), .ZN(n4961) );
  NOR2_X1 U6340 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4960) );
  NAND2_X1 U6341 ( .A1(n4961), .A2(n4960), .ZN(n4962) );
  INV_X4 U6342 ( .A(n5058), .ZN(n5534) );
  NOR2_X1 U6343 ( .A1(n8519), .A2(n5534), .ZN(n5344) );
  NAND2_X1 U6344 ( .A1(n5673), .A2(n4966), .ZN(n5057) );
  INV_X1 U6345 ( .A(SI_1_), .ZN(n9437) );
  MUX2_X1 U6346 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4710), .Z(n5065) );
  NAND2_X1 U6347 ( .A1(n5066), .A2(n5065), .ZN(n4968) );
  NAND2_X1 U6348 ( .A1(n4968), .A2(n4967), .ZN(n5072) );
  NAND2_X1 U6349 ( .A1(n5072), .A2(n5071), .ZN(n4970) );
  NAND2_X1 U6350 ( .A1(n4970), .A2(n4969), .ZN(n5092) );
  MUX2_X1 U6351 ( .A(n6291), .B(n6294), .S(n6292), .Z(n4971) );
  NAND2_X1 U6352 ( .A1(n5092), .A2(n5091), .ZN(n4974) );
  INV_X1 U6353 ( .A(n4971), .ZN(n4972) );
  NAND2_X1 U6354 ( .A1(n4974), .A2(n4973), .ZN(n5109) );
  MUX2_X1 U6355 ( .A(n6301), .B(n6297), .S(n6292), .Z(n4975) );
  NAND2_X1 U6356 ( .A1(n5109), .A2(n5108), .ZN(n4978) );
  INV_X1 U6357 ( .A(n4975), .ZN(n4976) );
  NAND2_X1 U6358 ( .A1(n4976), .A2(SI_4_), .ZN(n4977) );
  MUX2_X1 U6359 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6292), .Z(n4980) );
  NAND2_X1 U6360 ( .A1(n4980), .A2(SI_5_), .ZN(n4981) );
  MUX2_X1 U6361 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6292), .Z(n4982) );
  NAND2_X1 U6362 ( .A1(n4982), .A2(SI_6_), .ZN(n4983) );
  MUX2_X1 U6363 ( .A(n4984), .B(n6314), .S(n6292), .Z(n4985) );
  INV_X1 U6364 ( .A(n4985), .ZN(n4986) );
  INV_X1 U6365 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n4987) );
  MUX2_X1 U6366 ( .A(n4987), .B(n6325), .S(n6292), .Z(n4988) );
  INV_X1 U6367 ( .A(n4988), .ZN(n4989) );
  NAND2_X1 U6368 ( .A1(n4989), .A2(SI_8_), .ZN(n4990) );
  INV_X1 U6369 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n4993) );
  INV_X1 U6370 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n4992) );
  MUX2_X1 U6371 ( .A(n4993), .B(n4992), .S(n6292), .Z(n4994) );
  NAND2_X1 U6372 ( .A1(n4994), .A2(n9440), .ZN(n4997) );
  INV_X1 U6373 ( .A(n4994), .ZN(n4995) );
  NAND2_X1 U6374 ( .A1(n4995), .A2(SI_9_), .ZN(n4996) );
  INV_X1 U6375 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5000) );
  INV_X1 U6376 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n4999) );
  MUX2_X1 U6377 ( .A(n5000), .B(n4999), .S(n6292), .Z(n5001) );
  INV_X1 U6378 ( .A(SI_10_), .ZN(n9354) );
  INV_X1 U6379 ( .A(n5001), .ZN(n5002) );
  NAND2_X1 U6380 ( .A1(n5002), .A2(SI_10_), .ZN(n5003) );
  MUX2_X1 U6381 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6292), .Z(n5006) );
  INV_X1 U6382 ( .A(SI_11_), .ZN(n5005) );
  NAND2_X1 U6383 ( .A1(n5006), .A2(SI_11_), .ZN(n5007) );
  INV_X1 U6384 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5008) );
  INV_X1 U6385 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6424) );
  MUX2_X1 U6386 ( .A(n5008), .B(n6424), .S(n7589), .Z(n5010) );
  INV_X1 U6387 ( .A(SI_12_), .ZN(n5009) );
  INV_X1 U6388 ( .A(n5010), .ZN(n5011) );
  NAND2_X1 U6389 ( .A1(n5011), .A2(SI_12_), .ZN(n5012) );
  NAND2_X1 U6390 ( .A1(n5013), .A2(n5012), .ZN(n5243) );
  INV_X1 U6391 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6575) );
  INV_X1 U6392 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5014) );
  MUX2_X1 U6393 ( .A(n6575), .B(n5014), .S(n7589), .Z(n5015) );
  INV_X1 U6394 ( .A(SI_13_), .ZN(n9361) );
  NAND2_X1 U6395 ( .A1(n5015), .A2(n9361), .ZN(n5018) );
  INV_X1 U6396 ( .A(n5015), .ZN(n5016) );
  NAND2_X1 U6397 ( .A1(n5016), .A2(SI_13_), .ZN(n5017) );
  MUX2_X1 U6398 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7589), .Z(n5021) );
  INV_X1 U6399 ( .A(SI_14_), .ZN(n5020) );
  XNOR2_X1 U6400 ( .A(n5021), .B(n5020), .ZN(n5277) );
  INV_X1 U6401 ( .A(n5277), .ZN(n5022) );
  INV_X1 U6402 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6724) );
  INV_X1 U6403 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6722) );
  MUX2_X1 U6404 ( .A(n6724), .B(n6722), .S(n7589), .Z(n5023) );
  INV_X1 U6405 ( .A(SI_15_), .ZN(n9428) );
  NAND2_X1 U6406 ( .A1(n5023), .A2(n9428), .ZN(n5026) );
  INV_X1 U6407 ( .A(n5023), .ZN(n5024) );
  NAND2_X1 U6408 ( .A1(n5024), .A2(SI_15_), .ZN(n5025) );
  NAND2_X1 U6409 ( .A1(n5026), .A2(n5025), .ZN(n5313) );
  INV_X1 U6410 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5028) );
  INV_X1 U6411 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5027) );
  MUX2_X1 U6412 ( .A(n5028), .B(n5027), .S(n7589), .Z(n5029) );
  INV_X1 U6413 ( .A(SI_16_), .ZN(n9395) );
  NAND2_X1 U6414 ( .A1(n5029), .A2(n9395), .ZN(n5032) );
  INV_X1 U6415 ( .A(n5029), .ZN(n5030) );
  NAND2_X1 U6416 ( .A1(n5030), .A2(SI_16_), .ZN(n5031) );
  MUX2_X1 U6417 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n7589), .Z(n5035) );
  INV_X1 U6418 ( .A(SI_17_), .ZN(n5034) );
  XNOR2_X1 U6419 ( .A(n5035), .B(n5034), .ZN(n5327) );
  INV_X1 U6420 ( .A(n5327), .ZN(n5037) );
  NAND2_X1 U6421 ( .A1(n5035), .A2(SI_17_), .ZN(n5036) );
  MUX2_X1 U6422 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7589), .Z(n5348) );
  XNOR2_X1 U6423 ( .A(n5348), .B(SI_18_), .ZN(n5345) );
  XNOR2_X1 U6424 ( .A(n5347), .B(n5345), .ZN(n6956) );
  INV_X1 U6425 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5041) );
  INV_X2 U6426 ( .A(n5093), .ZN(n5484) );
  NAND2_X1 U6427 ( .A1(n6956), .A2(n5484), .ZN(n5048) );
  INV_X1 U6428 ( .A(n5044), .ZN(n5045) );
  NAND2_X1 U6429 ( .A1(n5045), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5046) );
  XNOR2_X1 U6430 ( .A(n5046), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8315) );
  AOI22_X1 U6431 ( .A1(n5353), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6338), .B2(
        n8315), .ZN(n5047) );
  NAND3_X1 U6432 ( .A1(n7806), .A2(n9982), .A3(n7284), .ZN(n5049) );
  NAND2_X1 U6433 ( .A1(n7802), .A2(n7643), .ZN(n6761) );
  NAND2_X2 U6434 ( .A1(n5049), .A2(n6761), .ZN(n5356) );
  XNOR2_X1 U6435 ( .A(n8511), .B(n4414), .ZN(n5343) );
  NAND2_X1 U6436 ( .A1(n4325), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U6437 ( .A1(n5416), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5052) );
  NAND2_X1 U6438 ( .A1(n5084), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5051) );
  NAND2_X1 U6439 ( .A1(n4337), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5050) );
  INV_X1 U6440 ( .A(n4913), .ZN(n8265) );
  INV_X1 U6441 ( .A(SI_0_), .ZN(n5055) );
  INV_X1 U6442 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5054) );
  OAI21_X1 U6443 ( .B1(n7589), .B2(n5055), .A(n5054), .ZN(n5056) );
  AND2_X1 U6444 ( .A1(n5057), .A2(n5056), .ZN(n8705) );
  NAND2_X1 U6445 ( .A1(n8265), .A2(n8139), .ZN(n6845) );
  INV_X1 U6446 ( .A(n6845), .ZN(n5059) );
  NAND2_X1 U6447 ( .A1(n5059), .A2(n5058), .ZN(n8135) );
  OR2_X1 U6448 ( .A1(n8139), .A2(n5356), .ZN(n5060) );
  AND2_X1 U6449 ( .A1(n8135), .A2(n5060), .ZN(n8189) );
  NAND2_X1 U6450 ( .A1(n4325), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5064) );
  NAND2_X1 U6451 ( .A1(n5084), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5063) );
  NAND2_X1 U6452 ( .A1(n5416), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5062) );
  NAND2_X1 U6453 ( .A1(n4337), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5061) );
  AND4_X2 U6454 ( .A1(n5064), .A2(n5063), .A3(n5062), .A4(n5061), .ZN(n8142)
         );
  INV_X1 U6455 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6298) );
  XNOR2_X1 U6456 ( .A(n5066), .B(n5065), .ZN(n6299) );
  INV_X1 U6457 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5068) );
  NAND2_X1 U6458 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5067) );
  XNOR2_X1 U6459 ( .A(n5068), .B(n5067), .ZN(n6477) );
  XNOR2_X1 U6460 ( .A(n8187), .B(n5356), .ZN(n5080) );
  OR2_X1 U6461 ( .A1(n5069), .A2(n4933), .ZN(n5070) );
  XNOR2_X1 U6462 ( .A(n5070), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6480) );
  INV_X1 U6463 ( .A(n6480), .ZN(n9516) );
  XNOR2_X1 U6464 ( .A(n5072), .B(n5071), .ZN(n6302) );
  OR2_X1 U6465 ( .A1(n5093), .A2(n6302), .ZN(n5073) );
  INV_X1 U6466 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5075) );
  NOR2_X1 U6467 ( .A1(n6633), .A2(n5534), .ZN(n5078) );
  INV_X1 U6468 ( .A(n5078), .ZN(n5076) );
  NAND2_X1 U6469 ( .A1(n8178), .A2(n5076), .ZN(n5079) );
  XNOR2_X1 U6470 ( .A(n8231), .B(n5356), .ZN(n5077) );
  NAND2_X1 U6471 ( .A1(n5078), .A2(n5077), .ZN(n5083) );
  INV_X1 U6472 ( .A(n5080), .ZN(n5081) );
  NAND2_X1 U6473 ( .A1(n5082), .A2(n5081), .ZN(n8232) );
  NAND2_X1 U6474 ( .A1(n4325), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5088) );
  INV_X1 U6475 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9368) );
  NAND2_X1 U6476 ( .A1(n5084), .A2(n9368), .ZN(n5087) );
  NAND2_X1 U6477 ( .A1(n5416), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U6478 ( .A1(n4337), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5085) );
  NOR2_X1 U6479 ( .A1(n6796), .A2(n5534), .ZN(n5095) );
  NAND2_X1 U6480 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5089), .ZN(n5090) );
  XNOR2_X1 U6481 ( .A(n5090), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6544) );
  INV_X1 U6482 ( .A(n6544), .ZN(n6290) );
  XNOR2_X1 U6483 ( .A(n5092), .B(n5091), .ZN(n6293) );
  OR2_X1 U6484 ( .A1(n7594), .A2(n6291), .ZN(n5094) );
  NAND2_X1 U6485 ( .A1(n5095), .A2(n5096), .ZN(n5112) );
  INV_X1 U6486 ( .A(n5096), .ZN(n6790) );
  NAND2_X1 U6487 ( .A1(n4337), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U6488 ( .A1(n7580), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5102) );
  NOR2_X1 U6489 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5099) );
  NOR2_X1 U6490 ( .A1(n5118), .A2(n5099), .ZN(n6772) );
  NAND2_X1 U6491 ( .A1(n5084), .A2(n6772), .ZN(n5101) );
  NAND2_X1 U6492 ( .A1(n5416), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5100) );
  OR2_X1 U6493 ( .A1(n9917), .A2(n5534), .ZN(n5116) );
  NAND2_X1 U6494 ( .A1(n5104), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5105) );
  MUX2_X1 U6495 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5105), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5107) );
  NAND2_X1 U6496 ( .A1(n5107), .A2(n5106), .ZN(n6475) );
  OR2_X1 U6497 ( .A1(n7594), .A2(n6301), .ZN(n5111) );
  XNOR2_X1 U6498 ( .A(n5109), .B(n5108), .ZN(n6300) );
  OR2_X1 U6499 ( .A1(n5093), .A2(n6300), .ZN(n5110) );
  OAI211_X1 U6500 ( .C1(n6466), .C2(n6475), .A(n5111), .B(n5110), .ZN(n6769)
         );
  XNOR2_X1 U6501 ( .A(n4414), .B(n6769), .ZN(n5115) );
  XNOR2_X1 U6502 ( .A(n5116), .B(n5115), .ZN(n6793) );
  INV_X1 U6503 ( .A(n5112), .ZN(n5113) );
  NOR2_X1 U6504 ( .A1(n6793), .A2(n5113), .ZN(n5114) );
  NAND2_X1 U6505 ( .A1(n5116), .A2(n5115), .ZN(n5117) );
  NAND2_X1 U6506 ( .A1(n6794), .A2(n5117), .ZN(n9910) );
  INV_X1 U6507 ( .A(n9910), .ZN(n5138) );
  NAND2_X1 U6508 ( .A1(n7580), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5126) );
  INV_X1 U6509 ( .A(n5145), .ZN(n5122) );
  INV_X1 U6510 ( .A(n5118), .ZN(n5120) );
  INV_X1 U6511 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5119) );
  NAND2_X1 U6512 ( .A1(n5120), .A2(n5119), .ZN(n5121) );
  NAND2_X1 U6513 ( .A1(n5122), .A2(n5121), .ZN(n9922) );
  INV_X1 U6514 ( .A(n9922), .ZN(n9959) );
  NAND2_X1 U6515 ( .A1(n5084), .A2(n9959), .ZN(n5125) );
  NAND2_X1 U6516 ( .A1(n5416), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5124) );
  NAND2_X1 U6517 ( .A1(n4337), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5123) );
  AND2_X1 U6518 ( .A1(n8261), .A2(n7604), .ZN(n5133) );
  NAND2_X1 U6519 ( .A1(n5106), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5127) );
  XNOR2_X1 U6520 ( .A(n5127), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6530) );
  INV_X1 U6521 ( .A(n6530), .ZN(n6303) );
  XNOR2_X1 U6522 ( .A(n5129), .B(n5128), .ZN(n6306) );
  OR2_X1 U6523 ( .A1(n5093), .A2(n6306), .ZN(n5131) );
  INV_X1 U6524 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6304) );
  OR2_X1 U6525 ( .A1(n7594), .A2(n6304), .ZN(n5130) );
  XNOR2_X1 U6526 ( .A(n9957), .B(n5132), .ZN(n5134) );
  NAND2_X1 U6527 ( .A1(n5133), .A2(n5134), .ZN(n5150) );
  INV_X1 U6528 ( .A(n5133), .ZN(n5135) );
  INV_X1 U6529 ( .A(n5134), .ZN(n6805) );
  NAND2_X1 U6530 ( .A1(n5135), .A2(n6805), .ZN(n5136) );
  NAND2_X1 U6531 ( .A1(n5150), .A2(n5136), .ZN(n9911) );
  INV_X1 U6532 ( .A(n9911), .ZN(n5137) );
  NAND2_X1 U6533 ( .A1(n5138), .A2(n5137), .ZN(n6804) );
  OR2_X1 U6534 ( .A1(n5139), .A2(n4933), .ZN(n5140) );
  XNOR2_X1 U6535 ( .A(n5140), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6505) );
  AOI22_X1 U6536 ( .A1(n5353), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6338), .B2(
        n6505), .ZN(n5144) );
  XNOR2_X1 U6537 ( .A(n5142), .B(n5141), .ZN(n6309) );
  OR2_X1 U6538 ( .A1(n6309), .A2(n5093), .ZN(n5143) );
  NAND2_X1 U6539 ( .A1(n5144), .A2(n5143), .ZN(n7175) );
  XNOR2_X1 U6540 ( .A(n7175), .B(n5132), .ZN(n5152) );
  NAND2_X1 U6541 ( .A1(n4315), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U6542 ( .A1(n7580), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5148) );
  OAI21_X1 U6543 ( .B1(n5145), .B2(P2_REG3_REG_6__SCAN_IN), .A(n5179), .ZN(
        n6811) );
  INV_X1 U6544 ( .A(n6811), .ZN(n7131) );
  NAND2_X1 U6545 ( .A1(n5084), .A2(n7131), .ZN(n5147) );
  NAND2_X1 U6546 ( .A1(n6326), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5146) );
  NAND4_X1 U6547 ( .A1(n5149), .A2(n5148), .A3(n5147), .A4(n5146), .ZN(n8260)
         );
  NAND2_X1 U6548 ( .A1(n8260), .A2(n7604), .ZN(n5153) );
  XNOR2_X1 U6549 ( .A(n5152), .B(n5153), .ZN(n6817) );
  AND2_X1 U6550 ( .A1(n6817), .A2(n5150), .ZN(n5151) );
  INV_X1 U6551 ( .A(n5152), .ZN(n5154) );
  NAND2_X1 U6552 ( .A1(n5154), .A2(n5153), .ZN(n5155) );
  XNOR2_X1 U6553 ( .A(n5157), .B(n5156), .ZN(n6315) );
  OR2_X1 U6554 ( .A1(n6315), .A2(n5093), .ZN(n5161) );
  NAND2_X1 U6555 ( .A1(n5139), .A2(n5158), .ZN(n5172) );
  NAND2_X1 U6556 ( .A1(n5172), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5159) );
  XNOR2_X1 U6557 ( .A(n5159), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6517) );
  AOI22_X1 U6558 ( .A1(n5353), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6338), .B2(
        n6517), .ZN(n5160) );
  XNOR2_X1 U6559 ( .A(n10011), .B(n4414), .ZN(n6973) );
  NAND2_X1 U6560 ( .A1(n4315), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U6561 ( .A1(n7580), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5164) );
  XNOR2_X1 U6562 ( .A(n5179), .B(P2_REG3_REG_7__SCAN_IN), .ZN(n7170) );
  NAND2_X1 U6563 ( .A1(n5084), .A2(n7170), .ZN(n5163) );
  NAND2_X1 U6564 ( .A1(n6326), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5162) );
  NAND4_X1 U6565 ( .A1(n5165), .A2(n5164), .A3(n5163), .A4(n5162), .ZN(n8259)
         );
  AND2_X1 U6566 ( .A1(n8259), .A2(n7604), .ZN(n5166) );
  NAND2_X1 U6567 ( .A1(n6973), .A2(n5166), .ZN(n6975) );
  INV_X1 U6568 ( .A(n6973), .ZN(n5168) );
  INV_X1 U6569 ( .A(n5166), .ZN(n5167) );
  NAND2_X1 U6570 ( .A1(n5168), .A2(n5167), .ZN(n5169) );
  NAND2_X1 U6571 ( .A1(n6975), .A2(n5169), .ZN(n6934) );
  XNOR2_X1 U6572 ( .A(n5171), .B(n5170), .ZN(n6322) );
  NAND2_X1 U6573 ( .A1(n6322), .A2(n5484), .ZN(n5178) );
  INV_X1 U6574 ( .A(n5211), .ZN(n5176) );
  NAND2_X1 U6575 ( .A1(n5173), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5174) );
  MUX2_X1 U6576 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5174), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5175) );
  AOI22_X1 U6577 ( .A1(n5353), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6338), .B2(
        n6572), .ZN(n5177) );
  XNOR2_X1 U6578 ( .A(n10017), .B(n4414), .ZN(n5201) );
  INV_X1 U6579 ( .A(n5201), .ZN(n5186) );
  NAND2_X1 U6580 ( .A1(n4315), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6581 ( .A1(n7580), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5184) );
  INV_X1 U6582 ( .A(n5179), .ZN(n5180) );
  AOI21_X1 U6583 ( .B1(n5180), .B2(P2_REG3_REG_7__SCAN_IN), .A(
        P2_REG3_REG_8__SCAN_IN), .ZN(n5181) );
  OR2_X1 U6584 ( .A1(n5181), .A2(n5193), .ZN(n6972) );
  INV_X1 U6585 ( .A(n6972), .ZN(n8573) );
  NAND2_X1 U6586 ( .A1(n5084), .A2(n8573), .ZN(n5183) );
  NAND2_X1 U6587 ( .A1(n6326), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5182) );
  NOR2_X1 U6588 ( .A1(n7218), .A2(n5534), .ZN(n5200) );
  NAND2_X1 U6589 ( .A1(n5186), .A2(n5200), .ZN(n5199) );
  AND2_X1 U6590 ( .A1(n6975), .A2(n5199), .ZN(n5187) );
  NAND2_X1 U6591 ( .A1(n6976), .A2(n5187), .ZN(n7069) );
  XNOR2_X1 U6592 ( .A(n5189), .B(n5188), .ZN(n6333) );
  NAND2_X1 U6593 ( .A1(n6333), .A2(n5484), .ZN(n5192) );
  OR2_X1 U6594 ( .A1(n5211), .A2(n4933), .ZN(n5190) );
  XNOR2_X1 U6595 ( .A(n5190), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6608) );
  AOI22_X1 U6596 ( .A1(n5353), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6338), .B2(
        n6608), .ZN(n5191) );
  XNOR2_X1 U6597 ( .A(n10027), .B(n4414), .ZN(n5205) );
  NAND2_X1 U6598 ( .A1(n4315), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6599 ( .A1(n7580), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5197) );
  OR2_X1 U6600 ( .A1(n5193), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5194) );
  AND2_X1 U6601 ( .A1(n5232), .A2(n5194), .ZN(n7234) );
  NAND2_X1 U6602 ( .A1(n5084), .A2(n7234), .ZN(n5196) );
  NAND2_X1 U6603 ( .A1(n6326), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5195) );
  OR2_X1 U6604 ( .A1(n7305), .A2(n5534), .ZN(n5206) );
  NAND2_X1 U6605 ( .A1(n5205), .A2(n5206), .ZN(n5203) );
  INV_X1 U6606 ( .A(n5199), .ZN(n5202) );
  XNOR2_X1 U6607 ( .A(n5201), .B(n5200), .ZN(n6977) );
  OR2_X1 U6608 ( .A1(n5202), .A2(n6977), .ZN(n7068) );
  AND2_X1 U6609 ( .A1(n5203), .A2(n7068), .ZN(n5204) );
  INV_X1 U6610 ( .A(n5205), .ZN(n7072) );
  INV_X1 U6611 ( .A(n5206), .ZN(n5207) );
  NAND2_X1 U6612 ( .A1(n7072), .A2(n5207), .ZN(n7066) );
  XNOR2_X1 U6613 ( .A(n5209), .B(n5208), .ZN(n6345) );
  NAND2_X1 U6614 ( .A1(n6345), .A2(n5484), .ZN(n5213) );
  NAND2_X1 U6615 ( .A1(n5211), .A2(n5210), .ZN(n5245) );
  NAND2_X1 U6616 ( .A1(n5245), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5226) );
  XNOR2_X1 U6617 ( .A(n5226), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6675) );
  AOI22_X1 U6618 ( .A1(n5353), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6338), .B2(
        n6675), .ZN(n5212) );
  NAND2_X1 U6619 ( .A1(n5213), .A2(n5212), .ZN(n9946) );
  XNOR2_X1 U6620 ( .A(n9946), .B(n5249), .ZN(n5218) );
  NAND2_X1 U6621 ( .A1(n4315), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U6622 ( .A1(n7580), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5216) );
  XNOR2_X1 U6623 ( .A(n5232), .B(P2_REG3_REG_10__SCAN_IN), .ZN(n9943) );
  NAND2_X1 U6624 ( .A1(n5084), .A2(n9943), .ZN(n5215) );
  NAND2_X1 U6625 ( .A1(n6326), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5214) );
  NOR2_X1 U6626 ( .A1(n7304), .A2(n5534), .ZN(n5219) );
  NAND2_X1 U6627 ( .A1(n5218), .A2(n5219), .ZN(n5222) );
  INV_X1 U6628 ( .A(n5218), .ZN(n7057) );
  INV_X1 U6629 ( .A(n5219), .ZN(n5220) );
  NAND2_X1 U6630 ( .A1(n7057), .A2(n5220), .ZN(n5221) );
  AND2_X1 U6631 ( .A1(n5222), .A2(n5221), .ZN(n6987) );
  XNOR2_X1 U6632 ( .A(n5224), .B(n5223), .ZN(n6349) );
  NAND2_X1 U6633 ( .A1(n6349), .A2(n5484), .ZN(n5230) );
  NAND2_X1 U6634 ( .A1(n5226), .A2(n5225), .ZN(n5227) );
  NAND2_X1 U6635 ( .A1(n5227), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5228) );
  XNOR2_X1 U6636 ( .A(n5228), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6859) );
  AOI22_X1 U6637 ( .A1(n5353), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6338), .B2(
        n6859), .ZN(n5229) );
  NAND2_X1 U6638 ( .A1(n5230), .A2(n5229), .ZN(n7347) );
  XNOR2_X1 U6639 ( .A(n7347), .B(n5249), .ZN(n9898) );
  NAND2_X1 U6640 ( .A1(n4315), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6641 ( .A1(n7580), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5236) );
  INV_X1 U6642 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6603) );
  INV_X1 U6643 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5231) );
  OAI21_X1 U6644 ( .B1(n5232), .B2(n6603), .A(n5231), .ZN(n5233) );
  AND2_X1 U6645 ( .A1(n5233), .A2(n5250), .ZN(n7313) );
  NAND2_X1 U6646 ( .A1(n5084), .A2(n7313), .ZN(n5235) );
  NAND2_X1 U6647 ( .A1(n6326), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5234) );
  NOR2_X1 U6648 ( .A1(n7355), .A2(n5534), .ZN(n5238) );
  NAND2_X1 U6649 ( .A1(n9898), .A2(n5238), .ZN(n5242) );
  INV_X1 U6650 ( .A(n9898), .ZN(n5240) );
  INV_X1 U6651 ( .A(n5238), .ZN(n5239) );
  NAND2_X1 U6652 ( .A1(n5240), .A2(n5239), .ZN(n5241) );
  AND2_X1 U6653 ( .A1(n5242), .A2(n5241), .ZN(n7055) );
  XNOR2_X1 U6654 ( .A(n5244), .B(n5243), .ZN(n6380) );
  NAND2_X1 U6655 ( .A1(n6380), .A2(n5484), .ZN(n5248) );
  NAND2_X1 U6656 ( .A1(n5263), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5246) );
  XNOR2_X1 U6657 ( .A(n5246), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6895) );
  AOI22_X1 U6658 ( .A1(n5353), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6338), .B2(
        n6895), .ZN(n5247) );
  XNOR2_X1 U6659 ( .A(n9901), .B(n5249), .ZN(n5256) );
  NAND2_X1 U6660 ( .A1(n4315), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5255) );
  NAND2_X1 U6661 ( .A1(n7580), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5254) );
  AND2_X1 U6662 ( .A1(n5250), .A2(n9374), .ZN(n5251) );
  OR2_X1 U6663 ( .A1(n5251), .A2(n5284), .ZN(n9907) );
  INV_X1 U6664 ( .A(n9907), .ZN(n7359) );
  NAND2_X1 U6665 ( .A1(n5084), .A2(n7359), .ZN(n5253) );
  NAND2_X1 U6666 ( .A1(n6326), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5252) );
  NOR2_X1 U6667 ( .A1(n7402), .A2(n5534), .ZN(n5257) );
  NAND2_X1 U6668 ( .A1(n5256), .A2(n5257), .ZN(n5260) );
  INV_X1 U6669 ( .A(n5256), .ZN(n7242) );
  INV_X1 U6670 ( .A(n5257), .ZN(n5258) );
  NAND2_X1 U6671 ( .A1(n7242), .A2(n5258), .ZN(n5259) );
  AND2_X1 U6672 ( .A1(n5260), .A2(n5259), .ZN(n9894) );
  NAND2_X1 U6673 ( .A1(n9903), .A2(n5260), .ZN(n5275) );
  XNOR2_X1 U6674 ( .A(n5262), .B(n5261), .ZN(n6441) );
  NAND2_X1 U6675 ( .A1(n6441), .A2(n5484), .ZN(n5265) );
  OAI21_X1 U6676 ( .B1(n5263), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5280) );
  XNOR2_X1 U6677 ( .A(n5280), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7012) );
  AOI22_X1 U6678 ( .A1(n5353), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6338), .B2(
        n7012), .ZN(n5264) );
  XNOR2_X1 U6679 ( .A(n7411), .B(n5249), .ZN(n5270) );
  NAND2_X1 U6680 ( .A1(n4315), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U6681 ( .A1(n7580), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5268) );
  INV_X1 U6682 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6892) );
  XNOR2_X1 U6683 ( .A(n5284), .B(n6892), .ZN(n7410) );
  NAND2_X1 U6684 ( .A1(n5084), .A2(n7410), .ZN(n5267) );
  NAND2_X1 U6685 ( .A1(n5416), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5266) );
  NOR2_X1 U6686 ( .A1(n7459), .A2(n5534), .ZN(n5271) );
  NAND2_X1 U6687 ( .A1(n5270), .A2(n5271), .ZN(n5276) );
  INV_X1 U6688 ( .A(n5270), .ZN(n5273) );
  INV_X1 U6689 ( .A(n5271), .ZN(n5272) );
  NAND2_X1 U6690 ( .A1(n5273), .A2(n5272), .ZN(n5274) );
  AND2_X1 U6691 ( .A1(n5276), .A2(n5274), .ZN(n7240) );
  XNOR2_X1 U6692 ( .A(n5278), .B(n5277), .ZN(n6623) );
  NAND2_X1 U6693 ( .A1(n6623), .A2(n5484), .ZN(n5283) );
  NAND2_X1 U6694 ( .A1(n5280), .A2(n5279), .ZN(n5281) );
  NAND2_X1 U6695 ( .A1(n5281), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5316) );
  XNOR2_X1 U6696 ( .A(n5316), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7291) );
  AOI22_X1 U6697 ( .A1(n7291), .A2(n6338), .B1(n5353), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5282) );
  XNOR2_X1 U6698 ( .A(n9536), .B(n5249), .ZN(n5293) );
  NAND2_X1 U6699 ( .A1(n7580), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5292) );
  INV_X1 U6700 ( .A(n5284), .ZN(n5286) );
  INV_X1 U6701 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5285) );
  OAI21_X1 U6702 ( .B1(n5286), .B2(n6892), .A(n5285), .ZN(n5287) );
  NAND2_X1 U6703 ( .A1(n5307), .A2(n5287), .ZN(n9539) );
  INV_X1 U6704 ( .A(n9539), .ZN(n5288) );
  NAND2_X1 U6705 ( .A1(n5084), .A2(n5288), .ZN(n5291) );
  NAND2_X1 U6706 ( .A1(n6326), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U6707 ( .A1(n4315), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5289) );
  NOR2_X1 U6708 ( .A1(n8092), .A2(n5534), .ZN(n5294) );
  XNOR2_X1 U6709 ( .A(n5293), .B(n5294), .ZN(n9532) );
  INV_X1 U6710 ( .A(n5293), .ZN(n5296) );
  INV_X1 U6711 ( .A(n5294), .ZN(n5295) );
  XNOR2_X1 U6712 ( .A(n5298), .B(n5297), .ZN(n6819) );
  NAND2_X1 U6713 ( .A1(n6819), .A2(n5484), .ZN(n5302) );
  OR2_X1 U6714 ( .A1(n5299), .A2(n4933), .ZN(n5300) );
  XNOR2_X1 U6715 ( .A(n5300), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8286) );
  AOI22_X1 U6716 ( .A1(n5353), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6338), .B2(
        n8286), .ZN(n5301) );
  XNOR2_X1 U6717 ( .A(n8660), .B(n5249), .ZN(n7484) );
  NAND2_X1 U6718 ( .A1(n4315), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6719 ( .A1(n7580), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5305) );
  XNOR2_X1 U6720 ( .A(n5333), .B(P2_REG3_REG_16__SCAN_IN), .ZN(n8543) );
  NAND2_X1 U6721 ( .A1(n5084), .A2(n8543), .ZN(n5304) );
  NAND2_X1 U6722 ( .A1(n6326), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5303) );
  NOR2_X1 U6723 ( .A1(n8520), .A2(n5534), .ZN(n7485) );
  NAND2_X1 U6724 ( .A1(n7580), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5312) );
  INV_X1 U6725 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9497) );
  NAND2_X1 U6726 ( .A1(n5307), .A2(n9497), .ZN(n5308) );
  AND2_X1 U6727 ( .A1(n5333), .A2(n5308), .ZN(n8552) );
  NAND2_X1 U6728 ( .A1(n5084), .A2(n8552), .ZN(n5311) );
  NAND2_X1 U6729 ( .A1(n6326), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5310) );
  NAND2_X1 U6730 ( .A1(n4315), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5309) );
  NAND4_X1 U6731 ( .A1(n5312), .A2(n5311), .A3(n5310), .A4(n5309), .ZN(n8255)
         );
  NAND2_X1 U6732 ( .A1(n8255), .A2(n7604), .ZN(n7482) );
  INV_X1 U6733 ( .A(n7482), .ZN(n5323) );
  XNOR2_X1 U6734 ( .A(n5314), .B(n5313), .ZN(n6721) );
  NAND2_X1 U6735 ( .A1(n5316), .A2(n5315), .ZN(n5317) );
  NAND2_X1 U6736 ( .A1(n5317), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5319) );
  INV_X1 U6737 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5318) );
  XNOR2_X1 U6738 ( .A(n5319), .B(n5318), .ZN(n7427) );
  OAI22_X1 U6739 ( .A1(n7427), .A2(n6466), .B1(n7594), .B2(n6724), .ZN(n5320)
         );
  INV_X1 U6740 ( .A(n5320), .ZN(n5321) );
  XNOR2_X1 U6741 ( .A(n8665), .B(n4414), .ZN(n7481) );
  INV_X1 U6742 ( .A(n7481), .ZN(n7470) );
  AOI22_X1 U6743 ( .A1(n7484), .A2(n7485), .B1(n5323), .B2(n7470), .ZN(n5326)
         );
  NAND2_X1 U6744 ( .A1(n7481), .A2(n7482), .ZN(n5322) );
  AOI21_X1 U6745 ( .B1(n7485), .B2(n5322), .A(n7484), .ZN(n5325) );
  NOR3_X1 U6746 ( .A1(n7470), .A2(n5323), .A3(n7485), .ZN(n5324) );
  XNOR2_X1 U6747 ( .A(n5328), .B(n5327), .ZN(n6884) );
  NAND2_X1 U6748 ( .A1(n6884), .A2(n5484), .ZN(n5332) );
  NAND2_X1 U6749 ( .A1(n5329), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5330) );
  XNOR2_X1 U6750 ( .A(n5330), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8300) );
  AOI22_X1 U6751 ( .A1(n5353), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6338), .B2(
        n8300), .ZN(n5331) );
  XNOR2_X1 U6752 ( .A(n8656), .B(n4414), .ZN(n7512) );
  NAND2_X1 U6753 ( .A1(n4315), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6754 ( .A1(n7580), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5338) );
  INV_X1 U6755 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7422) );
  INV_X1 U6756 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9435) );
  OAI21_X1 U6757 ( .B1(n5333), .B2(n7422), .A(n9435), .ZN(n5335) );
  AND2_X1 U6758 ( .A1(n5335), .A2(n5334), .ZN(n8525) );
  NAND2_X1 U6759 ( .A1(n5084), .A2(n8525), .ZN(n5337) );
  NAND2_X1 U6760 ( .A1(n6326), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5336) );
  OR2_X1 U6761 ( .A1(n8536), .A2(n5534), .ZN(n5340) );
  NOR2_X1 U6762 ( .A1(n7512), .A2(n5340), .ZN(n5341) );
  AOI21_X1 U6763 ( .B1(n7512), .B2(n5340), .A(n5341), .ZN(n7449) );
  INV_X1 U6764 ( .A(n5341), .ZN(n5342) );
  XNOR2_X1 U6765 ( .A(n5343), .B(n5344), .ZN(n7513) );
  INV_X1 U6766 ( .A(n5345), .ZN(n5346) );
  NAND2_X1 U6767 ( .A1(n5348), .A2(SI_18_), .ZN(n5349) );
  INV_X1 U6768 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7140) );
  INV_X1 U6769 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7138) );
  MUX2_X1 U6770 ( .A(n7140), .B(n7138), .S(n7589), .Z(n5350) );
  INV_X1 U6771 ( .A(SI_19_), .ZN(n9434) );
  NAND2_X1 U6772 ( .A1(n5350), .A2(n9434), .ZN(n5369) );
  INV_X1 U6773 ( .A(n5350), .ZN(n5351) );
  NAND2_X1 U6774 ( .A1(n5351), .A2(SI_19_), .ZN(n5352) );
  NAND2_X1 U6775 ( .A1(n5369), .A2(n5352), .ZN(n5367) );
  XNOR2_X1 U6776 ( .A(n5366), .B(n5367), .ZN(n7137) );
  NAND2_X1 U6777 ( .A1(n7137), .A2(n5484), .ZN(n5355) );
  AOI22_X1 U6778 ( .A1(n5353), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6338), .B2(
        n9962), .ZN(n5354) );
  XNOR2_X1 U6779 ( .A(n8645), .B(n5249), .ZN(n5365) );
  NAND2_X1 U6780 ( .A1(n7580), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5363) );
  NAND2_X1 U6781 ( .A1(n4315), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5362) );
  INV_X1 U6782 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5357) );
  NAND2_X1 U6783 ( .A1(n5358), .A2(n5357), .ZN(n5359) );
  AND2_X1 U6784 ( .A1(n5377), .A2(n5359), .ZN(n8495) );
  NAND2_X1 U6785 ( .A1(n5084), .A2(n8495), .ZN(n5361) );
  NAND2_X1 U6786 ( .A1(n5416), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5360) );
  NOR2_X1 U6787 ( .A1(n8505), .A2(n5534), .ZN(n5364) );
  NOR2_X1 U6788 ( .A1(n5365), .A2(n5364), .ZN(n7529) );
  NAND2_X1 U6789 ( .A1(n5365), .A2(n5364), .ZN(n7530) );
  INV_X1 U6790 ( .A(n5367), .ZN(n5368) );
  INV_X1 U6791 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7251) );
  INV_X1 U6792 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7298) );
  MUX2_X1 U6793 ( .A(n7251), .B(n7298), .S(n7589), .Z(n5372) );
  INV_X1 U6794 ( .A(SI_20_), .ZN(n5371) );
  NAND2_X1 U6795 ( .A1(n5372), .A2(n5371), .ZN(n5388) );
  INV_X1 U6796 ( .A(n5372), .ZN(n5373) );
  NAND2_X1 U6797 ( .A1(n5373), .A2(SI_20_), .ZN(n5374) );
  XNOR2_X1 U6798 ( .A(n5387), .B(n5386), .ZN(n7250) );
  NAND2_X1 U6799 ( .A1(n7250), .A2(n5484), .ZN(n5376) );
  OR2_X1 U6800 ( .A1(n7594), .A2(n7251), .ZN(n5375) );
  XNOR2_X1 U6801 ( .A(n8474), .B(n5249), .ZN(n5383) );
  NAND2_X1 U6802 ( .A1(n4315), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5382) );
  INV_X1 U6803 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9405) );
  NAND2_X1 U6804 ( .A1(n5377), .A2(n9405), .ZN(n5378) );
  AND2_X1 U6805 ( .A1(n5394), .A2(n5378), .ZN(n8472) );
  NAND2_X1 U6806 ( .A1(n5084), .A2(n8472), .ZN(n5381) );
  NAND2_X1 U6807 ( .A1(n7580), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U6808 ( .A1(n6326), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5379) );
  NOR2_X1 U6809 ( .A1(n8493), .A2(n5534), .ZN(n5385) );
  XNOR2_X1 U6810 ( .A(n5383), .B(n5385), .ZN(n8220) );
  INV_X1 U6811 ( .A(n5383), .ZN(n5384) );
  NAND2_X1 U6812 ( .A1(n5387), .A2(n5386), .ZN(n5389) );
  MUX2_X1 U6813 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7589), .Z(n5404) );
  INV_X1 U6814 ( .A(SI_21_), .ZN(n5390) );
  XNOR2_X1 U6815 ( .A(n5404), .B(n5390), .ZN(n5403) );
  XNOR2_X1 U6816 ( .A(n5407), .B(n5403), .ZN(n7267) );
  NAND2_X1 U6817 ( .A1(n7267), .A2(n5484), .ZN(n5392) );
  INV_X1 U6818 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7285) );
  OR2_X1 U6819 ( .A1(n7594), .A2(n7285), .ZN(n5391) );
  XNOR2_X1 U6820 ( .A(n8461), .B(n5249), .ZN(n5402) );
  NAND2_X1 U6821 ( .A1(n5393), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5414) );
  INV_X1 U6822 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9408) );
  NAND2_X1 U6823 ( .A1(n5394), .A2(n9408), .ZN(n5395) );
  NAND2_X1 U6824 ( .A1(n5414), .A2(n5395), .ZN(n8458) );
  OR2_X1 U6825 ( .A1(n8458), .A2(n5098), .ZN(n5400) );
  NAND2_X1 U6826 ( .A1(n7580), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6827 ( .A1(n4315), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5396) );
  AND2_X1 U6828 ( .A1(n5397), .A2(n5396), .ZN(n5399) );
  NAND2_X1 U6829 ( .A1(n6326), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5398) );
  INV_X1 U6830 ( .A(n8447), .ZN(n8481) );
  NAND2_X1 U6831 ( .A1(n8481), .A2(n7604), .ZN(n5401) );
  XNOR2_X1 U6832 ( .A(n5402), .B(n5401), .ZN(n8194) );
  INV_X1 U6833 ( .A(n5403), .ZN(n5406) );
  NAND2_X1 U6834 ( .A1(n5404), .A2(SI_21_), .ZN(n5405) );
  INV_X1 U6835 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8115) );
  INV_X1 U6836 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7346) );
  MUX2_X1 U6837 ( .A(n8115), .B(n7346), .S(n7589), .Z(n5408) );
  INV_X1 U6838 ( .A(SI_22_), .ZN(n9468) );
  NAND2_X1 U6839 ( .A1(n5408), .A2(n9468), .ZN(n5423) );
  INV_X1 U6840 ( .A(n5408), .ZN(n5409) );
  NAND2_X1 U6841 ( .A1(n5409), .A2(SI_22_), .ZN(n5410) );
  NAND2_X1 U6842 ( .A1(n5423), .A2(n5410), .ZN(n5424) );
  XNOR2_X1 U6843 ( .A(n5425), .B(n5424), .ZN(n7345) );
  NAND2_X1 U6844 ( .A1(n7345), .A2(n5484), .ZN(n5412) );
  OR2_X1 U6845 ( .A1(n7594), .A2(n8115), .ZN(n5411) );
  XNOR2_X1 U6846 ( .A(n8629), .B(n5249), .ZN(n5421) );
  INV_X1 U6847 ( .A(n5421), .ZN(n5413) );
  INV_X1 U6848 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9392) );
  NAND2_X1 U6849 ( .A1(n5414), .A2(n9392), .ZN(n5415) );
  AND2_X1 U6850 ( .A1(n5434), .A2(n5415), .ZN(n8439) );
  NAND2_X1 U6851 ( .A1(n8439), .A2(n5084), .ZN(n5419) );
  AOI22_X1 U6852 ( .A1(n4315), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n7580), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n5418) );
  NAND2_X1 U6853 ( .A1(n5416), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U6854 ( .A1(n8130), .A2(n5420), .ZN(n8134) );
  NAND2_X2 U6855 ( .A1(n8134), .A2(n4917), .ZN(n5440) );
  INV_X1 U6856 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7386) );
  INV_X1 U6857 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7383) );
  MUX2_X1 U6858 ( .A(n7386), .B(n7383), .S(n7589), .Z(n5426) );
  INV_X1 U6859 ( .A(SI_23_), .ZN(n9423) );
  NAND2_X1 U6860 ( .A1(n5426), .A2(n9423), .ZN(n5443) );
  INV_X1 U6861 ( .A(n5426), .ZN(n5427) );
  NAND2_X1 U6862 ( .A1(n5427), .A2(SI_23_), .ZN(n5428) );
  AND2_X1 U6863 ( .A1(n5443), .A2(n5428), .ZN(n5441) );
  NAND2_X1 U6864 ( .A1(n7384), .A2(n5484), .ZN(n5430) );
  OR2_X1 U6865 ( .A1(n7594), .A2(n7386), .ZN(n5429) );
  XNOR2_X1 U6866 ( .A(n8622), .B(n5249), .ZN(n5439) );
  NAND2_X1 U6867 ( .A1(n5432), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5449) );
  INV_X1 U6868 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U6869 ( .A1(n5434), .A2(n5433), .ZN(n5435) );
  NAND2_X1 U6870 ( .A1(n5449), .A2(n5435), .ZN(n8171) );
  OR2_X1 U6871 ( .A1(n8171), .A2(n5098), .ZN(n5438) );
  AOI22_X1 U6872 ( .A1(n4315), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n4325), .B2(
        P2_REG1_REG_23__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U6873 ( .A1(n6326), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5436) );
  INV_X1 U6874 ( .A(n8448), .ZN(n8252) );
  NAND2_X1 U6875 ( .A1(n8252), .A2(n7604), .ZN(n8167) );
  MUX2_X1 U6876 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n7589), .Z(n5463) );
  INV_X1 U6877 ( .A(SI_24_), .ZN(n5445) );
  XNOR2_X1 U6878 ( .A(n5463), .B(n5445), .ZN(n5462) );
  XNOR2_X1 U6879 ( .A(n5461), .B(n5462), .ZN(n7494) );
  NAND2_X1 U6880 ( .A1(n7494), .A2(n5484), .ZN(n5447) );
  INV_X1 U6881 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7495) );
  OR2_X1 U6882 ( .A1(n7594), .A2(n7495), .ZN(n5446) );
  XNOR2_X1 U6883 ( .A(n8617), .B(n5249), .ZN(n5457) );
  INV_X1 U6884 ( .A(n5457), .ZN(n5448) );
  INV_X1 U6885 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9346) );
  NAND2_X1 U6886 ( .A1(n5449), .A2(n9346), .ZN(n5450) );
  NAND2_X1 U6887 ( .A1(n5470), .A2(n5450), .ZN(n8408) );
  OR2_X1 U6888 ( .A1(n8408), .A2(n5098), .ZN(n5456) );
  INV_X1 U6889 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U6890 ( .A1(n7580), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U6891 ( .A1(n4315), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5451) );
  OAI211_X1 U6892 ( .C1(n5453), .C2(n7584), .A(n5452), .B(n5451), .ZN(n5454)
         );
  INV_X1 U6893 ( .A(n5454), .ZN(n5455) );
  NOR2_X1 U6894 ( .A1(n8392), .A2(n5534), .ZN(n8212) );
  NAND2_X1 U6895 ( .A1(n5458), .A2(n5457), .ZN(n5459) );
  NAND2_X1 U6896 ( .A1(n5463), .A2(SI_24_), .ZN(n5464) );
  INV_X1 U6897 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7525) );
  INV_X1 U6898 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7526) );
  MUX2_X1 U6899 ( .A(n7525), .B(n7526), .S(n7589), .Z(n5465) );
  INV_X1 U6900 ( .A(SI_25_), .ZN(n9393) );
  NAND2_X1 U6901 ( .A1(n5465), .A2(n9393), .ZN(n5478) );
  INV_X1 U6902 ( .A(n5465), .ZN(n5466) );
  NAND2_X1 U6903 ( .A1(n5466), .A2(SI_25_), .ZN(n5467) );
  NAND2_X1 U6904 ( .A1(n5478), .A2(n5467), .ZN(n5479) );
  NAND2_X1 U6905 ( .A1(n7523), .A2(n5484), .ZN(n5469) );
  OR2_X1 U6906 ( .A1(n7594), .A2(n7525), .ZN(n5468) );
  XNOR2_X1 U6907 ( .A(n8614), .B(n5249), .ZN(n8203) );
  INV_X1 U6908 ( .A(n8203), .ZN(n5477) );
  INV_X1 U6909 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8207) );
  NAND2_X1 U6910 ( .A1(n5470), .A2(n8207), .ZN(n5471) );
  AND2_X1 U6911 ( .A1(n5488), .A2(n5471), .ZN(n8397) );
  INV_X1 U6912 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U6913 ( .A1(n4315), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U6914 ( .A1(n7580), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5472) );
  OAI211_X1 U6915 ( .C1(n5474), .C2(n7584), .A(n5473), .B(n5472), .ZN(n5475)
         );
  AOI21_X1 U6916 ( .B1(n8397), .B2(n5084), .A(n5475), .ZN(n8415) );
  INV_X1 U6917 ( .A(n8415), .ZN(n8251) );
  NAND2_X1 U6918 ( .A1(n8251), .A2(n7604), .ZN(n8202) );
  INV_X1 U6919 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7551) );
  INV_X1 U6920 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7553) );
  MUX2_X1 U6921 ( .A(n7551), .B(n7553), .S(n7589), .Z(n5481) );
  INV_X1 U6922 ( .A(SI_26_), .ZN(n9412) );
  NAND2_X1 U6923 ( .A1(n5481), .A2(n9412), .ZN(n5501) );
  INV_X1 U6924 ( .A(n5481), .ZN(n5482) );
  NAND2_X1 U6925 ( .A1(n5482), .A2(SI_26_), .ZN(n5483) );
  AND2_X1 U6926 ( .A1(n5501), .A2(n5483), .ZN(n5499) );
  OR2_X1 U6927 ( .A1(n7594), .A2(n7551), .ZN(n5485) );
  NAND2_X1 U6928 ( .A1(n5487), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5526) );
  INV_X1 U6929 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9476) );
  NAND2_X1 U6930 ( .A1(n5488), .A2(n9476), .ZN(n5489) );
  AND2_X1 U6931 ( .A1(n5526), .A2(n5489), .ZN(n8382) );
  NAND2_X1 U6932 ( .A1(n8382), .A2(n5084), .ZN(n5495) );
  INV_X1 U6933 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U6934 ( .A1(n4315), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U6935 ( .A1(n7580), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5490) );
  OAI211_X1 U6936 ( .C1(n5492), .C2(n7584), .A(n5491), .B(n5490), .ZN(n5493)
         );
  INV_X1 U6937 ( .A(n5493), .ZN(n5494) );
  OR2_X1 U6938 ( .A1(n8393), .A2(n5534), .ZN(n5496) );
  AOI21_X1 U6939 ( .B1(n8157), .B2(n5496), .A(n5497), .ZN(n8241) );
  INV_X1 U6940 ( .A(n5497), .ZN(n5498) );
  NAND2_X1 U6941 ( .A1(n8158), .A2(n5498), .ZN(n5518) );
  NAND2_X1 U6942 ( .A1(n5500), .A2(n5499), .ZN(n5502) );
  INV_X1 U6943 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8703) );
  INV_X1 U6944 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n6179) );
  MUX2_X1 U6945 ( .A(n8703), .B(n6179), .S(n7589), .Z(n5503) );
  INV_X1 U6946 ( .A(SI_27_), .ZN(n9420) );
  NAND2_X1 U6947 ( .A1(n5503), .A2(n9420), .ZN(n5522) );
  INV_X1 U6948 ( .A(n5503), .ZN(n5504) );
  NAND2_X1 U6949 ( .A1(n5504), .A2(SI_27_), .ZN(n5505) );
  AND2_X1 U6950 ( .A1(n5522), .A2(n5505), .ZN(n5520) );
  OR2_X1 U6951 ( .A1(n7594), .A2(n8703), .ZN(n5506) );
  XNOR2_X1 U6952 ( .A(n8602), .B(n5249), .ZN(n5512) );
  XNOR2_X1 U6953 ( .A(n5526), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8363) );
  INV_X1 U6954 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U6955 ( .A1(n4315), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U6956 ( .A1(n7580), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5508) );
  OAI211_X1 U6957 ( .C1(n5510), .C2(n7584), .A(n5509), .B(n5508), .ZN(n5511)
         );
  AOI21_X1 U6958 ( .B1(n8363), .B2(n5084), .A(n5511), .ZN(n8242) );
  NOR2_X1 U6959 ( .A1(n8242), .A2(n5534), .ZN(n5513) );
  NAND2_X1 U6960 ( .A1(n5512), .A2(n5513), .ZN(n5519) );
  INV_X1 U6961 ( .A(n5512), .ZN(n5515) );
  INV_X1 U6962 ( .A(n5513), .ZN(n5514) );
  NAND2_X1 U6963 ( .A1(n5515), .A2(n5514), .ZN(n5516) );
  NAND2_X1 U6964 ( .A1(n5519), .A2(n5516), .ZN(n8159) );
  NAND2_X1 U6965 ( .A1(n5518), .A2(n5517), .ZN(n8160) );
  MUX2_X1 U6966 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7589), .Z(n7563) );
  INV_X1 U6967 ( .A(SI_28_), .ZN(n9441) );
  XNOR2_X1 U6968 ( .A(n7563), .B(n9441), .ZN(n7561) );
  INV_X1 U6969 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8699) );
  OR2_X1 U6970 ( .A1(n7594), .A2(n8699), .ZN(n5524) );
  INV_X1 U6971 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9469) );
  INV_X1 U6972 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5588) );
  OAI21_X1 U6973 ( .B1(n5526), .B2(n9469), .A(n5588), .ZN(n5527) );
  NAND2_X1 U6974 ( .A1(n8103), .A2(n5084), .ZN(n5533) );
  INV_X1 U6975 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U6976 ( .A1(n4315), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U6977 ( .A1(n7580), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5528) );
  OAI211_X1 U6978 ( .C1(n5530), .C2(n7584), .A(n5529), .B(n5528), .ZN(n5531)
         );
  INV_X1 U6979 ( .A(n5531), .ZN(n5532) );
  OR2_X1 U6980 ( .A1(n8368), .A2(n5534), .ZN(n5535) );
  XNOR2_X1 U6981 ( .A(n5535), .B(n5249), .ZN(n5572) );
  NOR3_X1 U6982 ( .A1(n8105), .A2(n10018), .A3(n5572), .ZN(n5536) );
  AOI21_X1 U6983 ( .B1(n8105), .B2(n5572), .A(n5536), .ZN(n5537) );
  NAND2_X1 U6984 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  NAND2_X1 U6985 ( .A1(n5540), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5564) );
  INV_X1 U6986 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U6987 ( .A1(n5564), .A2(n5563), .ZN(n5566) );
  NAND2_X1 U6988 ( .A1(n5566), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U6989 ( .A1(n5544), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5545) );
  XNOR2_X1 U6990 ( .A(n5545), .B(P2_IR_REG_26__SCAN_IN), .ZN(n5551) );
  INV_X1 U6991 ( .A(n5551), .ZN(n7552) );
  AND2_X1 U6992 ( .A1(n7496), .A2(n7552), .ZN(n9974) );
  NAND2_X1 U6993 ( .A1(n5546), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5547) );
  XNOR2_X1 U6994 ( .A(n5547), .B(P2_IR_REG_25__SCAN_IN), .ZN(n5562) );
  XOR2_X1 U6995 ( .A(n7496), .B(P2_B_REG_SCAN_IN), .Z(n5548) );
  INV_X1 U6996 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9975) );
  AND2_X1 U6997 ( .A1(n9971), .A2(n9975), .ZN(n5550) );
  INV_X1 U6998 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9977) );
  NOR2_X1 U6999 ( .A1(n5562), .A2(n5551), .ZN(n9978) );
  AOI21_X1 U7000 ( .B1(n9971), .B2(n9977), .A(n9978), .ZN(n6629) );
  NOR4_X1 U7001 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5555) );
  NOR4_X1 U7002 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5554) );
  NOR4_X1 U7003 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5553) );
  NOR4_X1 U7004 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5552) );
  NAND4_X1 U7005 ( .A1(n5555), .A2(n5554), .A3(n5553), .A4(n5552), .ZN(n5561)
         );
  NOR2_X1 U7006 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n5559) );
  NOR4_X1 U7007 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5558) );
  NOR4_X1 U7008 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5557) );
  NOR4_X1 U7009 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5556) );
  NAND4_X1 U7010 ( .A1(n5559), .A2(n5558), .A3(n5557), .A4(n5556), .ZN(n5560)
         );
  OAI21_X1 U7011 ( .B1(n5561), .B2(n5560), .A(n9971), .ZN(n6628) );
  AND2_X1 U7012 ( .A1(n6629), .A2(n6628), .ZN(n6757) );
  NAND2_X1 U7013 ( .A1(n6643), .A2(n6757), .ZN(n5583) );
  INV_X1 U7014 ( .A(n7802), .ZN(n7627) );
  NAND2_X1 U7015 ( .A1(n5583), .A2(n7627), .ZN(n5568) );
  INV_X1 U7016 ( .A(n5562), .ZN(n7524) );
  OR2_X1 U7017 ( .A1(n5564), .A2(n5563), .ZN(n5565) );
  NAND2_X1 U7018 ( .A1(n5566), .A2(n5565), .ZN(n6337) );
  AND2_X1 U7019 ( .A1(n9972), .A2(n10018), .ZN(n5567) );
  INV_X1 U7020 ( .A(n9972), .ZN(n5570) );
  NAND2_X1 U7021 ( .A1(n7815), .A2(n7643), .ZN(n6448) );
  NAND2_X1 U7022 ( .A1(n10048), .A2(n6448), .ZN(n5569) );
  OAI21_X1 U7023 ( .B1(n8105), .B2(n9913), .A(n9909), .ZN(n5574) );
  NAND3_X1 U7024 ( .A1(n8597), .A2(n10048), .A3(n5572), .ZN(n5571) );
  OAI21_X1 U7025 ( .B1(n8597), .B2(n5572), .A(n5571), .ZN(n5573) );
  NAND2_X1 U7026 ( .A1(n5583), .A2(n6759), .ZN(n8138) );
  OR2_X1 U7027 ( .A1(n7812), .A2(n6448), .ZN(n6627) );
  AND3_X1 U7028 ( .A1(n6449), .A2(n6337), .A3(n6627), .ZN(n5576) );
  NAND2_X1 U7029 ( .A1(n8138), .A2(n5576), .ZN(n5577) );
  NAND2_X1 U7030 ( .A1(n5577), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9923) );
  INV_X1 U7031 ( .A(n5578), .ZN(n8355) );
  INV_X1 U7032 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U7033 ( .A1(n4315), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U7034 ( .A1(n7580), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5579) );
  OAI211_X1 U7035 ( .C1(n5581), .C2(n7584), .A(n5580), .B(n5579), .ZN(n5582)
         );
  AOI21_X1 U7036 ( .B1(n8355), .B2(n5084), .A(n5582), .ZN(n8109) );
  INV_X1 U7037 ( .A(n5583), .ZN(n5585) );
  AND2_X1 U7038 ( .A1(n9972), .A2(n7812), .ZN(n5584) );
  INV_X1 U7039 ( .A(n5587), .ZN(n5591) );
  NAND2_X1 U7040 ( .A1(n9892), .A2(n8480), .ZN(n9915) );
  OAI22_X1 U7041 ( .A1(n8109), .A2(n9915), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5588), .ZN(n5589) );
  AOI21_X1 U7042 ( .B1(n8103), .B2(n8222), .A(n5589), .ZN(n5590) );
  INV_X1 U7043 ( .A(n5590), .ZN(n5593) );
  INV_X1 U7044 ( .A(n6448), .ZN(n6339) );
  NAND2_X1 U7045 ( .A1(n9892), .A2(n8478), .ZN(n9916) );
  NOR2_X1 U7046 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5600) );
  INV_X1 U7047 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7048 ( .A1(n5941), .A2(n5944), .ZN(n5602) );
  NOR2_X1 U7049 ( .A1(n5602), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5963) );
  AND2_X1 U7050 ( .A1(n5616), .A2(n5963), .ZN(n5603) );
  INV_X1 U7051 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U7052 ( .A1(n5610), .A2(n5609), .ZN(n5605) );
  NAND2_X1 U7053 ( .A1(n5605), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5607) );
  INV_X1 U7054 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7055 ( .A1(n5607), .A2(n5606), .ZN(n5653) );
  OR2_X1 U7056 ( .A1(n5607), .A2(n5606), .ZN(n5608) );
  NAND2_X1 U7057 ( .A1(n5653), .A2(n5608), .ZN(n6243) );
  NOR2_X1 U7058 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5614) );
  INV_X1 U7059 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5612) );
  INV_X1 U7060 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5615) );
  INV_X1 U7061 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U7062 ( .A1(n5628), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5621) );
  INV_X1 U7063 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U7064 ( .A1(n5621), .A2(n5627), .ZN(n5623) );
  NAND2_X1 U7065 ( .A1(n5623), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5619) );
  XNOR2_X1 U7066 ( .A(n5619), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6223) );
  INV_X1 U7067 ( .A(n5639), .ZN(n6238) );
  NAND2_X1 U7068 ( .A1(n6238), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5620) );
  XNOR2_X1 U7069 ( .A(n5620), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6220) );
  INV_X1 U7070 ( .A(n6220), .ZN(n7499) );
  OR2_X1 U7071 ( .A1(n5621), .A2(n5627), .ZN(n5622) );
  NOR2_X1 U7072 ( .A1(n7499), .A2(n7528), .ZN(n5624) );
  INV_X1 U7073 ( .A(n6354), .ZN(n5663) );
  XNOR2_X1 U7074 ( .A(n5625), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n6288) );
  INV_X1 U7075 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U7076 ( .A1(n5627), .A2(n5626), .ZN(n5630) );
  INV_X1 U7077 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5629) );
  NOR2_X1 U7078 ( .A1(n5630), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n5632) );
  AND2_X1 U7079 ( .A1(n5632), .A2(n5631), .ZN(n5636) );
  INV_X1 U7080 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5637) );
  MUX2_X1 U7081 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6288), .S(n6275), .Z(n6930) );
  AND2_X1 U7082 ( .A1(n5663), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n5635) );
  AND2_X1 U7083 ( .A1(n5637), .A2(n5636), .ZN(n5638) );
  NAND2_X1 U7084 ( .A1(n5641), .A2(n5642), .ZN(n9262) );
  XNOR2_X2 U7085 ( .A(n5640), .B(n9260), .ZN(n5645) );
  INV_X1 U7086 ( .A(n5645), .ZN(n5646) );
  INV_X4 U7087 ( .A(n6035), .ZN(n5992) );
  INV_X1 U7088 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5644) );
  OR2_X1 U7089 ( .A1(n5992), .A2(n5644), .ZN(n5652) );
  NAND2_X1 U7090 ( .A1(n6316), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5651) );
  INV_X1 U7091 ( .A(n6085), .ZN(n6107) );
  INV_X1 U7092 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5647) );
  OR2_X1 U7093 ( .A1(n6107), .A2(n5647), .ZN(n5650) );
  INV_X1 U7094 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9692) );
  OR2_X1 U7095 ( .A1(n5743), .A2(n9692), .ZN(n5649) );
  NAND2_X1 U7096 ( .A1(n5653), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5655) );
  XNOR2_X1 U7097 ( .A(n5655), .B(n5654), .ZN(n6241) );
  NAND2_X1 U7098 ( .A1(n5657), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5659) );
  XNOR2_X1 U7099 ( .A(n5659), .B(n5658), .ZN(n8000) );
  AND2_X1 U7100 ( .A1(n5656), .A2(n8000), .ZN(n6926) );
  NAND2_X1 U7101 ( .A1(n6241), .A2(n6926), .ZN(n5660) );
  NAND2_X1 U7102 ( .A1(n8827), .A2(n4319), .ZN(n5661) );
  NAND2_X1 U7103 ( .A1(n8827), .A2(n6199), .ZN(n5665) );
  AOI22_X1 U7104 ( .A1(n6930), .A2(n5696), .B1(n5663), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U7105 ( .A1(n5665), .A2(n5664), .ZN(n6662) );
  NAND2_X1 U7106 ( .A1(n6663), .A2(n6662), .ZN(n6661) );
  NAND2_X1 U7107 ( .A1(n8087), .A2(n8000), .ZN(n6688) );
  AND2_X2 U7108 ( .A1(n6688), .A2(n6687), .ZN(n5733) );
  INV_X1 U7109 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6693) );
  OR2_X1 U7110 ( .A1(n5992), .A2(n6693), .ZN(n5671) );
  NAND2_X1 U7111 ( .A1(n6316), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5670) );
  INV_X1 U7112 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5667) );
  OR2_X1 U7113 ( .A1(n5743), .A2(n5667), .ZN(n5669) );
  OR2_X1 U7114 ( .A1(n6107), .A2(n4603), .ZN(n5668) );
  NAND2_X1 U7115 ( .A1(n8825), .A2(n6199), .ZN(n5676) );
  INV_X1 U7116 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5672) );
  NAND2_X4 U7117 ( .A1(n6275), .A2(n5673), .ZN(n7877) );
  INV_X1 U7118 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U7119 ( .A1(n5676), .A2(n5675), .ZN(n5677) );
  XNOR2_X1 U7120 ( .A(n5677), .B(n5718), .ZN(n5681) );
  AND2_X1 U7121 ( .A1(n7835), .A2(n6093), .ZN(n5679) );
  AOI21_X1 U7122 ( .B1(n8825), .B2(n5678), .A(n5679), .ZN(n6726) );
  NAND2_X1 U7123 ( .A1(n6727), .A2(n6726), .ZN(n6725) );
  INV_X1 U7124 ( .A(n5680), .ZN(n5683) );
  INV_X1 U7125 ( .A(n5681), .ZN(n5682) );
  NAND2_X1 U7126 ( .A1(n5683), .A2(n5682), .ZN(n6729) );
  NAND2_X1 U7127 ( .A1(n6725), .A2(n6729), .ZN(n6715) );
  INV_X1 U7128 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5684) );
  OR2_X1 U7129 ( .A1(n4317), .A2(n6881), .ZN(n5689) );
  INV_X1 U7130 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5685) );
  OR2_X1 U7131 ( .A1(n6107), .A2(n5685), .ZN(n5688) );
  INV_X1 U7132 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n5686) );
  OR2_X1 U7133 ( .A1(n5992), .A2(n5686), .ZN(n5687) );
  NAND4_X2 U7134 ( .A1(n5690), .A2(n5689), .A3(n5688), .A4(n5687), .ZN(n8823)
         );
  NAND2_X1 U7135 ( .A1(n8823), .A2(n6199), .ZN(n5698) );
  OR2_X1 U7136 ( .A1(n5691), .A2(n5965), .ZN(n5693) );
  INV_X1 U7137 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5692) );
  NAND2_X1 U7138 ( .A1(n5693), .A2(n5692), .ZN(n5711) );
  OAI21_X1 U7139 ( .B1(n5693), .B2(n5692), .A(n5711), .ZN(n6393) );
  INV_X1 U7140 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6295) );
  OR2_X1 U7141 ( .A1(n7877), .A2(n6295), .ZN(n5695) );
  OR2_X1 U7142 ( .A1(n5806), .A2(n6302), .ZN(n5694) );
  OAI211_X1 U7143 ( .C1(n6275), .C2(n6393), .A(n5695), .B(n5694), .ZN(n6716)
         );
  NAND2_X1 U7144 ( .A1(n6716), .A2(n5696), .ZN(n5697) );
  NAND2_X1 U7145 ( .A1(n5698), .A2(n5697), .ZN(n5699) );
  XNOR2_X1 U7146 ( .A(n5699), .B(n5718), .ZN(n5701) );
  AND2_X1 U7147 ( .A1(n6716), .A2(n6199), .ZN(n5700) );
  AOI21_X1 U7148 ( .B1(n8823), .B2(n4319), .A(n5700), .ZN(n5702) );
  XNOR2_X1 U7149 ( .A(n5701), .B(n5702), .ZN(n6714) );
  NAND2_X1 U7150 ( .A1(n6715), .A2(n6714), .ZN(n5705) );
  INV_X1 U7151 ( .A(n5701), .ZN(n5703) );
  NAND2_X1 U7152 ( .A1(n5703), .A2(n5702), .ZN(n5704) );
  NAND2_X1 U7153 ( .A1(n5705), .A2(n5704), .ZN(n6615) );
  NAND2_X1 U7154 ( .A1(n6316), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5710) );
  INV_X4 U7155 ( .A(n6085), .ZN(n6369) );
  INV_X1 U7156 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5706) );
  OR2_X1 U7157 ( .A1(n6369), .A2(n5706), .ZN(n5709) );
  INV_X1 U7158 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6382) );
  OR2_X1 U7159 ( .A1(n4316), .A2(n6382), .ZN(n5708) );
  OR2_X1 U7160 ( .A1(n5992), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5707) );
  NAND4_X2 U7161 ( .A1(n5710), .A2(n5709), .A3(n5708), .A4(n5707), .ZN(n8822)
         );
  NAND2_X1 U7162 ( .A1(n8822), .A2(n6199), .ZN(n5717) );
  NAND2_X1 U7163 ( .A1(n5711), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5713) );
  INV_X1 U7164 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5712) );
  XNOR2_X1 U7165 ( .A(n5713), .B(n5712), .ZN(n6400) );
  OR2_X1 U7166 ( .A1(n5806), .A2(n6293), .ZN(n5714) );
  OAI211_X1 U7167 ( .C1(n6275), .C2(n6400), .A(n5715), .B(n5714), .ZN(n7027)
         );
  NAND2_X1 U7168 ( .A1(n7027), .A2(n5696), .ZN(n5716) );
  NAND2_X1 U7169 ( .A1(n5717), .A2(n5716), .ZN(n5719) );
  XNOR2_X1 U7170 ( .A(n5719), .B(n5718), .ZN(n5736) );
  AND2_X1 U7171 ( .A1(n7027), .A2(n6093), .ZN(n5720) );
  AOI21_X1 U7172 ( .B1(n8822), .B2(n4319), .A(n5720), .ZN(n5737) );
  XNOR2_X1 U7173 ( .A(n5736), .B(n5737), .ZN(n6616) );
  NAND2_X1 U7174 ( .A1(n6615), .A2(n6616), .ZN(n6649) );
  NAND2_X1 U7175 ( .A1(n6316), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5724) );
  INV_X1 U7176 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6960) );
  OR2_X1 U7177 ( .A1(n6369), .A2(n6960), .ZN(n5723) );
  XNOR2_X1 U7178 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6959) );
  OR2_X1 U7179 ( .A1(n5992), .A2(n6959), .ZN(n5722) );
  INV_X1 U7180 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6405) );
  OR2_X1 U7181 ( .A1(n4317), .A2(n6405), .ZN(n5721) );
  NAND2_X1 U7182 ( .A1(n8821), .A2(n6199), .ZN(n5732) );
  NAND2_X1 U7183 ( .A1(n5725), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5726) );
  MUX2_X1 U7184 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5726), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5728) );
  NAND2_X1 U7185 ( .A1(n5728), .A2(n5727), .ZN(n6406) );
  OR2_X1 U7186 ( .A1(n7877), .A2(n6297), .ZN(n5730) );
  OR2_X1 U7187 ( .A1(n5806), .A2(n6300), .ZN(n5729) );
  OAI211_X1 U7188 ( .C1(n6275), .C2(n6406), .A(n5730), .B(n5729), .ZN(n7038)
         );
  NAND2_X1 U7189 ( .A1(n7038), .A2(n5696), .ZN(n5731) );
  NAND2_X1 U7190 ( .A1(n5732), .A2(n5731), .ZN(n5734) );
  XNOR2_X1 U7191 ( .A(n5734), .B(n5733), .ZN(n6651) );
  AND2_X1 U7192 ( .A1(n7038), .A2(n6093), .ZN(n5735) );
  AOI21_X1 U7193 ( .B1(n8821), .B2(n5678), .A(n5735), .ZN(n6650) );
  NAND2_X1 U7194 ( .A1(n6651), .A2(n6650), .ZN(n5739) );
  INV_X1 U7195 ( .A(n5736), .ZN(n5738) );
  NAND2_X1 U7196 ( .A1(n5738), .A2(n5737), .ZN(n6648) );
  AND2_X1 U7197 ( .A1(n5739), .A2(n6648), .ZN(n5761) );
  NAND2_X1 U7198 ( .A1(n6649), .A2(n5761), .ZN(n5759) );
  INV_X1 U7199 ( .A(n6651), .ZN(n5741) );
  INV_X1 U7200 ( .A(n6650), .ZN(n5740) );
  NAND2_X1 U7201 ( .A1(n5741), .A2(n5740), .ZN(n5762) );
  AOI21_X1 U7202 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5742) );
  NOR2_X1 U7203 ( .A1(n5742), .A2(n5768), .ZN(n8751) );
  NAND2_X1 U7204 ( .A1(n6035), .A2(n8751), .ZN(n5751) );
  INV_X1 U7205 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5744) );
  OR2_X1 U7206 ( .A1(n4316), .A2(n5744), .ZN(n5750) );
  INV_X1 U7207 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5745) );
  OR2_X1 U7208 ( .A1(n5746), .A2(n5745), .ZN(n5749) );
  INV_X1 U7209 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5747) );
  OR2_X1 U7210 ( .A1(n6369), .A2(n5747), .ZN(n5748) );
  NAND4_X1 U7211 ( .A1(n5751), .A2(n5750), .A3(n5749), .A4(n5748), .ZN(n8820)
         );
  NAND2_X1 U7212 ( .A1(n8820), .A2(n6093), .ZN(n5756) );
  NAND2_X1 U7213 ( .A1(n5727), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5752) );
  XNOR2_X1 U7214 ( .A(n5752), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9742) );
  INV_X1 U7215 ( .A(n9742), .ZN(n6307) );
  OR2_X1 U7216 ( .A1(n5806), .A2(n6306), .ZN(n5754) );
  INV_X1 U7217 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6305) );
  OR2_X1 U7218 ( .A1(n7877), .A2(n6305), .ZN(n5753) );
  OAI211_X1 U7219 ( .C1(n6275), .C2(n6307), .A(n5754), .B(n5753), .ZN(n8750)
         );
  NAND2_X1 U7220 ( .A1(n8750), .A2(n5696), .ZN(n5755) );
  NAND2_X1 U7221 ( .A1(n5756), .A2(n5755), .ZN(n5757) );
  AND2_X1 U7222 ( .A1(n5762), .A2(n4340), .ZN(n5758) );
  AND2_X1 U7223 ( .A1(n6616), .A2(n5762), .ZN(n5760) );
  NAND2_X1 U7224 ( .A1(n6615), .A2(n5760), .ZN(n5765) );
  NAND2_X1 U7225 ( .A1(n5765), .A2(n5764), .ZN(n5766) );
  AND2_X1 U7226 ( .A1(n8750), .A2(n6093), .ZN(n5767) );
  AOI21_X1 U7227 ( .B1(n8820), .B2(n5678), .A(n5767), .ZN(n8748) );
  NAND2_X1 U7228 ( .A1(n6316), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5773) );
  INV_X1 U7229 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6411) );
  OR2_X1 U7230 ( .A1(n4316), .A2(n6411), .ZN(n5772) );
  OAI21_X1 U7231 ( .B1(n5768), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5784), .ZN(
        n7049) );
  OR2_X1 U7232 ( .A1(n5992), .A2(n7049), .ZN(n5771) );
  INV_X1 U7233 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5769) );
  OR2_X1 U7234 ( .A1(n6369), .A2(n5769), .ZN(n5770) );
  NAND4_X1 U7235 ( .A1(n5773), .A2(n5772), .A3(n5771), .A4(n5770), .ZN(n8819)
         );
  NAND2_X1 U7236 ( .A1(n8819), .A2(n6093), .ZN(n5779) );
  OR2_X1 U7237 ( .A1(n5774), .A2(n5965), .ZN(n5775) );
  XNOR2_X1 U7238 ( .A(n5775), .B(n5790), .ZN(n6410) );
  INV_X1 U7239 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6310) );
  OR2_X1 U7240 ( .A1(n7877), .A2(n6310), .ZN(n5777) );
  OR2_X1 U7241 ( .A1(n5806), .A2(n6309), .ZN(n5776) );
  NAND2_X1 U7242 ( .A1(n8123), .A2(n5696), .ZN(n5778) );
  NAND2_X1 U7243 ( .A1(n5779), .A2(n5778), .ZN(n5780) );
  XNOR2_X1 U7244 ( .A(n5780), .B(n5733), .ZN(n8117) );
  AND2_X1 U7245 ( .A1(n8123), .A2(n6093), .ZN(n5781) );
  AOI21_X1 U7246 ( .B1(n8819), .B2(n5678), .A(n5781), .ZN(n8116) );
  NAND2_X1 U7247 ( .A1(n6316), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5789) );
  INV_X1 U7248 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5782) );
  OR2_X1 U7249 ( .A1(n4316), .A2(n5782), .ZN(n5788) );
  AND2_X1 U7250 ( .A1(n5784), .A2(n5783), .ZN(n5785) );
  OR2_X1 U7251 ( .A1(n5785), .A2(n5800), .ZN(n7083) );
  OR2_X1 U7252 ( .A1(n5992), .A2(n7083), .ZN(n5787) );
  INV_X1 U7253 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7084) );
  OR2_X1 U7254 ( .A1(n6369), .A2(n7084), .ZN(n5786) );
  NAND4_X1 U7255 ( .A1(n5789), .A2(n5788), .A3(n5787), .A4(n5786), .ZN(n8818)
         );
  NAND2_X1 U7256 ( .A1(n8818), .A2(n6093), .ZN(n5795) );
  NAND2_X1 U7257 ( .A1(n5774), .A2(n5790), .ZN(n5807) );
  NAND2_X1 U7258 ( .A1(n5807), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5791) );
  XNOR2_X1 U7259 ( .A(n5791), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6429) );
  INV_X1 U7260 ( .A(n6429), .ZN(n6418) );
  OR2_X1 U7261 ( .A1(n6315), .A2(n5806), .ZN(n5793) );
  OR2_X1 U7262 ( .A1(n7877), .A2(n6314), .ZN(n5792) );
  NAND2_X1 U7263 ( .A1(n7102), .A2(n5696), .ZN(n5794) );
  NAND2_X1 U7264 ( .A1(n5795), .A2(n5794), .ZN(n5796) );
  XNOR2_X1 U7265 ( .A(n5796), .B(n5733), .ZN(n5798) );
  AOI22_X1 U7266 ( .A1(n8818), .A2(n5678), .B1(n6093), .B2(n7102), .ZN(n5797)
         );
  NAND2_X1 U7267 ( .A1(n5798), .A2(n5797), .ZN(n6278) );
  OR2_X1 U7268 ( .A1(n5798), .A2(n5797), .ZN(n6280) );
  NAND2_X1 U7269 ( .A1(n6200), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5805) );
  INV_X1 U7270 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5799) );
  OR2_X1 U7271 ( .A1(n5746), .A2(n5799), .ZN(n5804) );
  NAND2_X1 U7272 ( .A1(n5800), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5827) );
  OR2_X1 U7273 ( .A1(n5800), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U7274 ( .A1(n5827), .A2(n5801), .ZN(n7196) );
  OR2_X1 U7275 ( .A1(n5992), .A2(n7196), .ZN(n5803) );
  INV_X1 U7276 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6576) );
  OR2_X1 U7277 ( .A1(n6369), .A2(n6576), .ZN(n5802) );
  NAND4_X1 U7278 ( .A1(n5805), .A2(n5804), .A3(n5803), .A4(n5802), .ZN(n8817)
         );
  NAND2_X1 U7279 ( .A1(n8817), .A2(n5678), .ZN(n5814) );
  NAND2_X1 U7280 ( .A1(n6322), .A2(n5962), .ZN(n5812) );
  NAND2_X1 U7281 ( .A1(n5809), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5808) );
  MUX2_X1 U7282 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5808), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5810) );
  NAND2_X1 U7283 ( .A1(n5810), .A2(n5841), .ZN(n6577) );
  INV_X1 U7284 ( .A(n6577), .ZN(n6587) );
  AOI22_X1 U7285 ( .A1(n6030), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6029), .B2(
        n6587), .ZN(n5811) );
  NAND2_X1 U7286 ( .A1(n5812), .A2(n5811), .ZN(n7277) );
  NAND2_X1 U7287 ( .A1(n7277), .A2(n6093), .ZN(n5813) );
  NAND2_X1 U7288 ( .A1(n5814), .A2(n5813), .ZN(n5819) );
  NAND2_X1 U7289 ( .A1(n5818), .A2(n5819), .ZN(n7191) );
  NAND2_X1 U7290 ( .A1(n8817), .A2(n6093), .ZN(n5816) );
  NAND2_X1 U7291 ( .A1(n7277), .A2(n5696), .ZN(n5815) );
  NAND2_X1 U7292 ( .A1(n5816), .A2(n5815), .ZN(n5817) );
  XNOR2_X1 U7293 ( .A(n5817), .B(n5733), .ZN(n7194) );
  NAND2_X1 U7294 ( .A1(n7191), .A2(n7194), .ZN(n5822) );
  NAND2_X1 U7295 ( .A1(n6333), .A2(n5962), .ZN(n5825) );
  NAND2_X1 U7296 ( .A1(n5841), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5823) );
  XNOR2_X1 U7297 ( .A(n5823), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9769) );
  AOI22_X1 U7298 ( .A1(n6030), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6029), .B2(
        n9769), .ZN(n5824) );
  NAND2_X1 U7299 ( .A1(n7319), .A2(n5696), .ZN(n5835) );
  NAND2_X1 U7300 ( .A1(n6316), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U7301 ( .A1(n5827), .A2(n5826), .ZN(n5828) );
  NAND2_X1 U7302 ( .A1(n5848), .A2(n5828), .ZN(n7271) );
  OR2_X1 U7303 ( .A1(n5992), .A2(n7271), .ZN(n5832) );
  INV_X1 U7304 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7272) );
  OR2_X1 U7305 ( .A1(n6369), .A2(n7272), .ZN(n5831) );
  INV_X1 U7306 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5829) );
  OR2_X1 U7307 ( .A1(n4317), .A2(n5829), .ZN(n5830) );
  NAND4_X1 U7308 ( .A1(n5833), .A2(n5832), .A3(n5831), .A4(n5830), .ZN(n8816)
         );
  INV_X2 U7309 ( .A(n6217), .ZN(n6093) );
  NAND2_X1 U7310 ( .A1(n8816), .A2(n6093), .ZN(n5834) );
  NAND2_X1 U7311 ( .A1(n5835), .A2(n5834), .ZN(n5836) );
  XNOR2_X1 U7312 ( .A(n5836), .B(n5718), .ZN(n5837) );
  AOI22_X1 U7313 ( .A1(n7319), .A2(n6093), .B1(n5678), .B2(n8816), .ZN(n5838)
         );
  XNOR2_X1 U7314 ( .A(n5837), .B(n5838), .ZN(n7157) );
  INV_X1 U7315 ( .A(n5837), .ZN(n5839) );
  NAND2_X1 U7316 ( .A1(n5839), .A2(n5838), .ZN(n5840) );
  NAND2_X1 U7317 ( .A1(n6345), .A2(n5962), .ZN(n5846) );
  INV_X1 U7318 ( .A(n5841), .ZN(n5843) );
  INV_X1 U7319 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5842) );
  NAND2_X1 U7320 ( .A1(n5843), .A2(n5842), .ZN(n5861) );
  NAND2_X1 U7321 ( .A1(n5861), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5844) );
  XNOR2_X1 U7322 ( .A(n5844), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9782) );
  AOI22_X1 U7323 ( .A1(n6030), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6029), .B2(
        n9782), .ZN(n5845) );
  NAND2_X1 U7324 ( .A1(n9522), .A2(n5696), .ZN(n5855) );
  NAND2_X1 U7325 ( .A1(n6316), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5853) );
  INV_X1 U7326 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5847) );
  OR2_X1 U7327 ( .A1(n6369), .A2(n5847), .ZN(n5852) );
  INV_X1 U7328 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7209) );
  NAND2_X1 U7329 ( .A1(n5848), .A2(n7209), .ZN(n5849) );
  NAND2_X1 U7330 ( .A1(n5866), .A2(n5849), .ZN(n7210) );
  OR2_X1 U7331 ( .A1(n5992), .A2(n7210), .ZN(n5851) );
  INV_X1 U7332 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6584) );
  OR2_X1 U7333 ( .A1(n4317), .A2(n6584), .ZN(n5850) );
  NAND4_X1 U7334 ( .A1(n5853), .A2(n5852), .A3(n5851), .A4(n5850), .ZN(n9640)
         );
  NAND2_X1 U7335 ( .A1(n9640), .A2(n6093), .ZN(n5854) );
  NAND2_X1 U7336 ( .A1(n5855), .A2(n5854), .ZN(n5856) );
  XNOR2_X1 U7337 ( .A(n5856), .B(n5733), .ZN(n7206) );
  AND2_X1 U7338 ( .A1(n9640), .A2(n5678), .ZN(n5857) );
  AOI21_X1 U7339 ( .B1(n9522), .B2(n6093), .A(n5857), .ZN(n5858) );
  AND2_X1 U7340 ( .A1(n7206), .A2(n5858), .ZN(n5860) );
  INV_X1 U7341 ( .A(n7206), .ZN(n5859) );
  INV_X1 U7342 ( .A(n5858), .ZN(n7205) );
  NAND2_X1 U7343 ( .A1(n6349), .A2(n5962), .ZN(n5864) );
  OAI21_X1 U7344 ( .B1(n5861), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5862) );
  XNOR2_X1 U7345 ( .A(n5862), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6745) );
  AOI22_X1 U7346 ( .A1(n6030), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6029), .B2(
        n6745), .ZN(n5863) );
  NAND2_X1 U7347 ( .A1(n9650), .A2(n5696), .ZN(n5873) );
  NAND2_X1 U7348 ( .A1(n6316), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5871) );
  INV_X1 U7349 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9635) );
  OR2_X1 U7350 ( .A1(n6369), .A2(n9635), .ZN(n5870) );
  INV_X1 U7351 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5865) );
  AND2_X1 U7352 ( .A1(n5866), .A2(n5865), .ZN(n5867) );
  OR2_X1 U7353 ( .A1(n5867), .A2(n5888), .ZN(n9634) );
  OR2_X1 U7354 ( .A1(n5992), .A2(n9634), .ZN(n5869) );
  INV_X1 U7355 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6738) );
  OR2_X1 U7356 ( .A1(n4317), .A2(n6738), .ZN(n5868) );
  NAND4_X1 U7357 ( .A1(n5871), .A2(n5870), .A3(n5869), .A4(n5868), .ZN(n8815)
         );
  NAND2_X1 U7358 ( .A1(n8815), .A2(n6093), .ZN(n5872) );
  NAND2_X1 U7359 ( .A1(n5873), .A2(n5872), .ZN(n5874) );
  XNOR2_X1 U7360 ( .A(n5874), .B(n5718), .ZN(n5878) );
  AND2_X1 U7361 ( .A1(n8815), .A2(n5678), .ZN(n5875) );
  AOI21_X1 U7362 ( .B1(n9650), .B2(n6093), .A(n5875), .ZN(n5876) );
  XNOR2_X1 U7363 ( .A(n5878), .B(n5876), .ZN(n7334) );
  INV_X1 U7364 ( .A(n5876), .ZN(n5877) );
  NAND2_X1 U7365 ( .A1(n5878), .A2(n5877), .ZN(n5879) );
  NAND2_X1 U7366 ( .A1(n6380), .A2(n5962), .ZN(n5887) );
  NOR2_X1 U7367 ( .A1(n5881), .A2(n5965), .ZN(n5882) );
  MUX2_X1 U7368 ( .A(n5965), .B(n5882), .S(P1_IR_REG_12__SCAN_IN), .Z(n5885)
         );
  INV_X1 U7369 ( .A(n5884), .ZN(n5964) );
  OR2_X1 U7370 ( .A1(n5885), .A2(n5964), .ZN(n6832) );
  INV_X1 U7371 ( .A(n6832), .ZN(n6752) );
  AOI22_X1 U7372 ( .A1(n6030), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6029), .B2(
        n6752), .ZN(n5886) );
  NAND2_X1 U7373 ( .A1(n9237), .A2(n5696), .ZN(n5895) );
  NAND2_X1 U7374 ( .A1(n6316), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5893) );
  INV_X1 U7375 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6824) );
  OR2_X1 U7376 ( .A1(n4316), .A2(n6824), .ZN(n5892) );
  NAND2_X1 U7377 ( .A1(n5888), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5910) );
  OR2_X1 U7378 ( .A1(n5888), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5889) );
  NAND2_X1 U7379 ( .A1(n5910), .A2(n5889), .ZN(n7392) );
  OR2_X1 U7380 ( .A1(n5992), .A2(n7392), .ZN(n5891) );
  INV_X1 U7381 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6831) );
  OR2_X1 U7382 ( .A1(n6369), .A2(n6831), .ZN(n5890) );
  NAND4_X1 U7383 ( .A1(n5893), .A2(n5892), .A3(n5891), .A4(n5890), .ZN(n9639)
         );
  NAND2_X1 U7384 ( .A1(n9639), .A2(n6093), .ZN(n5894) );
  NAND2_X1 U7385 ( .A1(n5895), .A2(n5894), .ZN(n5896) );
  XNOR2_X1 U7386 ( .A(n5896), .B(n5733), .ZN(n5898) );
  AND2_X1 U7387 ( .A1(n9639), .A2(n5678), .ZN(n5897) );
  AOI21_X1 U7388 ( .B1(n9237), .B2(n6093), .A(n5897), .ZN(n5899) );
  NAND2_X1 U7389 ( .A1(n5898), .A2(n5899), .ZN(n5904) );
  INV_X1 U7390 ( .A(n5898), .ZN(n5901) );
  INV_X1 U7391 ( .A(n5899), .ZN(n5900) );
  NAND2_X1 U7392 ( .A1(n5901), .A2(n5900), .ZN(n5902) );
  NAND2_X1 U7393 ( .A1(n5904), .A2(n5902), .ZN(n7388) );
  INV_X1 U7394 ( .A(n7388), .ZN(n5903) );
  NAND2_X1 U7395 ( .A1(n6441), .A2(n5962), .ZN(n5907) );
  NAND2_X1 U7396 ( .A1(n5884), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5905) );
  XNOR2_X1 U7397 ( .A(n5905), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7256) );
  AOI22_X1 U7398 ( .A1(n6030), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6029), .B2(
        n7256), .ZN(n5906) );
  NAND2_X1 U7399 ( .A1(n9622), .A2(n5696), .ZN(n5917) );
  NAND2_X1 U7400 ( .A1(n6316), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5915) );
  INV_X1 U7401 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n5908) );
  OR2_X1 U7402 ( .A1(n4317), .A2(n5908), .ZN(n5914) );
  INV_X1 U7403 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7404 ( .A1(n5910), .A2(n5909), .ZN(n5911) );
  NAND2_X1 U7405 ( .A1(n5927), .A2(n5911), .ZN(n9609) );
  OR2_X1 U7406 ( .A1(n5992), .A2(n9609), .ZN(n5913) );
  INV_X1 U7407 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9610) );
  OR2_X1 U7408 ( .A1(n6369), .A2(n9610), .ZN(n5912) );
  NAND4_X1 U7409 ( .A1(n5915), .A2(n5914), .A3(n5913), .A4(n5912), .ZN(n8814)
         );
  NAND2_X1 U7410 ( .A1(n8814), .A2(n6093), .ZN(n5916) );
  NAND2_X1 U7411 ( .A1(n5917), .A2(n5916), .ZN(n5918) );
  XNOR2_X1 U7412 ( .A(n5918), .B(n5733), .ZN(n5920) );
  AND2_X1 U7413 ( .A1(n8814), .A2(n5678), .ZN(n5919) );
  AOI21_X1 U7414 ( .B1(n9622), .B2(n6093), .A(n5919), .ZN(n5921) );
  AND2_X1 U7415 ( .A1(n5920), .A2(n5921), .ZN(n7437) );
  INV_X1 U7416 ( .A(n5920), .ZN(n5923) );
  INV_X1 U7417 ( .A(n5921), .ZN(n5922) );
  NAND2_X1 U7418 ( .A1(n5923), .A2(n5922), .ZN(n7438) );
  NAND2_X1 U7419 ( .A1(n6623), .A2(n5962), .ZN(n5926) );
  OR2_X1 U7420 ( .A1(n5884), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7421 ( .A1(n5924), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5942) );
  XNOR2_X1 U7422 ( .A(n5942), .B(P1_IR_REG_14__SCAN_IN), .ZN(n8835) );
  AOI22_X1 U7423 ( .A1(n6030), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6029), .B2(
        n8835), .ZN(n5925) );
  NAND2_X1 U7424 ( .A1(n9232), .A2(n5696), .ZN(n5934) );
  NAND2_X1 U7425 ( .A1(n6316), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5932) );
  INV_X1 U7426 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7503) );
  OR2_X1 U7427 ( .A1(n6369), .A2(n7503), .ZN(n5931) );
  INV_X1 U7428 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7261) );
  AND2_X1 U7429 ( .A1(n5927), .A2(n7261), .ZN(n5928) );
  OR2_X1 U7430 ( .A1(n5928), .A2(n5950), .ZN(n7546) );
  OR2_X1 U7431 ( .A1(n5992), .A2(n7546), .ZN(n5930) );
  INV_X1 U7432 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7257) );
  OR2_X1 U7433 ( .A1(n4316), .A2(n7257), .ZN(n5929) );
  NAND4_X1 U7434 ( .A1(n5932), .A2(n5931), .A3(n5930), .A4(n5929), .ZN(n9616)
         );
  NAND2_X1 U7435 ( .A1(n9616), .A2(n6093), .ZN(n5933) );
  NAND2_X1 U7436 ( .A1(n5934), .A2(n5933), .ZN(n5935) );
  XNOR2_X1 U7437 ( .A(n5935), .B(n5718), .ZN(n5938) );
  NAND2_X1 U7438 ( .A1(n9232), .A2(n6199), .ZN(n5937) );
  NAND2_X1 U7439 ( .A1(n9616), .A2(n5678), .ZN(n5936) );
  NAND2_X1 U7440 ( .A1(n5937), .A2(n5936), .ZN(n7542) );
  NAND2_X1 U7441 ( .A1(n7540), .A2(n7542), .ZN(n5940) );
  NAND2_X1 U7442 ( .A1(n5939), .A2(n5938), .ZN(n7539) );
  NAND2_X1 U7443 ( .A1(n6721), .A2(n5962), .ZN(n5947) );
  NAND2_X1 U7444 ( .A1(n5942), .A2(n5941), .ZN(n5943) );
  NAND2_X1 U7445 ( .A1(n5943), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5945) );
  XNOR2_X1 U7446 ( .A(n5945), .B(n5944), .ZN(n8849) );
  INV_X1 U7447 ( .A(n8849), .ZN(n8838) );
  AOI22_X1 U7448 ( .A1(n6030), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6029), .B2(
        n8838), .ZN(n5946) );
  NAND2_X1 U7449 ( .A1(n9595), .A2(n5696), .ZN(n5957) );
  NAND2_X1 U7450 ( .A1(n6316), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5955) );
  INV_X1 U7451 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5948) );
  OR2_X1 U7452 ( .A1(n4317), .A2(n5948), .ZN(n5954) );
  INV_X1 U7453 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n5949) );
  OR2_X1 U7454 ( .A1(n6369), .A2(n5949), .ZN(n5953) );
  NOR2_X1 U7455 ( .A1(n5950), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5951) );
  OR2_X1 U7456 ( .A1(n5971), .A2(n5951), .ZN(n9592) );
  OR2_X1 U7457 ( .A1(n5992), .A2(n9592), .ZN(n5952) );
  NAND4_X1 U7458 ( .A1(n5955), .A2(n5954), .A3(n5953), .A4(n5952), .ZN(n8909)
         );
  NAND2_X1 U7459 ( .A1(n8909), .A2(n6093), .ZN(n5956) );
  NAND2_X1 U7460 ( .A1(n5957), .A2(n5956), .ZN(n5958) );
  XNOR2_X1 U7461 ( .A(n5958), .B(n5718), .ZN(n5961) );
  NAND2_X1 U7462 ( .A1(n9595), .A2(n6199), .ZN(n5960) );
  NAND2_X1 U7463 ( .A1(n8909), .A2(n5678), .ZN(n5959) );
  NAND2_X1 U7464 ( .A1(n5960), .A2(n5959), .ZN(n9574) );
  NAND2_X1 U7465 ( .A1(n6819), .A2(n5962), .ZN(n5969) );
  AND2_X1 U7466 ( .A1(n5964), .A2(n5963), .ZN(n5966) );
  OR2_X1 U7467 ( .A1(n5966), .A2(n5965), .ZN(n5967) );
  XNOR2_X1 U7468 ( .A(n5967), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8866) );
  AOI22_X1 U7469 ( .A1(n6030), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6029), .B2(
        n8866), .ZN(n5968) );
  NAND2_X1 U7470 ( .A1(n9227), .A2(n5696), .ZN(n5979) );
  NAND2_X1 U7471 ( .A1(n6316), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5977) );
  INV_X1 U7472 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5970) );
  OR2_X1 U7473 ( .A1(n6369), .A2(n5970), .ZN(n5976) );
  OR2_X1 U7474 ( .A1(n5971), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7475 ( .A1(n5990), .A2(n5972), .ZN(n8741) );
  OR2_X1 U7476 ( .A1(n5992), .A2(n8741), .ZN(n5975) );
  INV_X1 U7477 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n5973) );
  OR2_X1 U7478 ( .A1(n4316), .A2(n5973), .ZN(n5974) );
  NAND4_X1 U7479 ( .A1(n5977), .A2(n5976), .A3(n5975), .A4(n5974), .ZN(n8912)
         );
  NAND2_X1 U7480 ( .A1(n8912), .A2(n6093), .ZN(n5978) );
  NAND2_X1 U7481 ( .A1(n5979), .A2(n5978), .ZN(n5980) );
  XNOR2_X1 U7482 ( .A(n5980), .B(n5718), .ZN(n5982) );
  AND2_X1 U7483 ( .A1(n8912), .A2(n5678), .ZN(n5981) );
  AOI21_X1 U7484 ( .B1(n9227), .B2(n6199), .A(n5981), .ZN(n5983) );
  XNOR2_X1 U7485 ( .A(n5982), .B(n5983), .ZN(n8739) );
  INV_X1 U7486 ( .A(n5982), .ZN(n5984) );
  NAND2_X1 U7487 ( .A1(n5984), .A2(n5983), .ZN(n5985) );
  NAND2_X1 U7488 ( .A1(n8737), .A2(n5985), .ZN(n8757) );
  NAND2_X1 U7489 ( .A1(n6884), .A2(n5962), .ZN(n5988) );
  NAND2_X1 U7490 ( .A1(n5986), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6005) );
  XNOR2_X1 U7491 ( .A(n6005), .B(P1_IR_REG_17__SCAN_IN), .ZN(n8884) );
  AOI22_X1 U7492 ( .A1(n6030), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6029), .B2(
        n8884), .ZN(n5987) );
  NAND2_X1 U7493 ( .A1(n9222), .A2(n5696), .ZN(n5998) );
  NAND2_X1 U7494 ( .A1(n6316), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5996) );
  INV_X1 U7495 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n5989) );
  OR2_X1 U7496 ( .A1(n4316), .A2(n5989), .ZN(n5995) );
  INV_X1 U7497 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8760) );
  NAND2_X1 U7498 ( .A1(n5990), .A2(n8760), .ZN(n5991) );
  NAND2_X1 U7499 ( .A1(n6011), .A2(n5991), .ZN(n9127) );
  OR2_X1 U7500 ( .A1(n5992), .A2(n9127), .ZN(n5994) );
  INV_X1 U7501 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8861) );
  OR2_X1 U7502 ( .A1(n6369), .A2(n8861), .ZN(n5993) );
  NAND4_X1 U7503 ( .A1(n5996), .A2(n5995), .A3(n5994), .A4(n5993), .ZN(n8913)
         );
  NAND2_X1 U7504 ( .A1(n8913), .A2(n6093), .ZN(n5997) );
  NAND2_X1 U7505 ( .A1(n5998), .A2(n5997), .ZN(n5999) );
  XNOR2_X1 U7506 ( .A(n5999), .B(n5718), .ZN(n6001) );
  AND2_X1 U7507 ( .A1(n8913), .A2(n5678), .ZN(n6000) );
  AOI21_X1 U7508 ( .B1(n9222), .B2(n6093), .A(n6000), .ZN(n6002) );
  XNOR2_X1 U7509 ( .A(n6001), .B(n6002), .ZN(n8758) );
  NAND2_X1 U7510 ( .A1(n8757), .A2(n8758), .ZN(n8756) );
  INV_X1 U7511 ( .A(n6001), .ZN(n6003) );
  NAND2_X1 U7512 ( .A1(n6003), .A2(n6002), .ZN(n6004) );
  NAND2_X1 U7513 ( .A1(n8756), .A2(n6004), .ZN(n6024) );
  NAND2_X1 U7514 ( .A1(n6956), .A2(n5962), .ZN(n6009) );
  NAND2_X1 U7515 ( .A1(n6005), .A2(n4783), .ZN(n6006) );
  NAND2_X1 U7516 ( .A1(n6006), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6007) );
  XNOR2_X1 U7517 ( .A(n6007), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9788) );
  AOI22_X1 U7518 ( .A1(n6030), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6029), .B2(
        n9788), .ZN(n6008) );
  NAND2_X1 U7519 ( .A1(n9217), .A2(n5696), .ZN(n6020) );
  INV_X1 U7520 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6010) );
  AND2_X1 U7521 ( .A1(n6011), .A2(n6010), .ZN(n6012) );
  NOR2_X1 U7522 ( .A1(n6033), .A2(n6012), .ZN(n9118) );
  NAND2_X1 U7523 ( .A1(n6035), .A2(n9118), .ZN(n6018) );
  INV_X1 U7524 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n6013) );
  OR2_X1 U7525 ( .A1(n5746), .A2(n6013), .ZN(n6017) );
  INV_X1 U7526 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n6014) );
  OR2_X1 U7527 ( .A1(n6369), .A2(n6014), .ZN(n6016) );
  INV_X1 U7528 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8882) );
  OR2_X1 U7529 ( .A1(n4316), .A2(n8882), .ZN(n6015) );
  NAND4_X1 U7530 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .ZN(n9104)
         );
  NAND2_X1 U7531 ( .A1(n9104), .A2(n6093), .ZN(n6019) );
  NAND2_X1 U7532 ( .A1(n6020), .A2(n6019), .ZN(n6021) );
  XNOR2_X1 U7533 ( .A(n6021), .B(n5733), .ZN(n6025) );
  NAND2_X1 U7534 ( .A1(n6024), .A2(n6025), .ZN(n8790) );
  NAND2_X1 U7535 ( .A1(n9217), .A2(n6093), .ZN(n6023) );
  NAND2_X1 U7536 ( .A1(n9104), .A2(n5678), .ZN(n6022) );
  NAND2_X1 U7537 ( .A1(n6023), .A2(n6022), .ZN(n8793) );
  NAND2_X1 U7538 ( .A1(n8790), .A2(n8793), .ZN(n6028) );
  NAND2_X1 U7539 ( .A1(n7137), .A2(n5962), .ZN(n6032) );
  AOI22_X1 U7540 ( .A1(n6030), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9073), .B2(
        n6029), .ZN(n6031) );
  NAND2_X1 U7541 ( .A1(n9210), .A2(n5696), .ZN(n6043) );
  NAND2_X1 U7542 ( .A1(n6033), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6052) );
  OR2_X1 U7543 ( .A1(n6033), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6034) );
  AND2_X1 U7544 ( .A1(n6052), .A2(n6034), .ZN(n9097) );
  NAND2_X1 U7545 ( .A1(n9097), .A2(n6035), .ZN(n6041) );
  NAND2_X1 U7546 ( .A1(n6316), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6040) );
  INV_X1 U7547 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n6036) );
  OR2_X1 U7548 ( .A1(n4317), .A2(n6036), .ZN(n6039) );
  INV_X1 U7549 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n6037) );
  OR2_X1 U7550 ( .A1(n6369), .A2(n6037), .ZN(n6038) );
  NAND4_X1 U7551 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), .ZN(n9088)
         );
  NAND2_X1 U7552 ( .A1(n9088), .A2(n6093), .ZN(n6042) );
  NAND2_X1 U7553 ( .A1(n6043), .A2(n6042), .ZN(n6044) );
  XNOR2_X1 U7554 ( .A(n6044), .B(n5718), .ZN(n6046) );
  AND2_X1 U7555 ( .A1(n9088), .A2(n4319), .ZN(n6045) );
  AOI21_X1 U7556 ( .B1(n9210), .B2(n6093), .A(n6045), .ZN(n6047) );
  XNOR2_X1 U7557 ( .A(n6046), .B(n6047), .ZN(n8716) );
  INV_X1 U7558 ( .A(n6046), .ZN(n6048) );
  NAND2_X1 U7559 ( .A1(n6048), .A2(n6047), .ZN(n6049) );
  NAND2_X1 U7560 ( .A1(n7250), .A2(n5962), .ZN(n6051) );
  OR2_X1 U7561 ( .A1(n7877), .A2(n7298), .ZN(n6050) );
  NAND2_X1 U7562 ( .A1(n9205), .A2(n5696), .ZN(n6061) );
  INV_X1 U7563 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8775) );
  NAND2_X1 U7564 ( .A1(n6052), .A2(n8775), .ZN(n6053) );
  NAND2_X1 U7565 ( .A1(n6069), .A2(n6053), .ZN(n9081) );
  NOR2_X1 U7566 ( .A1(n9081), .A2(n5992), .ZN(n6059) );
  INV_X1 U7567 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7568 ( .A1(n6316), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6054) );
  OAI21_X1 U7569 ( .B1(n4317), .B2(n6055), .A(n6054), .ZN(n6058) );
  INV_X1 U7570 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n6056) );
  NOR2_X1 U7571 ( .A1(n6369), .A2(n6056), .ZN(n6057) );
  NAND2_X1 U7572 ( .A1(n9103), .A2(n6093), .ZN(n6060) );
  NAND2_X1 U7573 ( .A1(n6061), .A2(n6060), .ZN(n6062) );
  XNOR2_X1 U7574 ( .A(n6062), .B(n5718), .ZN(n6064) );
  AND2_X1 U7575 ( .A1(n9103), .A2(n5678), .ZN(n6063) );
  AOI21_X1 U7576 ( .B1(n9205), .B2(n6093), .A(n6063), .ZN(n6065) );
  XNOR2_X1 U7577 ( .A(n6064), .B(n6065), .ZN(n8774) );
  INV_X1 U7578 ( .A(n6064), .ZN(n6066) );
  NAND2_X1 U7579 ( .A1(n7267), .A2(n5962), .ZN(n6068) );
  INV_X1 U7580 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7268) );
  OR2_X1 U7581 ( .A1(n7877), .A2(n7268), .ZN(n6067) );
  NAND2_X1 U7582 ( .A1(n9202), .A2(n5696), .ZN(n6074) );
  INV_X1 U7583 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8724) );
  AND2_X1 U7584 ( .A1(n6069), .A2(n8724), .ZN(n6070) );
  OR2_X1 U7585 ( .A1(n6083), .A2(n6070), .ZN(n9072) );
  AOI22_X1 U7586 ( .A1(n6316), .A2(P1_REG0_REG_21__SCAN_IN), .B1(n6085), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7587 ( .A1(n6200), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6071) );
  OAI211_X1 U7588 ( .C1(n9072), .C2(n5992), .A(n6072), .B(n6071), .ZN(n9087)
         );
  NAND2_X1 U7589 ( .A1(n9087), .A2(n6093), .ZN(n6073) );
  NAND2_X1 U7590 ( .A1(n6074), .A2(n6073), .ZN(n6075) );
  XNOR2_X1 U7591 ( .A(n6075), .B(n5718), .ZN(n6077) );
  AND2_X1 U7592 ( .A1(n9087), .A2(n4319), .ZN(n6076) );
  AOI21_X1 U7593 ( .B1(n9202), .B2(n6093), .A(n6076), .ZN(n6078) );
  XNOR2_X1 U7594 ( .A(n6077), .B(n6078), .ZN(n8723) );
  INV_X1 U7595 ( .A(n6077), .ZN(n6079) );
  NAND2_X1 U7596 ( .A1(n6079), .A2(n6078), .ZN(n6080) );
  NAND2_X1 U7597 ( .A1(n7345), .A2(n5962), .ZN(n6082) );
  OR2_X1 U7598 ( .A1(n7877), .A2(n7346), .ZN(n6081) );
  OR2_X1 U7599 ( .A1(n6083), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7600 ( .A1(n6083), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7601 ( .A1(n6084), .A2(n6104), .ZN(n9057) );
  OR2_X1 U7602 ( .A1(n9057), .A2(n5992), .ZN(n6091) );
  INV_X1 U7603 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7604 ( .A1(n6085), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7605 ( .A1(n6316), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6086) );
  OAI211_X1 U7606 ( .C1(n4316), .C2(n6088), .A(n6087), .B(n6086), .ZN(n6089)
         );
  INV_X1 U7607 ( .A(n6089), .ZN(n6090) );
  NAND2_X1 U7608 ( .A1(n6091), .A2(n6090), .ZN(n9038) );
  AND2_X1 U7609 ( .A1(n9038), .A2(n5678), .ZN(n6092) );
  AOI21_X1 U7610 ( .B1(n9197), .B2(n6093), .A(n6092), .ZN(n6098) );
  NAND2_X1 U7611 ( .A1(n9197), .A2(n5696), .ZN(n6096) );
  NAND2_X1 U7612 ( .A1(n9038), .A2(n6093), .ZN(n6095) );
  NAND2_X1 U7613 ( .A1(n6096), .A2(n6095), .ZN(n6097) );
  XNOR2_X1 U7614 ( .A(n6097), .B(n5733), .ZN(n8783) );
  NAND2_X1 U7615 ( .A1(n8781), .A2(n8783), .ZN(n6100) );
  NAND2_X1 U7616 ( .A1(n7384), .A2(n5962), .ZN(n6102) );
  OR2_X1 U7617 ( .A1(n7877), .A2(n7383), .ZN(n6101) );
  NAND2_X1 U7618 ( .A1(n9192), .A2(n5696), .ZN(n6113) );
  NAND2_X1 U7619 ( .A1(n6200), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6111) );
  INV_X1 U7620 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n6103) );
  OR2_X1 U7621 ( .A1(n5746), .A2(n6103), .ZN(n6110) );
  OAI21_X1 U7622 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n6105), .A(n6125), .ZN(
        n9043) );
  OR2_X1 U7623 ( .A1(n5992), .A2(n9043), .ZN(n6109) );
  INV_X1 U7624 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6106) );
  OR2_X1 U7625 ( .A1(n6107), .A2(n6106), .ZN(n6108) );
  NAND4_X1 U7626 ( .A1(n6111), .A2(n6110), .A3(n6109), .A4(n6108), .ZN(n8919)
         );
  NAND2_X1 U7627 ( .A1(n8919), .A2(n6093), .ZN(n6112) );
  NAND2_X1 U7628 ( .A1(n6113), .A2(n6112), .ZN(n6114) );
  XNOR2_X1 U7629 ( .A(n6114), .B(n5733), .ZN(n6117) );
  AND2_X1 U7630 ( .A1(n8919), .A2(n4319), .ZN(n6116) );
  AOI21_X1 U7631 ( .B1(n9192), .B2(n6093), .A(n6116), .ZN(n8708) );
  NAND2_X1 U7632 ( .A1(n6118), .A2(n6117), .ZN(n8707) );
  NAND2_X1 U7633 ( .A1(n6119), .A2(n8707), .ZN(n8766) );
  NAND2_X1 U7634 ( .A1(n7494), .A2(n5962), .ZN(n6121) );
  INV_X1 U7635 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7497) );
  OR2_X1 U7636 ( .A1(n7877), .A2(n7497), .ZN(n6120) );
  NAND2_X1 U7637 ( .A1(n9187), .A2(n5696), .ZN(n6133) );
  NAND2_X1 U7638 ( .A1(n6316), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6131) );
  INV_X1 U7639 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6122) );
  OR2_X1 U7640 ( .A1(n4316), .A2(n6122), .ZN(n6130) );
  INV_X1 U7641 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7642 ( .A1(n6125), .A2(n6124), .ZN(n6126) );
  NAND2_X1 U7643 ( .A1(n6145), .A2(n6126), .ZN(n9028) );
  OR2_X1 U7644 ( .A1(n5992), .A2(n9028), .ZN(n6129) );
  INV_X1 U7645 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6127) );
  OR2_X1 U7646 ( .A1(n6369), .A2(n6127), .ZN(n6128) );
  NAND4_X1 U7647 ( .A1(n6131), .A2(n6130), .A3(n6129), .A4(n6128), .ZN(n9037)
         );
  NAND2_X1 U7648 ( .A1(n9037), .A2(n6093), .ZN(n6132) );
  NAND2_X1 U7649 ( .A1(n6133), .A2(n6132), .ZN(n6134) );
  XNOR2_X1 U7650 ( .A(n6134), .B(n5718), .ZN(n6136) );
  AND2_X1 U7651 ( .A1(n9037), .A2(n4319), .ZN(n6135) );
  AOI21_X1 U7652 ( .B1(n9187), .B2(n6093), .A(n6135), .ZN(n6137) );
  XNOR2_X1 U7653 ( .A(n6136), .B(n6137), .ZN(n8767) );
  INV_X1 U7654 ( .A(n6136), .ZN(n6138) );
  NAND2_X1 U7655 ( .A1(n6138), .A2(n6137), .ZN(n6139) );
  NAND2_X1 U7656 ( .A1(n7523), .A2(n5962), .ZN(n6141) );
  OR2_X1 U7657 ( .A1(n7877), .A2(n7526), .ZN(n6140) );
  NAND2_X1 U7658 ( .A1(n9180), .A2(n5696), .ZN(n6153) );
  NAND2_X1 U7659 ( .A1(n6316), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6151) );
  INV_X1 U7660 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6142) );
  OR2_X1 U7661 ( .A1(n4317), .A2(n6142), .ZN(n6150) );
  INV_X1 U7662 ( .A(n6145), .ZN(n6143) );
  NAND2_X1 U7663 ( .A1(n6143), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6164) );
  INV_X1 U7664 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7665 ( .A1(n6145), .A2(n6144), .ZN(n6146) );
  NAND2_X1 U7666 ( .A1(n6164), .A2(n6146), .ZN(n9007) );
  OR2_X1 U7667 ( .A1(n5992), .A2(n9007), .ZN(n6149) );
  INV_X1 U7668 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n6147) );
  OR2_X1 U7669 ( .A1(n6369), .A2(n6147), .ZN(n6148) );
  NAND4_X1 U7670 ( .A1(n6151), .A2(n6150), .A3(n6149), .A4(n6148), .ZN(n8998)
         );
  NAND2_X1 U7671 ( .A1(n8998), .A2(n6199), .ZN(n6152) );
  NAND2_X1 U7672 ( .A1(n6153), .A2(n6152), .ZN(n6154) );
  XNOR2_X1 U7673 ( .A(n6154), .B(n5718), .ZN(n6156) );
  AND2_X1 U7674 ( .A1(n8998), .A2(n5678), .ZN(n6155) );
  AOI21_X1 U7675 ( .B1(n9180), .B2(n6093), .A(n6155), .ZN(n6157) );
  XNOR2_X1 U7676 ( .A(n6156), .B(n6157), .ZN(n8731) );
  INV_X1 U7677 ( .A(n6156), .ZN(n6158) );
  OR2_X1 U7678 ( .A1(n7877), .A2(n7553), .ZN(n6159) );
  NAND2_X1 U7679 ( .A1(n9175), .A2(n5696), .ZN(n6172) );
  NAND2_X1 U7680 ( .A1(n6200), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6170) );
  INV_X1 U7681 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n6161) );
  OR2_X1 U7682 ( .A1(n5746), .A2(n6161), .ZN(n6169) );
  INV_X1 U7683 ( .A(n6164), .ZN(n6162) );
  INV_X1 U7684 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7685 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  NAND2_X1 U7686 ( .A1(n6204), .A2(n6165), .ZN(n8991) );
  INV_X1 U7687 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6166) );
  OR2_X1 U7688 ( .A1(n6369), .A2(n6166), .ZN(n6167) );
  NAND4_X1 U7689 ( .A1(n6170), .A2(n6169), .A3(n6168), .A4(n6167), .ZN(n9015)
         );
  NAND2_X1 U7690 ( .A1(n9015), .A2(n6199), .ZN(n6171) );
  NAND2_X1 U7691 ( .A1(n6172), .A2(n6171), .ZN(n6173) );
  XNOR2_X1 U7692 ( .A(n6173), .B(n5733), .ZN(n6178) );
  INV_X1 U7693 ( .A(n6178), .ZN(n6176) );
  AND2_X1 U7694 ( .A1(n9015), .A2(n4319), .ZN(n6174) );
  AOI21_X1 U7695 ( .B1(n9175), .B2(n6093), .A(n6174), .ZN(n6177) );
  INV_X1 U7696 ( .A(n6177), .ZN(n6175) );
  NAND2_X1 U7697 ( .A1(n6176), .A2(n6175), .ZN(n8803) );
  OR2_X1 U7698 ( .A1(n7877), .A2(n6179), .ZN(n6180) );
  NAND2_X1 U7699 ( .A1(n9172), .A2(n5696), .ZN(n6189) );
  NAND2_X1 U7700 ( .A1(n6316), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6187) );
  INV_X1 U7701 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6182) );
  OR2_X1 U7702 ( .A1(n4317), .A2(n6182), .ZN(n6186) );
  INV_X1 U7703 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6203) );
  XNOR2_X1 U7704 ( .A(n6204), .B(n6203), .ZN(n8146) );
  INV_X1 U7705 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6183) );
  OR2_X1 U7706 ( .A1(n6369), .A2(n6183), .ZN(n6184) );
  NAND4_X1 U7707 ( .A1(n6187), .A2(n6186), .A3(n6185), .A4(n6184), .ZN(n8997)
         );
  NAND2_X1 U7708 ( .A1(n8997), .A2(n6199), .ZN(n6188) );
  NAND2_X1 U7709 ( .A1(n6189), .A2(n6188), .ZN(n6190) );
  XNOR2_X1 U7710 ( .A(n6190), .B(n5733), .ZN(n6192) );
  AND2_X1 U7711 ( .A1(n8997), .A2(n4319), .ZN(n6191) );
  AOI21_X1 U7712 ( .B1(n9172), .B2(n6093), .A(n6191), .ZN(n6193) );
  NAND2_X1 U7713 ( .A1(n6192), .A2(n6193), .ZN(n6266) );
  INV_X1 U7714 ( .A(n6192), .ZN(n6195) );
  INV_X1 U7715 ( .A(n6193), .ZN(n6194) );
  NAND2_X1 U7716 ( .A1(n6195), .A2(n6194), .ZN(n6196) );
  NAND2_X1 U7717 ( .A1(n6266), .A2(n6196), .ZN(n8144) );
  NAND2_X1 U7718 ( .A1(n9271), .A2(n5962), .ZN(n6198) );
  INV_X1 U7719 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9273) );
  OR2_X1 U7720 ( .A1(n7877), .A2(n9273), .ZN(n6197) );
  NAND2_X1 U7721 ( .A1(n9166), .A2(n6199), .ZN(n6214) );
  NAND2_X1 U7722 ( .A1(n6200), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6212) );
  INV_X1 U7723 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6201) );
  OR2_X1 U7724 ( .A1(n5746), .A2(n6201), .ZN(n6211) );
  INV_X1 U7725 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6202) );
  OAI21_X1 U7726 ( .B1(n6204), .B2(n6203), .A(n6202), .ZN(n6207) );
  INV_X1 U7727 ( .A(n6204), .ZN(n6206) );
  AND2_X1 U7728 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6205) );
  NAND2_X1 U7729 ( .A1(n6206), .A2(n6205), .ZN(n8956) );
  NAND2_X1 U7730 ( .A1(n6207), .A2(n8956), .ZN(n8968) );
  OR2_X1 U7731 ( .A1(n5992), .A2(n8968), .ZN(n6210) );
  INV_X1 U7732 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n6208) );
  OR2_X1 U7733 ( .A1(n6369), .A2(n6208), .ZN(n6209) );
  OR2_X1 U7734 ( .A1(n4318), .A2(n8981), .ZN(n6213) );
  NAND2_X1 U7735 ( .A1(n6214), .A2(n6213), .ZN(n6215) );
  XNOR2_X1 U7736 ( .A(n6215), .B(n5733), .ZN(n6219) );
  NAND2_X1 U7737 ( .A1(n9166), .A2(n5696), .ZN(n6216) );
  OAI21_X1 U7738 ( .B1(n8981), .B2(n6217), .A(n6216), .ZN(n6218) );
  XNOR2_X1 U7739 ( .A(n6219), .B(n6218), .ZN(n6246) );
  INV_X1 U7740 ( .A(n6246), .ZN(n6267) );
  NAND2_X1 U7741 ( .A1(n7528), .A2(P1_B_REG_SCAN_IN), .ZN(n6221) );
  MUX2_X1 U7742 ( .A(n6221), .B(P1_B_REG_SCAN_IN), .S(n6220), .Z(n6222) );
  INV_X1 U7743 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6313) );
  INV_X1 U7744 ( .A(n6223), .ZN(n7555) );
  AND2_X1 U7745 ( .A1(n7555), .A2(n7499), .ZN(n6224) );
  AOI21_X1 U7746 ( .B1(n6443), .B2(n6313), .A(n6224), .ZN(n6700) );
  NOR2_X1 U7747 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n6228) );
  NOR4_X1 U7748 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6227) );
  NOR4_X1 U7749 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6226) );
  NOR4_X1 U7750 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6225) );
  NAND4_X1 U7751 ( .A1(n6228), .A2(n6227), .A3(n6226), .A4(n6225), .ZN(n6234)
         );
  NOR4_X1 U7752 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6232) );
  NOR4_X1 U7753 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6231) );
  NOR4_X1 U7754 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6230) );
  NOR4_X1 U7755 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6229) );
  NAND4_X1 U7756 ( .A1(n6232), .A2(n6231), .A3(n6230), .A4(n6229), .ZN(n6233)
         );
  OAI21_X1 U7757 ( .B1(n6234), .B2(n6233), .A(n6443), .ZN(n6698) );
  NAND2_X1 U7758 ( .A1(n6700), .A2(n6698), .ZN(n6865) );
  INV_X1 U7759 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6446) );
  NAND2_X1 U7760 ( .A1(n6443), .A2(n6446), .ZN(n6235) );
  NAND2_X1 U7761 ( .A1(n7555), .A2(n7528), .ZN(n6444) );
  NAND2_X1 U7762 ( .A1(n6235), .A2(n6444), .ZN(n6697) );
  OR2_X1 U7763 ( .A1(n6865), .A2(n6697), .ZN(n6659) );
  NAND2_X1 U7764 ( .A1(n6236), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6237) );
  MUX2_X1 U7765 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6237), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n6239) );
  NAND2_X1 U7766 ( .A1(n6239), .A2(n6238), .ZN(n7381) );
  NAND2_X1 U7767 ( .A1(n7381), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6273) );
  INV_X1 U7768 ( .A(n6273), .ZN(n6240) );
  NOR2_X1 U7769 ( .A1(n6659), .A2(n8084), .ZN(n6255) );
  NAND2_X1 U7770 ( .A1(n6242), .A2(n6243), .ZN(n6927) );
  NAND2_X1 U7771 ( .A1(n8087), .A2(n8072), .ZN(n7999) );
  AND2_X1 U7772 ( .A1(n9854), .A2(n7999), .ZN(n6244) );
  NAND2_X1 U7773 ( .A1(n6255), .A2(n6244), .ZN(n8812) );
  NAND3_X1 U7774 ( .A1(n6267), .A2(n9576), .A3(n6266), .ZN(n6245) );
  NAND2_X1 U7775 ( .A1(n8143), .A2(n6247), .ZN(n6271) );
  OR2_X1 U7776 ( .A1(n6927), .A2(n5656), .ZN(n6929) );
  INV_X1 U7777 ( .A(n6929), .ZN(n6248) );
  NAND3_X1 U7778 ( .A1(n6248), .A2(n6447), .A3(n6659), .ZN(n6252) );
  OR2_X1 U7779 ( .A1(n7999), .A2(n6926), .ZN(n6249) );
  AND2_X1 U7780 ( .A1(n6252), .A2(n6703), .ZN(n9570) );
  NAND2_X1 U7781 ( .A1(n9854), .A2(n6659), .ZN(n6250) );
  NAND4_X1 U7782 ( .A1(n6250), .A2(n6354), .A3(n7381), .A4(n6249), .ZN(n6251)
         );
  NAND2_X1 U7783 ( .A1(n6251), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6253) );
  OR2_X1 U7784 ( .A1(n6688), .A2(n6687), .ZN(n8085) );
  INV_X1 U7785 ( .A(n8085), .ZN(n6254) );
  AND2_X1 U7786 ( .A1(n6255), .A2(n6254), .ZN(n6257) );
  INV_X1 U7787 ( .A(n9711), .ZN(n9691) );
  AND2_X2 U7788 ( .A1(n6257), .A2(n9691), .ZN(n9564) );
  AOI22_X1 U7789 ( .A1(n9564), .A2(n8997), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6265) );
  INV_X1 U7790 ( .A(n6257), .ZN(n6258) );
  NAND2_X1 U7791 ( .A1(n6316), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6263) );
  INV_X1 U7792 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8957) );
  OR2_X1 U7793 ( .A1(n6369), .A2(n8957), .ZN(n6262) );
  OR2_X1 U7794 ( .A1(n5992), .A2(n8956), .ZN(n6261) );
  INV_X1 U7795 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6259) );
  OR2_X1 U7796 ( .A1(n4316), .A2(n6259), .ZN(n6260) );
  NAND4_X1 U7797 ( .A1(n6263), .A2(n6262), .A3(n6261), .A4(n6260), .ZN(n8974)
         );
  NAND2_X1 U7798 ( .A1(n8806), .A2(n8974), .ZN(n6264) );
  OAI211_X1 U7799 ( .C1(n9580), .C2(n8968), .A(n6265), .B(n6264), .ZN(n6269)
         );
  NOR3_X1 U7800 ( .A1(n6267), .A2(n8812), .A3(n6266), .ZN(n6268) );
  AOI211_X1 U7801 ( .C1(n8810), .C2(n9166), .A(n6269), .B(n6268), .ZN(n6270)
         );
  NAND3_X1 U7802 ( .A1(n6272), .A2(n6271), .A3(n6270), .ZN(P1_U3218) );
  OR2_X1 U7803 ( .A1(n6354), .A2(n6273), .ZN(n8824) );
  INV_X1 U7804 ( .A(n8824), .ZN(P1_U4006) );
  NAND2_X1 U7805 ( .A1(n7999), .A2(n6354), .ZN(n6274) );
  NAND2_X1 U7806 ( .A1(n6274), .A2(n7381), .ZN(n6357) );
  NAND2_X1 U7807 ( .A1(n6357), .A2(n6275), .ZN(n9685) );
  NAND2_X1 U7808 ( .A1(n9685), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U7809 ( .A(n9979), .ZN(n6276) );
  NOR2_X2 U7810 ( .A1(n6449), .A2(n6276), .ZN(P2_U3966) );
  AOI21_X1 U7811 ( .B1(n6280), .B2(n6278), .A(n6277), .ZN(n6279) );
  AOI211_X1 U7812 ( .C1(n4393), .C2(n6280), .A(n8812), .B(n6279), .ZN(n6287)
         );
  AND2_X1 U7813 ( .A1(n8810), .A2(n7102), .ZN(n6286) );
  NOR2_X1 U7814 ( .A1(n9580), .A2(n7083), .ZN(n6285) );
  INV_X1 U7815 ( .A(n8817), .ZN(n6283) );
  NAND2_X1 U7816 ( .A1(n9564), .A2(n8819), .ZN(n6282) );
  AND2_X1 U7817 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6415) );
  INV_X1 U7818 ( .A(n6415), .ZN(n6281) );
  OAI211_X1 U7819 ( .C1(n6283), .C2(n9568), .A(n6282), .B(n6281), .ZN(n6284)
         );
  OR4_X1 U7820 ( .A1(n6287), .A2(n6286), .A3(n6285), .A4(n6284), .ZN(P1_U3211)
         );
  XNOR2_X1 U7821 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U7822 ( .A(n6288), .ZN(n6289) );
  NAND2_X1 U7823 ( .A1(P1_STATE_REG_SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9686) );
  OAI21_X1 U7824 ( .B1(n6289), .B2(P1_STATE_REG_SCAN_IN), .A(n9686), .ZN(
        P1_U3353) );
  AND2_X1 U7825 ( .A1(n6292), .A2(P2_U3152), .ZN(n8690) );
  INV_X1 U7826 ( .A(n8690), .ZN(n8704) );
  OR2_X1 U7827 ( .A1(n6292), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8695) );
  OAI222_X1 U7828 ( .A1(n8704), .A2(n6291), .B1(n8695), .B2(n6293), .C1(
        P2_U3152), .C2(n6290), .ZN(P2_U3355) );
  AND2_X1 U7829 ( .A1(n7589), .A2(P1_U3084), .ZN(n9270) );
  INV_X2 U7830 ( .A(n9270), .ZN(n9277) );
  OAI222_X1 U7831 ( .A1(n4314), .A2(n6294), .B1(n9277), .B2(n6293), .C1(n6400), 
        .C2(P1_U3084), .ZN(P1_U3350) );
  OAI222_X1 U7832 ( .A1(n4314), .A2(n6295), .B1(n9277), .B2(n6302), .C1(n6393), 
        .C2(P1_U3084), .ZN(P1_U3351) );
  OAI222_X1 U7833 ( .A1(n4314), .A2(n6296), .B1(n9277), .B2(n6299), .C1(n6361), 
        .C2(P1_U3084), .ZN(P1_U3352) );
  OAI222_X1 U7834 ( .A1(n4314), .A2(n6297), .B1(n9277), .B2(n6300), .C1(n6406), 
        .C2(P1_U3084), .ZN(P1_U3349) );
  INV_X1 U7835 ( .A(n8695), .ZN(n8696) );
  INV_X1 U7836 ( .A(n8696), .ZN(n8702) );
  OAI222_X1 U7837 ( .A1(P2_U3152), .A2(n6477), .B1(n8702), .B2(n6299), .C1(
        n6298), .C2(n8704), .ZN(P2_U3357) );
  OAI222_X1 U7838 ( .A1(n8704), .A2(n6301), .B1(n8702), .B2(n6300), .C1(
        P2_U3152), .C2(n6475), .ZN(P2_U3354) );
  OAI222_X1 U7839 ( .A1(P2_U3152), .A2(n9516), .B1(n8702), .B2(n6302), .C1(
        n4422), .C2(n8704), .ZN(P2_U3356) );
  OAI222_X1 U7840 ( .A1(n8704), .A2(n6304), .B1(n8695), .B2(n6306), .C1(
        P2_U3152), .C2(n6303), .ZN(P2_U3353) );
  OAI222_X1 U7841 ( .A1(n6307), .A2(P1_U3084), .B1(n9277), .B2(n6306), .C1(
        n6305), .C2(n4314), .ZN(P1_U3348) );
  AOI22_X1 U7842 ( .A1(n6505), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n8690), .ZN(n6308) );
  OAI21_X1 U7843 ( .B1(n6309), .B2(n8695), .A(n6308), .ZN(P2_U3352) );
  OAI222_X1 U7844 ( .A1(n4314), .A2(n6310), .B1(n9277), .B2(n6309), .C1(n6410), 
        .C2(P1_U3084), .ZN(P1_U3347) );
  AOI22_X1 U7845 ( .A1(n6517), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n8690), .ZN(n6311) );
  OAI21_X1 U7846 ( .B1(n6315), .B2(n8695), .A(n6311), .ZN(P2_U3351) );
  NAND2_X1 U7847 ( .A1(n6700), .A2(n6447), .ZN(n6312) );
  OAI21_X1 U7848 ( .B1(n6313), .B2(n6447), .A(n6312), .ZN(P1_U3440) );
  OAI222_X1 U7849 ( .A1(n6418), .A2(P1_U3084), .B1(n9277), .B2(n6315), .C1(
        n6314), .C2(n4314), .ZN(P1_U3346) );
  INV_X1 U7850 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6321) );
  INV_X1 U7851 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U7852 ( .A1(n6316), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6318) );
  INV_X1 U7853 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8898) );
  OR2_X1 U7854 ( .A1(n6369), .A2(n8898), .ZN(n6317) );
  OAI211_X1 U7855 ( .C1(n4317), .C2(n6319), .A(n6318), .B(n6317), .ZN(n8896)
         );
  NAND2_X1 U7856 ( .A1(n8896), .A2(P1_U4006), .ZN(n6320) );
  OAI21_X1 U7857 ( .B1(P1_U4006), .B2(n6321), .A(n6320), .ZN(P1_U3586) );
  INV_X1 U7858 ( .A(n6322), .ZN(n6324) );
  AOI22_X1 U7859 ( .A1(n6572), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n8690), .ZN(n6323) );
  OAI21_X1 U7860 ( .B1(n6324), .B2(n8695), .A(n6323), .ZN(P2_U3350) );
  OAI222_X1 U7861 ( .A1(n4314), .A2(n6325), .B1(n9277), .B2(n6324), .C1(n6577), 
        .C2(P1_U3084), .ZN(P1_U3345) );
  INV_X1 U7862 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U7863 ( .A1(n7580), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6329) );
  NAND2_X1 U7864 ( .A1(n4315), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6328) );
  NAND2_X1 U7865 ( .A1(n6326), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6327) );
  AND3_X1 U7866 ( .A1(n6329), .A2(n6328), .A3(n6327), .ZN(n8331) );
  INV_X1 U7867 ( .A(n8331), .ZN(n6330) );
  NAND2_X1 U7868 ( .A1(n6330), .A2(P2_U3966), .ZN(n6331) );
  OAI21_X1 U7869 ( .B1(P2_U3966), .B2(n6332), .A(n6331), .ZN(P2_U3583) );
  INV_X1 U7870 ( .A(n6333), .ZN(n6336) );
  AOI22_X1 U7871 ( .A1(n6608), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n8690), .ZN(n6334) );
  OAI21_X1 U7872 ( .B1(n6336), .B2(n8695), .A(n6334), .ZN(P2_U3349) );
  AOI22_X1 U7874 ( .A1(n9769), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n4313), .ZN(n6335) );
  OAI21_X1 U7875 ( .B1(n6336), .B2(n9277), .A(n6335), .ZN(P1_U3344) );
  OAI21_X1 U7876 ( .B1(n9972), .B2(n7811), .A(n6338), .ZN(n6341) );
  NAND2_X1 U7877 ( .A1(n9972), .A2(n6339), .ZN(n6340) );
  INV_X1 U7878 ( .A(n8325), .ZN(n9926) );
  NOR2_X1 U7879 ( .A1(n9926), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X2 U7880 ( .A(P2_U3966), .ZN(n8264) );
  NAND2_X1 U7881 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n8264), .ZN(n6342) );
  OAI21_X1 U7882 ( .B1(n8092), .B2(n8264), .A(n6342), .ZN(P2_U3566) );
  NAND2_X1 U7883 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n8264), .ZN(n6343) );
  OAI21_X1 U7884 ( .B1(n7459), .B2(n8264), .A(n6343), .ZN(P2_U3565) );
  NAND2_X1 U7885 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n8264), .ZN(n6344) );
  OAI21_X1 U7886 ( .B1(n8536), .B2(n8264), .A(n6344), .ZN(P2_U3569) );
  INV_X1 U7887 ( .A(n6345), .ZN(n6348) );
  AOI22_X1 U7888 ( .A1(n9782), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n4313), .ZN(n6346) );
  OAI21_X1 U7889 ( .B1(n6348), .B2(n9277), .A(n6346), .ZN(P1_U3343) );
  AOI22_X1 U7890 ( .A1(n6675), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n8690), .ZN(n6347) );
  OAI21_X1 U7891 ( .B1(n6348), .B2(n8695), .A(n6347), .ZN(P2_U3348) );
  INV_X1 U7892 ( .A(n6745), .ZN(n6739) );
  INV_X1 U7893 ( .A(n6349), .ZN(n6351) );
  INV_X1 U7894 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6350) );
  OAI222_X1 U7895 ( .A1(P1_U3084), .A2(n6739), .B1(n9277), .B2(n6351), .C1(
        n6350), .C2(n4314), .ZN(P1_U3342) );
  INV_X1 U7896 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6352) );
  INV_X1 U7897 ( .A(n6859), .ZN(n6682) );
  OAI222_X1 U7898 ( .A1(n8704), .A2(n6352), .B1(n8702), .B2(n6351), .C1(n6682), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U7899 ( .A(n7381), .ZN(n6353) );
  NOR2_X1 U7900 ( .A1(n6354), .A2(n6353), .ZN(n9710) );
  INV_X1 U7901 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6366) );
  NOR2_X1 U7902 ( .A1(n6355), .A2(P1_U3084), .ZN(n9274) );
  AND2_X1 U7903 ( .A1(n6357), .A2(n9274), .ZN(n8887) );
  AND2_X1 U7904 ( .A1(n8887), .A2(n9711), .ZN(n9789) );
  INV_X1 U7905 ( .A(n6361), .ZN(n6392) );
  XNOR2_X1 U7906 ( .A(n6361), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n6359) );
  AND2_X1 U7907 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6358) );
  OR2_X1 U7908 ( .A1(n9711), .A2(P1_U3084), .ZN(n9688) );
  INV_X1 U7909 ( .A(n6355), .ZN(n9689) );
  NOR2_X1 U7910 ( .A1(n9688), .A2(n9689), .ZN(n6356) );
  NAND2_X1 U7911 ( .A1(n6357), .A2(n6356), .ZN(n9736) );
  INV_X1 U7912 ( .A(n9736), .ZN(n9797) );
  NAND2_X1 U7913 ( .A1(n6359), .A2(n6358), .ZN(n6385) );
  OAI211_X1 U7914 ( .C1(n6359), .C2(n6358), .A(n9797), .B(n6385), .ZN(n6360)
         );
  OAI21_X1 U7915 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6693), .A(n6360), .ZN(n6364) );
  NAND2_X1 U7916 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9708) );
  NOR2_X1 U7917 ( .A1(n6362), .A2(n9708), .ZN(n6391) );
  NAND2_X1 U7918 ( .A1(n8887), .A2(n9691), .ZN(n9775) );
  AOI211_X1 U7919 ( .C1(n9708), .C2(n6362), .A(n6391), .B(n9775), .ZN(n6363)
         );
  AOI211_X1 U7920 ( .C1(n9789), .C2(n6392), .A(n6364), .B(n6363), .ZN(n6365)
         );
  OAI21_X1 U7921 ( .B1(n9802), .B2(n6366), .A(n6365), .ZN(P1_U3242) );
  NAND2_X1 U7922 ( .A1(n6316), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6372) );
  INV_X1 U7923 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6367) );
  OR2_X1 U7924 ( .A1(n4316), .A2(n6367), .ZN(n6371) );
  INV_X1 U7925 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n6368) );
  OR2_X1 U7926 ( .A1(n6369), .A2(n6368), .ZN(n6370) );
  AND3_X1 U7927 ( .A1(n6372), .A2(n6371), .A3(n6370), .ZN(n8953) );
  INV_X1 U7928 ( .A(P1_U4006), .ZN(n8826) );
  NAND2_X1 U7929 ( .A1(n8826), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6373) );
  OAI21_X1 U7930 ( .B1(n8953), .B2(n8826), .A(n6373), .ZN(P1_U3585) );
  OAI211_X1 U7931 ( .C1(n8072), .C2(n9658), .A(n6703), .B(n6697), .ZN(n6866)
         );
  INV_X1 U7932 ( .A(n6700), .ZN(n6374) );
  NAND2_X1 U7933 ( .A1(n6374), .A2(n6698), .ZN(n6375) );
  INV_X2 U7934 ( .A(n9877), .ZN(n9879) );
  INV_X1 U7935 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6379) );
  INV_X1 U7936 ( .A(n6930), .ZN(n6666) );
  AND2_X1 U7937 ( .A1(n8827), .A2(n6666), .ZN(n7832) );
  NOR2_X1 U7938 ( .A1(n8827), .A2(n6666), .ZN(n6871) );
  OR2_X1 U7939 ( .A1(n7832), .A2(n6871), .ZN(n8038) );
  AND2_X1 U7940 ( .A1(n8085), .A2(n6927), .ZN(n6377) );
  AND2_X1 U7941 ( .A1(n8825), .A2(n9638), .ZN(n6376) );
  AOI21_X1 U7942 ( .B1(n8038), .B2(n6377), .A(n6376), .ZN(n6933) );
  OAI21_X1 U7943 ( .B1(n6927), .B2(n6666), .A(n6933), .ZN(n9242) );
  NAND2_X1 U7944 ( .A1(n9242), .A2(n9879), .ZN(n6378) );
  OAI21_X1 U7945 ( .B1(n9879), .B2(n6379), .A(n6378), .ZN(P1_U3454) );
  INV_X1 U7946 ( .A(n6380), .ZN(n6423) );
  AOI22_X1 U7947 ( .A1(n6895), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n8690), .ZN(n6381) );
  OAI21_X1 U7948 ( .B1(n6423), .B2(n8695), .A(n6381), .ZN(P2_U3346) );
  INV_X1 U7949 ( .A(n9802), .ZN(n9783) );
  INV_X1 U7950 ( .A(n9789), .ZN(n8873) );
  AND2_X1 U7951 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6619) );
  INV_X1 U7952 ( .A(n6619), .ZN(n6390) );
  OR2_X1 U7953 ( .A1(n6400), .A2(n6382), .ZN(n9724) );
  NAND2_X1 U7954 ( .A1(n6400), .A2(n6382), .ZN(n6383) );
  AND2_X1 U7955 ( .A1(n9724), .A2(n6383), .ZN(n6388) );
  XNOR2_X1 U7956 ( .A(n6393), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9701) );
  NAND2_X1 U7957 ( .A1(n6392), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6384) );
  NAND2_X1 U7958 ( .A1(n6385), .A2(n6384), .ZN(n9700) );
  NAND2_X1 U7959 ( .A1(n9701), .A2(n9700), .ZN(n9699) );
  INV_X1 U7960 ( .A(n6393), .ZN(n9715) );
  NAND2_X1 U7961 ( .A1(n9715), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U7962 ( .A1(n9699), .A2(n6386), .ZN(n6387) );
  AND2_X1 U7963 ( .A1(n6388), .A2(n6387), .ZN(n9727) );
  INV_X1 U7964 ( .A(n9727), .ZN(n6408) );
  OAI211_X1 U7965 ( .C1(n6388), .C2(n6387), .A(n9797), .B(n6408), .ZN(n6389)
         );
  OAI211_X1 U7966 ( .C1(n8873), .C2(n6400), .A(n6390), .B(n6389), .ZN(n6397)
         );
  AOI21_X1 U7967 ( .B1(n6392), .B2(P1_REG2_REG_1__SCAN_IN), .A(n6391), .ZN(
        n9706) );
  XOR2_X1 U7968 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6393), .Z(n9705) );
  NOR2_X1 U7969 ( .A1(n9706), .A2(n9705), .ZN(n9704) );
  AOI21_X1 U7970 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n9715), .A(n9704), .ZN(
        n6395) );
  XOR2_X1 U7971 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6400), .Z(n6394) );
  NOR2_X1 U7972 ( .A1(n6395), .A2(n6394), .ZN(n6401) );
  AOI211_X1 U7973 ( .C1(n6395), .C2(n6394), .A(n6401), .B(n9775), .ZN(n6396)
         );
  AOI211_X1 U7974 ( .C1(P1_ADDR_REG_3__SCAN_IN), .C2(n9783), .A(n6397), .B(
        n6396), .ZN(n6398) );
  INV_X1 U7975 ( .A(n6398), .ZN(P1_U3244) );
  INV_X1 U7976 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6422) );
  INV_X1 U7977 ( .A(n9775), .ZN(n9798) );
  INV_X1 U7978 ( .A(n6410), .ZN(n9749) );
  XNOR2_X1 U7979 ( .A(n9749), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n9754) );
  NOR2_X1 U7980 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9742), .ZN(n6399) );
  AOI21_X1 U7981 ( .B1(n9742), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6399), .ZN(
        n9744) );
  INV_X1 U7982 ( .A(n6406), .ZN(n9722) );
  INV_X1 U7983 ( .A(n6400), .ZN(n6402) );
  AOI21_X1 U7984 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n6402), .A(n6401), .ZN(
        n9720) );
  XNOR2_X1 U7985 ( .A(n6406), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9721) );
  NAND2_X1 U7986 ( .A1(n9720), .A2(n9721), .ZN(n9719) );
  OAI21_X1 U7987 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9722), .A(n9719), .ZN(
        n9745) );
  NAND2_X1 U7988 ( .A1(n9744), .A2(n9745), .ZN(n9743) );
  OAI21_X1 U7989 ( .B1(n9742), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9743), .ZN(
        n9753) );
  AOI22_X1 U7990 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6429), .B1(n6418), .B2(
        n7084), .ZN(n6403) );
  OAI21_X1 U7991 ( .B1(n6404), .B2(n6403), .A(n6425), .ZN(n6420) );
  AOI22_X1 U7992 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6429), .B1(n6418), .B2(
        n5782), .ZN(n6414) );
  XNOR2_X1 U7993 ( .A(n6410), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9751) );
  XNOR2_X1 U7994 ( .A(n6406), .B(n6405), .ZN(n9725) );
  INV_X1 U7995 ( .A(n9725), .ZN(n6407) );
  NAND3_X1 U7996 ( .A1(n6408), .A2(n6407), .A3(n9724), .ZN(n9729) );
  OAI21_X1 U7997 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9722), .A(n9729), .ZN(
        n9739) );
  NAND2_X1 U7998 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9742), .ZN(n6409) );
  OAI21_X1 U7999 ( .B1(n9742), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6409), .ZN(
        n9738) );
  NOR2_X1 U8000 ( .A1(n9739), .A2(n9738), .ZN(n9737) );
  AOI21_X1 U8001 ( .B1(n9742), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9737), .ZN(
        n9750) );
  AOI22_X1 U8002 ( .A1(n9751), .A2(n9750), .B1(n6411), .B2(n6410), .ZN(n6412)
         );
  INV_X1 U8003 ( .A(n6412), .ZN(n6413) );
  NAND2_X1 U8004 ( .A1(n6414), .A2(n6413), .ZN(n6430) );
  OAI21_X1 U8005 ( .B1(n6414), .B2(n6413), .A(n6430), .ZN(n6416) );
  AOI21_X1 U8006 ( .B1(n9797), .B2(n6416), .A(n6415), .ZN(n6417) );
  OAI21_X1 U8007 ( .B1(n8873), .B2(n6418), .A(n6417), .ZN(n6419) );
  AOI21_X1 U8008 ( .B1(n9798), .B2(n6420), .A(n6419), .ZN(n6421) );
  OAI21_X1 U8009 ( .B1(n9802), .B2(n6422), .A(n6421), .ZN(P1_U3248) );
  OAI222_X1 U8010 ( .A1(n4314), .A2(n6424), .B1(n9277), .B2(n6423), .C1(n6832), 
        .C2(P1_U3084), .ZN(P1_U3341) );
  INV_X1 U8011 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6439) );
  MUX2_X1 U8012 ( .A(n6576), .B(P1_REG2_REG_8__SCAN_IN), .S(n6577), .Z(n6426)
         );
  NAND2_X1 U8013 ( .A1(n6426), .A2(n6427), .ZN(n6579) );
  OAI21_X1 U8014 ( .B1(n6427), .B2(n6426), .A(n6579), .ZN(n6437) );
  INV_X1 U8015 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6428) );
  NOR2_X1 U8016 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6428), .ZN(n7195) );
  INV_X1 U8017 ( .A(n7195), .ZN(n6435) );
  INV_X1 U8018 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9884) );
  MUX2_X1 U8019 ( .A(n9884), .B(P1_REG1_REG_8__SCAN_IN), .S(n6577), .Z(n6433)
         );
  OR2_X1 U8020 ( .A1(n6429), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6431) );
  AND2_X1 U8021 ( .A1(n6431), .A2(n6430), .ZN(n6432) );
  NAND2_X1 U8022 ( .A1(n6433), .A2(n6432), .ZN(n6585) );
  OAI211_X1 U8023 ( .C1(n6433), .C2(n6432), .A(n9797), .B(n6585), .ZN(n6434)
         );
  OAI211_X1 U8024 ( .C1(n8873), .C2(n6577), .A(n6435), .B(n6434), .ZN(n6436)
         );
  AOI21_X1 U8025 ( .B1(n9798), .B2(n6437), .A(n6436), .ZN(n6438) );
  OAI21_X1 U8026 ( .B1(n9802), .B2(n6439), .A(n6438), .ZN(P1_U3249) );
  NAND2_X1 U8027 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n8264), .ZN(n6440) );
  OAI21_X1 U8028 ( .B1(n8393), .B2(n8264), .A(n6440), .ZN(P2_U3578) );
  INV_X1 U8029 ( .A(n6441), .ZN(n6574) );
  AOI22_X1 U8030 ( .A1(n7256), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n4313), .ZN(n6442) );
  OAI21_X1 U8031 ( .B1(n6574), .B2(n9277), .A(n6442), .ZN(P1_U3340) );
  NOR2_X1 U8032 ( .A1(n8084), .A2(n6443), .ZN(n9816) );
  OAI21_X1 U8033 ( .B1(n9834), .B2(P1_D_REG_1__SCAN_IN), .A(n6444), .ZN(n6445)
         );
  OAI21_X1 U8034 ( .B1(n6447), .B2(n6446), .A(n6445), .ZN(P1_U3441) );
  NAND2_X1 U8035 ( .A1(n9972), .A2(n6448), .ZN(n6452) );
  OR2_X1 U8036 ( .A1(n5587), .A2(P2_U3152), .ZN(n8697) );
  INV_X1 U8037 ( .A(n7811), .ZN(n7814) );
  OAI21_X1 U8038 ( .B1(n6449), .B2(n8697), .A(n7814), .ZN(n6450) );
  INV_X1 U8039 ( .A(n6450), .ZN(n6451) );
  NAND2_X1 U8040 ( .A1(n6452), .A2(n6451), .ZN(n6468) );
  NAND2_X1 U8041 ( .A1(n6468), .A2(n6466), .ZN(n6453) );
  NAND2_X1 U8042 ( .A1(n6453), .A2(n8264), .ZN(n6489) );
  NAND2_X1 U8043 ( .A1(n6489), .A2(n5587), .ZN(n9927) );
  INV_X1 U8044 ( .A(n9927), .ZN(n8291) );
  INV_X1 U8045 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n6473) );
  INV_X1 U8046 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10071) );
  MUX2_X1 U8047 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10071), .S(n6608), .Z(n6470)
         );
  XNOR2_X1 U8048 ( .A(n6475), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U8049 ( .A1(n6544), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6458) );
  XNOR2_X1 U8050 ( .A(n6477), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n8272) );
  AND2_X1 U8051 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n8271) );
  NAND2_X1 U8052 ( .A1(n8272), .A2(n8271), .ZN(n8270) );
  INV_X1 U8053 ( .A(n6477), .ZN(n8269) );
  NAND2_X1 U8054 ( .A1(n8269), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6454) );
  AND2_X1 U8055 ( .A1(n8270), .A2(n6454), .ZN(n9510) );
  NAND2_X1 U8056 ( .A1(n6480), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6455) );
  OAI21_X1 U8057 ( .B1(n6480), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6455), .ZN(
        n9509) );
  OR2_X1 U8058 ( .A1(n9510), .A2(n9509), .ZN(n9511) );
  AND2_X1 U8059 ( .A1(n9511), .A2(n6455), .ZN(n6534) );
  OR2_X1 U8060 ( .A1(n6544), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6456) );
  NAND2_X1 U8061 ( .A1(n6456), .A2(n6458), .ZN(n6533) );
  NOR2_X1 U8062 ( .A1(n6534), .A2(n6533), .ZN(n6532) );
  INV_X1 U8063 ( .A(n6532), .ZN(n6457) );
  NAND2_X1 U8064 ( .A1(n6458), .A2(n6457), .ZN(n6547) );
  NAND2_X1 U8065 ( .A1(n6546), .A2(n6547), .ZN(n6551) );
  INV_X1 U8066 ( .A(n6475), .ZN(n6560) );
  NAND2_X1 U8067 ( .A1(n6560), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U8068 ( .A1(n6551), .A2(n6459), .ZN(n6520) );
  OR2_X1 U8069 ( .A1(n6530), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6460) );
  NAND2_X1 U8070 ( .A1(n6530), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6461) );
  AND2_X1 U8071 ( .A1(n6460), .A2(n6461), .ZN(n6521) );
  NAND2_X1 U8072 ( .A1(n6520), .A2(n6521), .ZN(n6519) );
  NAND2_X1 U8073 ( .A1(n6519), .A2(n6461), .ZN(n6496) );
  INV_X1 U8074 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6462) );
  XNOR2_X1 U8075 ( .A(n6505), .B(n6462), .ZN(n6497) );
  NAND2_X1 U8076 ( .A1(n6496), .A2(n6497), .ZN(n6495) );
  NAND2_X1 U8077 ( .A1(n6505), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U8078 ( .A1(n6495), .A2(n6463), .ZN(n6508) );
  INV_X1 U8079 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10067) );
  MUX2_X1 U8080 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10067), .S(n6517), .Z(n6509)
         );
  NAND2_X1 U8081 ( .A1(n6508), .A2(n6509), .ZN(n6507) );
  NAND2_X1 U8082 ( .A1(n6517), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U8083 ( .A1(n6507), .A2(n6464), .ZN(n6563) );
  INV_X1 U8084 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10069) );
  MUX2_X1 U8085 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10069), .S(n6572), .Z(n6564)
         );
  NAND2_X1 U8086 ( .A1(n6563), .A2(n6564), .ZN(n6562) );
  NAND2_X1 U8087 ( .A1(n6572), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6465) );
  NAND2_X1 U8088 ( .A1(n6562), .A2(n6465), .ZN(n6469) );
  AND2_X1 U8089 ( .A1(n6466), .A2(n8701), .ZN(n6467) );
  NAND2_X1 U8090 ( .A1(n6469), .A2(n6470), .ZN(n6598) );
  OAI211_X1 U8091 ( .C1(n6470), .C2(n6469), .A(n9924), .B(n6598), .ZN(n6472)
         );
  NAND2_X1 U8092 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n6471) );
  OAI211_X1 U8093 ( .C1(n8325), .C2(n6473), .A(n6472), .B(n6471), .ZN(n6493)
         );
  INV_X1 U8094 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6474) );
  XNOR2_X1 U8095 ( .A(n6475), .B(n6474), .ZN(n6556) );
  NAND2_X1 U8096 ( .A1(n6480), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6476) );
  OAI21_X1 U8097 ( .B1(n6480), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6476), .ZN(
        n9505) );
  INV_X1 U8098 ( .A(n9505), .ZN(n6479) );
  XNOR2_X1 U8099 ( .A(n6477), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n8268) );
  AND2_X1 U8100 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n8267) );
  NAND2_X1 U8101 ( .A1(n8268), .A2(n8267), .ZN(n8266) );
  NAND2_X1 U8102 ( .A1(n8269), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U8103 ( .A1(n8266), .A2(n6478), .ZN(n9504) );
  AND2_X1 U8104 ( .A1(n6479), .A2(n9504), .ZN(n9508) );
  AOI21_X1 U8105 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n6480), .A(n9508), .ZN(
        n6541) );
  NAND2_X1 U8106 ( .A1(n6544), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6481) );
  OAI21_X1 U8107 ( .B1(n6544), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6481), .ZN(
        n6540) );
  NOR2_X1 U8108 ( .A1(n6541), .A2(n6540), .ZN(n6539) );
  NAND2_X1 U8109 ( .A1(n6530), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6482) );
  OAI21_X1 U8110 ( .B1(n6530), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6482), .ZN(
        n6526) );
  AOI21_X1 U8111 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n6530), .A(n6525), .ZN(
        n6502) );
  XNOR2_X1 U8112 ( .A(n6505), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n6501) );
  NOR2_X1 U8113 ( .A1(n6502), .A2(n6501), .ZN(n6500) );
  AOI21_X1 U8114 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n6505), .A(n6500), .ZN(
        n6514) );
  INV_X1 U8115 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6483) );
  MUX2_X1 U8116 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6483), .S(n6517), .Z(n6484)
         );
  INV_X1 U8117 ( .A(n6484), .ZN(n6513) );
  INV_X1 U8118 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6485) );
  MUX2_X1 U8119 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6485), .S(n6572), .Z(n6486)
         );
  INV_X1 U8120 ( .A(n6486), .ZN(n6568) );
  NAND2_X1 U8121 ( .A1(n6608), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6487) );
  OAI21_X1 U8122 ( .B1(n6608), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6487), .ZN(
        n6490) );
  NOR2_X1 U8123 ( .A1(n5587), .A2(n8701), .ZN(n6488) );
  NAND2_X1 U8124 ( .A1(n6489), .A2(n6488), .ZN(n9929) );
  NOR2_X1 U8125 ( .A1(n6491), .A2(n6490), .ZN(n6607) );
  AOI211_X1 U8126 ( .C1(n6491), .C2(n6490), .A(n9929), .B(n6607), .ZN(n6492)
         );
  AOI211_X1 U8127 ( .C1(n8291), .C2(n6608), .A(n6493), .B(n6492), .ZN(n6494)
         );
  INV_X1 U8128 ( .A(n6494), .ZN(P2_U3254) );
  INV_X1 U8129 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10119) );
  OAI211_X1 U8130 ( .C1(n6497), .C2(n6496), .A(n9924), .B(n6495), .ZN(n6499)
         );
  NAND2_X1 U8131 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n6498) );
  OAI211_X1 U8132 ( .C1(n8325), .C2(n10119), .A(n6499), .B(n6498), .ZN(n6504)
         );
  AOI211_X1 U8133 ( .C1(n6502), .C2(n6501), .A(n6500), .B(n9929), .ZN(n6503)
         );
  AOI211_X1 U8134 ( .C1(n8291), .C2(n6505), .A(n6504), .B(n6503), .ZN(n6506)
         );
  INV_X1 U8135 ( .A(n6506), .ZN(P2_U3251) );
  INV_X1 U8136 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10117) );
  OAI211_X1 U8137 ( .C1(n6509), .C2(n6508), .A(n9924), .B(n6507), .ZN(n6511)
         );
  NAND2_X1 U8138 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3152), .ZN(n6510) );
  OAI211_X1 U8139 ( .C1(n8325), .C2(n10117), .A(n6511), .B(n6510), .ZN(n6516)
         );
  AOI211_X1 U8140 ( .C1(n6514), .C2(n6513), .A(n6512), .B(n9929), .ZN(n6515)
         );
  AOI211_X1 U8141 ( .C1(n8291), .C2(n6517), .A(n6516), .B(n6515), .ZN(n6518)
         );
  INV_X1 U8142 ( .A(n6518), .ZN(P2_U3252) );
  INV_X1 U8143 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6524) );
  OAI211_X1 U8144 ( .C1(n6521), .C2(n6520), .A(n9924), .B(n6519), .ZN(n6523)
         );
  NAND2_X1 U8145 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n6522) );
  OAI211_X1 U8146 ( .C1(n8325), .C2(n6524), .A(n6523), .B(n6522), .ZN(n6529)
         );
  AOI211_X1 U8147 ( .C1(n6527), .C2(n6526), .A(n6525), .B(n9929), .ZN(n6528)
         );
  AOI211_X1 U8148 ( .C1(n8291), .C2(n6530), .A(n6529), .B(n6528), .ZN(n6531)
         );
  INV_X1 U8149 ( .A(n6531), .ZN(P2_U3250) );
  INV_X1 U8150 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6538) );
  AOI21_X1 U8151 ( .B1(n6534), .B2(n6533), .A(n6532), .ZN(n6535) );
  NAND2_X1 U8152 ( .A1(n9924), .A2(n6535), .ZN(n6537) );
  NAND2_X1 U8153 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3152), .ZN(n6536) );
  OAI211_X1 U8154 ( .C1(n8325), .C2(n6538), .A(n6537), .B(n6536), .ZN(n6543)
         );
  AOI211_X1 U8155 ( .C1(n6541), .C2(n6540), .A(n6539), .B(n9929), .ZN(n6542)
         );
  AOI211_X1 U8156 ( .C1(n8291), .C2(n6544), .A(n6543), .B(n6542), .ZN(n6545)
         );
  INV_X1 U8157 ( .A(n6545), .ZN(P2_U3248) );
  INV_X1 U8158 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6554) );
  INV_X1 U8159 ( .A(n6546), .ZN(n6549) );
  INV_X1 U8160 ( .A(n6547), .ZN(n6548) );
  NAND2_X1 U8161 ( .A1(n6549), .A2(n6548), .ZN(n6550) );
  NAND3_X1 U8162 ( .A1(n9924), .A2(n6551), .A3(n6550), .ZN(n6553) );
  NAND2_X1 U8163 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n6552) );
  OAI211_X1 U8164 ( .C1(n8325), .C2(n6554), .A(n6553), .B(n6552), .ZN(n6559)
         );
  AOI211_X1 U8165 ( .C1(n6557), .C2(n6556), .A(n6555), .B(n9929), .ZN(n6558)
         );
  AOI211_X1 U8166 ( .C1(n8291), .C2(n6560), .A(n6559), .B(n6558), .ZN(n6561)
         );
  INV_X1 U8167 ( .A(n6561), .ZN(P2_U3249) );
  INV_X1 U8168 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10111) );
  OAI211_X1 U8169 ( .C1(n6564), .C2(n6563), .A(n9924), .B(n6562), .ZN(n6566)
         );
  NAND2_X1 U8170 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n6565) );
  OAI211_X1 U8171 ( .C1(n8325), .C2(n10111), .A(n6566), .B(n6565), .ZN(n6571)
         );
  AOI211_X1 U8172 ( .C1(n6569), .C2(n6568), .A(n9929), .B(n6567), .ZN(n6570)
         );
  AOI211_X1 U8173 ( .C1(n8291), .C2(n6572), .A(n6571), .B(n6570), .ZN(n6573)
         );
  INV_X1 U8174 ( .A(n6573), .ZN(P2_U3253) );
  INV_X1 U8175 ( .A(n7012), .ZN(n6903) );
  OAI222_X1 U8176 ( .A1(n8704), .A2(n6575), .B1(n8702), .B2(n6574), .C1(n6903), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8177 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U8178 ( .A1(n6577), .A2(n6576), .ZN(n6578) );
  NAND2_X1 U8179 ( .A1(n6579), .A2(n6578), .ZN(n9765) );
  NAND2_X1 U8180 ( .A1(n9769), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6580) );
  OAI21_X1 U8181 ( .B1(n9769), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6580), .ZN(
        n9764) );
  NOR2_X1 U8182 ( .A1(n9765), .A2(n9764), .ZN(n9763) );
  XNOR2_X1 U8183 ( .A(n9782), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n9777) );
  NOR2_X1 U8184 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6745), .ZN(n6581) );
  AOI21_X1 U8185 ( .B1(n6745), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6581), .ZN(
        n6582) );
  OAI21_X1 U8186 ( .B1(n6583), .B2(n6582), .A(n6746), .ZN(n6594) );
  AOI22_X1 U8187 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n6745), .B1(n6739), .B2(
        n6738), .ZN(n6590) );
  MUX2_X1 U8188 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6584), .S(n9782), .Z(n9773)
         );
  INV_X1 U8189 ( .A(n6585), .ZN(n6586) );
  AOI21_X1 U8190 ( .B1(n6587), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6586), .ZN(
        n9762) );
  NOR2_X1 U8191 ( .A1(n9769), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6588) );
  AOI21_X1 U8192 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9769), .A(n6588), .ZN(
        n9761) );
  NAND2_X1 U8193 ( .A1(n9762), .A2(n9761), .ZN(n9760) );
  OAI21_X1 U8194 ( .B1(n9769), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9760), .ZN(
        n9774) );
  NAND2_X1 U8195 ( .A1(n9773), .A2(n9774), .ZN(n9772) );
  OAI21_X1 U8196 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n9782), .A(n9772), .ZN(
        n6589) );
  NAND2_X1 U8197 ( .A1(n6590), .A2(n6589), .ZN(n6736) );
  OAI21_X1 U8198 ( .B1(n6590), .B2(n6589), .A(n6736), .ZN(n6591) );
  AND2_X1 U8199 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7336) );
  AOI21_X1 U8200 ( .B1(n9797), .B2(n6591), .A(n7336), .ZN(n6592) );
  OAI21_X1 U8201 ( .B1(n8873), .B2(n6739), .A(n6592), .ZN(n6593) );
  AOI21_X1 U8202 ( .B1(n9798), .B2(n6594), .A(n6593), .ZN(n6595) );
  OAI21_X1 U8203 ( .B1(n9802), .B2(n6596), .A(n6595), .ZN(P1_U3252) );
  INV_X1 U8204 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U8205 ( .A1(n6608), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6597) );
  AND2_X1 U8206 ( .A1(n6598), .A2(n6597), .ZN(n6601) );
  INV_X1 U8207 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6599) );
  MUX2_X1 U8208 ( .A(n6599), .B(P2_REG1_REG_10__SCAN_IN), .S(n6675), .Z(n6600)
         );
  NOR2_X1 U8209 ( .A1(n6601), .A2(n6600), .ZN(n6668) );
  AOI21_X1 U8210 ( .B1(n6601), .B2(n6600), .A(n6668), .ZN(n6602) );
  NAND2_X1 U8211 ( .A1(n9924), .A2(n6602), .ZN(n6605) );
  NOR2_X1 U8212 ( .A1(n6603), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6990) );
  INV_X1 U8213 ( .A(n6990), .ZN(n6604) );
  OAI211_X1 U8214 ( .C1(n8325), .C2(n6606), .A(n6605), .B(n6604), .ZN(n6613)
         );
  NAND2_X1 U8215 ( .A1(n6675), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6609) );
  OAI21_X1 U8216 ( .B1(n6675), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6609), .ZN(
        n6610) );
  AOI211_X1 U8217 ( .C1(n6611), .C2(n6610), .A(n6674), .B(n9929), .ZN(n6612)
         );
  AOI211_X1 U8218 ( .C1(n8291), .C2(n6675), .A(n6613), .B(n6612), .ZN(n6614)
         );
  INV_X1 U8219 ( .A(n6614), .ZN(P2_U3255) );
  XOR2_X1 U8220 ( .A(n6615), .B(n6616), .Z(n6622) );
  INV_X1 U8221 ( .A(n9564), .ZN(n8761) );
  INV_X1 U8222 ( .A(n8823), .ZN(n6617) );
  NOR2_X1 U8223 ( .A1(n8761), .A2(n6617), .ZN(n6618) );
  AOI211_X1 U8224 ( .C1(n8806), .C2(n8821), .A(n6619), .B(n6618), .ZN(n6621)
         );
  INV_X1 U8225 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7028) );
  AOI22_X1 U8226 ( .A1(n7028), .A2(n8798), .B1(n8810), .B2(n7027), .ZN(n6620)
         );
  OAI211_X1 U8227 ( .C1(n6622), .C2(n8812), .A(n6621), .B(n6620), .ZN(P1_U3216) );
  INV_X1 U8228 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6624) );
  INV_X1 U8229 ( .A(n6623), .ZN(n6626) );
  INV_X1 U8230 ( .A(n7291), .ZN(n7010) );
  OAI222_X1 U8231 ( .A1(n8704), .A2(n6624), .B1(n8702), .B2(n6626), .C1(n7010), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8232 ( .A(n8835), .ZN(n8828) );
  INV_X1 U8233 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6625) );
  OAI222_X1 U8234 ( .A1(P1_U3084), .A2(n8828), .B1(n9277), .B2(n6626), .C1(
        n6625), .C2(n4314), .ZN(P1_U3339) );
  NAND3_X1 U8235 ( .A1(n6628), .A2(n8137), .A3(n6759), .ZN(n6630) );
  NOR2_X1 U8236 ( .A1(n6630), .A2(n6629), .ZN(n6644) );
  AND2_X2 U8237 ( .A1(n6644), .A2(n6643), .ZN(n10077) );
  INV_X1 U8238 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6642) );
  NAND2_X1 U8239 ( .A1(n8142), .A2(n8187), .ZN(n7658) );
  NAND2_X1 U8240 ( .A1(n7648), .A2(n7658), .ZN(n6840) );
  NAND2_X1 U8241 ( .A1(n6840), .A2(n6845), .ZN(n6632) );
  NAND2_X1 U8242 ( .A1(n8142), .A2(n9988), .ZN(n6631) );
  NAND2_X1 U8243 ( .A1(n6632), .A2(n6631), .ZN(n6778) );
  NAND2_X1 U8244 ( .A1(n6634), .A2(n6842), .ZN(n7660) );
  NAND2_X1 U8245 ( .A1(n7659), .A2(n7660), .ZN(n6637) );
  NAND2_X1 U8246 ( .A1(n6633), .A2(n6634), .ZN(n6635) );
  INV_X1 U8247 ( .A(n6796), .ZN(n8263) );
  INV_X1 U8248 ( .A(n8183), .ZN(n7112) );
  XNOR2_X1 U8249 ( .A(n6756), .B(n7664), .ZN(n7121) );
  XNOR2_X1 U8250 ( .A(n7815), .B(n6761), .ZN(n6636) );
  NAND2_X1 U8251 ( .A1(n6636), .A2(n8383), .ZN(n7406) );
  NAND3_X1 U8252 ( .A1(n8113), .A2(n9962), .A3(n7802), .ZN(n9551) );
  NAND2_X1 U8253 ( .A1(n7406), .A2(n9551), .ZN(n10054) );
  NAND2_X1 U8254 ( .A1(n6996), .A2(n7658), .ZN(n7642) );
  XNOR2_X1 U8255 ( .A(n6763), .B(n7664), .ZN(n6638) );
  NAND2_X1 U8256 ( .A1(n7627), .A2(n7643), .ZN(n7603) );
  INV_X1 U8257 ( .A(n9939), .ZN(n8483) );
  OAI22_X1 U8258 ( .A1(n6633), .A2(n8537), .B1(n9917), .B2(n8535), .ZN(n8182)
         );
  AOI21_X1 U8259 ( .B1(n6638), .B2(n8483), .A(n8182), .ZN(n7111) );
  OR2_X1 U8260 ( .A1(n8187), .A2(n8139), .ZN(n6846) );
  OR2_X1 U8261 ( .A1(n6781), .A2(n7112), .ZN(n6639) );
  AND2_X1 U8262 ( .A1(n6639), .A2(n6770), .ZN(n7114) );
  INV_X1 U8263 ( .A(n10049), .ZN(n10019) );
  AOI22_X1 U8264 ( .A1(n7114), .A2(n10019), .B1(n10018), .B2(n8183), .ZN(n6640) );
  OAI211_X1 U8265 ( .C1(n7121), .C2(n9983), .A(n7111), .B(n6640), .ZN(n6645)
         );
  NAND2_X1 U8266 ( .A1(n6645), .A2(n10077), .ZN(n6641) );
  OAI21_X1 U8267 ( .B1(n10077), .B2(n6642), .A(n6641), .ZN(P2_U3523) );
  INV_X1 U8268 ( .A(n6643), .ZN(n6758) );
  AND2_X2 U8269 ( .A1(n6644), .A2(n6758), .ZN(n10057) );
  INV_X1 U8270 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U8271 ( .A1(n6645), .A2(n10057), .ZN(n6646) );
  OAI21_X1 U8272 ( .B1(n10057), .B2(n6647), .A(n6646), .ZN(P2_U3460) );
  NAND2_X1 U8273 ( .A1(n6649), .A2(n6648), .ZN(n6653) );
  XNOR2_X1 U8274 ( .A(n6651), .B(n6650), .ZN(n6652) );
  XNOR2_X1 U8275 ( .A(n6653), .B(n6652), .ZN(n6658) );
  AND2_X1 U8276 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9731) );
  INV_X1 U8277 ( .A(n8820), .ZN(n6911) );
  NOR2_X1 U8278 ( .A1(n9568), .A2(n6911), .ZN(n6654) );
  AOI211_X1 U8279 ( .C1(n9564), .C2(n8822), .A(n9731), .B(n6654), .ZN(n6657)
         );
  INV_X1 U8280 ( .A(n6959), .ZN(n6655) );
  INV_X1 U8281 ( .A(n7038), .ZN(n6958) );
  AOI22_X1 U8282 ( .A1(n6655), .A2(n8798), .B1(n8810), .B2(n7038), .ZN(n6656)
         );
  OAI211_X1 U8283 ( .C1(n6658), .C2(n8812), .A(n6657), .B(n6656), .ZN(P1_U3228) );
  INV_X1 U8284 ( .A(n8810), .ZN(n8795) );
  INV_X1 U8285 ( .A(n6659), .ZN(n6660) );
  AOI21_X1 U8286 ( .B1(n6703), .B2(n6660), .A(n8810), .ZN(n6733) );
  NAND2_X1 U8287 ( .A1(n6733), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6665) );
  OAI21_X1 U8288 ( .B1(n6663), .B2(n6662), .A(n6661), .ZN(n9707) );
  AOI22_X1 U8289 ( .A1(n9707), .A2(n9576), .B1(n8806), .B2(n8825), .ZN(n6664)
         );
  OAI211_X1 U8290 ( .C1(n8795), .C2(n6666), .A(n6665), .B(n6664), .ZN(P1_U3230) );
  INV_X1 U8291 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n6667) );
  NOR2_X1 U8292 ( .A1(n8325), .A2(n6667), .ZN(n6673) );
  AOI21_X1 U8293 ( .B1(n6675), .B2(P2_REG1_REG_10__SCAN_IN), .A(n6668), .ZN(
        n6671) );
  INV_X1 U8294 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6669) );
  MUX2_X1 U8295 ( .A(n6669), .B(P2_REG1_REG_11__SCAN_IN), .S(n6859), .Z(n6670)
         );
  NOR2_X1 U8296 ( .A1(n6671), .A2(n6670), .ZN(n6851) );
  INV_X1 U8297 ( .A(n9924), .ZN(n9928) );
  AOI211_X1 U8298 ( .C1(n6671), .C2(n6670), .A(n6851), .B(n9928), .ZN(n6672)
         );
  AOI211_X1 U8299 ( .C1(P2_REG3_REG_11__SCAN_IN), .C2(P2_U3152), .A(n6673), 
        .B(n6672), .ZN(n6681) );
  NOR2_X1 U8300 ( .A1(n6859), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6676) );
  AOI21_X1 U8301 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n6859), .A(n6676), .ZN(
        n6677) );
  OAI21_X1 U8302 ( .B1(n6678), .B2(n6677), .A(n6858), .ZN(n6679) );
  INV_X1 U8303 ( .A(n9929), .ZN(n9925) );
  NAND2_X1 U8304 ( .A1(n6679), .A2(n9925), .ZN(n6680) );
  OAI211_X1 U8305 ( .C1(n9927), .C2(n6682), .A(n6681), .B(n6680), .ZN(P2_U3256) );
  NAND2_X1 U8306 ( .A1(n8826), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6683) );
  OAI21_X1 U8307 ( .B1(n8981), .B2(n8826), .A(n6683), .ZN(P1_U3583) );
  OR2_X1 U8308 ( .A1(n6242), .A2(n8000), .ZN(n6685) );
  OR2_X1 U8309 ( .A1(n6243), .A2(n5656), .ZN(n6684) );
  XNOR2_X1 U8310 ( .A(n8039), .B(n6871), .ZN(n6686) );
  OR2_X1 U8311 ( .A1(n7999), .A2(n9711), .ZN(n9585) );
  AOI222_X1 U8312 ( .A1(n9613), .A2(n6686), .B1(n8827), .B2(n9641), .C1(n8823), 
        .C2(n9638), .ZN(n6710) );
  INV_X1 U8313 ( .A(n6710), .ZN(n6696) );
  OR2_X1 U8314 ( .A1(n4771), .A2(n6688), .ZN(n6690) );
  NAND3_X1 U8315 ( .A1(n6242), .A2(n8072), .A3(n6926), .ZN(n6689) );
  NAND2_X1 U8316 ( .A1(n4771), .A2(n9073), .ZN(n6964) );
  AND2_X1 U8317 ( .A1(n8827), .A2(n6930), .ZN(n6691) );
  OAI21_X1 U8318 ( .B1(n6692), .B2(n6691), .A(n6868), .ZN(n6711) );
  AOI21_X1 U8319 ( .B1(n9864), .B2(n6964), .A(n6711), .ZN(n6695) );
  OAI22_X1 U8320 ( .A1(n9633), .A2(n6693), .B1(n6872), .B2(n6929), .ZN(n6694)
         );
  NOR3_X1 U8321 ( .A1(n6696), .A2(n6695), .A3(n6694), .ZN(n6707) );
  INV_X1 U8322 ( .A(n6697), .ZN(n6699) );
  NAND2_X1 U8323 ( .A1(n6699), .A2(n6698), .ZN(n6701) );
  NOR2_X1 U8324 ( .A1(n6701), .A2(n6700), .ZN(n6702) );
  NAND2_X1 U8325 ( .A1(n6703), .A2(n6702), .ZN(n6704) );
  NOR2_X1 U8326 ( .A1(n6704), .A2(n9073), .ZN(n9147) );
  INV_X1 U8327 ( .A(n9873), .ZN(n9860) );
  NAND2_X1 U8328 ( .A1(n7835), .A2(n6930), .ZN(n6705) );
  AND3_X1 U8329 ( .A1(n9860), .A2(n6878), .A3(n6705), .ZN(n6708) );
  AOI22_X1 U8330 ( .A1(n9147), .A2(n6708), .B1(n9149), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6706) );
  OAI21_X1 U8331 ( .B1(n6707), .B2(n9149), .A(n6706), .ZN(P1_U3290) );
  INV_X1 U8332 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6713) );
  NAND2_X1 U8333 ( .A1(n9864), .A2(n9658), .ZN(n9875) );
  AOI21_X1 U8334 ( .B1(n9563), .B2(n7835), .A(n6708), .ZN(n6709) );
  OAI211_X1 U8335 ( .C1(n9240), .C2(n6711), .A(n6710), .B(n6709), .ZN(n9241)
         );
  NAND2_X1 U8336 ( .A1(n9241), .A2(n9879), .ZN(n6712) );
  OAI21_X1 U8337 ( .B1(n9879), .B2(n6713), .A(n6712), .ZN(P1_U3457) );
  XOR2_X1 U8338 ( .A(n6715), .B(n6714), .Z(n6720) );
  INV_X1 U8339 ( .A(n6716), .ZN(n7831) );
  AOI22_X1 U8340 ( .A1(n8806), .A2(n8822), .B1(n9564), .B2(n8825), .ZN(n6717)
         );
  OAI21_X1 U8341 ( .B1(n7831), .B2(n8795), .A(n6717), .ZN(n6718) );
  AOI21_X1 U8342 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n6733), .A(n6718), .ZN(
        n6719) );
  OAI21_X1 U8343 ( .B1(n6720), .B2(n8812), .A(n6719), .ZN(P1_U3235) );
  INV_X1 U8344 ( .A(n6721), .ZN(n6723) );
  OAI222_X1 U8345 ( .A1(n8849), .A2(P1_U3084), .B1(n9277), .B2(n6723), .C1(
        n6722), .C2(n4314), .ZN(P1_U3338) );
  OAI222_X1 U8346 ( .A1(n8704), .A2(n6724), .B1(n8702), .B2(n6723), .C1(
        P2_U3152), .C2(n7427), .ZN(P2_U3343) );
  INV_X1 U8347 ( .A(n6725), .ZN(n6730) );
  AOI21_X1 U8348 ( .B1(n6727), .B2(n6729), .A(n6726), .ZN(n6728) );
  AOI21_X1 U8349 ( .B1(n6730), .B2(n6729), .A(n6728), .ZN(n6735) );
  AOI22_X1 U8350 ( .A1(n8806), .A2(n8823), .B1(n9564), .B2(n8827), .ZN(n6731)
         );
  OAI21_X1 U8351 ( .B1(n6872), .B2(n8795), .A(n6731), .ZN(n6732) );
  AOI21_X1 U8352 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6733), .A(n6732), .ZN(
        n6734) );
  OAI21_X1 U8353 ( .B1(n6735), .B2(n8812), .A(n6734), .ZN(P1_U3220) );
  INV_X1 U8354 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6754) );
  MUX2_X1 U8355 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6824), .S(n6832), .Z(n6741)
         );
  INV_X1 U8356 ( .A(n6736), .ZN(n6737) );
  AOI21_X1 U8357 ( .B1(n6739), .B2(n6738), .A(n6737), .ZN(n6740) );
  NOR2_X1 U8358 ( .A1(n6740), .A2(n6741), .ZN(n6823) );
  AOI21_X1 U8359 ( .B1(n6741), .B2(n6740), .A(n6823), .ZN(n6744) );
  INV_X1 U8360 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6742) );
  NOR2_X1 U8361 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6742), .ZN(n7390) );
  INV_X1 U8362 ( .A(n7390), .ZN(n6743) );
  OAI21_X1 U8363 ( .B1(n9736), .B2(n6744), .A(n6743), .ZN(n6751) );
  XNOR2_X1 U8364 ( .A(n6832), .B(n6831), .ZN(n6749) );
  OR2_X1 U8365 ( .A1(n6745), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6747) );
  NAND2_X1 U8366 ( .A1(n6747), .A2(n6746), .ZN(n6748) );
  AOI211_X1 U8367 ( .C1(n6749), .C2(n6748), .A(n6833), .B(n9775), .ZN(n6750)
         );
  AOI211_X1 U8368 ( .C1(n9789), .C2(n6752), .A(n6751), .B(n6750), .ZN(n6753)
         );
  OAI21_X1 U8369 ( .B1(n9802), .B2(n6754), .A(n6753), .ZN(P1_U3253) );
  NAND2_X1 U8370 ( .A1(n9917), .A2(n6769), .ZN(n7653) );
  INV_X1 U8371 ( .A(n9917), .ZN(n8262) );
  NAND2_X1 U8372 ( .A1(n8262), .A2(n9999), .ZN(n7124) );
  XNOR2_X1 U8373 ( .A(n6942), .B(n7608), .ZN(n10003) );
  INV_X1 U8374 ( .A(n10003), .ZN(n6777) );
  NAND3_X1 U8375 ( .A1(n6758), .A2(n8137), .A3(n6757), .ZN(n6768) );
  INV_X1 U8376 ( .A(n6759), .ZN(n6760) );
  NAND2_X1 U8377 ( .A1(n9972), .A2(n6760), .ZN(n7464) );
  OR2_X1 U8378 ( .A1(n6761), .A2(n8383), .ZN(n7231) );
  NAND2_X1 U8379 ( .A1(n7406), .A2(n7231), .ZN(n9967) );
  NAND2_X1 U8380 ( .A1(n9968), .A2(n9967), .ZN(n8565) );
  INV_X1 U8381 ( .A(n7608), .ZN(n6764) );
  NAND2_X1 U8382 ( .A1(n6764), .A2(n6765), .ZN(n7125) );
  OAI211_X1 U8383 ( .C1(n6765), .C2(n6764), .A(n8483), .B(n7125), .ZN(n6767)
         );
  AOI22_X1 U8384 ( .A1(n8263), .A2(n8478), .B1(n8480), .B2(n8261), .ZN(n6766)
         );
  NAND2_X1 U8385 ( .A1(n6767), .A2(n6766), .ZN(n10001) );
  NOR2_X1 U8386 ( .A1(n9982), .A2(n7802), .ZN(n9958) );
  NAND2_X1 U8387 ( .A1(n9968), .A2(n9958), .ZN(n8554) );
  INV_X1 U8388 ( .A(n6770), .ZN(n6771) );
  OAI21_X1 U8389 ( .B1(n6771), .B2(n9999), .A(n6945), .ZN(n10000) );
  INV_X1 U8390 ( .A(n6772), .ZN(n6795) );
  OAI22_X1 U8391 ( .A1(n8354), .A2(n10000), .B1(n6795), .B2(n7464), .ZN(n6773)
         );
  AOI21_X1 U8392 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n9944), .A(n6773), .ZN(
        n6774) );
  OAI21_X1 U8393 ( .B1(n9999), .B2(n8554), .A(n6774), .ZN(n6775) );
  AOI21_X1 U8394 ( .B1(n10001), .B2(n9968), .A(n6775), .ZN(n6776) );
  OAI21_X1 U8395 ( .B1(n6777), .B2(n8565), .A(n6776), .ZN(P2_U3292) );
  XNOR2_X1 U8396 ( .A(n6778), .B(n6637), .ZN(n9997) );
  INV_X1 U8397 ( .A(n9997), .ZN(n6788) );
  XOR2_X1 U8398 ( .A(n6637), .B(n6779), .Z(n6780) );
  OAI222_X1 U8399 ( .A1(n8537), .A2(n8142), .B1(n8535), .B2(n6796), .C1(n9939), 
        .C2(n6780), .ZN(n9995) );
  INV_X1 U8400 ( .A(n6846), .ZN(n6783) );
  INV_X1 U8401 ( .A(n6781), .ZN(n6782) );
  OAI21_X1 U8402 ( .B1(n6634), .B2(n6783), .A(n6782), .ZN(n9994) );
  OAI22_X1 U8403 ( .A1(n8354), .A2(n9994), .B1(n5075), .B2(n7464), .ZN(n6784)
         );
  AOI21_X1 U8404 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n9944), .A(n6784), .ZN(
        n6785) );
  OAI21_X1 U8405 ( .B1(n6634), .B2(n8554), .A(n6785), .ZN(n6786) );
  AOI21_X1 U8406 ( .B1(n9995), .B2(n9968), .A(n6786), .ZN(n6787) );
  OAI21_X1 U8407 ( .B1(n6788), .B2(n8565), .A(n6787), .ZN(P2_U3294) );
  INV_X1 U8408 ( .A(n6789), .ZN(n6792) );
  NAND2_X1 U8409 ( .A1(n9893), .A2(n7604), .ZN(n8179) );
  NOR3_X1 U8410 ( .A1(n8179), .A2(n6790), .A3(n6796), .ZN(n6791) );
  AOI21_X1 U8411 ( .B1(n6792), .B2(n9893), .A(n6791), .ZN(n6803) );
  INV_X1 U8412 ( .A(n6793), .ZN(n6802) );
  NOR2_X1 U8413 ( .A1(n6794), .A2(n9909), .ZN(n6800) );
  NOR2_X1 U8414 ( .A1(n9923), .A2(n6795), .ZN(n6799) );
  INV_X1 U8415 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9425) );
  OAI22_X1 U8416 ( .A1(n9913), .A2(n9999), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9425), .ZN(n6798) );
  INV_X1 U8417 ( .A(n8261), .ZN(n6941) );
  OAI22_X1 U8418 ( .A1(n6796), .A2(n9916), .B1(n9915), .B2(n6941), .ZN(n6797)
         );
  NOR4_X1 U8419 ( .A1(n6800), .A2(n6799), .A3(n6798), .A4(n6797), .ZN(n6801)
         );
  OAI21_X1 U8420 ( .B1(n6803), .B2(n6802), .A(n6801), .ZN(P2_U3232) );
  INV_X1 U8421 ( .A(n6804), .ZN(n9908) );
  NOR3_X1 U8422 ( .A1(n8179), .A2(n6805), .A3(n6941), .ZN(n6806) );
  AOI21_X1 U8423 ( .B1(n9908), .B2(n9893), .A(n6806), .ZN(n6818) );
  INV_X1 U8424 ( .A(n6807), .ZN(n6815) );
  INV_X1 U8425 ( .A(n7175), .ZN(n10005) );
  NAND2_X1 U8426 ( .A1(n8261), .A2(n8478), .ZN(n6809) );
  NAND2_X1 U8427 ( .A1(n8259), .A2(n8480), .ZN(n6808) );
  AND2_X1 U8428 ( .A1(n6809), .A2(n6808), .ZN(n7127) );
  INV_X1 U8429 ( .A(n7127), .ZN(n6810) );
  AOI22_X1 U8430 ( .A1(n9892), .A2(n6810), .B1(P2_REG3_REG_6__SCAN_IN), .B2(
        P2_U3152), .ZN(n6813) );
  OR2_X1 U8431 ( .A1(n9923), .A2(n6811), .ZN(n6812) );
  OAI211_X1 U8432 ( .C1(n10005), .C2(n9913), .A(n6813), .B(n6812), .ZN(n6814)
         );
  AOI21_X1 U8433 ( .B1(n6815), .B2(n9893), .A(n6814), .ZN(n6816) );
  OAI21_X1 U8434 ( .B1(n6818), .B2(n6817), .A(n6816), .ZN(P2_U3241) );
  INV_X1 U8435 ( .A(n6819), .ZN(n6822) );
  AOI22_X1 U8436 ( .A1(n8286), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8690), .ZN(n6820) );
  OAI21_X1 U8437 ( .B1(n6822), .B2(n8695), .A(n6820), .ZN(P2_U3342) );
  AOI22_X1 U8438 ( .A1(n8866), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n4313), .ZN(n6821) );
  OAI21_X1 U8439 ( .B1(n6822), .B2(n9277), .A(n6821), .ZN(P1_U3337) );
  INV_X1 U8440 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6839) );
  AOI21_X1 U8441 ( .B1(n6832), .B2(n6824), .A(n6823), .ZN(n6826) );
  MUX2_X1 U8442 ( .A(n5908), .B(P1_REG1_REG_13__SCAN_IN), .S(n7256), .Z(n6825)
         );
  NOR2_X1 U8443 ( .A1(n6826), .A2(n6825), .ZN(n7254) );
  AOI21_X1 U8444 ( .B1(n6826), .B2(n6825), .A(n7254), .ZN(n6827) );
  NAND2_X1 U8445 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7442) );
  OAI21_X1 U8446 ( .B1(n6827), .B2(n9736), .A(n7442), .ZN(n6828) );
  AOI21_X1 U8447 ( .B1(n7256), .B2(n9789), .A(n6828), .ZN(n6838) );
  OR2_X1 U8448 ( .A1(n7256), .A2(n9610), .ZN(n6830) );
  NAND2_X1 U8449 ( .A1(n7256), .A2(n9610), .ZN(n6829) );
  NAND2_X1 U8450 ( .A1(n6830), .A2(n6829), .ZN(n6836) );
  INV_X1 U8451 ( .A(n7252), .ZN(n6834) );
  OAI211_X1 U8452 ( .C1(n6836), .C2(n6835), .A(n9798), .B(n6834), .ZN(n6837)
         );
  OAI211_X1 U8453 ( .C1(n6839), .C2(n9802), .A(n6838), .B(n6837), .ZN(P1_U3254) );
  XNOR2_X1 U8454 ( .A(n6996), .B(n6840), .ZN(n6841) );
  NAND2_X1 U8455 ( .A1(n6841), .A2(n8483), .ZN(n6844) );
  AOI22_X1 U8456 ( .A1(n6842), .A2(n8480), .B1(n8478), .B2(n8265), .ZN(n6843)
         );
  NAND2_X1 U8457 ( .A1(n6844), .A2(n6843), .ZN(n9990) );
  INV_X1 U8458 ( .A(n9990), .ZN(n6850) );
  INV_X1 U8459 ( .A(n8565), .ZN(n8576) );
  XNOR2_X1 U8460 ( .A(n6840), .B(n6845), .ZN(n9992) );
  AOI22_X1 U8461 ( .A1(n8576), .A2(n9992), .B1(n9945), .B2(n8187), .ZN(n6849)
         );
  INV_X1 U8462 ( .A(n8139), .ZN(n9981) );
  OAI21_X1 U8463 ( .B1(n9988), .B2(n9981), .A(n6846), .ZN(n9989) );
  INV_X1 U8464 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9398) );
  OAI22_X1 U8465 ( .A1(n8354), .A2(n9989), .B1(n9398), .B2(n7464), .ZN(n6847)
         );
  AOI21_X1 U8466 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n9944), .A(n6847), .ZN(
        n6848) );
  OAI211_X1 U8467 ( .C1(n9944), .C2(n6850), .A(n6849), .B(n6848), .ZN(P2_U3295) );
  INV_X1 U8468 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6857) );
  AOI21_X1 U8469 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n6859), .A(n6851), .ZN(
        n6854) );
  INV_X1 U8470 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6852) );
  MUX2_X1 U8471 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6852), .S(n6895), .Z(n6853)
         );
  NAND2_X1 U8472 ( .A1(n6853), .A2(n6854), .ZN(n6897) );
  OAI21_X1 U8473 ( .B1(n6854), .B2(n6853), .A(n6897), .ZN(n6855) );
  NAND2_X1 U8474 ( .A1(n9924), .A2(n6855), .ZN(n6856) );
  NAND2_X1 U8475 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9889) );
  OAI211_X1 U8476 ( .C1(n8325), .C2(n6857), .A(n6856), .B(n9889), .ZN(n6863)
         );
  OAI21_X1 U8477 ( .B1(n6859), .B2(P2_REG2_REG_11__SCAN_IN), .A(n6858), .ZN(
        n6861) );
  XNOR2_X1 U8478 ( .A(n6895), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n6860) );
  NOR2_X1 U8479 ( .A1(n6861), .A2(n6860), .ZN(n6888) );
  AOI211_X1 U8480 ( .C1(n6861), .C2(n6860), .A(n9929), .B(n6888), .ZN(n6862)
         );
  AOI211_X1 U8481 ( .C1(n8291), .C2(n6895), .A(n6863), .B(n6862), .ZN(n6864)
         );
  INV_X1 U8482 ( .A(n6864), .ZN(P2_U3257) );
  INV_X2 U8483 ( .A(n9886), .ZN(n9888) );
  INV_X1 U8484 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6881) );
  NAND2_X1 U8485 ( .A1(n8825), .A2(n7835), .ZN(n6867) );
  INV_X1 U8486 ( .A(n6908), .ZN(n6869) );
  AOI21_X1 U8487 ( .B1(n8043), .B2(n6870), .A(n6869), .ZN(n7185) );
  NAND2_X1 U8488 ( .A1(n8039), .A2(n6871), .ZN(n6874) );
  OR2_X1 U8489 ( .A1(n8825), .A2(n6872), .ZN(n6873) );
  NAND2_X1 U8490 ( .A1(n6874), .A2(n6873), .ZN(n6913) );
  XNOR2_X1 U8491 ( .A(n6913), .B(n8043), .ZN(n6877) );
  AOI22_X1 U8492 ( .A1(n9638), .A2(n8822), .B1(n8825), .B2(n9641), .ZN(n6875)
         );
  OAI21_X1 U8493 ( .B1(n7185), .B2(n9864), .A(n6875), .ZN(n6876) );
  AOI21_X1 U8494 ( .B1(n9613), .B2(n6877), .A(n6876), .ZN(n7190) );
  AOI21_X1 U8495 ( .B1(n6716), .B2(n6878), .A(n7024), .ZN(n7188) );
  AOI22_X1 U8496 ( .A1(n7188), .A2(n9860), .B1(n9563), .B2(n6716), .ZN(n6879)
         );
  OAI211_X1 U8497 ( .C1(n7185), .C2(n9658), .A(n7190), .B(n6879), .ZN(n6882)
         );
  NAND2_X1 U8498 ( .A1(n6882), .A2(n9888), .ZN(n6880) );
  OAI21_X1 U8499 ( .B1(n9888), .B2(n6881), .A(n6880), .ZN(P1_U3525) );
  NAND2_X1 U8500 ( .A1(n6882), .A2(n9879), .ZN(n6883) );
  OAI21_X1 U8501 ( .B1(n9879), .B2(n5684), .A(n6883), .ZN(P1_U3460) );
  INV_X1 U8502 ( .A(n6884), .ZN(n6887) );
  AOI22_X1 U8503 ( .A1(n8884), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n4313), .ZN(n6885) );
  OAI21_X1 U8504 ( .B1(n6887), .B2(n9277), .A(n6885), .ZN(P1_U3336) );
  AOI22_X1 U8505 ( .A1(n8300), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n8690), .ZN(n6886) );
  OAI21_X1 U8506 ( .B1(n6887), .B2(n8695), .A(n6886), .ZN(P2_U3341) );
  AOI21_X1 U8507 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n6895), .A(n6888), .ZN(
        n6891) );
  INV_X1 U8508 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6889) );
  AOI22_X1 U8509 ( .A1(n7012), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n6889), .B2(
        n6903), .ZN(n6890) );
  NAND2_X1 U8510 ( .A1(n6891), .A2(n6890), .ZN(n7004) );
  OAI21_X1 U8511 ( .B1(n6891), .B2(n6890), .A(n7004), .ZN(n6905) );
  INV_X1 U8512 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6893) );
  OAI22_X1 U8513 ( .A1(n8325), .A2(n6893), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6892), .ZN(n6894) );
  INV_X1 U8514 ( .A(n6894), .ZN(n6902) );
  INV_X1 U8515 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9556) );
  AOI22_X1 U8516 ( .A1(n7012), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n9556), .B2(
        n6903), .ZN(n6899) );
  OR2_X1 U8517 ( .A1(n6895), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6896) );
  NAND2_X1 U8518 ( .A1(n6897), .A2(n6896), .ZN(n6898) );
  NAND2_X1 U8519 ( .A1(n6899), .A2(n6898), .ZN(n7011) );
  OAI21_X1 U8520 ( .B1(n6899), .B2(n6898), .A(n7011), .ZN(n6900) );
  NAND2_X1 U8521 ( .A1(n9924), .A2(n6900), .ZN(n6901) );
  OAI211_X1 U8522 ( .C1(n9927), .C2(n6903), .A(n6902), .B(n6901), .ZN(n6904)
         );
  AOI21_X1 U8523 ( .B1(n6905), .B2(n9925), .A(n6904), .ZN(n6906) );
  INV_X1 U8524 ( .A(n6906), .ZN(P2_U3258) );
  INV_X1 U8525 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6923) );
  OR2_X1 U8526 ( .A1(n8823), .A2(n6716), .ZN(n6907) );
  OR2_X1 U8527 ( .A1(n8822), .A2(n7027), .ZN(n6909) );
  NAND2_X1 U8528 ( .A1(n7018), .A2(n6909), .ZN(n6910) );
  OR2_X1 U8529 ( .A1(n8821), .A2(n6958), .ZN(n8009) );
  NAND2_X1 U8530 ( .A1(n8821), .A2(n6958), .ZN(n8002) );
  NAND2_X1 U8531 ( .A1(n8009), .A2(n8002), .ZN(n8037) );
  OAI21_X1 U8532 ( .B1(n6910), .B2(n8037), .A(n7040), .ZN(n6965) );
  INV_X1 U8533 ( .A(n6965), .ZN(n6921) );
  INV_X1 U8534 ( .A(n9864), .ZN(n9646) );
  INV_X1 U8535 ( .A(n8822), .ZN(n6912) );
  OAI22_X1 U8536 ( .A1(n6912), .A2(n9585), .B1(n6911), .B2(n9583), .ZN(n6919)
         );
  NAND2_X1 U8537 ( .A1(n6913), .A2(n8043), .ZN(n6915) );
  OR2_X1 U8538 ( .A1(n8823), .A2(n7831), .ZN(n6914) );
  INV_X1 U8539 ( .A(n7019), .ZN(n8044) );
  NAND2_X1 U8540 ( .A1(n8005), .A2(n8044), .ZN(n6916) );
  OR2_X1 U8541 ( .A1(n8822), .A2(n9835), .ZN(n8008) );
  NAND2_X1 U8542 ( .A1(n6916), .A2(n8008), .ZN(n7035) );
  XNOR2_X1 U8543 ( .A(n7035), .B(n8037), .ZN(n6917) );
  NOR2_X1 U8544 ( .A1(n6917), .A2(n9643), .ZN(n6918) );
  AOI211_X1 U8545 ( .C1(n9646), .C2(n6965), .A(n6919), .B(n6918), .ZN(n6968)
         );
  NAND2_X1 U8546 ( .A1(n7024), .A2(n9835), .ZN(n7026) );
  OR2_X1 U8547 ( .A1(n7026), .A2(n7038), .ZN(n7047) );
  INV_X1 U8548 ( .A(n7047), .ZN(n7143) );
  AOI21_X1 U8549 ( .B1(n7038), .B2(n7026), .A(n7143), .ZN(n6963) );
  AOI22_X1 U8550 ( .A1(n6963), .A2(n9860), .B1(n9563), .B2(n7038), .ZN(n6920)
         );
  OAI211_X1 U8551 ( .C1(n6921), .C2(n9658), .A(n6968), .B(n6920), .ZN(n6924)
         );
  NAND2_X1 U8552 ( .A1(n6924), .A2(n9879), .ZN(n6922) );
  OAI21_X1 U8553 ( .B1(n9879), .B2(n6923), .A(n6922), .ZN(P1_U3466) );
  NAND2_X1 U8554 ( .A1(n6924), .A2(n9888), .ZN(n6925) );
  OAI21_X1 U8555 ( .B1(n9888), .B2(n6405), .A(n6925), .ZN(P1_U3527) );
  INV_X1 U8556 ( .A(n6926), .ZN(n8082) );
  OR2_X1 U8557 ( .A1(n6927), .A2(n8082), .ZN(n6928) );
  OR2_X1 U8558 ( .A1(n9149), .A2(n6928), .ZN(n8960) );
  OAI21_X1 U8559 ( .B1(n9631), .B2(n9651), .A(n6930), .ZN(n6932) );
  INV_X1 U8560 ( .A(n9633), .ZN(n9593) );
  AOI22_X1 U8561 ( .A1(n9647), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9593), .ZN(n6931) );
  OAI211_X1 U8562 ( .C1(n9647), .C2(n6933), .A(n6932), .B(n6931), .ZN(P1_U3291) );
  INV_X1 U8563 ( .A(n6976), .ZN(n6974) );
  AOI211_X1 U8564 ( .C1(n6935), .C2(n6934), .A(n9909), .B(n6974), .ZN(n6936)
         );
  INV_X1 U8565 ( .A(n6936), .ZN(n6940) );
  INV_X1 U8566 ( .A(n8260), .ZN(n9914) );
  NOR2_X1 U8567 ( .A1(n9916), .A2(n9914), .ZN(n6938) );
  INV_X1 U8568 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9410) );
  OAI22_X1 U8569 ( .A1(n9915), .A2(n7218), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9410), .ZN(n6937) );
  AOI211_X1 U8570 ( .C1(n8222), .C2(n7170), .A(n6938), .B(n6937), .ZN(n6939)
         );
  OAI211_X1 U8571 ( .C1(n10011), .C2(n9913), .A(n6940), .B(n6939), .ZN(
        P2_U3215) );
  INV_X1 U8572 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6952) );
  NAND2_X1 U8573 ( .A1(n6941), .A2(n9957), .ZN(n7656) );
  NAND2_X1 U8574 ( .A1(n8261), .A2(n9912), .ZN(n7667) );
  NAND2_X1 U8575 ( .A1(n7656), .A2(n7667), .ZN(n7611) );
  NAND2_X1 U8576 ( .A1(n6942), .A2(n7608), .ZN(n6944) );
  NAND2_X1 U8577 ( .A1(n9917), .A2(n9999), .ZN(n6943) );
  NAND2_X1 U8578 ( .A1(n6944), .A2(n6943), .ZN(n7122) );
  XOR2_X1 U8579 ( .A(n7611), .B(n7122), .Z(n9955) );
  NAND2_X1 U8580 ( .A1(n6945), .A2(n9957), .ZN(n6946) );
  NAND2_X1 U8581 ( .A1(n6946), .A2(n10019), .ZN(n6947) );
  NOR2_X1 U8582 ( .A1(n7130), .A2(n6947), .ZN(n9956) );
  NAND2_X1 U8583 ( .A1(n7125), .A2(n7124), .ZN(n6948) );
  XOR2_X1 U8584 ( .A(n7611), .B(n6948), .Z(n6949) );
  OAI222_X1 U8585 ( .A1(n8535), .A2(n9914), .B1(n8537), .B2(n9917), .C1(n9939), 
        .C2(n6949), .ZN(n9964) );
  AOI211_X1 U8586 ( .C1(n10018), .C2(n9957), .A(n9956), .B(n9964), .ZN(n6950)
         );
  OAI21_X1 U8587 ( .B1(n9983), .B2(n9955), .A(n6950), .ZN(n6953) );
  NAND2_X1 U8588 ( .A1(n6953), .A2(n10077), .ZN(n6951) );
  OAI21_X1 U8589 ( .B1(n10077), .B2(n6952), .A(n6951), .ZN(P2_U3525) );
  INV_X1 U8590 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6955) );
  NAND2_X1 U8591 ( .A1(n6953), .A2(n10057), .ZN(n6954) );
  OAI21_X1 U8592 ( .B1(n10057), .B2(n6955), .A(n6954), .ZN(P2_U3466) );
  INV_X1 U8593 ( .A(n6956), .ZN(n7002) );
  AOI22_X1 U8594 ( .A1(n8315), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8690), .ZN(n6957) );
  OAI21_X1 U8595 ( .B1(n7002), .B2(n8695), .A(n6957), .ZN(P2_U3340) );
  NOR2_X1 U8596 ( .A1(n9152), .A2(n6958), .ZN(n6962) );
  OAI22_X1 U8597 ( .A1(n9128), .A2(n6960), .B1(n6959), .B2(n9633), .ZN(n6961)
         );
  AOI211_X1 U8598 ( .C1(n6963), .C2(n9631), .A(n6962), .B(n6961), .ZN(n6967)
         );
  NOR2_X1 U8599 ( .A1(n9647), .A2(n6964), .ZN(n9632) );
  NAND2_X1 U8600 ( .A1(n6965), .A2(n9632), .ZN(n6966) );
  OAI211_X1 U8601 ( .C1(n6968), .C2(n9149), .A(n6967), .B(n6966), .ZN(P1_U3287) );
  OR2_X1 U8602 ( .A1(n7305), .A2(n8535), .ZN(n6970) );
  NAND2_X1 U8603 ( .A1(n8259), .A2(n8478), .ZN(n6969) );
  NAND2_X1 U8604 ( .A1(n6970), .A2(n6969), .ZN(n8571) );
  AOI22_X1 U8605 ( .A1(n9892), .A2(n8571), .B1(P2_REG3_REG_8__SCAN_IN), .B2(
        P2_U3152), .ZN(n6971) );
  OAI21_X1 U8606 ( .B1(n6972), .B2(n9923), .A(n6971), .ZN(n6983) );
  INV_X1 U8607 ( .A(n8179), .ZN(n9897) );
  NAND3_X1 U8608 ( .A1(n9897), .A2(n6973), .A3(n8259), .ZN(n6981) );
  OAI21_X1 U8609 ( .B1(n6974), .B2(n6977), .A(n9893), .ZN(n6980) );
  NAND2_X1 U8610 ( .A1(n6976), .A2(n6975), .ZN(n6978) );
  AND2_X1 U8611 ( .A1(n6978), .A2(n6977), .ZN(n6979) );
  AOI21_X1 U8612 ( .B1(n6981), .B2(n6980), .A(n6979), .ZN(n6982) );
  AOI211_X1 U8613 ( .C1(n9902), .C2(n10017), .A(n6983), .B(n6982), .ZN(n6984)
         );
  INV_X1 U8614 ( .A(n6984), .ZN(P2_U3223) );
  INV_X1 U8615 ( .A(n9946), .ZN(n10034) );
  OAI211_X1 U8616 ( .C1(n6987), .C2(n6985), .A(n7056), .B(n9893), .ZN(n6995)
         );
  INV_X1 U8617 ( .A(n9943), .ZN(n6992) );
  OR2_X1 U8618 ( .A1(n7305), .A2(n8537), .ZN(n6989) );
  OR2_X1 U8619 ( .A1(n7355), .A2(n8535), .ZN(n6988) );
  NAND2_X1 U8620 ( .A1(n6989), .A2(n6988), .ZN(n9941) );
  AOI21_X1 U8621 ( .B1(n9892), .B2(n9941), .A(n6990), .ZN(n6991) );
  OAI21_X1 U8622 ( .B1(n9923), .B2(n6992), .A(n6991), .ZN(n6993) );
  INV_X1 U8623 ( .A(n6993), .ZN(n6994) );
  OAI211_X1 U8624 ( .C1(n10034), .C2(n9913), .A(n6995), .B(n6994), .ZN(
        P2_U3219) );
  NAND2_X1 U8625 ( .A1(n8265), .A2(n9981), .ZN(n7644) );
  NAND2_X1 U8626 ( .A1(n6996), .A2(n7644), .ZN(n7607) );
  INV_X1 U8627 ( .A(n7607), .ZN(n9984) );
  AOI22_X1 U8628 ( .A1(n7607), .A2(n8483), .B1(n8480), .B2(n6997), .ZN(n9980)
         );
  INV_X1 U8629 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9422) );
  OAI22_X1 U8630 ( .A1(n9944), .A2(n9980), .B1(n9422), .B2(n7464), .ZN(n6998)
         );
  AOI21_X1 U8631 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n9944), .A(n6998), .ZN(
        n7000) );
  OAI21_X1 U8632 ( .B1(n9945), .B2(n9951), .A(n8139), .ZN(n6999) );
  OAI211_X1 U8633 ( .C1(n9984), .C2(n8565), .A(n7000), .B(n6999), .ZN(P2_U3296) );
  INV_X1 U8634 ( .A(n9788), .ZN(n8881) );
  INV_X1 U8635 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7001) );
  OAI222_X1 U8636 ( .A1(n8881), .A2(P1_U3084), .B1(n9277), .B2(n7002), .C1(
        n7001), .C2(n4314), .ZN(P1_U3335) );
  NOR2_X1 U8637 ( .A1(n7291), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7003) );
  AOI21_X1 U8638 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7291), .A(n7003), .ZN(
        n7006) );
  OAI21_X1 U8639 ( .B1(n7006), .B2(n7005), .A(n7286), .ZN(n7009) );
  NAND2_X1 U8640 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n9529) );
  NAND2_X1 U8641 ( .A1(n9926), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7007) );
  OAI211_X1 U8642 ( .C1(n9927), .C2(n7010), .A(n9529), .B(n7007), .ZN(n7008)
         );
  AOI21_X1 U8643 ( .B1(n7009), .B2(n9925), .A(n7008), .ZN(n7017) );
  INV_X1 U8644 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9550) );
  AOI22_X1 U8645 ( .A1(n7291), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n9550), .B2(
        n7010), .ZN(n7014) );
  OAI21_X1 U8646 ( .B1(n7012), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7011), .ZN(
        n7013) );
  NAND2_X1 U8647 ( .A1(n7014), .A2(n7013), .ZN(n7290) );
  OAI21_X1 U8648 ( .B1(n7014), .B2(n7013), .A(n7290), .ZN(n7015) );
  NAND2_X1 U8649 ( .A1(n7015), .A2(n9924), .ZN(n7016) );
  NAND2_X1 U8650 ( .A1(n7017), .A2(n7016), .ZN(P2_U3259) );
  XNOR2_X1 U8651 ( .A(n8005), .B(n7019), .ZN(n7023) );
  OAI21_X1 U8652 ( .B1(n7020), .B2(n7019), .A(n7018), .ZN(n9839) );
  NAND2_X1 U8653 ( .A1(n9839), .A2(n9646), .ZN(n7022) );
  AOI22_X1 U8654 ( .A1(n9641), .A2(n8823), .B1(n8821), .B2(n9638), .ZN(n7021)
         );
  OAI211_X1 U8655 ( .C1(n9643), .C2(n7023), .A(n7022), .B(n7021), .ZN(n9837)
         );
  INV_X1 U8656 ( .A(n9837), .ZN(n7033) );
  OR2_X1 U8657 ( .A1(n7024), .A2(n9835), .ZN(n7025) );
  NAND2_X1 U8658 ( .A1(n7026), .A2(n7025), .ZN(n9836) );
  NAND2_X1 U8659 ( .A1(n9651), .A2(n7027), .ZN(n7030) );
  AOI22_X1 U8660 ( .A1(n9647), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9593), .B2(
        n7028), .ZN(n7029) );
  OAI211_X1 U8661 ( .C1(n9836), .C2(n8960), .A(n7030), .B(n7029), .ZN(n7031)
         );
  AOI21_X1 U8662 ( .B1(n9839), .B2(n9632), .A(n7031), .ZN(n7032) );
  OAI21_X1 U8663 ( .B1(n7033), .B2(n9149), .A(n7032), .ZN(P1_U3288) );
  INV_X1 U8664 ( .A(n8009), .ZN(n7034) );
  NAND2_X1 U8665 ( .A1(n7898), .A2(n8002), .ZN(n7892) );
  NAND2_X1 U8666 ( .A1(n8820), .A2(n9842), .ZN(n7897) );
  NAND2_X1 U8667 ( .A1(n7899), .A2(n7897), .ZN(n7144) );
  NOR2_X1 U8668 ( .A1(n7892), .A2(n7144), .ZN(n7146) );
  INV_X1 U8669 ( .A(n7899), .ZN(n7036) );
  NOR2_X1 U8670 ( .A1(n7146), .A2(n7036), .ZN(n7037) );
  NAND2_X1 U8671 ( .A1(n8819), .A2(n9846), .ZN(n7902) );
  INV_X1 U8672 ( .A(n7042), .ZN(n7900) );
  XNOR2_X1 U8673 ( .A(n7037), .B(n7900), .ZN(n7046) );
  OR2_X1 U8674 ( .A1(n8821), .A2(n7038), .ZN(n7039) );
  INV_X1 U8675 ( .A(n7144), .ZN(n8041) );
  NAND2_X1 U8676 ( .A1(n8820), .A2(n8750), .ZN(n7041) );
  NAND2_X1 U8677 ( .A1(n7043), .A2(n7042), .ZN(n7090) );
  OAI21_X1 U8678 ( .B1(n7043), .B2(n7042), .A(n7090), .ZN(n9850) );
  NAND2_X1 U8679 ( .A1(n9850), .A2(n9646), .ZN(n7045) );
  AOI22_X1 U8680 ( .A1(n9641), .A2(n8820), .B1(n8818), .B2(n9638), .ZN(n7044)
         );
  OAI211_X1 U8681 ( .C1(n7046), .C2(n9643), .A(n7045), .B(n7044), .ZN(n9848)
         );
  INV_X1 U8682 ( .A(n9848), .ZN(n7054) );
  NOR2_X1 U8683 ( .A1(n7141), .A2(n9846), .ZN(n7048) );
  OR2_X1 U8684 ( .A1(n7085), .A2(n7048), .ZN(n9847) );
  INV_X1 U8685 ( .A(n7049), .ZN(n8124) );
  AOI22_X1 U8686 ( .A1(n9647), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n8124), .B2(
        n9593), .ZN(n7051) );
  NAND2_X1 U8687 ( .A1(n9651), .A2(n8123), .ZN(n7050) );
  OAI211_X1 U8688 ( .C1(n9847), .C2(n8960), .A(n7051), .B(n7050), .ZN(n7052)
         );
  AOI21_X1 U8689 ( .B1(n9850), .B2(n9632), .A(n7052), .ZN(n7053) );
  OAI21_X1 U8690 ( .B1(n7054), .B2(n9149), .A(n7053), .ZN(P1_U3285) );
  INV_X1 U8691 ( .A(n7347), .ZN(n10042) );
  AOI21_X1 U8692 ( .B1(n7056), .B2(n4743), .A(n9909), .ZN(n7060) );
  NOR3_X1 U8693 ( .A1(n7057), .A2(n7304), .A3(n8179), .ZN(n7059) );
  OAI21_X1 U8694 ( .B1(n7060), .B2(n7059), .A(n7058), .ZN(n7064) );
  NOR2_X1 U8695 ( .A1(n9916), .A2(n7304), .ZN(n7062) );
  OAI22_X1 U8696 ( .A1(n9915), .A2(n7402), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5231), .ZN(n7061) );
  AOI211_X1 U8697 ( .C1(n8222), .C2(n7313), .A(n7062), .B(n7061), .ZN(n7063)
         );
  OAI211_X1 U8698 ( .C1(n10042), .C2(n9913), .A(n7064), .B(n7063), .ZN(
        P2_U3238) );
  INV_X1 U8699 ( .A(n6985), .ZN(n7073) );
  INV_X1 U8700 ( .A(n7065), .ZN(n7067) );
  NAND2_X1 U8701 ( .A1(n7067), .A2(n7066), .ZN(n7071) );
  AND2_X1 U8702 ( .A1(n7069), .A2(n7068), .ZN(n7070) );
  AOI22_X1 U8703 ( .A1(n7073), .A2(n7072), .B1(n7071), .B2(n7070), .ZN(n7079)
         );
  INV_X1 U8704 ( .A(n9916), .ZN(n8228) );
  AOI22_X1 U8705 ( .A1(n8228), .A2(n4814), .B1(P2_REG3_REG_9__SCAN_IN), .B2(
        P2_U3152), .ZN(n7075) );
  NAND2_X1 U8706 ( .A1(n8222), .A2(n7234), .ZN(n7074) );
  OAI211_X1 U8707 ( .C1(n7304), .C2(n9915), .A(n7075), .B(n7074), .ZN(n7077)
         );
  NOR3_X1 U8708 ( .A1(n6985), .A2(n7305), .A3(n8179), .ZN(n7076) );
  AOI211_X1 U8709 ( .C1(n9902), .C2(n10027), .A(n7077), .B(n7076), .ZN(n7078)
         );
  OAI21_X1 U8710 ( .B1(n7079), .B2(n9909), .A(n7078), .ZN(P2_U3233) );
  NAND2_X1 U8711 ( .A1(n8040), .A2(n7899), .ZN(n8010) );
  INV_X1 U8712 ( .A(n8010), .ZN(n7080) );
  NAND2_X1 U8713 ( .A1(n7902), .A2(n7897), .ZN(n7081) );
  NAND2_X1 U8714 ( .A1(n7081), .A2(n8040), .ZN(n7829) );
  INV_X1 U8715 ( .A(n7102), .ZN(n9855) );
  NAND2_X1 U8716 ( .A1(n8818), .A2(n9855), .ZN(n8003) );
  XNOR2_X1 U8717 ( .A(n7837), .B(n7095), .ZN(n7082) );
  AOI222_X1 U8718 ( .A1(n9613), .A2(n7082), .B1(n8817), .B2(n9638), .C1(n8819), 
        .C2(n9641), .ZN(n9853) );
  OAI22_X1 U8719 ( .A1(n9128), .A2(n7084), .B1(n7083), .B2(n9633), .ZN(n7088)
         );
  OAI211_X1 U8720 ( .C1(n7085), .C2(n9855), .A(n9860), .B(n7105), .ZN(n9852)
         );
  INV_X1 U8721 ( .A(n9147), .ZN(n7086) );
  NOR2_X1 U8722 ( .A1(n9852), .A2(n7086), .ZN(n7087) );
  AOI211_X1 U8723 ( .C1(n9651), .C2(n7102), .A(n7088), .B(n7087), .ZN(n7094)
         );
  OR2_X1 U8724 ( .A1(n8819), .A2(n8123), .ZN(n7089) );
  NAND2_X1 U8725 ( .A1(n7090), .A2(n7089), .ZN(n7091) );
  OAI21_X1 U8726 ( .B1(n7091), .B2(n7095), .A(n7104), .ZN(n9857) );
  NAND2_X1 U8727 ( .A1(n5718), .A2(n8085), .ZN(n7092) );
  INV_X1 U8728 ( .A(n9156), .ZN(n7280) );
  NAND2_X1 U8729 ( .A1(n9857), .A2(n7280), .ZN(n7093) );
  OAI211_X1 U8730 ( .C1(n9853), .C2(n9149), .A(n7094), .B(n7093), .ZN(P1_U3284) );
  INV_X1 U8731 ( .A(n7095), .ZN(n7096) );
  NAND2_X1 U8732 ( .A1(n7097), .A2(n7904), .ZN(n7099) );
  INV_X1 U8733 ( .A(n7277), .ZN(n7106) );
  OR2_X1 U8734 ( .A1(n8817), .A2(n7106), .ZN(n7913) );
  NAND2_X1 U8735 ( .A1(n7106), .A2(n8817), .ZN(n7916) );
  INV_X1 U8736 ( .A(n8051), .ZN(n7098) );
  AOI21_X1 U8737 ( .B1(n7099), .B2(n7098), .A(n9643), .ZN(n7101) );
  OR2_X2 U8738 ( .A1(n7099), .A2(n7098), .ZN(n7269) );
  INV_X1 U8739 ( .A(n8816), .ZN(n7326) );
  INV_X1 U8740 ( .A(n8818), .ZN(n8121) );
  OAI22_X1 U8741 ( .A1(n7326), .A2(n9583), .B1(n8121), .B2(n9585), .ZN(n7100)
         );
  AOI21_X1 U8742 ( .B1(n7101), .B2(n7269), .A(n7100), .ZN(n9863) );
  OR2_X1 U8743 ( .A1(n8818), .A2(n7102), .ZN(n7103) );
  XNOR2_X1 U8744 ( .A(n7276), .B(n8051), .ZN(n9865) );
  INV_X1 U8745 ( .A(n9865), .ZN(n9867) );
  NAND2_X1 U8746 ( .A1(n9867), .A2(n7280), .ZN(n7110) );
  AOI21_X1 U8747 ( .B1(n7277), .B2(n7105), .A(n4390), .ZN(n9861) );
  NOR2_X1 U8748 ( .A1(n9152), .A2(n7106), .ZN(n7108) );
  OAI22_X1 U8749 ( .A1(n9128), .A2(n6576), .B1(n7196), .B2(n9633), .ZN(n7107)
         );
  AOI211_X1 U8750 ( .C1(n9861), .C2(n9631), .A(n7108), .B(n7107), .ZN(n7109)
         );
  OAI211_X1 U8751 ( .C1(n9647), .C2(n9863), .A(n7110), .B(n7109), .ZN(P1_U3283) );
  NOR2_X1 U8752 ( .A1(n7111), .A2(n9944), .ZN(n7119) );
  NOR2_X1 U8753 ( .A1(n8554), .A2(n7112), .ZN(n7118) );
  INV_X1 U8754 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7113) );
  NOR2_X1 U8755 ( .A1(n9968), .A2(n7113), .ZN(n7117) );
  INV_X1 U8756 ( .A(n7114), .ZN(n7115) );
  OAI22_X1 U8757 ( .A1(n8354), .A2(n7115), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n7464), .ZN(n7116) );
  NOR4_X1 U8758 ( .A1(n7119), .A2(n7118), .A3(n7117), .A4(n7116), .ZN(n7120)
         );
  OAI21_X1 U8759 ( .B1(n7121), .B2(n8565), .A(n7120), .ZN(P2_U3293) );
  NAND2_X1 U8760 ( .A1(n8261), .A2(n9957), .ZN(n7123) );
  XNOR2_X1 U8761 ( .A(n8260), .B(n7175), .ZN(n7173) );
  XNOR2_X1 U8762 ( .A(n7168), .B(n7173), .ZN(n10009) );
  INV_X1 U8763 ( .A(n10009), .ZN(n7136) );
  AND2_X1 U8764 ( .A1(n7124), .A2(n7667), .ZN(n7669) );
  NAND2_X1 U8765 ( .A1(n7125), .A2(n7669), .ZN(n7126) );
  NAND2_X1 U8766 ( .A1(n7126), .A2(n7656), .ZN(n7174) );
  INV_X1 U8767 ( .A(n7173), .ZN(n7612) );
  XNOR2_X1 U8768 ( .A(n7174), .B(n7612), .ZN(n7128) );
  OAI21_X1 U8769 ( .B1(n7128), .B2(n9939), .A(n7127), .ZN(n10007) );
  INV_X1 U8770 ( .A(n7169), .ZN(n7129) );
  OAI21_X1 U8771 ( .B1(n10005), .B2(n7130), .A(n7129), .ZN(n10006) );
  AOI22_X1 U8772 ( .A1(n9944), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n7131), .B2(
        n9960), .ZN(n7133) );
  NAND2_X1 U8773 ( .A1(n9945), .A2(n7175), .ZN(n7132) );
  OAI211_X1 U8774 ( .C1(n10006), .C2(n8354), .A(n7133), .B(n7132), .ZN(n7134)
         );
  AOI21_X1 U8775 ( .B1(n10007), .B2(n9968), .A(n7134), .ZN(n7135) );
  OAI21_X1 U8776 ( .B1(n7136), .B2(n8565), .A(n7135), .ZN(P2_U3290) );
  INV_X1 U8777 ( .A(n7137), .ZN(n7139) );
  OAI222_X1 U8778 ( .A1(n8000), .A2(P1_U3084), .B1(n9277), .B2(n7139), .C1(
        n7138), .C2(n4314), .ZN(P1_U3334) );
  OAI222_X1 U8779 ( .A1(n8704), .A2(n7140), .B1(n8702), .B2(n7139), .C1(n8383), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  INV_X1 U8780 ( .A(n7141), .ZN(n7142) );
  OAI211_X1 U8781 ( .C1(n9842), .C2(n7143), .A(n7142), .B(n9860), .ZN(n9841)
         );
  NOR2_X1 U8782 ( .A1(n9841), .A2(n9073), .ZN(n7149) );
  AND2_X1 U8783 ( .A1(n7892), .A2(n7144), .ZN(n7145) );
  OAI21_X1 U8784 ( .B1(n7146), .B2(n7145), .A(n9613), .ZN(n7148) );
  AOI22_X1 U8785 ( .A1(n9641), .A2(n8821), .B1(n8819), .B2(n9638), .ZN(n7147)
         );
  NAND2_X1 U8786 ( .A1(n7148), .A2(n7147), .ZN(n9843) );
  AOI211_X1 U8787 ( .C1(n9593), .C2(n8751), .A(n7149), .B(n9843), .ZN(n7155)
         );
  INV_X1 U8788 ( .A(n7150), .ZN(n7151) );
  AOI21_X1 U8789 ( .B1(n8041), .B2(n7152), .A(n7151), .ZN(n9845) );
  OAI22_X1 U8790 ( .A1(n9842), .A2(n9152), .B1(n9128), .B2(n5747), .ZN(n7153)
         );
  AOI21_X1 U8791 ( .B1(n9845), .B2(n7280), .A(n7153), .ZN(n7154) );
  OAI21_X1 U8792 ( .B1(n7155), .B2(n9149), .A(n7154), .ZN(P1_U3286) );
  XNOR2_X1 U8793 ( .A(n7156), .B(n7157), .ZN(n7164) );
  AND2_X1 U8794 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9767) );
  AOI21_X1 U8795 ( .B1(n9564), .B2(n8817), .A(n9767), .ZN(n7162) );
  AND2_X1 U8796 ( .A1(n7319), .A2(n9563), .ZN(n9869) );
  NAND2_X1 U8797 ( .A1(n9869), .A2(n9570), .ZN(n7161) );
  INV_X1 U8798 ( .A(n7271), .ZN(n7158) );
  NAND2_X1 U8799 ( .A1(n8798), .A2(n7158), .ZN(n7160) );
  NAND2_X1 U8800 ( .A1(n8806), .A2(n9640), .ZN(n7159) );
  NAND4_X1 U8801 ( .A1(n7162), .A2(n7161), .A3(n7160), .A4(n7159), .ZN(n7163)
         );
  AOI21_X1 U8802 ( .B1(n7164), .B2(n9576), .A(n7163), .ZN(n7165) );
  INV_X1 U8803 ( .A(n7165), .ZN(P1_U3229) );
  AND2_X1 U8804 ( .A1(n8260), .A2(n7175), .ZN(n7167) );
  NAND2_X1 U8805 ( .A1(n9914), .A2(n10005), .ZN(n7166) );
  NAND2_X1 U8806 ( .A1(n10011), .A2(n8259), .ZN(n7683) );
  INV_X1 U8807 ( .A(n8259), .ZN(n7222) );
  INV_X1 U8808 ( .A(n10011), .ZN(n7171) );
  NAND2_X1 U8809 ( .A1(n7222), .A2(n7171), .ZN(n7682) );
  NAND2_X1 U8810 ( .A1(n7683), .A2(n7682), .ZN(n7680) );
  XNOR2_X1 U8811 ( .A(n7221), .B(n7680), .ZN(n10015) );
  NAND2_X1 U8812 ( .A1(n7169), .A2(n10011), .ZN(n8579) );
  OAI21_X1 U8813 ( .B1(n7169), .B2(n10011), .A(n8579), .ZN(n10012) );
  AOI22_X1 U8814 ( .A1(n9945), .A2(n7171), .B1(n9960), .B2(n7170), .ZN(n7172)
         );
  OAI21_X1 U8815 ( .B1(n10012), .B2(n8354), .A(n7172), .ZN(n7181) );
  NAND2_X1 U8816 ( .A1(n9914), .A2(n7175), .ZN(n7679) );
  INV_X1 U8817 ( .A(n7220), .ZN(n8568) );
  AOI211_X1 U8818 ( .C1(n7680), .C2(n7177), .A(n9939), .B(n8568), .ZN(n7179)
         );
  OAI22_X1 U8819 ( .A1(n9914), .A2(n8537), .B1(n7218), .B2(n8535), .ZN(n7178)
         );
  OR2_X1 U8820 ( .A1(n7179), .A2(n7178), .ZN(n10013) );
  MUX2_X1 U8821 ( .A(n10013), .B(P2_REG2_REG_7__SCAN_IN), .S(n9944), .Z(n7180)
         );
  AOI211_X1 U8822 ( .C1(n8576), .C2(n10015), .A(n7181), .B(n7180), .ZN(n7182)
         );
  INV_X1 U8823 ( .A(n7182), .ZN(P2_U3289) );
  AOI22_X1 U8824 ( .A1(n9647), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9593), .ZN(n7183) );
  OAI21_X1 U8825 ( .B1(n9152), .B2(n7831), .A(n7183), .ZN(n7187) );
  INV_X1 U8826 ( .A(n9632), .ZN(n7184) );
  NOR2_X1 U8827 ( .A1(n7185), .A2(n7184), .ZN(n7186) );
  AOI211_X1 U8828 ( .C1(n7188), .C2(n9631), .A(n7187), .B(n7186), .ZN(n7189)
         );
  OAI21_X1 U8829 ( .B1(n9647), .B2(n7190), .A(n7189), .ZN(P1_U3289) );
  NAND2_X1 U8830 ( .A1(n7192), .A2(n7191), .ZN(n7193) );
  XOR2_X1 U8831 ( .A(n7194), .B(n7193), .Z(n7203) );
  AOI21_X1 U8832 ( .B1(n8806), .B2(n8816), .A(n7195), .ZN(n7201) );
  AND2_X1 U8833 ( .A1(n9563), .A2(n7277), .ZN(n9859) );
  NAND2_X1 U8834 ( .A1(n9570), .A2(n9859), .ZN(n7200) );
  INV_X1 U8835 ( .A(n7196), .ZN(n7197) );
  NAND2_X1 U8836 ( .A1(n8798), .A2(n7197), .ZN(n7199) );
  NAND2_X1 U8837 ( .A1(n9564), .A2(n8818), .ZN(n7198) );
  NAND4_X1 U8838 ( .A1(n7201), .A2(n7200), .A3(n7199), .A4(n7198), .ZN(n7202)
         );
  AOI21_X1 U8839 ( .B1(n7203), .B2(n9576), .A(n7202), .ZN(n7204) );
  INV_X1 U8840 ( .A(n7204), .ZN(P1_U3219) );
  XNOR2_X1 U8841 ( .A(n7206), .B(n7205), .ZN(n7207) );
  XNOR2_X1 U8842 ( .A(n7208), .B(n7207), .ZN(n7216) );
  NOR2_X1 U8843 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7209), .ZN(n9780) );
  AOI21_X1 U8844 ( .B1(n9564), .B2(n8816), .A(n9780), .ZN(n7214) );
  NAND2_X1 U8845 ( .A1(n8810), .A2(n9522), .ZN(n7213) );
  INV_X1 U8846 ( .A(n7210), .ZN(n7328) );
  NAND2_X1 U8847 ( .A1(n8798), .A2(n7328), .ZN(n7212) );
  NAND2_X1 U8848 ( .A1(n8806), .A2(n8815), .ZN(n7211) );
  NAND4_X1 U8849 ( .A1(n7214), .A2(n7213), .A3(n7212), .A4(n7211), .ZN(n7215)
         );
  AOI21_X1 U8850 ( .B1(n7216), .B2(n9576), .A(n7215), .ZN(n7217) );
  INV_X1 U8851 ( .A(n7217), .ZN(P1_U3215) );
  NAND2_X1 U8852 ( .A1(n10017), .A2(n7218), .ZN(n7686) );
  INV_X1 U8853 ( .A(n7683), .ZN(n8567) );
  NOR2_X1 U8854 ( .A1(n8566), .A2(n8567), .ZN(n7219) );
  NAND2_X1 U8855 ( .A1(n8569), .A2(n7686), .ZN(n7301) );
  OR2_X1 U8856 ( .A1(n10027), .A2(n7305), .ZN(n7698) );
  NAND2_X1 U8857 ( .A1(n10027), .A2(n7305), .ZN(n7690) );
  NAND2_X1 U8858 ( .A1(n7698), .A2(n7690), .ZN(n7300) );
  XNOR2_X1 U8859 ( .A(n7301), .B(n7300), .ZN(n7230) );
  NAND2_X1 U8860 ( .A1(n7221), .A2(n7680), .ZN(n7224) );
  NAND2_X1 U8861 ( .A1(n10011), .A2(n7222), .ZN(n7223) );
  NAND2_X1 U8862 ( .A1(n7224), .A2(n7223), .ZN(n8574) );
  INV_X1 U8863 ( .A(n8574), .ZN(n7225) );
  NAND2_X1 U8864 ( .A1(n10017), .A2(n4814), .ZN(n7226) );
  OAI21_X1 U8865 ( .B1(n7227), .B2(n7300), .A(n7306), .ZN(n10032) );
  INV_X1 U8866 ( .A(n7406), .ZN(n9942) );
  NAND2_X1 U8867 ( .A1(n10032), .A2(n9942), .ZN(n7229) );
  INV_X1 U8868 ( .A(n7304), .ZN(n8257) );
  AOI22_X1 U8869 ( .A1(n8478), .A2(n4814), .B1(n8257), .B2(n8480), .ZN(n7228)
         );
  OAI211_X1 U8870 ( .C1(n9939), .C2(n7230), .A(n7229), .B(n7228), .ZN(n10030)
         );
  INV_X1 U8871 ( .A(n10030), .ZN(n7239) );
  INV_X1 U8872 ( .A(n7231), .ZN(n7232) );
  AND2_X1 U8873 ( .A1(n9968), .A2(n7232), .ZN(n9952) );
  AND2_X1 U8874 ( .A1(n8577), .A2(n10027), .ZN(n7233) );
  OR2_X1 U8875 ( .A1(n7233), .A2(n9949), .ZN(n10029) );
  AOI22_X1 U8876 ( .A1(n9944), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7234), .B2(
        n9960), .ZN(n7236) );
  NAND2_X1 U8877 ( .A1(n9945), .A2(n10027), .ZN(n7235) );
  OAI211_X1 U8878 ( .C1(n10029), .C2(n8354), .A(n7236), .B(n7235), .ZN(n7237)
         );
  AOI21_X1 U8879 ( .B1(n10032), .B2(n9952), .A(n7237), .ZN(n7238) );
  OAI21_X1 U8880 ( .B1(n7239), .B2(n9944), .A(n7238), .ZN(P2_U3287) );
  INV_X1 U8881 ( .A(n7240), .ZN(n7241) );
  AOI21_X1 U8882 ( .B1(n9903), .B2(n7241), .A(n9909), .ZN(n7245) );
  NOR3_X1 U8883 ( .A1(n7242), .A2(n7402), .A3(n8179), .ZN(n7244) );
  OAI21_X1 U8884 ( .B1(n7245), .B2(n7244), .A(n7243), .ZN(n7249) );
  NOR2_X1 U8885 ( .A1(n9916), .A2(n7402), .ZN(n7247) );
  OAI22_X1 U8886 ( .A1(n9915), .A2(n8092), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6892), .ZN(n7246) );
  AOI211_X1 U8887 ( .C1(n8222), .C2(n7410), .A(n7247), .B(n7246), .ZN(n7248)
         );
  OAI211_X1 U8888 ( .C1(n4706), .C2(n9913), .A(n7249), .B(n7248), .ZN(P2_U3236) );
  INV_X1 U8889 ( .A(n7250), .ZN(n7299) );
  OAI222_X1 U8890 ( .A1(n8704), .A2(n7251), .B1(P2_U3152), .B2(n7802), .C1(
        n8695), .C2(n7299), .ZN(P2_U3338) );
  XNOR2_X1 U8891 ( .A(n8828), .B(n8829), .ZN(n7253) );
  NOR2_X1 U8892 ( .A1(n7503), .A2(n7253), .ZN(n8830) );
  AOI211_X1 U8893 ( .C1(n7253), .C2(n7503), .A(n8830), .B(n9775), .ZN(n7265)
         );
  INV_X1 U8894 ( .A(n7254), .ZN(n7255) );
  OAI21_X1 U8895 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n7256), .A(n7255), .ZN(
        n7259) );
  MUX2_X1 U8896 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7257), .S(n8835), .Z(n7258)
         );
  NAND2_X1 U8897 ( .A1(n7258), .A2(n7259), .ZN(n8834) );
  OAI21_X1 U8898 ( .B1(n7259), .B2(n7258), .A(n8834), .ZN(n7260) );
  NAND2_X1 U8899 ( .A1(n7260), .A2(n9797), .ZN(n7263) );
  NOR2_X1 U8900 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7261), .ZN(n7544) );
  INV_X1 U8901 ( .A(n7544), .ZN(n7262) );
  OAI211_X1 U8902 ( .C1(n8873), .C2(n8828), .A(n7263), .B(n7262), .ZN(n7264)
         );
  AOI211_X1 U8903 ( .C1(P1_ADDR_REG_14__SCAN_IN), .C2(n9783), .A(n7265), .B(
        n7264), .ZN(n7266) );
  INV_X1 U8904 ( .A(n7266), .ZN(P1_U3255) );
  INV_X1 U8905 ( .A(n7267), .ZN(n7283) );
  OAI222_X1 U8906 ( .A1(P1_U3084), .A2(n6243), .B1(n9277), .B2(n7283), .C1(
        n7268), .C2(n4314), .ZN(P1_U3332) );
  OR2_X1 U8907 ( .A1(n7326), .A2(n7319), .ZN(n7855) );
  NAND2_X1 U8908 ( .A1(n7319), .A2(n7326), .ZN(n7914) );
  AND2_X1 U8909 ( .A1(n7855), .A2(n7914), .ZN(n8050) );
  XOR2_X1 U8910 ( .A(n8050), .B(n7371), .Z(n7270) );
  AOI222_X1 U8911 ( .A1(n9613), .A2(n7270), .B1(n9640), .B2(n9638), .C1(n8817), 
        .C2(n9641), .ZN(n9871) );
  OAI22_X1 U8912 ( .A1(n9128), .A2(n7272), .B1(n7271), .B2(n9633), .ZN(n7275)
         );
  INV_X1 U8913 ( .A(n7319), .ZN(n7273) );
  OAI21_X1 U8914 ( .B1(n4390), .B2(n7273), .A(n7327), .ZN(n9872) );
  NOR2_X1 U8915 ( .A1(n9872), .A2(n8960), .ZN(n7274) );
  AOI211_X1 U8916 ( .C1(n9651), .C2(n7319), .A(n7275), .B(n7274), .ZN(n7282)
         );
  NAND2_X1 U8917 ( .A1(n8817), .A2(n7277), .ZN(n7278) );
  NAND2_X1 U8918 ( .A1(n7279), .A2(n7278), .ZN(n7321) );
  XNOR2_X1 U8919 ( .A(n7321), .B(n8050), .ZN(n9876) );
  NAND2_X1 U8920 ( .A1(n9876), .A2(n7280), .ZN(n7281) );
  OAI211_X1 U8921 ( .C1(n9871), .C2(n9149), .A(n7282), .B(n7281), .ZN(P1_U3282) );
  OAI222_X1 U8922 ( .A1(n8704), .A2(n7285), .B1(P2_U3152), .B2(n7284), .C1(
        n8702), .C2(n7283), .ZN(P2_U3337) );
  INV_X1 U8923 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7287) );
  NAND2_X1 U8924 ( .A1(n7288), .A2(n7287), .ZN(n7428) );
  OAI21_X1 U8925 ( .B1(n7288), .B2(n7287), .A(n7428), .ZN(n7296) );
  NOR2_X1 U8926 ( .A1(n9497), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7477) );
  AOI21_X1 U8927 ( .B1(n9926), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7477), .ZN(
        n7289) );
  OAI21_X1 U8928 ( .B1(n7427), .B2(n9927), .A(n7289), .ZN(n7295) );
  OAI21_X1 U8929 ( .B1(n7291), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7290), .ZN(
        n7417) );
  XNOR2_X1 U8930 ( .A(n7417), .B(n7427), .ZN(n7293) );
  INV_X1 U8931 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7292) );
  NOR2_X1 U8932 ( .A1(n7292), .A2(n7293), .ZN(n7418) );
  AOI211_X1 U8933 ( .C1(n7293), .C2(n7292), .A(n7418), .B(n9928), .ZN(n7294)
         );
  AOI211_X1 U8934 ( .C1(n9925), .C2(n7296), .A(n7295), .B(n7294), .ZN(n7297)
         );
  INV_X1 U8935 ( .A(n7297), .ZN(P2_U3260) );
  OAI222_X1 U8936 ( .A1(P1_U3084), .A2(n5656), .B1(n9277), .B2(n7299), .C1(
        n7298), .C2(n4314), .ZN(P1_U3333) );
  OR2_X1 U8937 ( .A1(n7347), .A2(n7355), .ZN(n7697) );
  NAND2_X1 U8938 ( .A1(n7347), .A2(n7355), .ZN(n7706) );
  NAND2_X1 U8939 ( .A1(n7697), .A2(n7706), .ZN(n7618) );
  INV_X1 U8940 ( .A(n7300), .ZN(n7615) );
  NAND2_X1 U8941 ( .A1(n7301), .A2(n7615), .ZN(n7302) );
  NAND2_X1 U8942 ( .A1(n9946), .A2(n7304), .ZN(n7695) );
  XOR2_X1 U8943 ( .A(n7618), .B(n7352), .Z(n7303) );
  OAI222_X1 U8944 ( .A1(n8535), .A2(n7402), .B1(n8537), .B2(n7304), .C1(n9939), 
        .C2(n7303), .ZN(n10044) );
  INV_X1 U8945 ( .A(n10044), .ZN(n7318) );
  INV_X1 U8946 ( .A(n7305), .ZN(n8258) );
  INV_X1 U8947 ( .A(n9935), .ZN(n7308) );
  INV_X1 U8948 ( .A(n7614), .ZN(n7307) );
  NAND2_X1 U8949 ( .A1(n7308), .A2(n7307), .ZN(n7310) );
  NAND2_X1 U8950 ( .A1(n9946), .A2(n8257), .ZN(n7309) );
  NAND2_X1 U8951 ( .A1(n7310), .A2(n7309), .ZN(n7311) );
  OAI21_X1 U8952 ( .B1(n7311), .B2(n7618), .A(n7350), .ZN(n7312) );
  INV_X1 U8953 ( .A(n7312), .ZN(n10046) );
  XNOR2_X1 U8954 ( .A(n9947), .B(n10042), .ZN(n10043) );
  AOI22_X1 U8955 ( .A1(n9944), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7313), .B2(
        n9960), .ZN(n7315) );
  NAND2_X1 U8956 ( .A1(n7347), .A2(n9945), .ZN(n7314) );
  OAI211_X1 U8957 ( .C1(n10043), .C2(n8354), .A(n7315), .B(n7314), .ZN(n7316)
         );
  AOI21_X1 U8958 ( .B1(n10046), .B2(n8576), .A(n7316), .ZN(n7317) );
  OAI21_X1 U8959 ( .B1(n7318), .B2(n9944), .A(n7317), .ZN(P2_U3285) );
  AND2_X1 U8960 ( .A1(n7319), .A2(n8816), .ZN(n7320) );
  INV_X1 U8961 ( .A(n9640), .ZN(n7322) );
  NAND2_X1 U8962 ( .A1(n9522), .A2(n7322), .ZN(n7918) );
  NAND2_X1 U8963 ( .A1(n7922), .A2(n7918), .ZN(n7365) );
  INV_X1 U8964 ( .A(n7365), .ZN(n8052) );
  XNOR2_X1 U8965 ( .A(n7366), .B(n8052), .ZN(n9524) );
  INV_X1 U8966 ( .A(n8815), .ZN(n7373) );
  INV_X1 U8967 ( .A(n7855), .ZN(n7323) );
  OAI21_X1 U8968 ( .B1(n7371), .B2(n7323), .A(n7914), .ZN(n7324) );
  XNOR2_X1 U8969 ( .A(n7324), .B(n7365), .ZN(n7325) );
  OAI222_X1 U8970 ( .A1(n9585), .A2(n7326), .B1(n9583), .B2(n7373), .C1(n7325), 
        .C2(n9643), .ZN(n9520) );
  INV_X1 U8971 ( .A(n9522), .ZN(n7331) );
  AOI211_X1 U8972 ( .C1(n9522), .C2(n7327), .A(n9873), .B(n9627), .ZN(n9521)
         );
  NAND2_X1 U8973 ( .A1(n9521), .A2(n9147), .ZN(n7330) );
  AOI22_X1 U8974 ( .A1(n9647), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7328), .B2(
        n9593), .ZN(n7329) );
  OAI211_X1 U8975 ( .C1(n7331), .C2(n9152), .A(n7330), .B(n7329), .ZN(n7332)
         );
  AOI21_X1 U8976 ( .B1(n9520), .B2(n9128), .A(n7332), .ZN(n7333) );
  OAI21_X1 U8977 ( .B1(n9524), .B2(n9156), .A(n7333), .ZN(P1_U3281) );
  XOR2_X1 U8978 ( .A(n7335), .B(n7334), .Z(n7343) );
  AOI21_X1 U8979 ( .B1(n8806), .B2(n9639), .A(n7336), .ZN(n7341) );
  NAND2_X1 U8980 ( .A1(n9650), .A2(n8810), .ZN(n7340) );
  INV_X1 U8981 ( .A(n9634), .ZN(n7337) );
  NAND2_X1 U8982 ( .A1(n8798), .A2(n7337), .ZN(n7339) );
  NAND2_X1 U8983 ( .A1(n9564), .A2(n9640), .ZN(n7338) );
  NAND4_X1 U8984 ( .A1(n7341), .A2(n7340), .A3(n7339), .A4(n7338), .ZN(n7342)
         );
  AOI21_X1 U8985 ( .B1(n7343), .B2(n9576), .A(n7342), .ZN(n7344) );
  INV_X1 U8986 ( .A(n7344), .ZN(P1_U3234) );
  INV_X1 U8987 ( .A(n7345), .ZN(n8114) );
  OAI222_X1 U8988 ( .A1(n6242), .A2(P1_U3084), .B1(n9277), .B2(n8114), .C1(
        n7346), .C2(n4314), .ZN(P1_U3331) );
  INV_X1 U8989 ( .A(n7355), .ZN(n9896) );
  NAND2_X1 U8990 ( .A1(n7347), .A2(n9896), .ZN(n7348) );
  AND2_X1 U8991 ( .A1(n7350), .A2(n7348), .ZN(n7351) );
  NAND2_X1 U8992 ( .A1(n9901), .A2(n7402), .ZN(n7709) );
  NAND2_X1 U8993 ( .A1(n7710), .A2(n7709), .ZN(n7694) );
  AND2_X1 U8994 ( .A1(n7694), .A2(n7348), .ZN(n7349) );
  OAI21_X1 U8995 ( .B1(n7351), .B2(n7694), .A(n7397), .ZN(n10053) );
  INV_X1 U8996 ( .A(n10053), .ZN(n7364) );
  INV_X1 U8997 ( .A(n7697), .ZN(n7708) );
  OAI21_X1 U8998 ( .B1(n7352), .B2(n7708), .A(n7706), .ZN(n7354) );
  INV_X1 U8999 ( .A(n7401), .ZN(n7353) );
  AOI211_X1 U9000 ( .C1(n7694), .C2(n7354), .A(n9939), .B(n7353), .ZN(n7358)
         );
  OR2_X1 U9001 ( .A1(n7355), .A2(n8537), .ZN(n7357) );
  OR2_X1 U9002 ( .A1(n7459), .A2(n8535), .ZN(n7356) );
  NAND2_X1 U9003 ( .A1(n7357), .A2(n7356), .ZN(n9891) );
  OR2_X1 U9004 ( .A1(n7358), .A2(n9891), .ZN(n10051) );
  OAI21_X1 U9005 ( .B1(n4391), .B2(n4707), .A(n7408), .ZN(n10050) );
  AOI22_X1 U9006 ( .A1(n9944), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7359), .B2(
        n9960), .ZN(n7361) );
  NAND2_X1 U9007 ( .A1(n9901), .A2(n9945), .ZN(n7360) );
  OAI211_X1 U9008 ( .C1(n10050), .C2(n8354), .A(n7361), .B(n7360), .ZN(n7362)
         );
  AOI21_X1 U9009 ( .B1(n10051), .B2(n9968), .A(n7362), .ZN(n7363) );
  OAI21_X1 U9010 ( .B1(n7364), .B2(n8565), .A(n7363), .ZN(P2_U3284) );
  NAND2_X1 U9011 ( .A1(n7366), .A2(n7365), .ZN(n7368) );
  OR2_X1 U9012 ( .A1(n9522), .A2(n9640), .ZN(n7367) );
  NAND2_X1 U9013 ( .A1(n9650), .A2(n8815), .ZN(n7369) );
  INV_X1 U9014 ( .A(n9639), .ZN(n7370) );
  NAND2_X1 U9015 ( .A1(n9237), .A2(n7370), .ZN(n7919) );
  NAND2_X1 U9016 ( .A1(n7911), .A2(n7919), .ZN(n8054) );
  XNOR2_X1 U9017 ( .A(n7501), .B(n8054), .ZN(n9239) );
  NAND2_X1 U9018 ( .A1(n7922), .A2(n7855), .ZN(n7920) );
  NAND2_X1 U9019 ( .A1(n7918), .A2(n7914), .ZN(n7908) );
  NAND2_X1 U9020 ( .A1(n7908), .A2(n7922), .ZN(n7843) );
  AND2_X1 U9021 ( .A1(n9650), .A2(n7373), .ZN(n7841) );
  OR2_X1 U9022 ( .A1(n9650), .A2(n7373), .ZN(n7851) );
  XOR2_X1 U9023 ( .A(n8054), .B(n7506), .Z(n7372) );
  OAI222_X1 U9024 ( .A1(n9583), .A2(n7509), .B1(n9585), .B2(n7373), .C1(n9643), 
        .C2(n7372), .ZN(n9235) );
  INV_X1 U9025 ( .A(n9237), .ZN(n7378) );
  INV_X1 U9026 ( .A(n9650), .ZN(n9671) );
  NAND2_X1 U9027 ( .A1(n9627), .A2(n9671), .ZN(n9629) );
  INV_X1 U9028 ( .A(n9605), .ZN(n7374) );
  AOI211_X1 U9029 ( .C1(n9237), .C2(n9629), .A(n9873), .B(n7374), .ZN(n9236)
         );
  NAND2_X1 U9030 ( .A1(n9236), .A2(n9147), .ZN(n7377) );
  INV_X1 U9031 ( .A(n7392), .ZN(n7375) );
  AOI22_X1 U9032 ( .A1(n9647), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7375), .B2(
        n9593), .ZN(n7376) );
  OAI211_X1 U9033 ( .C1(n7378), .C2(n9152), .A(n7377), .B(n7376), .ZN(n7379)
         );
  AOI21_X1 U9034 ( .B1(n9235), .B2(n9128), .A(n7379), .ZN(n7380) );
  OAI21_X1 U9035 ( .B1(n9239), .B2(n9156), .A(n7380), .ZN(P1_U3279) );
  NAND2_X1 U9036 ( .A1(n7384), .A2(n9270), .ZN(n7382) );
  NOR2_X1 U9037 ( .A1(n7381), .A2(P1_U3084), .ZN(n8081) );
  INV_X1 U9038 ( .A(n8081), .ZN(n8086) );
  OAI211_X1 U9039 ( .C1(n7383), .C2(n4314), .A(n7382), .B(n8086), .ZN(P1_U3330) );
  NAND2_X1 U9040 ( .A1(n7384), .A2(n8696), .ZN(n7385) );
  OAI211_X1 U9041 ( .C1(n7386), .C2(n8704), .A(n7385), .B(n7814), .ZN(P2_U3335) );
  AOI21_X1 U9042 ( .B1(n7388), .B2(n7387), .A(n4394), .ZN(n7395) );
  NOR2_X1 U9043 ( .A1(n9568), .A2(n7509), .ZN(n7389) );
  AOI211_X1 U9044 ( .C1(n9564), .C2(n8815), .A(n7390), .B(n7389), .ZN(n7391)
         );
  OAI21_X1 U9045 ( .B1(n9580), .B2(n7392), .A(n7391), .ZN(n7393) );
  AOI21_X1 U9046 ( .B1(n8810), .B2(n9237), .A(n7393), .ZN(n7394) );
  OAI21_X1 U9047 ( .B1(n7395), .B2(n8812), .A(n7394), .ZN(P1_U3222) );
  INV_X1 U9048 ( .A(n7402), .ZN(n8256) );
  OR2_X1 U9049 ( .A1(n9901), .A2(n8256), .ZN(n7396) );
  OR2_X1 U9050 ( .A1(n7411), .A2(n7459), .ZN(n7719) );
  NAND2_X1 U9051 ( .A1(n7411), .A2(n7459), .ZN(n7718) );
  NAND2_X1 U9052 ( .A1(n7399), .A2(n7716), .ZN(n7400) );
  NAND2_X1 U9053 ( .A1(n7455), .A2(n7400), .ZN(n7407) );
  OAI21_X1 U9054 ( .B1(n7716), .B2(n4389), .A(n7457), .ZN(n7404) );
  OAI22_X1 U9055 ( .A1(n7402), .A2(n8537), .B1(n8092), .B2(n8535), .ZN(n7403)
         );
  AOI21_X1 U9056 ( .B1(n7404), .B2(n8483), .A(n7403), .ZN(n7405) );
  OAI21_X1 U9057 ( .B1(n7407), .B2(n7406), .A(n7405), .ZN(n9553) );
  INV_X1 U9058 ( .A(n9553), .ZN(n7416) );
  INV_X1 U9059 ( .A(n7407), .ZN(n9555) );
  NAND2_X1 U9060 ( .A1(n7408), .A2(n7411), .ZN(n7409) );
  NAND2_X1 U9061 ( .A1(n8101), .A2(n7409), .ZN(n9552) );
  AOI22_X1 U9062 ( .A1(n9944), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7410), .B2(
        n9960), .ZN(n7413) );
  NAND2_X1 U9063 ( .A1(n7411), .A2(n9945), .ZN(n7412) );
  OAI211_X1 U9064 ( .C1(n9552), .C2(n8354), .A(n7413), .B(n7412), .ZN(n7414)
         );
  AOI21_X1 U9065 ( .B1(n9555), .B2(n9952), .A(n7414), .ZN(n7415) );
  OAI21_X1 U9066 ( .B1(n7416), .B2(n9944), .A(n7415), .ZN(P2_U3283) );
  NOR2_X1 U9067 ( .A1(n7427), .A2(n7417), .ZN(n7419) );
  NOR2_X1 U9068 ( .A1(n7419), .A2(n7418), .ZN(n7421) );
  XOR2_X1 U9069 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8286), .Z(n7420) );
  NAND2_X1 U9070 ( .A1(n7420), .A2(n7421), .ZN(n8277) );
  OAI21_X1 U9071 ( .B1(n7421), .B2(n7420), .A(n8277), .ZN(n7435) );
  INV_X1 U9072 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7425) );
  NAND2_X1 U9073 ( .A1(n8291), .A2(n8286), .ZN(n7424) );
  NOR2_X1 U9074 ( .A1(n7422), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7488) );
  INV_X1 U9075 ( .A(n7488), .ZN(n7423) );
  OAI211_X1 U9076 ( .C1(n8325), .C2(n7425), .A(n7424), .B(n7423), .ZN(n7434)
         );
  NAND2_X1 U9077 ( .A1(n7427), .A2(n7426), .ZN(n7429) );
  NAND2_X1 U9078 ( .A1(n7429), .A2(n7428), .ZN(n7432) );
  NAND2_X1 U9079 ( .A1(n8286), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7430) );
  OAI21_X1 U9080 ( .B1(n8286), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7430), .ZN(
        n7431) );
  AOI211_X1 U9081 ( .C1(n7432), .C2(n7431), .A(n8285), .B(n9929), .ZN(n7433)
         );
  AOI211_X1 U9082 ( .C1(n7435), .C2(n9924), .A(n7434), .B(n7433), .ZN(n7436)
         );
  INV_X1 U9083 ( .A(n7436), .ZN(P2_U3261) );
  INV_X1 U9084 ( .A(n7437), .ZN(n7439) );
  NAND2_X1 U9085 ( .A1(n7439), .A2(n7438), .ZN(n7440) );
  XNOR2_X1 U9086 ( .A(n7441), .B(n7440), .ZN(n7448) );
  INV_X1 U9087 ( .A(n7442), .ZN(n7444) );
  INV_X1 U9088 ( .A(n9616), .ZN(n9586) );
  NOR2_X1 U9089 ( .A1(n9568), .A2(n9586), .ZN(n7443) );
  AOI211_X1 U9090 ( .C1(n9564), .C2(n9639), .A(n7444), .B(n7443), .ZN(n7445)
         );
  OAI21_X1 U9091 ( .B1(n9580), .B2(n9609), .A(n7445), .ZN(n7446) );
  AOI21_X1 U9092 ( .B1(n8810), .B2(n9622), .A(n7446), .ZN(n7447) );
  OAI21_X1 U9093 ( .B1(n7448), .B2(n8812), .A(n7447), .ZN(P1_U3232) );
  INV_X1 U9094 ( .A(n8656), .ZN(n8528) );
  OAI211_X1 U9095 ( .C1(n7450), .C2(n7449), .A(n7514), .B(n9893), .ZN(n7454)
         );
  INV_X1 U9096 ( .A(n9915), .ZN(n8229) );
  INV_X1 U9097 ( .A(n8519), .ZN(n8253) );
  AOI22_X1 U9098 ( .A1(n8229), .A2(n8253), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n7451) );
  OAI21_X1 U9099 ( .B1(n8520), .B2(n9916), .A(n7451), .ZN(n7452) );
  AOI21_X1 U9100 ( .B1(n8525), .B2(n8222), .A(n7452), .ZN(n7453) );
  OAI211_X1 U9101 ( .C1(n8528), .C2(n9913), .A(n7454), .B(n7453), .ZN(P2_U3230) );
  NAND2_X1 U9102 ( .A1(n9536), .A2(n8092), .ZN(n7724) );
  NAND2_X1 U9103 ( .A1(n7455), .A2(n4915), .ZN(n7456) );
  AOI21_X1 U9104 ( .B1(n7721), .B2(n7456), .A(n4320), .ZN(n9544) );
  NAND2_X1 U9105 ( .A1(n7458), .A2(n7721), .ZN(n7556) );
  OAI211_X1 U9106 ( .C1(n7458), .C2(n7721), .A(n7556), .B(n8483), .ZN(n7463)
         );
  OR2_X1 U9107 ( .A1(n7459), .A2(n8537), .ZN(n7461) );
  NAND2_X1 U9108 ( .A1(n8255), .A2(n8480), .ZN(n7460) );
  NAND2_X1 U9109 ( .A1(n7461), .A2(n7460), .ZN(n9531) );
  INV_X1 U9110 ( .A(n9531), .ZN(n7462) );
  NAND2_X1 U9111 ( .A1(n7463), .A2(n7462), .ZN(n9548) );
  XNOR2_X1 U9112 ( .A(n8101), .B(n9536), .ZN(n9546) );
  INV_X1 U9113 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7465) );
  OAI22_X1 U9114 ( .A1(n9968), .A2(n7465), .B1(n9539), .B2(n7464), .ZN(n7466)
         );
  AOI21_X1 U9115 ( .B1(n9536), .B2(n9945), .A(n7466), .ZN(n7467) );
  OAI21_X1 U9116 ( .B1(n9546), .B2(n8354), .A(n7467), .ZN(n7468) );
  AOI21_X1 U9117 ( .B1(n9548), .B2(n9968), .A(n7468), .ZN(n7469) );
  OAI21_X1 U9118 ( .B1(n9544), .B2(n8565), .A(n7469), .ZN(P2_U3282) );
  INV_X1 U9119 ( .A(n8665), .ZN(n8555) );
  NAND2_X1 U9120 ( .A1(n9897), .A2(n8255), .ZN(n7472) );
  NAND2_X1 U9121 ( .A1(n9893), .A2(n7482), .ZN(n7471) );
  XNOR2_X1 U9122 ( .A(n7480), .B(n7470), .ZN(n7483) );
  MUX2_X1 U9123 ( .A(n7472), .B(n7471), .S(n7483), .Z(n7479) );
  OR2_X1 U9124 ( .A1(n8520), .A2(n8535), .ZN(n7474) );
  OR2_X1 U9125 ( .A1(n8092), .A2(n8537), .ZN(n7473) );
  NAND2_X1 U9126 ( .A1(n7474), .A2(n7473), .ZN(n8559) );
  INV_X1 U9127 ( .A(n8552), .ZN(n7475) );
  NOR2_X1 U9128 ( .A1(n9923), .A2(n7475), .ZN(n7476) );
  AOI211_X1 U9129 ( .C1(n9892), .C2(n8559), .A(n7477), .B(n7476), .ZN(n7478)
         );
  OAI211_X1 U9130 ( .C1(n8555), .C2(n9913), .A(n7479), .B(n7478), .ZN(P2_U3243) );
  AOI22_X1 U9131 ( .A1(n7483), .A2(n7482), .B1(n7481), .B2(n7480), .ZN(n7487)
         );
  XOR2_X1 U9132 ( .A(n7485), .B(n7484), .Z(n7486) );
  XNOR2_X1 U9133 ( .A(n7487), .B(n7486), .ZN(n7493) );
  AOI21_X1 U9134 ( .B1(n8228), .B2(n8255), .A(n7488), .ZN(n7490) );
  NAND2_X1 U9135 ( .A1(n8222), .A2(n8543), .ZN(n7489) );
  OAI211_X1 U9136 ( .C1(n8536), .C2(n9915), .A(n7490), .B(n7489), .ZN(n7491)
         );
  AOI21_X1 U9137 ( .B1(n8660), .B2(n9902), .A(n7491), .ZN(n7492) );
  OAI21_X1 U9138 ( .B1(n7493), .B2(n9909), .A(n7492), .ZN(P2_U3228) );
  INV_X1 U9139 ( .A(n7494), .ZN(n7498) );
  OAI222_X1 U9140 ( .A1(P2_U3152), .A2(n7496), .B1(n8702), .B2(n7498), .C1(
        n7495), .C2(n8704), .ZN(P2_U3334) );
  OAI222_X1 U9141 ( .A1(n7499), .A2(P1_U3084), .B1(n9277), .B2(n7498), .C1(
        n7497), .C2(n4314), .ZN(P1_U3329) );
  XNOR2_X1 U9142 ( .A(n9232), .B(n9616), .ZN(n8930) );
  AND2_X1 U9143 ( .A1(n9237), .A2(n9639), .ZN(n7500) );
  INV_X1 U9144 ( .A(n9622), .ZN(n9665) );
  XOR2_X1 U9145 ( .A(n8930), .B(n8905), .Z(n9234) );
  INV_X1 U9146 ( .A(n9606), .ZN(n7502) );
  INV_X1 U9147 ( .A(n9232), .ZN(n8906) );
  AOI211_X1 U9148 ( .C1(n9232), .C2(n7502), .A(n9873), .B(n9599), .ZN(n9231)
         );
  NOR2_X1 U9149 ( .A1(n8906), .A2(n9152), .ZN(n7505) );
  OAI22_X1 U9150 ( .A1(n9128), .A2(n7503), .B1(n7546), .B2(n9633), .ZN(n7504)
         );
  AOI211_X1 U9151 ( .C1(n9231), .C2(n9147), .A(n7505), .B(n7504), .ZN(n7511)
         );
  INV_X1 U9152 ( .A(n8909), .ZN(n9143) );
  INV_X1 U9153 ( .A(n7911), .ZN(n7926) );
  OR2_X1 U9154 ( .A1(n9622), .A2(n7509), .ZN(n7849) );
  NAND2_X1 U9155 ( .A1(n9622), .A2(n7509), .ZN(n7840) );
  INV_X1 U9156 ( .A(n7840), .ZN(n7507) );
  XNOR2_X1 U9157 ( .A(n8931), .B(n8930), .ZN(n7508) );
  OAI222_X1 U9158 ( .A1(n9585), .A2(n7509), .B1(n9583), .B2(n9143), .C1(n9643), 
        .C2(n7508), .ZN(n9230) );
  NAND2_X1 U9159 ( .A1(n9230), .A2(n9128), .ZN(n7510) );
  OAI211_X1 U9160 ( .C1(n9234), .C2(n9156), .A(n7511), .B(n7510), .ZN(P1_U3277) );
  NOR3_X1 U9161 ( .A1(n7512), .A2(n8536), .A3(n8179), .ZN(n7518) );
  AOI21_X1 U9162 ( .B1(n7514), .B2(n7513), .A(n9909), .ZN(n7517) );
  INV_X1 U9163 ( .A(n7515), .ZN(n7516) );
  OAI21_X1 U9164 ( .B1(n7518), .B2(n7517), .A(n7516), .ZN(n7522) );
  INV_X1 U9165 ( .A(n8505), .ZN(n8479) );
  NAND2_X1 U9166 ( .A1(n8229), .A2(n8479), .ZN(n7519) );
  NAND2_X1 U9167 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8302) );
  OAI211_X1 U9168 ( .C1(n8536), .C2(n9916), .A(n7519), .B(n8302), .ZN(n7520)
         );
  AOI21_X1 U9169 ( .B1(n8508), .B2(n8222), .A(n7520), .ZN(n7521) );
  OAI211_X1 U9170 ( .C1(n8511), .C2(n9913), .A(n7522), .B(n7521), .ZN(P2_U3240) );
  INV_X1 U9171 ( .A(n7523), .ZN(n7527) );
  OAI222_X1 U9172 ( .A1(n8704), .A2(n7525), .B1(n8702), .B2(n7527), .C1(
        P2_U3152), .C2(n7524), .ZN(P2_U3333) );
  OAI222_X1 U9173 ( .A1(P1_U3084), .A2(n7528), .B1(n9277), .B2(n7527), .C1(
        n7526), .C2(n4314), .ZN(P1_U3328) );
  INV_X1 U9174 ( .A(n7529), .ZN(n7531) );
  NAND2_X1 U9175 ( .A1(n7531), .A2(n7530), .ZN(n7532) );
  XNOR2_X1 U9176 ( .A(n4398), .B(n7532), .ZN(n7538) );
  NAND2_X1 U9177 ( .A1(n8228), .A2(n8253), .ZN(n7534) );
  NAND2_X1 U9178 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8324) );
  OAI211_X1 U9179 ( .C1(n8493), .C2(n9915), .A(n7534), .B(n8324), .ZN(n7536)
         );
  NOR2_X1 U9180 ( .A1(n4716), .A2(n9913), .ZN(n7535) );
  AOI211_X1 U9181 ( .C1(n8222), .C2(n8495), .A(n7536), .B(n7535), .ZN(n7537)
         );
  OAI21_X1 U9182 ( .B1(n7538), .B2(n9909), .A(n7537), .ZN(P2_U3221) );
  NAND2_X1 U9183 ( .A1(n7540), .A2(n7539), .ZN(n7541) );
  XOR2_X1 U9184 ( .A(n7542), .B(n7541), .Z(n7549) );
  NOR2_X1 U9185 ( .A1(n9568), .A2(n9143), .ZN(n7543) );
  AOI211_X1 U9186 ( .C1(n9564), .C2(n8814), .A(n7544), .B(n7543), .ZN(n7545)
         );
  OAI21_X1 U9187 ( .B1(n9580), .B2(n7546), .A(n7545), .ZN(n7547) );
  AOI21_X1 U9188 ( .B1(n8810), .B2(n9232), .A(n7547), .ZN(n7548) );
  OAI21_X1 U9189 ( .B1(n7549), .B2(n8812), .A(n7548), .ZN(P1_U3213) );
  INV_X1 U9190 ( .A(n7550), .ZN(n7554) );
  OAI222_X1 U9191 ( .A1(P2_U3152), .A2(n7552), .B1(n8702), .B2(n7554), .C1(
        n7551), .C2(n8704), .ZN(P2_U3332) );
  OAI222_X1 U9192 ( .A1(n7555), .A2(P1_U3084), .B1(n9277), .B2(n7554), .C1(
        n7553), .C2(n4314), .ZN(P1_U3327) );
  INV_X1 U9193 ( .A(n8255), .ZN(n8538) );
  INV_X1 U9194 ( .A(n7731), .ZN(n7558) );
  NAND2_X1 U9195 ( .A1(n8660), .A2(n8520), .ZN(n7732) );
  NAND2_X1 U9196 ( .A1(n8656), .A2(n8536), .ZN(n7639) );
  NAND2_X1 U9197 ( .A1(n7641), .A2(n7639), .ZN(n8516) );
  OR2_X1 U9198 ( .A1(n8649), .A2(n8519), .ZN(n7738) );
  NAND2_X1 U9199 ( .A1(n8649), .A2(n8519), .ZN(n7740) );
  NAND2_X1 U9200 ( .A1(n7738), .A2(n7740), .ZN(n8502) );
  INV_X1 U9201 ( .A(n7740), .ZN(n7559) );
  OR2_X1 U9202 ( .A1(n8645), .A2(n8505), .ZN(n7739) );
  NAND2_X1 U9203 ( .A1(n8645), .A2(n8505), .ZN(n7741) );
  INV_X1 U9204 ( .A(n7741), .ZN(n8475) );
  NAND2_X1 U9205 ( .A1(n8638), .A2(n8493), .ZN(n7750) );
  INV_X1 U9206 ( .A(n7742), .ZN(n7751) );
  OR2_X1 U9207 ( .A1(n8093), .A2(n8447), .ZN(n7759) );
  NAND2_X1 U9208 ( .A1(n8093), .A2(n8447), .ZN(n8444) );
  NAND2_X1 U9209 ( .A1(n8629), .A2(n8196), .ZN(n7745) );
  NAND2_X1 U9210 ( .A1(n7754), .A2(n7745), .ZN(n8098) );
  NAND2_X1 U9211 ( .A1(n8462), .A2(n4916), .ZN(n8442) );
  NAND2_X1 U9212 ( .A1(n8442), .A2(n7754), .ZN(n8422) );
  AND2_X1 U9213 ( .A1(n8622), .A2(n8448), .ZN(n8414) );
  NAND2_X1 U9214 ( .A1(n8617), .A2(n8392), .ZN(n7765) );
  NAND2_X1 U9215 ( .A1(n8614), .A2(n8415), .ZN(n7635) );
  NAND2_X1 U9216 ( .A1(n8608), .A2(n8393), .ZN(n7771) );
  NAND2_X1 U9217 ( .A1(n8602), .A2(n8242), .ZN(n7629) );
  INV_X1 U9218 ( .A(n7633), .ZN(n7560) );
  NAND2_X1 U9219 ( .A1(n8597), .A2(n8368), .ZN(n7630) );
  NAND2_X1 U9220 ( .A1(n7775), .A2(n7630), .ZN(n8340) );
  INV_X1 U9221 ( .A(n7563), .ZN(n7564) );
  NAND2_X1 U9222 ( .A1(n7564), .A2(n9441), .ZN(n7565) );
  MUX2_X1 U9223 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n7589), .Z(n7572) );
  INV_X1 U9224 ( .A(SI_29_), .ZN(n9362) );
  XNOR2_X1 U9225 ( .A(n7572), .B(n9362), .ZN(n7570) );
  NAND2_X1 U9226 ( .A1(n8692), .A2(n5484), .ZN(n7568) );
  INV_X1 U9227 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8693) );
  OR2_X1 U9228 ( .A1(n7594), .A2(n8693), .ZN(n7567) );
  NAND2_X1 U9229 ( .A1(n8327), .A2(n8109), .ZN(n7782) );
  NAND2_X1 U9230 ( .A1(n7569), .A2(n7780), .ZN(n7599) );
  INV_X1 U9231 ( .A(n7572), .ZN(n7573) );
  INV_X1 U9232 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8153) );
  INV_X1 U9233 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8155) );
  MUX2_X1 U9234 ( .A(n8153), .B(n8155), .S(n7589), .Z(n7575) );
  INV_X1 U9235 ( .A(SI_30_), .ZN(n7574) );
  NAND2_X1 U9236 ( .A1(n7575), .A2(n7574), .ZN(n7587) );
  INV_X1 U9237 ( .A(n7575), .ZN(n7576) );
  NAND2_X1 U9238 ( .A1(n7576), .A2(SI_30_), .ZN(n7577) );
  AND2_X1 U9239 ( .A1(n7587), .A2(n7577), .ZN(n7585) );
  NAND2_X1 U9240 ( .A1(n8152), .A2(n5484), .ZN(n7579) );
  OR2_X1 U9241 ( .A1(n7594), .A2(n8153), .ZN(n7578) );
  INV_X1 U9242 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n7583) );
  NAND2_X1 U9243 ( .A1(n4315), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7582) );
  NAND2_X1 U9244 ( .A1(n7580), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7581) );
  OAI211_X1 U9245 ( .C1(n7584), .C2(n7583), .A(n7582), .B(n7581), .ZN(n8347)
         );
  INV_X1 U9246 ( .A(n8347), .ZN(n7597) );
  NOR2_X1 U9247 ( .A1(n8587), .A2(n7597), .ZN(n7606) );
  MUX2_X1 U9248 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7589), .Z(n7591) );
  INV_X1 U9249 ( .A(SI_31_), .ZN(n7590) );
  XNOR2_X1 U9250 ( .A(n7591), .B(n7590), .ZN(n7592) );
  NAND2_X1 U9251 ( .A1(n8687), .A2(n5484), .ZN(n7596) );
  OR2_X1 U9252 ( .A1(n7594), .A2(n6321), .ZN(n7595) );
  NAND2_X1 U9253 ( .A1(n8587), .A2(n7597), .ZN(n7787) );
  OAI21_X1 U9254 ( .B1(n7599), .B2(n7606), .A(n7792), .ZN(n7601) );
  INV_X1 U9255 ( .A(n8587), .ZN(n8339) );
  NAND2_X1 U9256 ( .A1(n8331), .A2(n7643), .ZN(n7598) );
  AOI21_X1 U9257 ( .B1(n7599), .B2(n8339), .A(n7598), .ZN(n7600) );
  OAI21_X1 U9258 ( .B1(n7601), .B2(n7600), .A(n7799), .ZN(n7602) );
  XNOR2_X1 U9259 ( .A(n7602), .B(n9962), .ZN(n7605) );
  INV_X1 U9260 ( .A(n7792), .ZN(n7625) );
  INV_X1 U9261 ( .A(n7606), .ZN(n7788) );
  NOR3_X1 U9262 ( .A1(n6637), .A2(n7608), .A3(n7607), .ZN(n7610) );
  INV_X1 U9263 ( .A(n6840), .ZN(n7609) );
  NAND4_X1 U9264 ( .A1(n7610), .A2(n7627), .A3(n7664), .A4(n7609), .ZN(n7613)
         );
  NOR4_X1 U9265 ( .A1(n7613), .A2(n7612), .A3(n7680), .A4(n7611), .ZN(n7616)
         );
  NAND4_X1 U9266 ( .A1(n7616), .A2(n8575), .A3(n7615), .A4(n7614), .ZN(n7617)
         );
  NOR4_X1 U9267 ( .A1(n7398), .A2(n7694), .A3(n7618), .A4(n7617), .ZN(n7619)
         );
  NAND4_X1 U9268 ( .A1(n8532), .A2(n7721), .A3(n7619), .A4(n8557), .ZN(n7620)
         );
  NOR4_X1 U9269 ( .A1(n8490), .A2(n8516), .A3(n8502), .A4(n7620), .ZN(n7621)
         );
  NAND4_X1 U9270 ( .A1(n8443), .A2(n4564), .A3(n8463), .A4(n7621), .ZN(n7622)
         );
  NOR4_X1 U9271 ( .A1(n8389), .A2(n8413), .A3(n8432), .A4(n7622), .ZN(n7623)
         );
  NAND4_X1 U9272 ( .A1(n8107), .A2(n8100), .A3(n7623), .A4(n4581), .ZN(n7624)
         );
  XNOR2_X1 U9273 ( .A(n7626), .B(n9962), .ZN(n7628) );
  OAI22_X1 U9274 ( .A1(n7628), .A2(n7643), .B1(n7627), .B2(n7806), .ZN(n7804)
         );
  AND2_X1 U9275 ( .A1(n7630), .A2(n7629), .ZN(n7632) );
  NAND2_X1 U9276 ( .A1(n7643), .A2(n9962), .ZN(n7631) );
  MUX2_X1 U9277 ( .A(n7633), .B(n7632), .S(n7797), .Z(n7777) );
  OR2_X1 U9278 ( .A1(n8608), .A2(n8393), .ZN(n7770) );
  NAND2_X1 U9279 ( .A1(n7770), .A2(n7634), .ZN(n7637) );
  INV_X1 U9280 ( .A(n7635), .ZN(n7636) );
  OAI21_X1 U9281 ( .B1(n8448), .B2(n8622), .A(n8405), .ZN(n7638) );
  NAND2_X1 U9282 ( .A1(n7638), .A2(n7791), .ZN(n7763) );
  INV_X1 U9283 ( .A(n8432), .ZN(n8425) );
  MUX2_X1 U9284 ( .A(n7745), .B(n7754), .S(n7797), .Z(n7762) );
  AND2_X1 U9285 ( .A1(n7740), .A2(n7639), .ZN(n7640) );
  MUX2_X1 U9286 ( .A(n7641), .B(n7640), .S(n7791), .Z(n7737) );
  AND2_X1 U9287 ( .A1(n7648), .A2(n7644), .ZN(n7647) );
  AND2_X1 U9288 ( .A1(n7644), .A2(n7643), .ZN(n7645) );
  NOR2_X1 U9289 ( .A1(n7642), .A2(n7645), .ZN(n7646) );
  MUX2_X1 U9290 ( .A(n7647), .B(n7646), .S(n7797), .Z(n7662) );
  NAND2_X1 U9291 ( .A1(n7648), .A2(n7660), .ZN(n7649) );
  OAI211_X1 U9292 ( .C1(n7662), .C2(n7649), .A(n7797), .B(n7659), .ZN(n7652)
         );
  NAND2_X1 U9293 ( .A1(n7653), .A2(n7650), .ZN(n7651) );
  AOI21_X1 U9294 ( .B1(n7652), .B2(n7664), .A(n7651), .ZN(n7657) );
  INV_X1 U9295 ( .A(n7669), .ZN(n7655) );
  NAND2_X1 U9296 ( .A1(n7656), .A2(n7653), .ZN(n7654) );
  MUX2_X1 U9297 ( .A(n7655), .B(n7654), .S(n7791), .Z(n7663) );
  OAI211_X1 U9298 ( .C1(n7657), .C2(n7663), .A(n7656), .B(n7679), .ZN(n7678)
         );
  NAND2_X1 U9299 ( .A1(n7659), .A2(n7658), .ZN(n7661) );
  OAI21_X1 U9300 ( .B1(n7662), .B2(n7661), .A(n7660), .ZN(n7665) );
  INV_X1 U9301 ( .A(n7663), .ZN(n7672) );
  NAND3_X1 U9302 ( .A1(n7665), .A2(n7664), .A3(n7672), .ZN(n7666) );
  AND2_X1 U9303 ( .A1(n10005), .A2(n8260), .ZN(n7673) );
  AOI21_X1 U9304 ( .B1(n7666), .B2(n7791), .A(n7673), .ZN(n7677) );
  INV_X1 U9305 ( .A(n7667), .ZN(n7671) );
  NAND2_X1 U9306 ( .A1(n7669), .A2(n7668), .ZN(n7670) );
  INV_X1 U9307 ( .A(n7673), .ZN(n7674) );
  AOI21_X1 U9308 ( .B1(n7675), .B2(n7674), .A(n7797), .ZN(n7676) );
  NOR2_X1 U9309 ( .A1(n7679), .A2(n7797), .ZN(n7681) );
  MUX2_X1 U9310 ( .A(n7683), .B(n7682), .S(n7797), .Z(n7684) );
  NAND3_X1 U9311 ( .A1(n7685), .A2(n8575), .A3(n7684), .ZN(n7689) );
  MUX2_X1 U9312 ( .A(n7687), .B(n7686), .S(n7791), .Z(n7688) );
  NAND3_X1 U9313 ( .A1(n7689), .A2(n7690), .A3(n7688), .ZN(n7693) );
  NAND2_X1 U9314 ( .A1(n7695), .A2(n7690), .ZN(n7691) );
  NAND2_X1 U9315 ( .A1(n7691), .A2(n7797), .ZN(n7692) );
  NAND4_X1 U9316 ( .A1(n7693), .A2(n7696), .A3(n7698), .A4(n7692), .ZN(n7705)
         );
  INV_X1 U9317 ( .A(n7694), .ZN(n7704) );
  NAND2_X1 U9318 ( .A1(n7706), .A2(n7695), .ZN(n7701) );
  INV_X1 U9319 ( .A(n7695), .ZN(n7699) );
  OAI211_X1 U9320 ( .C1(n7699), .C2(n7698), .A(n7697), .B(n7696), .ZN(n7700)
         );
  MUX2_X1 U9321 ( .A(n7701), .B(n7700), .S(n7797), .Z(n7702) );
  INV_X1 U9322 ( .A(n7702), .ZN(n7703) );
  NAND3_X1 U9323 ( .A1(n7705), .A2(n7704), .A3(n7703), .ZN(n7715) );
  NAND2_X1 U9324 ( .A1(n7709), .A2(n7706), .ZN(n7707) );
  NAND2_X1 U9325 ( .A1(n7707), .A2(n7710), .ZN(n7713) );
  NAND2_X1 U9326 ( .A1(n7709), .A2(n7708), .ZN(n7711) );
  AND2_X1 U9327 ( .A1(n7711), .A2(n7710), .ZN(n7712) );
  MUX2_X1 U9328 ( .A(n7713), .B(n7712), .S(n7791), .Z(n7714) );
  NAND2_X1 U9329 ( .A1(n7715), .A2(n7714), .ZN(n7717) );
  NAND2_X1 U9330 ( .A1(n7717), .A2(n7716), .ZN(n7722) );
  MUX2_X1 U9331 ( .A(n7719), .B(n7718), .S(n7797), .Z(n7720) );
  MUX2_X1 U9332 ( .A(n7724), .B(n7723), .S(n7797), .Z(n7725) );
  NAND3_X1 U9333 ( .A1(n7726), .A2(n8557), .A3(n7725), .ZN(n7730) );
  OR2_X1 U9334 ( .A1(n8665), .A2(n7797), .ZN(n7728) );
  NAND2_X1 U9335 ( .A1(n8665), .A2(n7797), .ZN(n7727) );
  MUX2_X1 U9336 ( .A(n7728), .B(n7727), .S(n8538), .Z(n7729) );
  NAND3_X1 U9337 ( .A1(n7730), .A2(n8532), .A3(n7729), .ZN(n7734) );
  MUX2_X1 U9338 ( .A(n7732), .B(n7731), .S(n7797), .Z(n7733) );
  NAND2_X1 U9339 ( .A1(n7734), .A2(n7733), .ZN(n7735) );
  INV_X1 U9340 ( .A(n8516), .ZN(n8514) );
  NAND2_X1 U9341 ( .A1(n7735), .A2(n8514), .ZN(n7736) );
  NAND2_X1 U9342 ( .A1(n7737), .A2(n7736), .ZN(n7749) );
  NAND2_X1 U9343 ( .A1(n7739), .A2(n7738), .ZN(n7747) );
  AOI21_X1 U9344 ( .B1(n7749), .B2(n7740), .A(n7747), .ZN(n7744) );
  NAND2_X1 U9345 ( .A1(n7750), .A2(n7741), .ZN(n7743) );
  OAI211_X1 U9346 ( .C1(n7744), .C2(n7743), .A(n7742), .B(n7759), .ZN(n7746)
         );
  NAND3_X1 U9347 ( .A1(n7746), .A2(n7745), .A3(n7797), .ZN(n7757) );
  INV_X1 U9348 ( .A(n7757), .ZN(n7760) );
  INV_X1 U9349 ( .A(n8444), .ZN(n7756) );
  INV_X1 U9350 ( .A(n7747), .ZN(n7748) );
  AOI21_X1 U9351 ( .B1(n7749), .B2(n7748), .A(n8475), .ZN(n7752) );
  OAI211_X1 U9352 ( .C1(n7752), .C2(n7751), .A(n7750), .B(n8444), .ZN(n7753)
         );
  NAND3_X1 U9353 ( .A1(n7754), .A2(n7753), .A3(n7791), .ZN(n7755) );
  OAI21_X1 U9354 ( .B1(n7757), .B2(n7756), .A(n7755), .ZN(n7758) );
  OAI21_X1 U9355 ( .B1(n7760), .B2(n7759), .A(n7758), .ZN(n7761) );
  AOI21_X1 U9356 ( .B1(n7765), .B2(n4813), .A(n7791), .ZN(n7764) );
  AOI21_X1 U9357 ( .B1(n7766), .B2(n7765), .A(n7764), .ZN(n7769) );
  OAI21_X1 U9358 ( .B1(n7791), .B2(n7767), .A(n8099), .ZN(n7768) );
  NOR2_X1 U9359 ( .A1(n7769), .A2(n7768), .ZN(n7773) );
  MUX2_X1 U9360 ( .A(n7771), .B(n7770), .S(n7797), .Z(n7772) );
  OAI211_X1 U9361 ( .C1(n7774), .C2(n7773), .A(n8100), .B(n7772), .ZN(n7776)
         );
  INV_X1 U9362 ( .A(n8368), .ZN(n8349) );
  NAND2_X1 U9363 ( .A1(n7786), .A2(n8349), .ZN(n7779) );
  INV_X1 U9364 ( .A(n7782), .ZN(n7778) );
  AOI21_X1 U9365 ( .B1(n7779), .B2(n7780), .A(n7778), .ZN(n7785) );
  NAND2_X1 U9366 ( .A1(n7786), .A2(n8597), .ZN(n7783) );
  INV_X1 U9367 ( .A(n7780), .ZN(n7781) );
  AOI21_X1 U9368 ( .B1(n7783), .B2(n7782), .A(n7781), .ZN(n7784) );
  MUX2_X1 U9369 ( .A(n7785), .B(n7784), .S(n7797), .Z(n7796) );
  NOR2_X1 U9370 ( .A1(n8597), .A2(n8349), .ZN(n8342) );
  NAND3_X1 U9371 ( .A1(n7786), .A2(n8343), .A3(n8342), .ZN(n7789) );
  NAND3_X1 U9372 ( .A1(n7789), .A2(n7788), .A3(n7787), .ZN(n7795) );
  INV_X1 U9373 ( .A(n7790), .ZN(n7793) );
  OAI21_X1 U9374 ( .B1(n7796), .B2(n7795), .A(n7794), .ZN(n7801) );
  MUX2_X1 U9375 ( .A(n7799), .B(n7798), .S(n7797), .Z(n7800) );
  NAND2_X1 U9376 ( .A1(n7801), .A2(n7800), .ZN(n7803) );
  NAND2_X1 U9377 ( .A1(n7803), .A2(n7802), .ZN(n7805) );
  NAND2_X1 U9378 ( .A1(n7804), .A2(n7805), .ZN(n7809) );
  INV_X1 U9379 ( .A(n7805), .ZN(n7807) );
  NAND3_X1 U9380 ( .A1(n7807), .A2(n7806), .A3(n9982), .ZN(n7808) );
  INV_X1 U9381 ( .A(n8701), .ZN(n8328) );
  NAND4_X1 U9382 ( .A1(n9972), .A2(n8328), .A3(n7812), .A4(n8478), .ZN(n7813)
         );
  OAI211_X1 U9383 ( .C1(n7815), .C2(n7814), .A(n7813), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7816) );
  NAND2_X1 U9384 ( .A1(n8692), .A2(n5962), .ZN(n7818) );
  INV_X1 U9385 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9267) );
  OR2_X1 U9386 ( .A1(n7877), .A2(n9267), .ZN(n7817) );
  INV_X1 U9387 ( .A(n7982), .ZN(n8948) );
  AOI21_X1 U9388 ( .B1(n8955), .B2(n8974), .A(n8948), .ZN(n8023) );
  NAND2_X1 U9389 ( .A1(n9166), .A2(n8981), .ZN(n7983) );
  INV_X1 U9390 ( .A(n8997), .ZN(n8927) );
  NAND2_X1 U9391 ( .A1(n9175), .A2(n8982), .ZN(n8945) );
  INV_X1 U9392 ( .A(n8945), .ZN(n7819) );
  NAND2_X1 U9393 ( .A1(n8947), .A2(n7819), .ZN(n7820) );
  NAND3_X1 U9394 ( .A1(n7983), .A2(n7980), .A3(n7820), .ZN(n7822) );
  INV_X1 U9395 ( .A(n8974), .ZN(n7821) );
  AOI22_X1 U9396 ( .A1(n8023), .A2(n7822), .B1(n7821), .B2(n9162), .ZN(n8026)
         );
  INV_X1 U9397 ( .A(n8023), .ZN(n7872) );
  INV_X1 U9398 ( .A(n9037), .ZN(n8923) );
  NAND2_X1 U9399 ( .A1(n9187), .A2(n8923), .ZN(n9011) );
  OR2_X1 U9400 ( .A1(n9187), .A2(n8923), .ZN(n7958) );
  AND2_X1 U9401 ( .A1(n7958), .A2(n8942), .ZN(n7963) );
  NOR2_X1 U9402 ( .A1(n8944), .A2(n7963), .ZN(n7824) );
  NOR2_X1 U9403 ( .A1(n9175), .A2(n8982), .ZN(n8946) );
  INV_X1 U9404 ( .A(n8943), .ZN(n7823) );
  OR3_X1 U9405 ( .A1(n7824), .A2(n8946), .A3(n7823), .ZN(n8001) );
  INV_X1 U9406 ( .A(n9088), .ZN(n9116) );
  NAND2_X1 U9407 ( .A1(n9210), .A2(n9116), .ZN(n8937) );
  INV_X1 U9408 ( .A(n9104), .ZN(n9134) );
  NAND2_X1 U9409 ( .A1(n9217), .A2(n9134), .ZN(n8935) );
  AND2_X1 U9410 ( .A1(n8937), .A2(n8935), .ZN(n7951) );
  OR2_X1 U9411 ( .A1(n9217), .A2(n9134), .ZN(n8035) );
  INV_X1 U9412 ( .A(n8913), .ZN(n9144) );
  OR2_X1 U9413 ( .A1(n9222), .A2(n9144), .ZN(n9110) );
  NAND2_X1 U9414 ( .A1(n8035), .A2(n9110), .ZN(n8934) );
  OR2_X1 U9415 ( .A1(n9210), .A2(n9116), .ZN(n8034) );
  INV_X1 U9416 ( .A(n8034), .ZN(n7825) );
  INV_X1 U9417 ( .A(n9087), .ZN(n9054) );
  INV_X1 U9418 ( .A(n9103), .ZN(n9069) );
  NAND2_X1 U9419 ( .A1(n8033), .A2(n8938), .ZN(n7961) );
  AOI211_X1 U9420 ( .C1(n7951), .C2(n8934), .A(n7825), .B(n7961), .ZN(n7827)
         );
  INV_X1 U9421 ( .A(n9038), .ZN(n9070) );
  NAND2_X1 U9422 ( .A1(n9197), .A2(n9070), .ZN(n8061) );
  NAND2_X1 U9423 ( .A1(n9202), .A2(n9054), .ZN(n9049) );
  NAND2_X1 U9424 ( .A1(n8061), .A2(n9049), .ZN(n8941) );
  AND2_X1 U9425 ( .A1(n9205), .A2(n9069), .ZN(n8939) );
  AND2_X1 U9426 ( .A1(n8033), .A2(n8939), .ZN(n7826) );
  OR2_X1 U9427 ( .A1(n8941), .A2(n7826), .ZN(n7955) );
  OAI21_X1 U9428 ( .B1(n7827), .B2(n7955), .A(n8940), .ZN(n8019) );
  INV_X1 U9429 ( .A(n8019), .ZN(n7870) );
  NAND2_X1 U9430 ( .A1(n8822), .A2(n9835), .ZN(n7828) );
  AND2_X1 U9431 ( .A1(n7829), .A2(n7828), .ZN(n8004) );
  INV_X1 U9432 ( .A(n8004), .ZN(n7839) );
  INV_X1 U9433 ( .A(n8825), .ZN(n7836) );
  INV_X1 U9434 ( .A(n8002), .ZN(n7830) );
  AOI211_X1 U9435 ( .C1(n7831), .C2(n8823), .A(n6243), .B(n7830), .ZN(n7834)
         );
  INV_X1 U9436 ( .A(n7832), .ZN(n7833) );
  OAI211_X1 U9437 ( .C1(n7836), .C2(n7835), .A(n7834), .B(n7833), .ZN(n7838)
         );
  OAI21_X1 U9438 ( .B1(n7839), .B2(n7838), .A(n7837), .ZN(n7847) );
  NAND2_X1 U9439 ( .A1(n9595), .A2(n9143), .ZN(n8932) );
  INV_X1 U9440 ( .A(n8932), .ZN(n9139) );
  NAND2_X1 U9441 ( .A1(n9222), .A2(n9144), .ZN(n9112) );
  AND2_X1 U9442 ( .A1(n8935), .A2(n9112), .ZN(n8936) );
  INV_X1 U9443 ( .A(n8912), .ZN(n9584) );
  NAND2_X1 U9444 ( .A1(n9227), .A2(n9584), .ZN(n7942) );
  NAND2_X1 U9445 ( .A1(n8936), .A2(n7942), .ZN(n7848) );
  NAND2_X1 U9446 ( .A1(n9232), .A2(n9586), .ZN(n7927) );
  AND2_X1 U9447 ( .A1(n7927), .A2(n7840), .ZN(n7924) );
  INV_X1 U9448 ( .A(n7841), .ZN(n7842) );
  AND2_X1 U9449 ( .A1(n7919), .A2(n7842), .ZN(n7925) );
  INV_X1 U9450 ( .A(n7925), .ZN(n7844) );
  NOR2_X1 U9451 ( .A1(n7844), .A2(n4688), .ZN(n7854) );
  NAND3_X1 U9452 ( .A1(n7854), .A2(n7913), .A3(n7904), .ZN(n7845) );
  NOR3_X1 U9453 ( .A1(n7848), .A2(n4440), .A3(n7845), .ZN(n8014) );
  INV_X1 U9454 ( .A(n8014), .ZN(n7846) );
  AOI211_X1 U9455 ( .C1(n8003), .C2(n7847), .A(n9139), .B(n7846), .ZN(n7867)
         );
  INV_X1 U9456 ( .A(n7848), .ZN(n7863) );
  NOR2_X1 U9457 ( .A1(n9232), .A2(n9586), .ZN(n8929) );
  INV_X1 U9458 ( .A(n7849), .ZN(n7850) );
  OR2_X1 U9459 ( .A1(n8929), .A2(n7850), .ZN(n7928) );
  NAND2_X1 U9460 ( .A1(n7911), .A2(n7851), .ZN(n7852) );
  AND2_X1 U9461 ( .A1(n7852), .A2(n7919), .ZN(n7853) );
  NOR2_X1 U9462 ( .A1(n7928), .A2(n7853), .ZN(n7933) );
  INV_X1 U9463 ( .A(n7933), .ZN(n7860) );
  INV_X1 U9464 ( .A(n7854), .ZN(n7858) );
  NAND2_X1 U9465 ( .A1(n7855), .A2(n7916), .ZN(n7910) );
  INV_X1 U9466 ( .A(n7910), .ZN(n7856) );
  AND2_X1 U9467 ( .A1(n7922), .A2(n7856), .ZN(n7857) );
  NOR2_X1 U9468 ( .A1(n7858), .A2(n7857), .ZN(n7859) );
  OR2_X1 U9469 ( .A1(n7924), .A2(n8929), .ZN(n7930) );
  OAI211_X1 U9470 ( .C1(n7860), .C2(n7859), .A(n8932), .B(n7930), .ZN(n7861)
         );
  OR2_X1 U9471 ( .A1(n9227), .A2(n9584), .ZN(n7941) );
  OR2_X1 U9472 ( .A1(n9595), .A2(n9143), .ZN(n7935) );
  NAND3_X1 U9473 ( .A1(n7861), .A2(n7941), .A3(n7935), .ZN(n7862) );
  NAND2_X1 U9474 ( .A1(n7863), .A2(n7862), .ZN(n8017) );
  INV_X1 U9475 ( .A(n8017), .ZN(n7866) );
  INV_X1 U9476 ( .A(n7955), .ZN(n7864) );
  NAND2_X1 U9477 ( .A1(n7864), .A2(n8937), .ZN(n8015) );
  INV_X1 U9478 ( .A(n8015), .ZN(n7865) );
  OAI21_X1 U9479 ( .B1(n7867), .B2(n7866), .A(n7865), .ZN(n7869) );
  NAND2_X1 U9480 ( .A1(n9192), .A2(n9055), .ZN(n8032) );
  INV_X1 U9481 ( .A(n8032), .ZN(n7888) );
  NOR2_X1 U9482 ( .A1(n8944), .A2(n7888), .ZN(n8018) );
  INV_X1 U9483 ( .A(n8018), .ZN(n7868) );
  AOI21_X1 U9484 ( .B1(n7870), .B2(n7869), .A(n7868), .ZN(n7871) );
  OR4_X1 U9485 ( .A1(n7872), .A2(n8001), .A3(n8978), .A4(n7871), .ZN(n7876) );
  NAND2_X1 U9486 ( .A1(n8152), .A2(n5962), .ZN(n7874) );
  OR2_X1 U9487 ( .A1(n7877), .A2(n8155), .ZN(n7873) );
  INV_X1 U9488 ( .A(n8068), .ZN(n7875) );
  AOI21_X1 U9489 ( .B1(n8026), .B2(n7876), .A(n7875), .ZN(n7883) );
  NAND2_X1 U9490 ( .A1(n8687), .A2(n5962), .ZN(n7879) );
  OR2_X1 U9491 ( .A1(n7877), .A2(n6332), .ZN(n7878) );
  INV_X1 U9492 ( .A(n8896), .ZN(n7884) );
  NOR2_X1 U9493 ( .A1(n9157), .A2(n7884), .ZN(n8027) );
  INV_X1 U9494 ( .A(n8027), .ZN(n7881) );
  NAND2_X1 U9495 ( .A1(n8901), .A2(n8953), .ZN(n7880) );
  NAND2_X1 U9496 ( .A1(n7881), .A2(n7880), .ZN(n8071) );
  AND2_X1 U9497 ( .A1(n9157), .A2(n7884), .ZN(n8070) );
  INV_X1 U9498 ( .A(n8070), .ZN(n7882) );
  OAI21_X1 U9499 ( .B1(n7883), .B2(n8071), .A(n7882), .ZN(n8080) );
  NOR2_X1 U9500 ( .A1(n8080), .A2(n8000), .ZN(n8079) );
  OR2_X1 U9501 ( .A1(n8953), .A2(n7884), .ZN(n7885) );
  NAND2_X1 U9502 ( .A1(n8901), .A2(n7885), .ZN(n8025) );
  INV_X1 U9503 ( .A(n8942), .ZN(n7886) );
  NAND2_X1 U9504 ( .A1(n9011), .A2(n7886), .ZN(n7887) );
  AND2_X1 U9505 ( .A1(n8943), .A2(n7887), .ZN(n7891) );
  AND2_X1 U9506 ( .A1(n7958), .A2(n7888), .ZN(n7889) );
  NOR2_X1 U9507 ( .A1(n8944), .A2(n7889), .ZN(n7890) );
  INV_X1 U9508 ( .A(n7995), .ZN(n7988) );
  NAND2_X1 U9509 ( .A1(n7892), .A2(n7899), .ZN(n7894) );
  NAND2_X1 U9510 ( .A1(n7904), .A2(n8040), .ZN(n7893) );
  AOI21_X1 U9511 ( .B1(n7894), .B2(n7897), .A(n7893), .ZN(n7896) );
  INV_X1 U9512 ( .A(n7904), .ZN(n8047) );
  OAI211_X1 U9513 ( .C1(n8047), .C2(n7902), .A(n7995), .B(n8003), .ZN(n7895)
         );
  OR2_X1 U9514 ( .A1(n7896), .A2(n7895), .ZN(n7907) );
  AND2_X1 U9515 ( .A1(n7897), .A2(n8002), .ZN(n8006) );
  NAND2_X1 U9516 ( .A1(n7898), .A2(n8006), .ZN(n7901) );
  NAND3_X1 U9517 ( .A1(n7901), .A2(n7900), .A3(n7899), .ZN(n7903) );
  AND2_X1 U9518 ( .A1(n8003), .A2(n7902), .ZN(n8045) );
  NAND2_X1 U9519 ( .A1(n7903), .A2(n8045), .ZN(n7905) );
  NAND4_X1 U9520 ( .A1(n7905), .A2(n7988), .A3(n7904), .A4(n7913), .ZN(n7906)
         );
  NAND2_X1 U9521 ( .A1(n7907), .A2(n7906), .ZN(n7917) );
  INV_X1 U9522 ( .A(n7908), .ZN(n7909) );
  OAI21_X1 U9523 ( .B1(n7917), .B2(n7910), .A(n7909), .ZN(n7912) );
  NAND2_X1 U9524 ( .A1(n7914), .A2(n7913), .ZN(n7915) );
  AOI21_X1 U9525 ( .B1(n7917), .B2(n7916), .A(n7915), .ZN(n7921) );
  XNOR2_X1 U9526 ( .A(n9650), .B(n8815), .ZN(n9625) );
  OAI21_X1 U9527 ( .B1(n7922), .B2(n7995), .A(n9625), .ZN(n7923) );
  NAND2_X1 U9528 ( .A1(n7928), .A2(n7927), .ZN(n7929) );
  MUX2_X1 U9529 ( .A(n7930), .B(n7929), .S(n7988), .Z(n7931) );
  AND2_X1 U9530 ( .A1(n7931), .A2(n9588), .ZN(n7937) );
  AOI21_X1 U9531 ( .B1(n7932), .B2(n7937), .A(n9139), .ZN(n7940) );
  NAND2_X1 U9532 ( .A1(n7934), .A2(n7933), .ZN(n7938) );
  INV_X1 U9533 ( .A(n7935), .ZN(n7936) );
  AOI21_X1 U9534 ( .B1(n7938), .B2(n7937), .A(n7936), .ZN(n7939) );
  NAND2_X1 U9535 ( .A1(n7941), .A2(n7942), .ZN(n9137) );
  NAND2_X1 U9536 ( .A1(n9110), .A2(n9112), .ZN(n8036) );
  INV_X1 U9537 ( .A(n7941), .ZN(n7943) );
  INV_X1 U9538 ( .A(n7942), .ZN(n8933) );
  MUX2_X1 U9539 ( .A(n7943), .B(n8933), .S(n7995), .Z(n7944) );
  NOR2_X1 U9540 ( .A1(n8036), .A2(n7944), .ZN(n7945) );
  INV_X1 U9541 ( .A(n8934), .ZN(n7946) );
  MUX2_X1 U9542 ( .A(n8936), .B(n7946), .S(n7995), .Z(n7947) );
  AND2_X1 U9543 ( .A1(n8034), .A2(n8035), .ZN(n7949) );
  OR2_X1 U9544 ( .A1(n8939), .A2(n4673), .ZN(n7948) );
  AOI21_X1 U9545 ( .B1(n7952), .B2(n7949), .A(n7948), .ZN(n7954) );
  NAND2_X1 U9546 ( .A1(n8938), .A2(n8034), .ZN(n7950) );
  AOI21_X1 U9547 ( .B1(n7952), .B2(n7951), .A(n7950), .ZN(n7953) );
  MUX2_X1 U9548 ( .A(n7954), .B(n7953), .S(n7995), .Z(n7962) );
  AOI21_X1 U9549 ( .B1(n7962), .B2(n8033), .A(n7955), .ZN(n7957) );
  NAND2_X1 U9550 ( .A1(n8940), .A2(n7995), .ZN(n7956) );
  OAI211_X1 U9551 ( .C1(n7957), .C2(n7956), .A(n8032), .B(n9011), .ZN(n7959)
         );
  NAND2_X1 U9552 ( .A1(n7959), .A2(n7958), .ZN(n7967) );
  INV_X1 U9553 ( .A(n8941), .ZN(n7960) );
  OAI21_X1 U9554 ( .B1(n7962), .B2(n7961), .A(n7960), .ZN(n7964) );
  NAND3_X1 U9555 ( .A1(n7964), .A2(n7963), .A3(n8940), .ZN(n7965) );
  NAND2_X1 U9556 ( .A1(n7965), .A2(n7988), .ZN(n7966) );
  NAND2_X1 U9557 ( .A1(n7967), .A2(n7966), .ZN(n7968) );
  NAND2_X1 U9558 ( .A1(n9175), .A2(n8943), .ZN(n7970) );
  NAND2_X1 U9559 ( .A1(n7980), .A2(n7970), .ZN(n7973) );
  NAND2_X1 U9560 ( .A1(n8031), .A2(n9015), .ZN(n7971) );
  NAND2_X1 U9561 ( .A1(n8947), .A2(n7971), .ZN(n7972) );
  MUX2_X1 U9562 ( .A(n7973), .B(n7972), .S(n7995), .Z(n7974) );
  NAND2_X1 U9563 ( .A1(n8943), .A2(n8982), .ZN(n7975) );
  NAND2_X1 U9564 ( .A1(n8945), .A2(n7975), .ZN(n7978) );
  NOR2_X1 U9565 ( .A1(n8031), .A2(n9015), .ZN(n7976) );
  NOR2_X1 U9566 ( .A1(n7976), .A2(n9175), .ZN(n7977) );
  MUX2_X1 U9567 ( .A(n7978), .B(n7977), .S(n7995), .Z(n7979) );
  MUX2_X1 U9568 ( .A(n8947), .B(n7980), .S(n7995), .Z(n7981) );
  MUX2_X1 U9569 ( .A(n7983), .B(n7982), .S(n7995), .Z(n7984) );
  NOR3_X1 U9570 ( .A1(n7993), .A2(n9162), .A3(n8974), .ZN(n7992) );
  NAND2_X1 U9571 ( .A1(n8068), .A2(n8896), .ZN(n7986) );
  NAND2_X1 U9572 ( .A1(n7986), .A2(n9157), .ZN(n8028) );
  NAND2_X1 U9573 ( .A1(n8974), .A2(n7995), .ZN(n7987) );
  OAI211_X1 U9574 ( .C1(n8955), .C2(n7995), .A(n8028), .B(n7987), .ZN(n7991)
         );
  INV_X1 U9575 ( .A(n7993), .ZN(n7990) );
  NAND2_X1 U9576 ( .A1(n8974), .A2(n7988), .ZN(n7989) );
  OAI22_X1 U9577 ( .A1(n7992), .A2(n7991), .B1(n7990), .B2(n7989), .ZN(n7997)
         );
  INV_X1 U9578 ( .A(n8028), .ZN(n7996) );
  NAND3_X1 U9579 ( .A1(n8028), .A2(n7993), .A3(n9162), .ZN(n7994) );
  OAI21_X1 U9580 ( .B1(n8000), .B2(n7999), .A(n7998), .ZN(n8077) );
  INV_X1 U9581 ( .A(n8001), .ZN(n8022) );
  NAND4_X1 U9582 ( .A1(n8005), .A2(n8004), .A3(n8003), .A4(n8002), .ZN(n8013)
         );
  INV_X1 U9583 ( .A(n8006), .ZN(n8007) );
  AOI21_X1 U9584 ( .B1(n8009), .B2(n8008), .A(n8007), .ZN(n8011) );
  OAI21_X1 U9585 ( .B1(n8011), .B2(n8010), .A(n8045), .ZN(n8012) );
  NAND4_X1 U9586 ( .A1(n8014), .A2(n8932), .A3(n8013), .A4(n8012), .ZN(n8016)
         );
  AOI21_X1 U9587 ( .B1(n8017), .B2(n8016), .A(n8015), .ZN(n8020) );
  OAI21_X1 U9588 ( .B1(n8020), .B2(n8019), .A(n8018), .ZN(n8021) );
  NAND4_X1 U9589 ( .A1(n8023), .A2(n8022), .A3(n8947), .A4(n8021), .ZN(n8024)
         );
  NAND3_X1 U9590 ( .A1(n8026), .A2(n8025), .A3(n8024), .ZN(n8029) );
  AOI211_X1 U9591 ( .C1(n8029), .C2(n8028), .A(n6243), .B(n8027), .ZN(n8030)
         );
  NOR2_X1 U9592 ( .A1(n8030), .A2(n9073), .ZN(n8075) );
  XNOR2_X1 U9593 ( .A(n9175), .B(n8982), .ZN(n8995) );
  INV_X1 U9594 ( .A(n9013), .ZN(n8065) );
  INV_X1 U9595 ( .A(n9067), .ZN(n8060) );
  NAND2_X1 U9596 ( .A1(n8035), .A2(n8935), .ZN(n9113) );
  INV_X1 U9597 ( .A(n8036), .ZN(n9131) );
  NOR2_X1 U9598 ( .A1(n8038), .A2(n8037), .ZN(n8042) );
  NAND4_X1 U9599 ( .A1(n8042), .A2(n8041), .A3(n8040), .A4(n8039), .ZN(n8049)
         );
  NAND2_X1 U9600 ( .A1(n8044), .A2(n8043), .ZN(n8048) );
  INV_X1 U9601 ( .A(n8045), .ZN(n8046) );
  NOR4_X1 U9602 ( .A1(n8049), .A2(n8048), .A3(n8047), .A4(n8046), .ZN(n8053)
         );
  NAND4_X1 U9603 ( .A1(n8053), .A2(n8052), .A3(n8051), .A4(n8050), .ZN(n8055)
         );
  NOR2_X1 U9604 ( .A1(n8055), .A2(n8054), .ZN(n8056) );
  AND4_X1 U9605 ( .A1(n9588), .A2(n9611), .A3(n8056), .A4(n9625), .ZN(n8057)
         );
  NAND4_X1 U9606 ( .A1(n9131), .A2(n4842), .A3(n8057), .A4(n8930), .ZN(n8058)
         );
  NOR2_X1 U9607 ( .A1(n9113), .A2(n8058), .ZN(n8059) );
  NAND4_X1 U9608 ( .A1(n8060), .A2(n9101), .A3(n9085), .A4(n8059), .ZN(n8062)
         );
  NAND2_X1 U9609 ( .A1(n8940), .A2(n8061), .ZN(n9051) );
  NOR2_X1 U9610 ( .A1(n8062), .A2(n9051), .ZN(n8064) );
  INV_X1 U9611 ( .A(n9023), .ZN(n8063) );
  NAND4_X1 U9612 ( .A1(n8065), .A2(n9035), .A3(n8064), .A4(n8063), .ZN(n8066)
         );
  NOR3_X1 U9613 ( .A1(n8978), .A2(n8995), .A3(n8066), .ZN(n8067) );
  NAND4_X1 U9614 ( .A1(n8068), .A2(n8949), .A3(n8067), .A4(n8950), .ZN(n8069)
         );
  NOR3_X1 U9615 ( .A1(n8071), .A2(n8070), .A3(n8069), .ZN(n8073) );
  NOR2_X1 U9616 ( .A1(n8073), .A2(n8072), .ZN(n8074) );
  MUX2_X1 U9617 ( .A(n8075), .B(n9073), .S(n8074), .Z(n8076) );
  INV_X1 U9618 ( .A(n8080), .ZN(n8083) );
  OAI21_X1 U9619 ( .B1(n8083), .B2(n8082), .A(n8081), .ZN(n8090) );
  NOR4_X1 U9620 ( .A1(n8085), .A2(n8084), .A3(n6355), .A4(n9711), .ZN(n8089)
         );
  OAI21_X1 U9621 ( .B1(n8087), .B2(n8086), .A(P1_B_REG_SCAN_IN), .ZN(n8088) );
  INV_X1 U9622 ( .A(n8622), .ZN(n8430) );
  INV_X1 U9623 ( .A(n8520), .ZN(n8254) );
  INV_X1 U9624 ( .A(n9536), .ZN(n9545) );
  INV_X1 U9625 ( .A(n8493), .ZN(n8465) );
  NAND2_X1 U9626 ( .A1(n8454), .A2(n8094), .ZN(n8095) );
  OAI21_X1 U9627 ( .B1(n8481), .B2(n8093), .A(n8095), .ZN(n8436) );
  INV_X1 U9628 ( .A(n8629), .ZN(n8441) );
  AOI21_X1 U9629 ( .B1(n8436), .B2(n8098), .A(n8097), .ZN(n8433) );
  NAND2_X1 U9630 ( .A1(n8433), .A2(n8432), .ZN(n8624) );
  INV_X1 U9631 ( .A(n8242), .ZN(n8250) );
  XNOR2_X1 U9632 ( .A(n8341), .B(n8107), .ZN(n8601) );
  INV_X1 U9633 ( .A(n8614), .ZN(n8400) );
  NOR2_X1 U9634 ( .A1(n8101), .A2(n9536), .ZN(n8549) );
  INV_X1 U9635 ( .A(n8660), .ZN(n8546) );
  NAND2_X1 U9636 ( .A1(n8471), .A2(n8461), .ZN(n8455) );
  INV_X1 U9637 ( .A(n8362), .ZN(n8102) );
  AOI21_X1 U9638 ( .B1(n8597), .B2(n8102), .A(n8353), .ZN(n8598) );
  AOI22_X1 U9639 ( .A1(n8103), .A2(n9960), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9944), .ZN(n8104) );
  OAI21_X1 U9640 ( .B1(n8105), .B2(n8554), .A(n8104), .ZN(n8106) );
  AOI21_X1 U9641 ( .B1(n8598), .B2(n9951), .A(n8106), .ZN(n8112) );
  XNOR2_X1 U9642 ( .A(n8108), .B(n8107), .ZN(n8110) );
  INV_X1 U9643 ( .A(n8109), .ZN(n8249) );
  AOI222_X1 U9644 ( .A1(n8483), .A2(n8110), .B1(n8250), .B2(n8478), .C1(n8249), 
        .C2(n8480), .ZN(n8600) );
  OR2_X1 U9645 ( .A1(n8600), .A2(n9944), .ZN(n8111) );
  OAI211_X1 U9646 ( .C1(n8601), .C2(n8565), .A(n8112), .B(n8111), .ZN(P2_U3268) );
  OAI222_X1 U9647 ( .A1(n8704), .A2(n8115), .B1(n8702), .B2(n8114), .C1(n8113), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  XNOR2_X1 U9648 ( .A(n8117), .B(n8116), .ZN(n8118) );
  XNOR2_X1 U9649 ( .A(n8119), .B(n8118), .ZN(n8127) );
  INV_X1 U9650 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n8120) );
  NOR2_X1 U9651 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8120), .ZN(n9756) );
  NOR2_X1 U9652 ( .A1(n9568), .A2(n8121), .ZN(n8122) );
  AOI211_X1 U9653 ( .C1(n9564), .C2(n8820), .A(n9756), .B(n8122), .ZN(n8126)
         );
  AOI22_X1 U9654 ( .A1(n8124), .A2(n8798), .B1(n8810), .B2(n8123), .ZN(n8125)
         );
  OAI211_X1 U9655 ( .C1(n8127), .C2(n8812), .A(n8126), .B(n8125), .ZN(P1_U3237) );
  AOI22_X1 U9656 ( .A1(n8229), .A2(n8252), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8129) );
  NAND2_X1 U9657 ( .A1(n8222), .A2(n8439), .ZN(n8128) );
  OAI211_X1 U9658 ( .C1(n8447), .C2(n9916), .A(n8129), .B(n8128), .ZN(n8132)
         );
  NOR3_X1 U9659 ( .A1(n8130), .A2(n8196), .A3(n8179), .ZN(n8131) );
  AOI211_X1 U9660 ( .C1(n9902), .C2(n8629), .A(n8132), .B(n8131), .ZN(n8133)
         );
  OAI21_X1 U9661 ( .B1(n8134), .B2(n9909), .A(n8133), .ZN(P2_U3237) );
  OAI22_X1 U9662 ( .A1(n8179), .A2(n4913), .B1(n9981), .B2(n9909), .ZN(n8136)
         );
  NAND2_X1 U9663 ( .A1(n8136), .A2(n8135), .ZN(n8141) );
  NAND2_X1 U9664 ( .A1(n8138), .A2(n8137), .ZN(n8230) );
  AOI22_X1 U9665 ( .A1(n9902), .A2(n8139), .B1(n8230), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n8140) );
  OAI211_X1 U9666 ( .C1(n8142), .C2(n9915), .A(n8141), .B(n8140), .ZN(P2_U3234) );
  AOI21_X1 U9667 ( .B1(n8145), .B2(n8144), .A(n8143), .ZN(n8151) );
  AOI22_X1 U9668 ( .A1(n9564), .A2(n9015), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8148) );
  INV_X1 U9669 ( .A(n8146), .ZN(n8984) );
  NAND2_X1 U9670 ( .A1(n8798), .A2(n8984), .ZN(n8147) );
  OAI211_X1 U9671 ( .C1(n8981), .C2(n9568), .A(n8148), .B(n8147), .ZN(n8149)
         );
  AOI21_X1 U9672 ( .B1(n9172), .B2(n8810), .A(n8149), .ZN(n8150) );
  OAI21_X1 U9673 ( .B1(n8151), .B2(n8812), .A(n8150), .ZN(P1_U3212) );
  INV_X1 U9674 ( .A(n8152), .ZN(n8156) );
  OAI222_X1 U9675 ( .A1(n9277), .A2(n8156), .B1(n5645), .B2(P1_U3084), .C1(
        n8155), .C2(n4314), .ZN(P1_U3323) );
  NOR3_X1 U9676 ( .A1(n8157), .A2(n8393), .A3(n8179), .ZN(n8162) );
  AOI21_X1 U9677 ( .B1(n8158), .B2(n8159), .A(n9909), .ZN(n8161) );
  OAI21_X1 U9678 ( .B1(n8162), .B2(n8161), .A(n8160), .ZN(n8166) );
  NOR2_X1 U9679 ( .A1(n8393), .A2(n9916), .ZN(n8164) );
  OAI22_X1 U9680 ( .A1(n8368), .A2(n9915), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9469), .ZN(n8163) );
  AOI211_X1 U9681 ( .C1(n8222), .C2(n8363), .A(n8164), .B(n8163), .ZN(n8165)
         );
  OAI211_X1 U9682 ( .C1(n4900), .C2(n9913), .A(n8166), .B(n8165), .ZN(P2_U3216) );
  NAND2_X1 U9683 ( .A1(n8167), .A2(n9893), .ZN(n8170) );
  NAND2_X1 U9684 ( .A1(n9897), .A2(n8252), .ZN(n8169) );
  MUX2_X1 U9685 ( .A(n8170), .B(n8169), .S(n8168), .Z(n8175) );
  INV_X1 U9686 ( .A(n8171), .ZN(n8428) );
  AOI22_X1 U9687 ( .A1(n8228), .A2(n8096), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8172) );
  OAI21_X1 U9688 ( .B1(n8392), .B2(n9915), .A(n8172), .ZN(n8173) );
  AOI21_X1 U9689 ( .B1(n8428), .B2(n8222), .A(n8173), .ZN(n8174) );
  OAI211_X1 U9690 ( .C1(n8430), .C2(n9913), .A(n8175), .B(n8174), .ZN(P2_U3218) );
  INV_X1 U9691 ( .A(n8176), .ZN(n8177) );
  AOI21_X1 U9692 ( .B1(n8234), .B2(n8177), .A(n9909), .ZN(n8181) );
  NOR3_X1 U9693 ( .A1(n8179), .A2(n8178), .A3(n6633), .ZN(n8180) );
  OAI21_X1 U9694 ( .B1(n8181), .B2(n8180), .A(n6789), .ZN(n8186) );
  AOI22_X1 U9695 ( .A1(n9902), .A2(n8183), .B1(n9892), .B2(n8182), .ZN(n8185)
         );
  MUX2_X1 U9696 ( .A(P2_STATE_REG_SCAN_IN), .B(n9923), .S(n9368), .Z(n8184) );
  NAND3_X1 U9697 ( .A1(n8186), .A2(n8185), .A3(n8184), .ZN(P2_U3220) );
  AOI22_X1 U9698 ( .A1(n8228), .A2(n8265), .B1(n8229), .B2(n6842), .ZN(n8193)
         );
  AOI22_X1 U9699 ( .A1(n9902), .A2(n8187), .B1(n8230), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n8192) );
  OAI21_X1 U9700 ( .B1(n8189), .B2(n8188), .A(n8233), .ZN(n8190) );
  NAND2_X1 U9701 ( .A1(n8190), .A2(n9893), .ZN(n8191) );
  NAND3_X1 U9702 ( .A1(n8193), .A2(n8192), .A3(n8191), .ZN(P2_U3224) );
  XNOR2_X1 U9703 ( .A(n8195), .B(n8194), .ZN(n8201) );
  OAI22_X1 U9704 ( .A1(n9915), .A2(n8196), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9408), .ZN(n8197) );
  AOI21_X1 U9705 ( .B1(n8228), .B2(n8465), .A(n8197), .ZN(n8198) );
  OAI21_X1 U9706 ( .B1(n8458), .B2(n9923), .A(n8198), .ZN(n8199) );
  AOI21_X1 U9707 ( .B1(n8093), .B2(n9902), .A(n8199), .ZN(n8200) );
  OAI21_X1 U9708 ( .B1(n8201), .B2(n9909), .A(n8200), .ZN(P2_U3225) );
  XNOR2_X1 U9709 ( .A(n8203), .B(n8202), .ZN(n8204) );
  XNOR2_X1 U9710 ( .A(n8205), .B(n8204), .ZN(n8206) );
  NAND2_X1 U9711 ( .A1(n8206), .A2(n9893), .ZN(n8211) );
  OAI22_X1 U9712 ( .A1(n9916), .A2(n8392), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8207), .ZN(n8209) );
  NOR2_X1 U9713 ( .A1(n8393), .A2(n9915), .ZN(n8208) );
  AOI211_X1 U9714 ( .C1(n8222), .C2(n8397), .A(n8209), .B(n8208), .ZN(n8210)
         );
  OAI211_X1 U9715 ( .C1(n8400), .C2(n9913), .A(n8211), .B(n8210), .ZN(P2_U3227) );
  NAND2_X1 U9716 ( .A1(n9897), .A2(n4459), .ZN(n8215) );
  OR2_X1 U9717 ( .A1(n8212), .A2(n9909), .ZN(n8214) );
  MUX2_X1 U9718 ( .A(n8215), .B(n8214), .S(n8213), .Z(n8219) );
  NOR2_X1 U9719 ( .A1(n9923), .A2(n8408), .ZN(n8217) );
  OAI22_X1 U9720 ( .A1(n9916), .A2(n8448), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9346), .ZN(n8216) );
  AOI211_X1 U9721 ( .C1(n8229), .C2(n8251), .A(n8217), .B(n8216), .ZN(n8218)
         );
  OAI211_X1 U9722 ( .C1(n8411), .C2(n9913), .A(n8219), .B(n8218), .ZN(P2_U3231) );
  XNOR2_X1 U9723 ( .A(n8221), .B(n8220), .ZN(n8227) );
  AOI22_X1 U9724 ( .A1(n8229), .A2(n8481), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8224) );
  NAND2_X1 U9725 ( .A1(n8222), .A2(n8472), .ZN(n8223) );
  OAI211_X1 U9726 ( .C1(n8505), .C2(n9916), .A(n8224), .B(n8223), .ZN(n8225)
         );
  AOI21_X1 U9727 ( .B1(n8638), .B2(n9902), .A(n8225), .ZN(n8226) );
  OAI21_X1 U9728 ( .B1(n8227), .B2(n9909), .A(n8226), .ZN(P2_U3235) );
  AOI22_X1 U9729 ( .A1(n8229), .A2(n8263), .B1(n8228), .B2(n6997), .ZN(n8239)
         );
  AOI22_X1 U9730 ( .A1(n9902), .A2(n8231), .B1(n8230), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n8238) );
  AND2_X1 U9731 ( .A1(n8233), .A2(n8232), .ZN(n8236) );
  OAI211_X1 U9732 ( .C1(n8236), .C2(n8235), .A(n8234), .B(n9893), .ZN(n8237)
         );
  NAND3_X1 U9733 ( .A1(n8239), .A2(n8238), .A3(n8237), .ZN(P2_U3239) );
  OAI211_X1 U9734 ( .C1(n8240), .C2(n8241), .A(n8158), .B(n9893), .ZN(n8248)
         );
  OR2_X1 U9735 ( .A1(n8242), .A2(n8535), .ZN(n8244) );
  OR2_X1 U9736 ( .A1(n8415), .A2(n8537), .ZN(n8243) );
  NAND2_X1 U9737 ( .A1(n8244), .A2(n8243), .ZN(n8378) );
  INV_X1 U9738 ( .A(n8382), .ZN(n8245) );
  OAI22_X1 U9739 ( .A1(n8245), .A2(n9923), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9476), .ZN(n8246) );
  AOI21_X1 U9740 ( .B1(n8378), .B2(n9892), .A(n8246), .ZN(n8247) );
  OAI211_X1 U9741 ( .C1(n8375), .C2(n9913), .A(n8248), .B(n8247), .ZN(P2_U3242) );
  MUX2_X1 U9742 ( .A(n8347), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8264), .Z(
        P2_U3582) );
  MUX2_X1 U9743 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8249), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U9744 ( .A(n8349), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8264), .Z(
        P2_U3580) );
  MUX2_X1 U9745 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8250), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9746 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8251), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U9747 ( .A(n4459), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8264), .Z(
        P2_U3576) );
  MUX2_X1 U9748 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8252), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U9749 ( .A(n8096), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8264), .Z(
        P2_U3574) );
  MUX2_X1 U9750 ( .A(n8481), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8264), .Z(
        P2_U3573) );
  MUX2_X1 U9751 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8465), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9752 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8479), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9753 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8253), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9754 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8254), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9755 ( .A(n8255), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8264), .Z(
        P2_U3567) );
  MUX2_X1 U9756 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8256), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9757 ( .A(n9896), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8264), .Z(
        P2_U3563) );
  MUX2_X1 U9758 ( .A(n8257), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8264), .Z(
        P2_U3562) );
  MUX2_X1 U9759 ( .A(n8258), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8264), .Z(
        P2_U3561) );
  MUX2_X1 U9760 ( .A(n4814), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8264), .Z(
        P2_U3560) );
  MUX2_X1 U9761 ( .A(n8259), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8264), .Z(
        P2_U3559) );
  MUX2_X1 U9762 ( .A(n8260), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8264), .Z(
        P2_U3558) );
  MUX2_X1 U9763 ( .A(n8261), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8264), .Z(
        P2_U3557) );
  MUX2_X1 U9764 ( .A(n8262), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8264), .Z(
        P2_U3556) );
  MUX2_X1 U9765 ( .A(n8263), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8264), .Z(
        P2_U3555) );
  MUX2_X1 U9766 ( .A(n6842), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8264), .Z(
        P2_U3554) );
  MUX2_X1 U9767 ( .A(n6997), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8264), .Z(
        P2_U3553) );
  MUX2_X1 U9768 ( .A(n8265), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8264), .Z(
        P2_U3552) );
  OAI211_X1 U9769 ( .C1(n8268), .C2(n8267), .A(n9925), .B(n8266), .ZN(n8276)
         );
  AOI22_X1 U9770 ( .A1(n9926), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n8275) );
  NAND2_X1 U9771 ( .A1(n8291), .A2(n8269), .ZN(n8274) );
  OAI211_X1 U9772 ( .C1(n8272), .C2(n8271), .A(n9924), .B(n8270), .ZN(n8273)
         );
  NAND4_X1 U9773 ( .A1(n8276), .A2(n8275), .A3(n8274), .A4(n8273), .ZN(
        P2_U3246) );
  INV_X1 U9774 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8284) );
  XNOR2_X1 U9775 ( .A(n8300), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8280) );
  OR2_X1 U9776 ( .A1(n8286), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8278) );
  NAND2_X1 U9777 ( .A1(n8278), .A2(n8277), .ZN(n8279) );
  NOR2_X1 U9778 ( .A1(n8280), .A2(n8279), .ZN(n8299) );
  AOI21_X1 U9779 ( .B1(n8280), .B2(n8279), .A(n8299), .ZN(n8281) );
  NAND2_X1 U9780 ( .A1(n9924), .A2(n8281), .ZN(n8283) );
  NAND2_X1 U9781 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3152), .ZN(n8282) );
  OAI211_X1 U9782 ( .C1(n8325), .C2(n8284), .A(n8283), .B(n8282), .ZN(n8290)
         );
  NAND2_X1 U9783 ( .A1(n8300), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8295) );
  OAI21_X1 U9784 ( .B1(n8300), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8295), .ZN(
        n8287) );
  AOI211_X1 U9785 ( .C1(n8288), .C2(n8287), .A(n8293), .B(n9929), .ZN(n8289)
         );
  AOI211_X1 U9786 ( .C1(n8291), .C2(n8300), .A(n8290), .B(n8289), .ZN(n8292)
         );
  INV_X1 U9787 ( .A(n8292), .ZN(P2_U3262) );
  INV_X1 U9788 ( .A(n8315), .ZN(n8305) );
  NAND2_X1 U9789 ( .A1(n8295), .A2(n8294), .ZN(n8310) );
  XNOR2_X1 U9790 ( .A(n8305), .B(n8310), .ZN(n8297) );
  INV_X1 U9791 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8296) );
  NAND2_X1 U9792 ( .A1(n8297), .A2(n8296), .ZN(n8311) );
  OAI21_X1 U9793 ( .B1(n8297), .B2(n8296), .A(n8311), .ZN(n8308) );
  INV_X1 U9794 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8304) );
  INV_X1 U9795 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8298) );
  XNOR2_X1 U9796 ( .A(n8315), .B(n8298), .ZN(n8318) );
  AOI21_X1 U9797 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8300), .A(n8299), .ZN(
        n8317) );
  XNOR2_X1 U9798 ( .A(n8318), .B(n8317), .ZN(n8301) );
  NAND2_X1 U9799 ( .A1(n9924), .A2(n8301), .ZN(n8303) );
  OAI211_X1 U9800 ( .C1(n8325), .C2(n8304), .A(n8303), .B(n8302), .ZN(n8307)
         );
  NOR2_X1 U9801 ( .A1(n9927), .A2(n8305), .ZN(n8306) );
  AOI211_X1 U9802 ( .C1(n9925), .C2(n8308), .A(n8307), .B(n8306), .ZN(n8309)
         );
  INV_X1 U9803 ( .A(n8309), .ZN(P2_U3263) );
  INV_X1 U9804 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8326) );
  INV_X1 U9805 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8314) );
  OR2_X1 U9806 ( .A1(n8315), .A2(n8310), .ZN(n8312) );
  NAND2_X1 U9807 ( .A1(n8312), .A2(n8311), .ZN(n8313) );
  XNOR2_X1 U9808 ( .A(n8314), .B(n8313), .ZN(n8323) );
  INV_X1 U9809 ( .A(n8323), .ZN(n8321) );
  NOR2_X1 U9810 ( .A1(n8315), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8316) );
  AOI21_X1 U9811 ( .B1(n8318), .B2(n8317), .A(n8316), .ZN(n8319) );
  XNOR2_X1 U9812 ( .A(n8319), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U9813 ( .A1(n9924), .A2(n8322), .ZN(n8320) );
  AND2_X1 U9814 ( .A1(n8328), .A2(P2_B_REG_SCAN_IN), .ZN(n8329) );
  NOR2_X1 U9815 ( .A1(n8535), .A2(n8329), .ZN(n8348) );
  INV_X1 U9816 ( .A(n8348), .ZN(n8330) );
  NOR2_X1 U9817 ( .A1(n8331), .A2(n8330), .ZN(n9541) );
  INV_X1 U9818 ( .A(n9541), .ZN(n8332) );
  NOR2_X1 U9819 ( .A1(n9944), .A2(n8332), .ZN(n8336) );
  AOI21_X1 U9820 ( .B1(n9944), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8336), .ZN(
        n8334) );
  NAND2_X1 U9821 ( .A1(n9542), .A2(n9945), .ZN(n8333) );
  OAI211_X1 U9822 ( .C1(n9540), .C2(n8354), .A(n8334), .B(n8333), .ZN(P2_U3265) );
  INV_X1 U9823 ( .A(n8352), .ZN(n8335) );
  NOR2_X1 U9824 ( .A1(n8339), .A2(n8335), .ZN(n8585) );
  OR3_X1 U9825 ( .A1(n8585), .A2(n8584), .A3(n8354), .ZN(n8338) );
  AOI21_X1 U9826 ( .B1(n9944), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8336), .ZN(
        n8337) );
  OAI211_X1 U9827 ( .C1(n8339), .C2(n8554), .A(n8338), .B(n8337), .ZN(P2_U3266) );
  XNOR2_X1 U9828 ( .A(n8344), .B(n8346), .ZN(n8590) );
  INV_X1 U9829 ( .A(n8590), .ZN(n8360) );
  XOR2_X1 U9830 ( .A(n8346), .B(n8345), .Z(n8351) );
  AOI22_X1 U9831 ( .A1(n8349), .A2(n8478), .B1(n8348), .B2(n8347), .ZN(n8350)
         );
  OAI21_X1 U9832 ( .B1(n8591), .B2(n8353), .A(n8352), .ZN(n8592) );
  NOR2_X1 U9833 ( .A1(n8592), .A2(n8354), .ZN(n8358) );
  AOI22_X1 U9834 ( .A1(P2_REG2_REG_29__SCAN_IN), .A2(n9944), .B1(n8355), .B2(
        n9960), .ZN(n8356) );
  OAI21_X1 U9835 ( .B1(n8591), .B2(n8554), .A(n8356), .ZN(n8357) );
  AOI211_X1 U9836 ( .C1(n8594), .C2(n9968), .A(n8358), .B(n8357), .ZN(n8359)
         );
  OAI21_X1 U9837 ( .B1(n8360), .B2(n8565), .A(n8359), .ZN(P2_U3267) );
  XNOR2_X1 U9838 ( .A(n8361), .B(n8367), .ZN(n8606) );
  AOI21_X1 U9839 ( .B1(n8602), .B2(n8380), .A(n8362), .ZN(n8603) );
  AOI22_X1 U9840 ( .A1(n8363), .A2(n9960), .B1(n9944), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8364) );
  OAI21_X1 U9841 ( .B1(n4900), .B2(n8554), .A(n8364), .ZN(n8372) );
  AOI211_X1 U9842 ( .C1(n8367), .C2(n8366), .A(n9939), .B(n8365), .ZN(n8370)
         );
  OAI22_X1 U9843 ( .A1(n8368), .A2(n8535), .B1(n8393), .B2(n8537), .ZN(n8369)
         );
  NOR2_X1 U9844 ( .A1(n8370), .A2(n8369), .ZN(n8605) );
  NOR2_X1 U9845 ( .A1(n8605), .A2(n9944), .ZN(n8371) );
  AOI211_X1 U9846 ( .C1(n9951), .C2(n8603), .A(n8372), .B(n8371), .ZN(n8373)
         );
  OAI21_X1 U9847 ( .B1(n8606), .B2(n8565), .A(n8373), .ZN(P2_U3269) );
  XNOR2_X1 U9848 ( .A(n8374), .B(n4581), .ZN(n8611) );
  NOR2_X1 U9849 ( .A1(n8375), .A2(n8554), .ZN(n8386) );
  XNOR2_X1 U9850 ( .A(n8377), .B(n8376), .ZN(n8379) );
  INV_X1 U9851 ( .A(n8380), .ZN(n8381) );
  AOI211_X1 U9852 ( .C1(n8608), .C2(n8394), .A(n10049), .B(n8381), .ZN(n8607)
         );
  AOI22_X1 U9853 ( .A1(n8607), .A2(n8383), .B1(n9960), .B2(n8382), .ZN(n8384)
         );
  AOI21_X1 U9854 ( .B1(n8610), .B2(n8384), .A(n9944), .ZN(n8385) );
  AOI211_X1 U9855 ( .C1(n9944), .C2(P2_REG2_REG_26__SCAN_IN), .A(n8386), .B(
        n8385), .ZN(n8387) );
  OAI21_X1 U9856 ( .B1(n8565), .B2(n8611), .A(n8387), .ZN(P2_U3270) );
  XNOR2_X1 U9857 ( .A(n8388), .B(n8389), .ZN(n8616) );
  XNOR2_X1 U9858 ( .A(n8390), .B(n8389), .ZN(n8391) );
  OAI222_X1 U9859 ( .A1(n8535), .A2(n8393), .B1(n8537), .B2(n8392), .C1(n9939), 
        .C2(n8391), .ZN(n8612) );
  INV_X1 U9860 ( .A(n8406), .ZN(n8396) );
  INV_X1 U9861 ( .A(n8394), .ZN(n8395) );
  AOI211_X1 U9862 ( .C1(n8614), .C2(n8396), .A(n10049), .B(n8395), .ZN(n8613)
         );
  NOR2_X1 U9863 ( .A1(n9944), .A2(n9962), .ZN(n8524) );
  NAND2_X1 U9864 ( .A1(n8613), .A2(n8524), .ZN(n8399) );
  AOI22_X1 U9865 ( .A1(n9944), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8397), .B2(
        n9960), .ZN(n8398) );
  OAI211_X1 U9866 ( .C1(n8400), .C2(n8554), .A(n8399), .B(n8398), .ZN(n8401)
         );
  AOI21_X1 U9867 ( .B1(n8612), .B2(n9968), .A(n8401), .ZN(n8402) );
  OAI21_X1 U9868 ( .B1(n8616), .B2(n8565), .A(n8402), .ZN(P2_U3271) );
  AOI21_X1 U9869 ( .B1(n8405), .B2(n8404), .A(n8403), .ZN(n8621) );
  INV_X1 U9870 ( .A(n8427), .ZN(n8407) );
  AOI21_X1 U9871 ( .B1(n8617), .B2(n8407), .A(n8406), .ZN(n8618) );
  INV_X1 U9872 ( .A(n8408), .ZN(n8409) );
  AOI22_X1 U9873 ( .A1(n9944), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8409), .B2(
        n9960), .ZN(n8410) );
  OAI21_X1 U9874 ( .B1(n8411), .B2(n8554), .A(n8410), .ZN(n8420) );
  NOR2_X1 U9875 ( .A1(n8412), .A2(n9939), .ZN(n8418) );
  OAI21_X1 U9876 ( .B1(n8423), .B2(n8414), .A(n8413), .ZN(n8417) );
  OAI22_X1 U9877 ( .A1(n8415), .A2(n8535), .B1(n8448), .B2(n8537), .ZN(n8416)
         );
  AOI21_X1 U9878 ( .B1(n8418), .B2(n8417), .A(n8416), .ZN(n8620) );
  NOR2_X1 U9879 ( .A1(n8620), .A2(n9944), .ZN(n8419) );
  AOI211_X1 U9880 ( .C1(n8618), .C2(n9951), .A(n8420), .B(n8419), .ZN(n8421)
         );
  OAI21_X1 U9881 ( .B1(n8621), .B2(n8565), .A(n8421), .ZN(P2_U3272) );
  INV_X1 U9882 ( .A(n8423), .ZN(n8424) );
  OAI21_X1 U9883 ( .B1(n4805), .B2(n8425), .A(n8424), .ZN(n8426) );
  AOI222_X1 U9884 ( .A1(n8483), .A2(n8426), .B1(n8096), .B2(n8478), .C1(n4459), 
        .C2(n8480), .ZN(n8628) );
  AOI21_X1 U9885 ( .B1(n8622), .B2(n8437), .A(n8427), .ZN(n8623) );
  AOI22_X1 U9886 ( .A1(n9944), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8428), .B2(
        n9960), .ZN(n8429) );
  OAI21_X1 U9887 ( .B1(n8430), .B2(n8554), .A(n8429), .ZN(n8431) );
  AOI21_X1 U9888 ( .B1(n8623), .B2(n9951), .A(n8431), .ZN(n8435) );
  OR2_X1 U9889 ( .A1(n8433), .A2(n8432), .ZN(n8625) );
  NAND3_X1 U9890 ( .A1(n8625), .A2(n8624), .A3(n8576), .ZN(n8434) );
  OAI211_X1 U9891 ( .C1(n8628), .C2(n9944), .A(n8435), .B(n8434), .ZN(P2_U3273) );
  XNOR2_X1 U9892 ( .A(n8436), .B(n8443), .ZN(n8633) );
  INV_X1 U9893 ( .A(n8437), .ZN(n8438) );
  AOI21_X1 U9894 ( .B1(n8629), .B2(n8455), .A(n8438), .ZN(n8630) );
  AOI22_X1 U9895 ( .A1(n9944), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8439), .B2(
        n9960), .ZN(n8440) );
  OAI21_X1 U9896 ( .B1(n8441), .B2(n8554), .A(n8440), .ZN(n8452) );
  INV_X1 U9897 ( .A(n8442), .ZN(n8446) );
  AOI21_X1 U9898 ( .B1(n8462), .B2(n8444), .A(n8443), .ZN(n8445) );
  NOR3_X1 U9899 ( .A1(n8446), .A2(n8445), .A3(n9939), .ZN(n8450) );
  OAI22_X1 U9900 ( .A1(n8448), .A2(n8535), .B1(n8447), .B2(n8537), .ZN(n8449)
         );
  NOR2_X1 U9901 ( .A1(n8450), .A2(n8449), .ZN(n8632) );
  NOR2_X1 U9902 ( .A1(n8632), .A2(n9944), .ZN(n8451) );
  AOI211_X1 U9903 ( .C1(n8630), .C2(n9951), .A(n8452), .B(n8451), .ZN(n8453)
         );
  OAI21_X1 U9904 ( .B1(n8633), .B2(n8565), .A(n8453), .ZN(P2_U3274) );
  XNOR2_X1 U9905 ( .A(n8454), .B(n8463), .ZN(n8637) );
  INV_X1 U9906 ( .A(n8471), .ZN(n8457) );
  INV_X1 U9907 ( .A(n8455), .ZN(n8456) );
  AOI21_X1 U9908 ( .B1(n8093), .B2(n8457), .A(n8456), .ZN(n8634) );
  INV_X1 U9909 ( .A(n8458), .ZN(n8459) );
  AOI22_X1 U9910 ( .A1(n9944), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8459), .B2(
        n9960), .ZN(n8460) );
  OAI21_X1 U9911 ( .B1(n8461), .B2(n8554), .A(n8460), .ZN(n8468) );
  OAI21_X1 U9912 ( .B1(n8464), .B2(n8463), .A(n8462), .ZN(n8466) );
  AOI222_X1 U9913 ( .A1(n8483), .A2(n8466), .B1(n8096), .B2(n8480), .C1(n8465), 
        .C2(n8478), .ZN(n8636) );
  NOR2_X1 U9914 ( .A1(n8636), .A2(n9944), .ZN(n8467) );
  AOI211_X1 U9915 ( .C1(n8634), .C2(n9951), .A(n8468), .B(n8467), .ZN(n8469)
         );
  OAI21_X1 U9916 ( .B1(n8565), .B2(n8637), .A(n8469), .ZN(P2_U3275) );
  XNOR2_X1 U9917 ( .A(n8470), .B(n8476), .ZN(n8642) );
  AOI21_X1 U9918 ( .B1(n8638), .B2(n4718), .A(n8471), .ZN(n8639) );
  AOI22_X1 U9919 ( .A1(n9944), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8472), .B2(
        n9960), .ZN(n8473) );
  OAI21_X1 U9920 ( .B1(n8474), .B2(n8554), .A(n8473), .ZN(n8485) );
  NOR2_X1 U9921 ( .A1(n8489), .A2(n8475), .ZN(n8477) );
  XNOR2_X1 U9922 ( .A(n8477), .B(n8476), .ZN(n8482) );
  AOI222_X1 U9923 ( .A1(n8483), .A2(n8482), .B1(n8481), .B2(n8480), .C1(n8479), 
        .C2(n8478), .ZN(n8641) );
  NOR2_X1 U9924 ( .A1(n8641), .A2(n9944), .ZN(n8484) );
  AOI211_X1 U9925 ( .C1(n8639), .C2(n9951), .A(n8485), .B(n8484), .ZN(n8486)
         );
  OAI21_X1 U9926 ( .B1(n8565), .B2(n8642), .A(n8486), .ZN(P2_U3276) );
  XNOR2_X1 U9927 ( .A(n8488), .B(n8487), .ZN(n8647) );
  AOI21_X1 U9928 ( .B1(n8491), .B2(n8490), .A(n8489), .ZN(n8492) );
  OAI222_X1 U9929 ( .A1(n8535), .A2(n8493), .B1(n8537), .B2(n8519), .C1(n9939), 
        .C2(n8492), .ZN(n8643) );
  AOI211_X1 U9930 ( .C1(n8645), .C2(n8506), .A(n10049), .B(n8494), .ZN(n8644)
         );
  NAND2_X1 U9931 ( .A1(n8644), .A2(n8524), .ZN(n8497) );
  AOI22_X1 U9932 ( .A1(n9944), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8495), .B2(
        n9960), .ZN(n8496) );
  OAI211_X1 U9933 ( .C1(n4716), .C2(n8554), .A(n8497), .B(n8496), .ZN(n8498)
         );
  AOI21_X1 U9934 ( .B1(n8643), .B2(n9968), .A(n8498), .ZN(n8499) );
  OAI21_X1 U9935 ( .B1(n8565), .B2(n8647), .A(n8499), .ZN(P2_U3277) );
  XNOR2_X1 U9936 ( .A(n8500), .B(n8502), .ZN(n8653) );
  AOI21_X1 U9937 ( .B1(n8503), .B2(n8502), .A(n8501), .ZN(n8504) );
  OAI222_X1 U9938 ( .A1(n8537), .A2(n8536), .B1(n8535), .B2(n8505), .C1(n9939), 
        .C2(n8504), .ZN(n8648) );
  INV_X1 U9939 ( .A(n8506), .ZN(n8507) );
  AOI21_X1 U9940 ( .B1(n8649), .B2(n8521), .A(n8507), .ZN(n8650) );
  NAND2_X1 U9941 ( .A1(n8650), .A2(n9951), .ZN(n8510) );
  AOI22_X1 U9942 ( .A1(n9944), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8508), .B2(
        n9960), .ZN(n8509) );
  OAI211_X1 U9943 ( .C1(n8511), .C2(n8554), .A(n8510), .B(n8509), .ZN(n8512)
         );
  AOI21_X1 U9944 ( .B1(n8648), .B2(n9968), .A(n8512), .ZN(n8513) );
  OAI21_X1 U9945 ( .B1(n8653), .B2(n8565), .A(n8513), .ZN(P2_U3278) );
  XNOR2_X1 U9946 ( .A(n8515), .B(n8514), .ZN(n8658) );
  XNOR2_X1 U9947 ( .A(n8517), .B(n8516), .ZN(n8518) );
  OAI222_X1 U9948 ( .A1(n8537), .A2(n8520), .B1(n8535), .B2(n8519), .C1(n8518), 
        .C2(n9939), .ZN(n8654) );
  INV_X1 U9949 ( .A(n8541), .ZN(n8523) );
  INV_X1 U9950 ( .A(n8521), .ZN(n8522) );
  AOI211_X1 U9951 ( .C1(n8656), .C2(n8523), .A(n10049), .B(n8522), .ZN(n8655)
         );
  NAND2_X1 U9952 ( .A1(n8655), .A2(n8524), .ZN(n8527) );
  AOI22_X1 U9953 ( .A1(n9944), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8525), .B2(
        n9960), .ZN(n8526) );
  OAI211_X1 U9954 ( .C1(n8528), .C2(n8554), .A(n8527), .B(n8526), .ZN(n8529)
         );
  AOI21_X1 U9955 ( .B1(n8654), .B2(n9968), .A(n8529), .ZN(n8530) );
  OAI21_X1 U9956 ( .B1(n8658), .B2(n8565), .A(n8530), .ZN(P2_U3279) );
  AOI21_X1 U9957 ( .B1(n8532), .B2(n8531), .A(n4388), .ZN(n8659) );
  XNOR2_X1 U9958 ( .A(n8533), .B(n8532), .ZN(n8534) );
  NOR2_X1 U9959 ( .A1(n8534), .A2(n9939), .ZN(n8540) );
  OAI22_X1 U9960 ( .A1(n8538), .A2(n8537), .B1(n8536), .B2(n8535), .ZN(n8539)
         );
  AOI211_X1 U9961 ( .C1(n8659), .C2(n9942), .A(n8540), .B(n8539), .ZN(n8663)
         );
  INV_X1 U9962 ( .A(n8550), .ZN(n8542) );
  AOI21_X1 U9963 ( .B1(n8660), .B2(n8542), .A(n8541), .ZN(n8661) );
  NAND2_X1 U9964 ( .A1(n8661), .A2(n9951), .ZN(n8545) );
  AOI22_X1 U9965 ( .A1(n9944), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8543), .B2(
        n9960), .ZN(n8544) );
  OAI211_X1 U9966 ( .C1(n8546), .C2(n8554), .A(n8545), .B(n8544), .ZN(n8547)
         );
  AOI21_X1 U9967 ( .B1(n8659), .B2(n9952), .A(n8547), .ZN(n8548) );
  OAI21_X1 U9968 ( .B1(n8663), .B2(n9944), .A(n8548), .ZN(P2_U3280) );
  XOR2_X1 U9969 ( .A(n8557), .B(n4386), .Z(n8669) );
  INV_X1 U9970 ( .A(n8549), .ZN(n8551) );
  AOI21_X1 U9971 ( .B1(n8665), .B2(n8551), .A(n8550), .ZN(n8666) );
  AOI22_X1 U9972 ( .A1(n9944), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8552), .B2(
        n9960), .ZN(n8553) );
  OAI21_X1 U9973 ( .B1(n8555), .B2(n8554), .A(n8553), .ZN(n8563) );
  INV_X1 U9974 ( .A(n8556), .ZN(n8558) );
  AOI21_X1 U9975 ( .B1(n8558), .B2(n4909), .A(n9939), .ZN(n8561) );
  AOI21_X1 U9976 ( .B1(n8561), .B2(n8560), .A(n8559), .ZN(n8668) );
  NOR2_X1 U9977 ( .A1(n8668), .A2(n9944), .ZN(n8562) );
  AOI211_X1 U9978 ( .C1(n8666), .C2(n9951), .A(n8563), .B(n8562), .ZN(n8564)
         );
  OAI21_X1 U9979 ( .B1(n8565), .B2(n8669), .A(n8564), .ZN(P2_U3281) );
  OAI21_X1 U9980 ( .B1(n8568), .B2(n8567), .A(n8566), .ZN(n8570) );
  AOI21_X1 U9981 ( .B1(n8570), .B2(n8569), .A(n9939), .ZN(n8572) );
  NOR2_X1 U9982 ( .A1(n8572), .A2(n8571), .ZN(n10025) );
  MUX2_X1 U9983 ( .A(n6485), .B(n10025), .S(n9968), .Z(n8583) );
  AOI22_X1 U9984 ( .A1(n9945), .A2(n10017), .B1(n8573), .B2(n9960), .ZN(n8582)
         );
  NAND2_X1 U9985 ( .A1(n8574), .A2(n8575), .ZN(n10021) );
  NAND3_X1 U9986 ( .A1(n10022), .A2(n10021), .A3(n8576), .ZN(n8581) );
  INV_X1 U9987 ( .A(n8577), .ZN(n8578) );
  AOI21_X1 U9988 ( .B1(n10017), .B2(n8579), .A(n8578), .ZN(n10020) );
  NAND2_X1 U9989 ( .A1(n10020), .A2(n9951), .ZN(n8580) );
  NAND4_X1 U9990 ( .A1(n8583), .A2(n8582), .A3(n8581), .A4(n8580), .ZN(
        P2_U3288) );
  INV_X1 U9991 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8588) );
  NOR3_X1 U9992 ( .A1(n8585), .A2(n8584), .A3(n10049), .ZN(n8586) );
  AOI211_X1 U9993 ( .C1(n10018), .C2(n8587), .A(n9541), .B(n8586), .ZN(n8670)
         );
  MUX2_X1 U9994 ( .A(n8588), .B(n8670), .S(n10077), .Z(n8589) );
  INV_X1 U9995 ( .A(n8589), .ZN(P2_U3550) );
  NAND2_X1 U9996 ( .A1(n8590), .A2(n10054), .ZN(n8596) );
  OAI22_X1 U9997 ( .A1(n8592), .A2(n10049), .B1(n8591), .B2(n10048), .ZN(n8593) );
  NOR2_X1 U9998 ( .A1(n8594), .A2(n8593), .ZN(n8595) );
  NAND2_X1 U9999 ( .A1(n8596), .A2(n8595), .ZN(n8672) );
  MUX2_X1 U10000 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8672), .S(n10077), .Z(
        P2_U3549) );
  AOI22_X1 U10001 ( .A1(n8598), .A2(n10019), .B1(n10018), .B2(n8597), .ZN(
        n8599) );
  OAI211_X1 U10002 ( .C1(n8601), .C2(n9983), .A(n8600), .B(n8599), .ZN(n8673)
         );
  MUX2_X1 U10003 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8673), .S(n10077), .Z(
        P2_U3548) );
  AOI22_X1 U10004 ( .A1(n8603), .A2(n10019), .B1(n10018), .B2(n8602), .ZN(
        n8604) );
  OAI211_X1 U10005 ( .C1(n8606), .C2(n9983), .A(n8605), .B(n8604), .ZN(n8674)
         );
  MUX2_X1 U10006 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8674), .S(n10077), .Z(
        P2_U3547) );
  AOI21_X1 U10007 ( .B1(n10018), .B2(n8608), .A(n8607), .ZN(n8609) );
  OAI211_X1 U10008 ( .C1(n8611), .C2(n9983), .A(n8610), .B(n8609), .ZN(n8675)
         );
  MUX2_X1 U10009 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8675), .S(n10077), .Z(
        P2_U3546) );
  AOI211_X1 U10010 ( .C1(n10018), .C2(n8614), .A(n8613), .B(n8612), .ZN(n8615)
         );
  OAI21_X1 U10011 ( .B1(n9983), .B2(n8616), .A(n8615), .ZN(n8676) );
  MUX2_X1 U10012 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8676), .S(n10077), .Z(
        P2_U3545) );
  AOI22_X1 U10013 ( .A1(n8618), .A2(n10019), .B1(n10018), .B2(n8617), .ZN(
        n8619) );
  OAI211_X1 U10014 ( .C1(n8621), .C2(n9983), .A(n8620), .B(n8619), .ZN(n8677)
         );
  MUX2_X1 U10015 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8677), .S(n10077), .Z(
        P2_U3544) );
  AOI22_X1 U10016 ( .A1(n8623), .A2(n10019), .B1(n10018), .B2(n8622), .ZN(
        n8627) );
  NAND3_X1 U10017 ( .A1(n8625), .A2(n8624), .A3(n10054), .ZN(n8626) );
  NAND3_X1 U10018 ( .A1(n8628), .A2(n8627), .A3(n8626), .ZN(n8678) );
  MUX2_X1 U10019 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8678), .S(n10077), .Z(
        P2_U3543) );
  AOI22_X1 U10020 ( .A1(n8630), .A2(n10019), .B1(n10018), .B2(n8629), .ZN(
        n8631) );
  OAI211_X1 U10021 ( .C1(n8633), .C2(n9983), .A(n8632), .B(n8631), .ZN(n8679)
         );
  MUX2_X1 U10022 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8679), .S(n10077), .Z(
        P2_U3542) );
  AOI22_X1 U10023 ( .A1(n8634), .A2(n10019), .B1(n10018), .B2(n8093), .ZN(
        n8635) );
  OAI211_X1 U10024 ( .C1(n8637), .C2(n9983), .A(n8636), .B(n8635), .ZN(n8680)
         );
  MUX2_X1 U10025 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8680), .S(n10077), .Z(
        P2_U3541) );
  AOI22_X1 U10026 ( .A1(n8639), .A2(n10019), .B1(n10018), .B2(n8638), .ZN(
        n8640) );
  OAI211_X1 U10027 ( .C1(n8642), .C2(n9983), .A(n8641), .B(n8640), .ZN(n8681)
         );
  MUX2_X1 U10028 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8681), .S(n10077), .Z(
        P2_U3540) );
  AOI211_X1 U10029 ( .C1(n10018), .C2(n8645), .A(n8644), .B(n8643), .ZN(n8646)
         );
  OAI21_X1 U10030 ( .B1(n9983), .B2(n8647), .A(n8646), .ZN(n8682) );
  MUX2_X1 U10031 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8682), .S(n10077), .Z(
        P2_U3539) );
  INV_X1 U10032 ( .A(n8648), .ZN(n8652) );
  AOI22_X1 U10033 ( .A1(n8650), .A2(n10019), .B1(n10018), .B2(n8649), .ZN(
        n8651) );
  OAI211_X1 U10034 ( .C1(n8653), .C2(n9983), .A(n8652), .B(n8651), .ZN(n8683)
         );
  MUX2_X1 U10035 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8683), .S(n10077), .Z(
        P2_U3538) );
  AOI211_X1 U10036 ( .C1(n10018), .C2(n8656), .A(n8655), .B(n8654), .ZN(n8657)
         );
  OAI21_X1 U10037 ( .B1(n8658), .B2(n9983), .A(n8657), .ZN(n8684) );
  MUX2_X1 U10038 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8684), .S(n10077), .Z(
        P2_U3537) );
  INV_X1 U10039 ( .A(n8659), .ZN(n8664) );
  AOI22_X1 U10040 ( .A1(n8661), .A2(n10019), .B1(n10018), .B2(n8660), .ZN(
        n8662) );
  OAI211_X1 U10041 ( .C1(n9551), .C2(n8664), .A(n8663), .B(n8662), .ZN(n8685)
         );
  MUX2_X1 U10042 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8685), .S(n10077), .Z(
        P2_U3536) );
  AOI22_X1 U10043 ( .A1(n8666), .A2(n10019), .B1(n10018), .B2(n8665), .ZN(
        n8667) );
  OAI211_X1 U10044 ( .C1(n8669), .C2(n9983), .A(n8668), .B(n8667), .ZN(n8686)
         );
  MUX2_X1 U10045 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8686), .S(n10077), .Z(
        P2_U3535) );
  MUX2_X1 U10046 ( .A(n7583), .B(n8670), .S(n10057), .Z(n8671) );
  INV_X1 U10047 ( .A(n8671), .ZN(P2_U3518) );
  MUX2_X1 U10048 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8672), .S(n10057), .Z(
        P2_U3517) );
  MUX2_X1 U10049 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8673), .S(n10057), .Z(
        P2_U3516) );
  MUX2_X1 U10050 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8674), .S(n10057), .Z(
        P2_U3515) );
  MUX2_X1 U10051 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8675), .S(n10057), .Z(
        P2_U3514) );
  MUX2_X1 U10052 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8676), .S(n10057), .Z(
        P2_U3513) );
  MUX2_X1 U10053 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8677), .S(n10057), .Z(
        P2_U3512) );
  MUX2_X1 U10054 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8678), .S(n10057), .Z(
        P2_U3511) );
  MUX2_X1 U10055 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8679), .S(n10057), .Z(
        P2_U3510) );
  MUX2_X1 U10056 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8680), .S(n10057), .Z(
        P2_U3509) );
  MUX2_X1 U10057 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8681), .S(n10057), .Z(
        P2_U3508) );
  MUX2_X1 U10058 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8682), .S(n10057), .Z(
        P2_U3507) );
  MUX2_X1 U10059 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8683), .S(n10057), .Z(
        P2_U3505) );
  MUX2_X1 U10060 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8684), .S(n10057), .Z(
        P2_U3502) );
  MUX2_X1 U10061 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8685), .S(n10057), .Z(
        P2_U3499) );
  MUX2_X1 U10062 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8686), .S(n10057), .Z(
        P2_U3496) );
  INV_X1 U10063 ( .A(n8687), .ZN(n9265) );
  NOR4_X1 U10064 ( .A1(n8688), .A2(P2_IR_REG_30__SCAN_IN), .A3(n4933), .A4(
        P2_U3152), .ZN(n8689) );
  AOI21_X1 U10065 ( .B1(n8690), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8689), .ZN(
        n8691) );
  OAI21_X1 U10066 ( .B1(n9265), .B2(n8695), .A(n8691), .ZN(P2_U3327) );
  INV_X1 U10067 ( .A(n8692), .ZN(n9269) );
  OAI222_X1 U10068 ( .A1(n8695), .A2(n9269), .B1(P2_U3152), .B2(n8694), .C1(
        n8693), .C2(n8704), .ZN(P2_U3329) );
  NAND2_X1 U10069 ( .A1(n9271), .A2(n8696), .ZN(n8698) );
  OAI211_X1 U10070 ( .C1(n8704), .C2(n8699), .A(n8698), .B(n8697), .ZN(
        P2_U3330) );
  INV_X1 U10071 ( .A(n8700), .ZN(n9278) );
  OAI222_X1 U10072 ( .A1(n8704), .A2(n8703), .B1(n8702), .B2(n9278), .C1(n8701), .C2(P2_U3152), .ZN(P2_U3331) );
  MUX2_X1 U10073 ( .A(n8705), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10074 ( .A1(n8706), .A2(n8707), .ZN(n8709) );
  XNOR2_X1 U10075 ( .A(n8709), .B(n8708), .ZN(n8714) );
  AOI22_X1 U10076 ( .A1(n8806), .A2(n9037), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8711) );
  NAND2_X1 U10077 ( .A1(n9564), .A2(n9038), .ZN(n8710) );
  OAI211_X1 U10078 ( .C1(n9580), .C2(n9043), .A(n8711), .B(n8710), .ZN(n8712)
         );
  AOI21_X1 U10079 ( .B1(n9192), .B2(n8810), .A(n8712), .ZN(n8713) );
  OAI21_X1 U10080 ( .B1(n8714), .B2(n8812), .A(n8713), .ZN(P1_U3214) );
  NAND2_X1 U10081 ( .A1(n8717), .A2(n9576), .ZN(n8721) );
  NAND2_X1 U10082 ( .A1(n9564), .A2(n9104), .ZN(n8718) );
  NAND2_X1 U10083 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8877) );
  OAI211_X1 U10084 ( .C1(n9069), .C2(n9568), .A(n8718), .B(n8877), .ZN(n8719)
         );
  AOI21_X1 U10085 ( .B1(n9097), .B2(n8798), .A(n8719), .ZN(n8720) );
  OAI211_X1 U10086 ( .C1(n9099), .C2(n8795), .A(n8721), .B(n8720), .ZN(
        P1_U3217) );
  XOR2_X1 U10087 ( .A(n8722), .B(n8723), .Z(n8729) );
  OAI22_X1 U10088 ( .A1(n9070), .A2(n9568), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8724), .ZN(n8725) );
  AOI21_X1 U10089 ( .B1(n9564), .B2(n9103), .A(n8725), .ZN(n8726) );
  OAI21_X1 U10090 ( .B1(n9580), .B2(n9072), .A(n8726), .ZN(n8727) );
  AOI21_X1 U10091 ( .B1(n9202), .B2(n8810), .A(n8727), .ZN(n8728) );
  OAI21_X1 U10092 ( .B1(n8729), .B2(n8812), .A(n8728), .ZN(P1_U3221) );
  XOR2_X1 U10093 ( .A(n8731), .B(n8730), .Z(n8736) );
  AOI22_X1 U10094 ( .A1(n8806), .A2(n9015), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8733) );
  NAND2_X1 U10095 ( .A1(n9564), .A2(n9037), .ZN(n8732) );
  OAI211_X1 U10096 ( .C1(n9580), .C2(n9007), .A(n8733), .B(n8732), .ZN(n8734)
         );
  AOI21_X1 U10097 ( .B1(n9180), .B2(n8810), .A(n8734), .ZN(n8735) );
  OAI21_X1 U10098 ( .B1(n8736), .B2(n8812), .A(n8735), .ZN(P1_U3223) );
  INV_X1 U10099 ( .A(n9227), .ZN(n9153) );
  OAI21_X1 U10100 ( .B1(n8739), .B2(n8738), .A(n8737), .ZN(n8740) );
  NAND2_X1 U10101 ( .A1(n8740), .A2(n9576), .ZN(n8745) );
  INV_X1 U10102 ( .A(n8741), .ZN(n9148) );
  AOI22_X1 U10103 ( .A1(n9564), .A2(n8909), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n8742) );
  OAI21_X1 U10104 ( .B1(n9144), .B2(n9568), .A(n8742), .ZN(n8743) );
  AOI21_X1 U10105 ( .B1(n9148), .B2(n8798), .A(n8743), .ZN(n8744) );
  OAI211_X1 U10106 ( .C1(n9153), .C2(n8795), .A(n8745), .B(n8744), .ZN(
        P1_U3224) );
  OAI21_X1 U10107 ( .B1(n8748), .B2(n8746), .A(n8747), .ZN(n8749) );
  NAND2_X1 U10108 ( .A1(n8749), .A2(n9576), .ZN(n8755) );
  AND2_X1 U10109 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9741) );
  AOI21_X1 U10110 ( .B1(n9564), .B2(n8821), .A(n9741), .ZN(n8754) );
  AOI22_X1 U10111 ( .A1(n8751), .A2(n8798), .B1(n8810), .B2(n8750), .ZN(n8753)
         );
  NAND2_X1 U10112 ( .A1(n8806), .A2(n8819), .ZN(n8752) );
  NAND4_X1 U10113 ( .A1(n8755), .A2(n8754), .A3(n8753), .A4(n8752), .ZN(
        P1_U3225) );
  INV_X1 U10114 ( .A(n9222), .ZN(n9126) );
  OAI21_X1 U10115 ( .B1(n8758), .B2(n8757), .A(n8756), .ZN(n8759) );
  NAND2_X1 U10116 ( .A1(n8759), .A2(n9576), .ZN(n8765) );
  NOR2_X1 U10117 ( .A1(n9580), .A2(n9127), .ZN(n8763) );
  OAI22_X1 U10118 ( .A1(n8761), .A2(n9584), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8760), .ZN(n8762) );
  AOI211_X1 U10119 ( .C1(n8806), .C2(n9104), .A(n8763), .B(n8762), .ZN(n8764)
         );
  OAI211_X1 U10120 ( .C1(n9126), .C2(n8795), .A(n8765), .B(n8764), .ZN(
        P1_U3226) );
  XOR2_X1 U10121 ( .A(n8767), .B(n8766), .Z(n8772) );
  AOI22_X1 U10122 ( .A1(n8806), .A2(n8998), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8769) );
  NAND2_X1 U10123 ( .A1(n9564), .A2(n8919), .ZN(n8768) );
  OAI211_X1 U10124 ( .C1(n9580), .C2(n9028), .A(n8769), .B(n8768), .ZN(n8770)
         );
  AOI21_X1 U10125 ( .B1(n9187), .B2(n8810), .A(n8770), .ZN(n8771) );
  OAI21_X1 U10126 ( .B1(n8772), .B2(n8812), .A(n8771), .ZN(P1_U3227) );
  XOR2_X1 U10127 ( .A(n8773), .B(n8774), .Z(n8780) );
  OAI22_X1 U10128 ( .A1(n9054), .A2(n9568), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8775), .ZN(n8776) );
  AOI21_X1 U10129 ( .B1(n9564), .B2(n9088), .A(n8776), .ZN(n8777) );
  OAI21_X1 U10130 ( .B1(n9580), .B2(n9081), .A(n8777), .ZN(n8778) );
  AOI21_X1 U10131 ( .B1(n9205), .B2(n8810), .A(n8778), .ZN(n8779) );
  OAI21_X1 U10132 ( .B1(n8780), .B2(n8812), .A(n8779), .ZN(P1_U3231) );
  NAND2_X1 U10133 ( .A1(n8781), .A2(n8782), .ZN(n8784) );
  XNOR2_X1 U10134 ( .A(n8784), .B(n8783), .ZN(n8789) );
  AOI22_X1 U10135 ( .A1(n8806), .A2(n8919), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8786) );
  NAND2_X1 U10136 ( .A1(n9564), .A2(n9087), .ZN(n8785) );
  OAI211_X1 U10137 ( .C1(n9580), .C2(n9057), .A(n8786), .B(n8785), .ZN(n8787)
         );
  AOI21_X1 U10138 ( .B1(n9197), .B2(n8810), .A(n8787), .ZN(n8788) );
  OAI21_X1 U10139 ( .B1(n8789), .B2(n8812), .A(n8788), .ZN(P1_U3233) );
  NAND2_X1 U10140 ( .A1(n8791), .A2(n8790), .ZN(n8792) );
  XOR2_X1 U10141 ( .A(n8793), .B(n8792), .Z(n8800) );
  NAND2_X1 U10142 ( .A1(n9564), .A2(n8913), .ZN(n8794) );
  NAND2_X1 U10143 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9786) );
  OAI211_X1 U10144 ( .C1(n9116), .C2(n9568), .A(n8794), .B(n9786), .ZN(n8797)
         );
  INV_X1 U10145 ( .A(n9217), .ZN(n9121) );
  NOR2_X1 U10146 ( .A1(n9121), .A2(n8795), .ZN(n8796) );
  AOI211_X1 U10147 ( .C1(n9118), .C2(n8798), .A(n8797), .B(n8796), .ZN(n8799)
         );
  OAI21_X1 U10148 ( .B1(n8800), .B2(n8812), .A(n8799), .ZN(P1_U3236) );
  INV_X1 U10149 ( .A(n8802), .ZN(n8804) );
  NAND2_X1 U10150 ( .A1(n8804), .A2(n8803), .ZN(n8805) );
  XNOR2_X1 U10151 ( .A(n8801), .B(n8805), .ZN(n8813) );
  AOI22_X1 U10152 ( .A1(n9564), .A2(n8998), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8808) );
  NAND2_X1 U10153 ( .A1(n8806), .A2(n8997), .ZN(n8807) );
  OAI211_X1 U10154 ( .C1(n9580), .C2(n8991), .A(n8808), .B(n8807), .ZN(n8809)
         );
  AOI21_X1 U10155 ( .B1(n9175), .B2(n8810), .A(n8809), .ZN(n8811) );
  OAI21_X1 U10156 ( .B1(n8813), .B2(n8812), .A(n8811), .ZN(P1_U3238) );
  MUX2_X1 U10157 ( .A(n8974), .B(P1_DATAO_REG_29__SCAN_IN), .S(n8826), .Z(
        P1_U3584) );
  MUX2_X1 U10158 ( .A(n8997), .B(P1_DATAO_REG_27__SCAN_IN), .S(n8824), .Z(
        P1_U3582) );
  MUX2_X1 U10159 ( .A(n9015), .B(P1_DATAO_REG_26__SCAN_IN), .S(n8826), .Z(
        P1_U3581) );
  MUX2_X1 U10160 ( .A(n8998), .B(P1_DATAO_REG_25__SCAN_IN), .S(n8824), .Z(
        P1_U3580) );
  MUX2_X1 U10161 ( .A(n9037), .B(P1_DATAO_REG_24__SCAN_IN), .S(n8824), .Z(
        P1_U3579) );
  MUX2_X1 U10162 ( .A(n8919), .B(P1_DATAO_REG_23__SCAN_IN), .S(n8826), .Z(
        P1_U3578) );
  MUX2_X1 U10163 ( .A(n9038), .B(P1_DATAO_REG_22__SCAN_IN), .S(n8824), .Z(
        P1_U3577) );
  MUX2_X1 U10164 ( .A(n9087), .B(P1_DATAO_REG_21__SCAN_IN), .S(n8824), .Z(
        P1_U3576) );
  MUX2_X1 U10165 ( .A(n9103), .B(P1_DATAO_REG_20__SCAN_IN), .S(n8826), .Z(
        P1_U3575) );
  MUX2_X1 U10166 ( .A(n9088), .B(P1_DATAO_REG_19__SCAN_IN), .S(n8826), .Z(
        P1_U3574) );
  MUX2_X1 U10167 ( .A(n9104), .B(P1_DATAO_REG_18__SCAN_IN), .S(n8824), .Z(
        P1_U3573) );
  MUX2_X1 U10168 ( .A(n8913), .B(P1_DATAO_REG_17__SCAN_IN), .S(n8826), .Z(
        P1_U3572) );
  MUX2_X1 U10169 ( .A(n8912), .B(P1_DATAO_REG_16__SCAN_IN), .S(n8824), .Z(
        P1_U3571) );
  MUX2_X1 U10170 ( .A(n8909), .B(P1_DATAO_REG_15__SCAN_IN), .S(n8824), .Z(
        P1_U3570) );
  MUX2_X1 U10171 ( .A(n9616), .B(P1_DATAO_REG_14__SCAN_IN), .S(n8824), .Z(
        P1_U3569) );
  MUX2_X1 U10172 ( .A(n8814), .B(P1_DATAO_REG_13__SCAN_IN), .S(n8824), .Z(
        P1_U3568) );
  MUX2_X1 U10173 ( .A(n9639), .B(P1_DATAO_REG_12__SCAN_IN), .S(n8824), .Z(
        P1_U3567) );
  MUX2_X1 U10174 ( .A(n8815), .B(P1_DATAO_REG_11__SCAN_IN), .S(n8826), .Z(
        P1_U3566) );
  MUX2_X1 U10175 ( .A(n9640), .B(P1_DATAO_REG_10__SCAN_IN), .S(n8824), .Z(
        P1_U3565) );
  MUX2_X1 U10176 ( .A(n8816), .B(P1_DATAO_REG_9__SCAN_IN), .S(n8826), .Z(
        P1_U3564) );
  MUX2_X1 U10177 ( .A(n8817), .B(P1_DATAO_REG_8__SCAN_IN), .S(n8826), .Z(
        P1_U3563) );
  MUX2_X1 U10178 ( .A(n8818), .B(P1_DATAO_REG_7__SCAN_IN), .S(n8826), .Z(
        P1_U3562) );
  MUX2_X1 U10179 ( .A(n8819), .B(P1_DATAO_REG_6__SCAN_IN), .S(n8826), .Z(
        P1_U3561) );
  MUX2_X1 U10180 ( .A(n8820), .B(P1_DATAO_REG_5__SCAN_IN), .S(n8826), .Z(
        P1_U3560) );
  MUX2_X1 U10181 ( .A(n8821), .B(P1_DATAO_REG_4__SCAN_IN), .S(n8824), .Z(
        P1_U3559) );
  MUX2_X1 U10182 ( .A(n8822), .B(P1_DATAO_REG_3__SCAN_IN), .S(n8826), .Z(
        P1_U3558) );
  MUX2_X1 U10183 ( .A(n8823), .B(P1_DATAO_REG_2__SCAN_IN), .S(n8826), .Z(
        P1_U3557) );
  MUX2_X1 U10184 ( .A(n8825), .B(P1_DATAO_REG_1__SCAN_IN), .S(n8824), .Z(
        P1_U3556) );
  MUX2_X1 U10185 ( .A(n8827), .B(P1_DATAO_REG_0__SCAN_IN), .S(n8826), .Z(
        P1_U3555) );
  INV_X1 U10186 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n8841) );
  NOR2_X1 U10187 ( .A1(n8829), .A2(n8828), .ZN(n8831) );
  NOR2_X1 U10188 ( .A1(n8831), .A2(n8830), .ZN(n8842) );
  XNOR2_X1 U10189 ( .A(n8842), .B(n8849), .ZN(n8832) );
  NOR2_X1 U10190 ( .A1(n5949), .A2(n8832), .ZN(n8843) );
  AOI211_X1 U10191 ( .C1(n8832), .C2(n5949), .A(n8843), .B(n9775), .ZN(n8833)
         );
  INV_X1 U10192 ( .A(n8833), .ZN(n8840) );
  AND2_X1 U10193 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9565) );
  OAI21_X1 U10194 ( .B1(n8835), .B2(P1_REG1_REG_14__SCAN_IN), .A(n8834), .ZN(
        n8848) );
  XNOR2_X1 U10195 ( .A(n8849), .B(n8848), .ZN(n8836) );
  NOR2_X1 U10196 ( .A1(n5948), .A2(n8836), .ZN(n8850) );
  AOI211_X1 U10197 ( .C1(n8836), .C2(n5948), .A(n8850), .B(n9736), .ZN(n8837)
         );
  AOI211_X1 U10198 ( .C1(n9789), .C2(n8838), .A(n9565), .B(n8837), .ZN(n8839)
         );
  OAI211_X1 U10199 ( .C1(n9802), .C2(n8841), .A(n8840), .B(n8839), .ZN(
        P1_U3256) );
  NOR2_X1 U10200 ( .A1(n8842), .A2(n8849), .ZN(n8844) );
  NAND2_X1 U10201 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n8866), .ZN(n8845) );
  OAI21_X1 U10202 ( .B1(n8866), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8845), .ZN(
        n8846) );
  AOI211_X1 U10203 ( .C1(n8847), .C2(n8846), .A(n8860), .B(n9775), .ZN(n8859)
         );
  NOR2_X1 U10204 ( .A1(n8849), .A2(n8848), .ZN(n8851) );
  NOR2_X1 U10205 ( .A1(n8851), .A2(n8850), .ZN(n8853) );
  XNOR2_X1 U10206 ( .A(n8866), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n8852) );
  NOR2_X1 U10207 ( .A1(n8853), .A2(n8852), .ZN(n8865) );
  AOI211_X1 U10208 ( .C1(n8853), .C2(n8852), .A(n8865), .B(n9736), .ZN(n8858)
         );
  INV_X1 U10209 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n8856) );
  NAND2_X1 U10210 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n8855) );
  NAND2_X1 U10211 ( .A1(n9789), .A2(n8866), .ZN(n8854) );
  OAI211_X1 U10212 ( .C1(n9802), .C2(n8856), .A(n8855), .B(n8854), .ZN(n8857)
         );
  OR3_X1 U10213 ( .A1(n8859), .A2(n8858), .A3(n8857), .ZN(P1_U3257) );
  NOR2_X1 U10214 ( .A1(n8884), .A2(n8861), .ZN(n8862) );
  AOI21_X1 U10215 ( .B1(n8861), .B2(n8884), .A(n8862), .ZN(n8863) );
  AOI211_X1 U10216 ( .C1(n8864), .C2(n8863), .A(n8878), .B(n9775), .ZN(n8875)
         );
  INV_X1 U10217 ( .A(n8884), .ZN(n8872) );
  AOI21_X1 U10218 ( .B1(n8866), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8865), .ZN(
        n8868) );
  XNOR2_X1 U10219 ( .A(n8884), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n8867) );
  NOR2_X1 U10220 ( .A1(n8868), .A2(n8867), .ZN(n8883) );
  AOI211_X1 U10221 ( .C1(n8868), .C2(n8867), .A(n8883), .B(n9736), .ZN(n8869)
         );
  INV_X1 U10222 ( .A(n8869), .ZN(n8871) );
  NAND2_X1 U10223 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n8870) );
  OAI211_X1 U10224 ( .C1(n8873), .C2(n8872), .A(n8871), .B(n8870), .ZN(n8874)
         );
  AOI211_X1 U10225 ( .C1(P1_ADDR_REG_17__SCAN_IN), .C2(n9783), .A(n8875), .B(
        n8874), .ZN(n8876) );
  INV_X1 U10226 ( .A(n8876), .ZN(P1_U3258) );
  INV_X1 U10227 ( .A(n8877), .ZN(n8892) );
  AOI21_X1 U10228 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n8884), .A(n8878), .ZN(
        n9792) );
  NAND2_X1 U10229 ( .A1(n9788), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8879) );
  OAI21_X1 U10230 ( .B1(n9788), .B2(P1_REG2_REG_18__SCAN_IN), .A(n8879), .ZN(
        n9791) );
  NOR2_X1 U10231 ( .A1(n9792), .A2(n9791), .ZN(n9790) );
  AOI21_X1 U10232 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9788), .A(n9790), .ZN(
        n8880) );
  XNOR2_X1 U10233 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n8880), .ZN(n8891) );
  INV_X1 U10234 ( .A(n8891), .ZN(n8886) );
  AOI22_X1 U10235 ( .A1(n9788), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n8882), .B2(
        n8881), .ZN(n9795) );
  AOI21_X1 U10236 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n8884), .A(n8883), .ZN(
        n9794) );
  NAND2_X1 U10237 ( .A1(n9795), .A2(n9794), .ZN(n9793) );
  OAI21_X1 U10238 ( .B1(n9788), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9793), .ZN(
        n8885) );
  XOR2_X1 U10239 ( .A(n8885), .B(P1_REG1_REG_19__SCAN_IN), .Z(n8888) );
  INV_X1 U10240 ( .A(n8887), .ZN(n8890) );
  AOI21_X1 U10241 ( .B1(n8888), .B2(n9797), .A(n9789), .ZN(n8889) );
  INV_X1 U10242 ( .A(n9595), .ZN(n9598) );
  NAND2_X1 U10243 ( .A1(n9117), .A2(n9099), .ZN(n9094) );
  NOR2_X1 U10244 ( .A1(n4326), .A2(n8901), .ZN(n8893) );
  XOR2_X1 U10245 ( .A(n9157), .B(n8893), .Z(n9159) );
  INV_X1 U10246 ( .A(P1_B_REG_SCAN_IN), .ZN(n8894) );
  NOR2_X1 U10247 ( .A1(n6355), .A2(n8894), .ZN(n8895) );
  OR2_X1 U10248 ( .A1(n9583), .A2(n8895), .ZN(n8954) );
  INV_X1 U10249 ( .A(n8954), .ZN(n8897) );
  NAND2_X1 U10250 ( .A1(n8897), .A2(n8896), .ZN(n9654) );
  NOR2_X1 U10251 ( .A1(n9647), .A2(n9654), .ZN(n8902) );
  NOR2_X1 U10252 ( .A1(n9128), .A2(n8898), .ZN(n8899) );
  AOI211_X1 U10253 ( .C1(n9157), .C2(n9651), .A(n8902), .B(n8899), .ZN(n8900)
         );
  OAI21_X1 U10254 ( .B1(n9159), .B2(n8960), .A(n8900), .ZN(P1_U3261) );
  INV_X1 U10255 ( .A(n8901), .ZN(n9655) );
  XOR2_X1 U10256 ( .A(n8901), .B(n4326), .Z(n9657) );
  NAND2_X1 U10257 ( .A1(n9657), .A2(n9631), .ZN(n8904) );
  AOI21_X1 U10258 ( .B1(n9149), .B2(P1_REG2_REG_30__SCAN_IN), .A(n8902), .ZN(
        n8903) );
  OAI211_X1 U10259 ( .C1(n9655), .C2(n9152), .A(n8904), .B(n8903), .ZN(
        P1_U3262) );
  NOR2_X1 U10260 ( .A1(n9232), .A2(n9616), .ZN(n8907) );
  NAND2_X1 U10261 ( .A1(n9587), .A2(n8910), .ZN(n8911) );
  NOR2_X1 U10262 ( .A1(n9222), .A2(n8913), .ZN(n8914) );
  NAND2_X1 U10263 ( .A1(n9210), .A2(n9088), .ZN(n8915) );
  OAI21_X1 U10264 ( .B1(n9103), .B2(n9205), .A(n9078), .ZN(n8916) );
  INV_X1 U10265 ( .A(n9205), .ZN(n9084) );
  NAND2_X1 U10266 ( .A1(n9197), .A2(n9038), .ZN(n8918) );
  INV_X1 U10267 ( .A(n9197), .ZN(n9061) );
  OAI22_X2 U10268 ( .A1(n8922), .A2(n8921), .B1(n9055), .B2(n8920), .ZN(n9020)
         );
  NOR2_X1 U10269 ( .A1(n8924), .A2(n8923), .ZN(n8925) );
  NAND2_X1 U10270 ( .A1(n8965), .A2(n8972), .ZN(n8964) );
  OAI21_X1 U10271 ( .B1(n8981), .B2(n8971), .A(n8964), .ZN(n8928) );
  XNOR2_X1 U10272 ( .A(n8928), .B(n8950), .ZN(n9160) );
  INV_X1 U10273 ( .A(n9160), .ZN(n8963) );
  AOI21_X1 U10274 ( .B1(n8931), .B2(n8930), .A(n8929), .ZN(n9582) );
  NAND2_X1 U10275 ( .A1(n9582), .A2(n9588), .ZN(n9581) );
  OAI21_X1 U10276 ( .B1(n8979), .B2(n8978), .A(n8947), .ZN(n8973) );
  AOI21_X1 U10277 ( .B1(n8973), .B2(n8949), .A(n8948), .ZN(n8952) );
  INV_X1 U10278 ( .A(n8950), .ZN(n8951) );
  OAI21_X1 U10279 ( .B1(n8966), .B2(n8955), .A(n4326), .ZN(n9161) );
  OAI22_X1 U10280 ( .A1(n9128), .A2(n8957), .B1(n8956), .B2(n9633), .ZN(n8958)
         );
  AOI21_X1 U10281 ( .B1(n9162), .B2(n9651), .A(n8958), .ZN(n8959) );
  OAI21_X1 U10282 ( .B1(n9161), .B2(n8960), .A(n8959), .ZN(n8961) );
  AOI21_X1 U10283 ( .B1(n9164), .B2(n9128), .A(n8961), .ZN(n8962) );
  OAI21_X1 U10284 ( .B1(n8963), .B2(n9156), .A(n8962), .ZN(P1_U3355) );
  OAI21_X1 U10285 ( .B1(n8965), .B2(n8972), .A(n8964), .ZN(n9169) );
  INV_X1 U10286 ( .A(n8983), .ZN(n8967) );
  AOI211_X1 U10287 ( .C1(n9166), .C2(n8967), .A(n9873), .B(n8966), .ZN(n9165)
         );
  INV_X1 U10288 ( .A(n8968), .ZN(n8969) );
  AOI22_X1 U10289 ( .A1(n9647), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n8969), .B2(
        n9593), .ZN(n8970) );
  OAI21_X1 U10290 ( .B1(n8971), .B2(n9152), .A(n8970), .ZN(n8976) );
  XNOR2_X1 U10291 ( .A(n8973), .B(n8972), .ZN(n8975) );
  XOR2_X1 U10292 ( .A(n8978), .B(n8977), .Z(n9174) );
  XNOR2_X1 U10293 ( .A(n8979), .B(n8978), .ZN(n8980) );
  OAI222_X1 U10294 ( .A1(n9585), .A2(n8982), .B1(n9583), .B2(n8981), .C1(n8980), .C2(n9643), .ZN(n9170) );
  AOI211_X1 U10295 ( .C1(n9172), .C2(n8990), .A(n9873), .B(n8983), .ZN(n9171)
         );
  NAND2_X1 U10296 ( .A1(n9171), .A2(n9147), .ZN(n8986) );
  AOI22_X1 U10297 ( .A1(n9149), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n8984), .B2(
        n9593), .ZN(n8985) );
  OAI211_X1 U10298 ( .C1(n4584), .C2(n9152), .A(n8986), .B(n8985), .ZN(n8987)
         );
  AOI21_X1 U10299 ( .B1(n9170), .B2(n9128), .A(n8987), .ZN(n8988) );
  OAI21_X1 U10300 ( .B1(n9174), .B2(n9156), .A(n8988), .ZN(P1_U3264) );
  XNOR2_X1 U10301 ( .A(n8989), .B(n8995), .ZN(n9179) );
  AOI21_X1 U10302 ( .B1(n9175), .B2(n9004), .A(n4585), .ZN(n9176) );
  INV_X1 U10303 ( .A(n9175), .ZN(n8994) );
  INV_X1 U10304 ( .A(n8991), .ZN(n8992) );
  AOI22_X1 U10305 ( .A1(n9149), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n8992), .B2(
        n9593), .ZN(n8993) );
  OAI21_X1 U10306 ( .B1(n8994), .B2(n9152), .A(n8993), .ZN(n9001) );
  XNOR2_X1 U10307 ( .A(n8996), .B(n8995), .ZN(n8999) );
  AOI222_X1 U10308 ( .A1(n9613), .A2(n8999), .B1(n8998), .B2(n9641), .C1(n8997), .C2(n9638), .ZN(n9178) );
  NOR2_X1 U10309 ( .A1(n9178), .A2(n9647), .ZN(n9000) );
  AOI211_X1 U10310 ( .C1(n9176), .C2(n9631), .A(n9001), .B(n9000), .ZN(n9002)
         );
  OAI21_X1 U10311 ( .B1(n9179), .B2(n9156), .A(n9002), .ZN(P1_U3265) );
  XOR2_X1 U10312 ( .A(n9013), .B(n9003), .Z(n9184) );
  INV_X1 U10313 ( .A(n9026), .ZN(n9006) );
  INV_X1 U10314 ( .A(n9004), .ZN(n9005) );
  AOI21_X1 U10315 ( .B1(n9180), .B2(n9006), .A(n9005), .ZN(n9181) );
  INV_X1 U10316 ( .A(n9007), .ZN(n9008) );
  AOI22_X1 U10317 ( .A1(n9149), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9008), .B2(
        n9593), .ZN(n9009) );
  OAI21_X1 U10318 ( .B1(n9010), .B2(n9152), .A(n9009), .ZN(n9018) );
  INV_X1 U10319 ( .A(n9011), .ZN(n9012) );
  NOR2_X1 U10320 ( .A1(n9021), .A2(n9012), .ZN(n9014) );
  XNOR2_X1 U10321 ( .A(n9014), .B(n9013), .ZN(n9016) );
  AOI222_X1 U10322 ( .A1(n9613), .A2(n9016), .B1(n9015), .B2(n9638), .C1(n9037), .C2(n9641), .ZN(n9183) );
  NOR2_X1 U10323 ( .A1(n9183), .A2(n9647), .ZN(n9017) );
  AOI211_X1 U10324 ( .C1(n9181), .C2(n9631), .A(n9018), .B(n9017), .ZN(n9019)
         );
  OAI21_X1 U10325 ( .B1(n9184), .B2(n9156), .A(n9019), .ZN(P1_U3266) );
  XNOR2_X1 U10326 ( .A(n9020), .B(n9023), .ZN(n9189) );
  AOI22_X1 U10327 ( .A1(n9187), .A2(n9651), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9647), .ZN(n9032) );
  AOI21_X1 U10328 ( .B1(n9023), .B2(n9022), .A(n9021), .ZN(n9024) );
  OAI222_X1 U10329 ( .A1(n9585), .A2(n9055), .B1(n9583), .B2(n9025), .C1(n9643), .C2(n9024), .ZN(n9185) );
  INV_X1 U10330 ( .A(n9041), .ZN(n9027) );
  AOI211_X1 U10331 ( .C1(n9187), .C2(n9027), .A(n9873), .B(n9026), .ZN(n9186)
         );
  INV_X1 U10332 ( .A(n9186), .ZN(n9029) );
  OAI22_X1 U10333 ( .A1(n9029), .A2(n9073), .B1(n9633), .B2(n9028), .ZN(n9030)
         );
  OAI21_X1 U10334 ( .B1(n9185), .B2(n9030), .A(n9128), .ZN(n9031) );
  OAI211_X1 U10335 ( .C1(n9189), .C2(n9156), .A(n9032), .B(n9031), .ZN(
        P1_U3267) );
  XOR2_X1 U10336 ( .A(n9035), .B(n9033), .Z(n9194) );
  AOI22_X1 U10337 ( .A1(n9192), .A2(n9651), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9149), .ZN(n9047) );
  OAI211_X1 U10338 ( .C1(n9036), .C2(n9035), .A(n9034), .B(n9613), .ZN(n9040)
         );
  AOI22_X1 U10339 ( .A1(n9038), .A2(n9641), .B1(n9638), .B2(n9037), .ZN(n9039)
         );
  NAND2_X1 U10340 ( .A1(n9040), .A2(n9039), .ZN(n9190) );
  INV_X1 U10341 ( .A(n9056), .ZN(n9042) );
  AOI211_X1 U10342 ( .C1(n9192), .C2(n9042), .A(n9873), .B(n9041), .ZN(n9191)
         );
  INV_X1 U10343 ( .A(n9191), .ZN(n9044) );
  OAI22_X1 U10344 ( .A1(n9044), .A2(n9073), .B1(n9633), .B2(n9043), .ZN(n9045)
         );
  OAI21_X1 U10345 ( .B1(n9190), .B2(n9045), .A(n9128), .ZN(n9046) );
  OAI211_X1 U10346 ( .C1(n9194), .C2(n9156), .A(n9047), .B(n9046), .ZN(
        P1_U3268) );
  XOR2_X1 U10347 ( .A(n9048), .B(n9051), .Z(n9199) );
  INV_X1 U10348 ( .A(n9065), .ZN(n9050) );
  NAND2_X1 U10349 ( .A1(n9050), .A2(n9049), .ZN(n9052) );
  XNOR2_X1 U10350 ( .A(n9052), .B(n9051), .ZN(n9053) );
  OAI222_X1 U10351 ( .A1(n9583), .A2(n9055), .B1(n9585), .B2(n9054), .C1(n9053), .C2(n9643), .ZN(n9195) );
  AOI211_X1 U10352 ( .C1(n9197), .C2(n9071), .A(n9873), .B(n9056), .ZN(n9196)
         );
  NAND2_X1 U10353 ( .A1(n9196), .A2(n9147), .ZN(n9060) );
  INV_X1 U10354 ( .A(n9057), .ZN(n9058) );
  AOI22_X1 U10355 ( .A1(n9149), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9058), .B2(
        n9593), .ZN(n9059) );
  OAI211_X1 U10356 ( .C1(n9061), .C2(n9152), .A(n9060), .B(n9059), .ZN(n9062)
         );
  AOI21_X1 U10357 ( .B1(n9195), .B2(n9128), .A(n9062), .ZN(n9063) );
  OAI21_X1 U10358 ( .B1(n9199), .B2(n9156), .A(n9063), .ZN(P1_U3269) );
  XNOR2_X1 U10359 ( .A(n9064), .B(n9067), .ZN(n9204) );
  AOI22_X1 U10360 ( .A1(n9202), .A2(n9651), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9647), .ZN(n9077) );
  AOI21_X1 U10361 ( .B1(n9067), .B2(n9066), .A(n9065), .ZN(n9068) );
  OAI222_X1 U10362 ( .A1(n9583), .A2(n9070), .B1(n9585), .B2(n9069), .C1(n9643), .C2(n9068), .ZN(n9200) );
  AOI211_X1 U10363 ( .C1(n9202), .C2(n9079), .A(n9873), .B(n4591), .ZN(n9201)
         );
  INV_X1 U10364 ( .A(n9201), .ZN(n9074) );
  OAI22_X1 U10365 ( .A1(n9074), .A2(n9073), .B1(n9633), .B2(n9072), .ZN(n9075)
         );
  OAI21_X1 U10366 ( .B1(n9200), .B2(n9075), .A(n9128), .ZN(n9076) );
  OAI211_X1 U10367 ( .C1(n9204), .C2(n9156), .A(n9077), .B(n9076), .ZN(
        P1_U3270) );
  XOR2_X1 U10368 ( .A(n9078), .B(n9085), .Z(n9209) );
  INV_X1 U10369 ( .A(n9079), .ZN(n9080) );
  AOI21_X1 U10370 ( .B1(n9205), .B2(n9094), .A(n9080), .ZN(n9206) );
  INV_X1 U10371 ( .A(n9081), .ZN(n9082) );
  AOI22_X1 U10372 ( .A1(n9149), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9082), .B2(
        n9593), .ZN(n9083) );
  OAI21_X1 U10373 ( .B1(n9084), .B2(n9152), .A(n9083), .ZN(n9091) );
  XNOR2_X1 U10374 ( .A(n9086), .B(n9085), .ZN(n9089) );
  AOI222_X1 U10375 ( .A1(n9613), .A2(n9089), .B1(n9088), .B2(n9641), .C1(n9087), .C2(n9638), .ZN(n9208) );
  NOR2_X1 U10376 ( .A1(n9208), .A2(n9647), .ZN(n9090) );
  AOI211_X1 U10377 ( .C1(n9206), .C2(n9631), .A(n9091), .B(n9090), .ZN(n9092)
         );
  OAI21_X1 U10378 ( .B1(n9209), .B2(n9156), .A(n9092), .ZN(P1_U3271) );
  XNOR2_X1 U10379 ( .A(n9093), .B(n9101), .ZN(n9214) );
  INV_X1 U10380 ( .A(n9117), .ZN(n9096) );
  INV_X1 U10381 ( .A(n9094), .ZN(n9095) );
  AOI21_X1 U10382 ( .B1(n9210), .B2(n9096), .A(n9095), .ZN(n9211) );
  AOI22_X1 U10383 ( .A1(n9149), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9097), .B2(
        n9593), .ZN(n9098) );
  OAI21_X1 U10384 ( .B1(n9099), .B2(n9152), .A(n9098), .ZN(n9107) );
  OAI21_X1 U10385 ( .B1(n9102), .B2(n9101), .A(n9100), .ZN(n9105) );
  AOI222_X1 U10386 ( .A1(n9613), .A2(n9105), .B1(n9104), .B2(n9641), .C1(n9103), .C2(n9638), .ZN(n9213) );
  NOR2_X1 U10387 ( .A1(n9213), .A2(n9647), .ZN(n9106) );
  AOI211_X1 U10388 ( .C1(n9211), .C2(n9631), .A(n9107), .B(n9106), .ZN(n9108)
         );
  OAI21_X1 U10389 ( .B1(n9156), .B2(n9214), .A(n9108), .ZN(P1_U3272) );
  XNOR2_X1 U10390 ( .A(n9109), .B(n9113), .ZN(n9219) );
  INV_X1 U10391 ( .A(n9110), .ZN(n9111) );
  AOI21_X1 U10392 ( .B1(n9132), .B2(n9112), .A(n9111), .ZN(n9114) );
  XNOR2_X1 U10393 ( .A(n9114), .B(n9113), .ZN(n9115) );
  OAI222_X1 U10394 ( .A1(n9583), .A2(n9116), .B1(n9585), .B2(n9144), .C1(n9643), .C2(n9115), .ZN(n9215) );
  AOI211_X1 U10395 ( .C1(n9217), .C2(n4588), .A(n9873), .B(n9117), .ZN(n9216)
         );
  NAND2_X1 U10396 ( .A1(n9216), .A2(n9147), .ZN(n9120) );
  AOI22_X1 U10397 ( .A1(n9149), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9118), .B2(
        n9593), .ZN(n9119) );
  OAI211_X1 U10398 ( .C1(n9121), .C2(n9152), .A(n9120), .B(n9119), .ZN(n9122)
         );
  AOI21_X1 U10399 ( .B1(n9215), .B2(n9128), .A(n9122), .ZN(n9123) );
  OAI21_X1 U10400 ( .B1(n9219), .B2(n9156), .A(n9123), .ZN(P1_U3273) );
  XNOR2_X1 U10401 ( .A(n9124), .B(n9131), .ZN(n9224) );
  AOI211_X1 U10402 ( .C1(n9222), .C2(n9145), .A(n9873), .B(n9125), .ZN(n9221)
         );
  NOR2_X1 U10403 ( .A1(n9126), .A2(n9152), .ZN(n9130) );
  OAI22_X1 U10404 ( .A1(n9128), .A2(n8861), .B1(n9127), .B2(n9633), .ZN(n9129)
         );
  AOI211_X1 U10405 ( .C1(n9221), .C2(n9147), .A(n9130), .B(n9129), .ZN(n9136)
         );
  XNOR2_X1 U10406 ( .A(n9132), .B(n9131), .ZN(n9133) );
  OAI222_X1 U10407 ( .A1(n9583), .A2(n9134), .B1(n9585), .B2(n9584), .C1(n9133), .C2(n9643), .ZN(n9220) );
  NAND2_X1 U10408 ( .A1(n9220), .A2(n9128), .ZN(n9135) );
  OAI211_X1 U10409 ( .C1(n9224), .C2(n9156), .A(n9136), .B(n9135), .ZN(
        P1_U3274) );
  XNOR2_X1 U10410 ( .A(n9138), .B(n9137), .ZN(n9229) );
  NOR2_X1 U10411 ( .A1(n4842), .A2(n9139), .ZN(n9141) );
  AOI21_X1 U10412 ( .B1(n9141), .B2(n9581), .A(n9140), .ZN(n9142) );
  OAI222_X1 U10413 ( .A1(n9583), .A2(n9144), .B1(n9585), .B2(n9143), .C1(n9643), .C2(n9142), .ZN(n9225) );
  INV_X1 U10414 ( .A(n9145), .ZN(n9146) );
  AOI211_X1 U10415 ( .C1(n9227), .C2(n9597), .A(n9873), .B(n9146), .ZN(n9226)
         );
  NAND2_X1 U10416 ( .A1(n9226), .A2(n9147), .ZN(n9151) );
  AOI22_X1 U10417 ( .A1(n9149), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9148), .B2(
        n9593), .ZN(n9150) );
  OAI211_X1 U10418 ( .C1(n9153), .C2(n9152), .A(n9151), .B(n9150), .ZN(n9154)
         );
  AOI21_X1 U10419 ( .B1(n9225), .B2(n9128), .A(n9154), .ZN(n9155) );
  OAI21_X1 U10420 ( .B1(n9229), .B2(n9156), .A(n9155), .ZN(P1_U3275) );
  NAND2_X1 U10421 ( .A1(n9157), .A2(n9563), .ZN(n9158) );
  OAI211_X1 U10422 ( .C1(n9159), .C2(n9873), .A(n9654), .B(n9158), .ZN(n9243)
         );
  MUX2_X1 U10423 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9243), .S(n9888), .Z(
        P1_U3554) );
  MUX2_X1 U10424 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9244), .S(n9888), .Z(
        P1_U3552) );
  AOI21_X1 U10425 ( .B1(n9563), .B2(n9166), .A(n9165), .ZN(n9167) );
  OAI211_X1 U10426 ( .C1(n9169), .C2(n9240), .A(n9168), .B(n9167), .ZN(n9245)
         );
  MUX2_X1 U10427 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9245), .S(n9888), .Z(
        P1_U3551) );
  AOI211_X1 U10428 ( .C1(n9563), .C2(n9172), .A(n9171), .B(n9170), .ZN(n9173)
         );
  OAI21_X1 U10429 ( .B1(n9174), .B2(n9240), .A(n9173), .ZN(n9246) );
  MUX2_X1 U10430 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9246), .S(n9888), .Z(
        P1_U3550) );
  AOI22_X1 U10431 ( .A1(n9176), .A2(n9860), .B1(n9563), .B2(n9175), .ZN(n9177)
         );
  OAI211_X1 U10432 ( .C1(n9179), .C2(n9240), .A(n9178), .B(n9177), .ZN(n9247)
         );
  MUX2_X1 U10433 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9247), .S(n9888), .Z(
        P1_U3549) );
  AOI22_X1 U10434 ( .A1(n9181), .A2(n9860), .B1(n9563), .B2(n9180), .ZN(n9182)
         );
  OAI211_X1 U10435 ( .C1(n9184), .C2(n9240), .A(n9183), .B(n9182), .ZN(n9248)
         );
  MUX2_X1 U10436 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9248), .S(n9888), .Z(
        P1_U3548) );
  AOI211_X1 U10437 ( .C1(n9563), .C2(n9187), .A(n9186), .B(n9185), .ZN(n9188)
         );
  OAI21_X1 U10438 ( .B1(n9189), .B2(n9240), .A(n9188), .ZN(n9249) );
  MUX2_X1 U10439 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9249), .S(n9888), .Z(
        P1_U3547) );
  AOI211_X1 U10440 ( .C1(n9563), .C2(n9192), .A(n9191), .B(n9190), .ZN(n9193)
         );
  OAI21_X1 U10441 ( .B1(n9194), .B2(n9240), .A(n9193), .ZN(n9250) );
  MUX2_X1 U10442 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9250), .S(n9888), .Z(
        P1_U3546) );
  AOI211_X1 U10443 ( .C1(n9563), .C2(n9197), .A(n9196), .B(n9195), .ZN(n9198)
         );
  OAI21_X1 U10444 ( .B1(n9199), .B2(n9240), .A(n9198), .ZN(n9251) );
  MUX2_X1 U10445 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9251), .S(n9888), .Z(
        P1_U3545) );
  AOI211_X1 U10446 ( .C1(n9563), .C2(n9202), .A(n9201), .B(n9200), .ZN(n9203)
         );
  OAI21_X1 U10447 ( .B1(n9204), .B2(n9240), .A(n9203), .ZN(n9252) );
  MUX2_X1 U10448 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9252), .S(n9888), .Z(
        P1_U3544) );
  AOI22_X1 U10449 ( .A1(n9206), .A2(n9860), .B1(n9563), .B2(n9205), .ZN(n9207)
         );
  OAI211_X1 U10450 ( .C1(n9209), .C2(n9240), .A(n9208), .B(n9207), .ZN(n9253)
         );
  MUX2_X1 U10451 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9253), .S(n9888), .Z(
        P1_U3543) );
  AOI22_X1 U10452 ( .A1(n9211), .A2(n9860), .B1(n9563), .B2(n9210), .ZN(n9212)
         );
  OAI211_X1 U10453 ( .C1(n9214), .C2(n9240), .A(n9213), .B(n9212), .ZN(n9254)
         );
  MUX2_X1 U10454 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9254), .S(n9888), .Z(
        P1_U3542) );
  AOI211_X1 U10455 ( .C1(n9563), .C2(n9217), .A(n9216), .B(n9215), .ZN(n9218)
         );
  OAI21_X1 U10456 ( .B1(n9219), .B2(n9240), .A(n9218), .ZN(n9255) );
  MUX2_X1 U10457 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9255), .S(n9888), .Z(
        P1_U3541) );
  AOI211_X1 U10458 ( .C1(n9563), .C2(n9222), .A(n9221), .B(n9220), .ZN(n9223)
         );
  OAI21_X1 U10459 ( .B1(n9224), .B2(n9240), .A(n9223), .ZN(n9256) );
  MUX2_X1 U10460 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9256), .S(n9888), .Z(
        P1_U3540) );
  AOI211_X1 U10461 ( .C1(n9563), .C2(n9227), .A(n9226), .B(n9225), .ZN(n9228)
         );
  OAI21_X1 U10462 ( .B1(n9240), .B2(n9229), .A(n9228), .ZN(n9257) );
  MUX2_X1 U10463 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9257), .S(n9888), .Z(
        P1_U3539) );
  AOI211_X1 U10464 ( .C1(n9563), .C2(n9232), .A(n9231), .B(n9230), .ZN(n9233)
         );
  OAI21_X1 U10465 ( .B1(n9240), .B2(n9234), .A(n9233), .ZN(n9258) );
  MUX2_X1 U10466 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9258), .S(n9888), .Z(
        P1_U3537) );
  AOI211_X1 U10467 ( .C1(n9563), .C2(n9237), .A(n9236), .B(n9235), .ZN(n9238)
         );
  OAI21_X1 U10468 ( .B1(n9240), .B2(n9239), .A(n9238), .ZN(n9259) );
  MUX2_X1 U10469 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9259), .S(n9888), .Z(
        P1_U3535) );
  MUX2_X1 U10470 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9241), .S(n9888), .Z(
        P1_U3524) );
  MUX2_X1 U10471 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9242), .S(n9888), .Z(
        P1_U3523) );
  MUX2_X1 U10472 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9243), .S(n9879), .Z(
        P1_U3522) );
  MUX2_X1 U10473 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9244), .S(n9879), .Z(
        P1_U3520) );
  MUX2_X1 U10474 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9245), .S(n9879), .Z(
        P1_U3519) );
  MUX2_X1 U10475 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9246), .S(n9879), .Z(
        P1_U3518) );
  MUX2_X1 U10476 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9247), .S(n9879), .Z(
        P1_U3517) );
  MUX2_X1 U10477 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9248), .S(n9879), .Z(
        P1_U3516) );
  MUX2_X1 U10478 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9249), .S(n9879), .Z(
        P1_U3515) );
  MUX2_X1 U10479 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9250), .S(n9879), .Z(
        P1_U3514) );
  MUX2_X1 U10480 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9251), .S(n9879), .Z(
        P1_U3513) );
  MUX2_X1 U10481 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9252), .S(n9879), .Z(
        P1_U3512) );
  MUX2_X1 U10482 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9253), .S(n9879), .Z(
        P1_U3511) );
  MUX2_X1 U10483 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9254), .S(n9879), .Z(
        P1_U3510) );
  MUX2_X1 U10484 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9255), .S(n9879), .Z(
        P1_U3508) );
  MUX2_X1 U10485 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9256), .S(n9879), .Z(
        P1_U3505) );
  MUX2_X1 U10486 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9257), .S(n9879), .Z(
        P1_U3502) );
  MUX2_X1 U10487 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9258), .S(n9879), .Z(
        P1_U3496) );
  MUX2_X1 U10488 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9259), .S(n9879), .Z(
        P1_U3490) );
  NAND3_X1 U10489 ( .A1(n9260), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9261) );
  OAI22_X1 U10490 ( .A1(n9262), .A2(n9261), .B1(n6332), .B2(n4314), .ZN(n9263)
         );
  INV_X1 U10491 ( .A(n9263), .ZN(n9264) );
  OAI21_X1 U10492 ( .B1(n9265), .B2(n9277), .A(n9264), .ZN(P1_U3322) );
  OAI222_X1 U10493 ( .A1(n9277), .A2(n9269), .B1(n9268), .B2(P1_U3084), .C1(
        n9267), .C2(n4314), .ZN(P1_U3324) );
  NAND2_X1 U10494 ( .A1(n9271), .A2(n9270), .ZN(n9272) );
  OAI211_X1 U10495 ( .C1(n4314), .C2(n9273), .A(n9272), .B(n9688), .ZN(
        P1_U3325) );
  AOI21_X1 U10496 ( .B1(n4313), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n9274), .ZN(
        n9276) );
  OAI21_X1 U10497 ( .B1(n9278), .B2(n9277), .A(n9276), .ZN(P1_U3326) );
  INV_X1 U10498 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10115) );
  NOR2_X1 U10499 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9279) );
  AOI21_X1 U10500 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9279), .ZN(n10084) );
  NOR2_X1 U10501 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9280) );
  AOI21_X1 U10502 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9280), .ZN(n10087) );
  NOR2_X1 U10503 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9281) );
  AOI21_X1 U10504 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9281), .ZN(n10090) );
  NOR2_X1 U10505 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9282) );
  AOI21_X1 U10506 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9282), .ZN(n10093) );
  NOR2_X1 U10507 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9283) );
  AOI21_X1 U10508 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9283), .ZN(n10096) );
  INV_X1 U10509 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10123) );
  NOR2_X1 U10510 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9290) );
  XNOR2_X1 U10511 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10128) );
  NAND2_X1 U10512 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9288) );
  XOR2_X1 U10513 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10126) );
  NAND2_X1 U10514 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9286) );
  XOR2_X1 U10515 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10110) );
  AOI21_X1 U10516 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10078) );
  INV_X1 U10517 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9284) );
  NAND3_X1 U10518 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10080) );
  OAI21_X1 U10519 ( .B1(n10078), .B2(n9284), .A(n10080), .ZN(n10109) );
  NAND2_X1 U10520 ( .A1(n10110), .A2(n10109), .ZN(n9285) );
  NAND2_X1 U10521 ( .A1(n9286), .A2(n9285), .ZN(n10125) );
  NAND2_X1 U10522 ( .A1(n10126), .A2(n10125), .ZN(n9287) );
  NAND2_X1 U10523 ( .A1(n9288), .A2(n9287), .ZN(n10127) );
  NOR2_X1 U10524 ( .A1(n10128), .A2(n10127), .ZN(n9289) );
  NAND2_X1 U10525 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10122), .ZN(n9291) );
  NOR2_X1 U10526 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10122), .ZN(n10121) );
  AOI21_X1 U10527 ( .B1(n10123), .B2(n9291), .A(n10121), .ZN(n9292) );
  NAND2_X1 U10528 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n9292), .ZN(n9294) );
  XOR2_X1 U10529 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n9292), .Z(n10120) );
  NAND2_X1 U10530 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10120), .ZN(n9293) );
  NAND2_X1 U10531 ( .A1(n9294), .A2(n9293), .ZN(n9295) );
  NAND2_X1 U10532 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9295), .ZN(n9297) );
  XOR2_X1 U10533 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9295), .Z(n10118) );
  NAND2_X1 U10534 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10118), .ZN(n9296) );
  NAND2_X1 U10535 ( .A1(n9297), .A2(n9296), .ZN(n9298) );
  NAND2_X1 U10536 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9298), .ZN(n9300) );
  XOR2_X1 U10537 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9298), .Z(n10112) );
  NAND2_X1 U10538 ( .A1(n10112), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n9299) );
  NAND2_X1 U10539 ( .A1(n9300), .A2(n9299), .ZN(n9301) );
  AND2_X1 U10540 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9301), .ZN(n9302) );
  XNOR2_X1 U10541 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9301), .ZN(n10108) );
  INV_X1 U10542 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10107) );
  NOR2_X1 U10543 ( .A1(n10108), .A2(n10107), .ZN(n10106) );
  NAND2_X1 U10544 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9303) );
  OAI21_X1 U10545 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9303), .ZN(n10104) );
  AOI21_X1 U10546 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10103), .ZN(n10102) );
  NAND2_X1 U10547 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9304) );
  OAI21_X1 U10548 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9304), .ZN(n10101) );
  NOR2_X1 U10549 ( .A1(n10102), .A2(n10101), .ZN(n10100) );
  AOI21_X1 U10550 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10100), .ZN(n10099) );
  NOR2_X1 U10551 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9305) );
  AOI21_X1 U10552 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9305), .ZN(n10098) );
  NAND2_X1 U10553 ( .A1(n10099), .A2(n10098), .ZN(n10097) );
  OAI21_X1 U10554 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10097), .ZN(n10095) );
  NAND2_X1 U10555 ( .A1(n10096), .A2(n10095), .ZN(n10094) );
  OAI21_X1 U10556 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10094), .ZN(n10092) );
  NAND2_X1 U10557 ( .A1(n10093), .A2(n10092), .ZN(n10091) );
  OAI21_X1 U10558 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10091), .ZN(n10089) );
  NAND2_X1 U10559 ( .A1(n10090), .A2(n10089), .ZN(n10088) );
  OAI21_X1 U10560 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10088), .ZN(n10086) );
  NAND2_X1 U10561 ( .A1(n10087), .A2(n10086), .ZN(n10085) );
  OAI21_X1 U10562 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10085), .ZN(n10083) );
  NAND2_X1 U10563 ( .A1(n10084), .A2(n10083), .ZN(n10082) );
  OAI21_X1 U10564 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10082), .ZN(n10114) );
  NOR2_X1 U10565 ( .A1(n10115), .A2(n10114), .ZN(n9306) );
  NAND2_X1 U10566 ( .A1(n10115), .A2(n10114), .ZN(n10113) );
  OAI21_X1 U10567 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n9306), .A(n10113), .ZN(
        n9499) );
  AOI22_X1 U10568 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_f55), .B1(
        SI_12_), .B2(keyinput_f20), .ZN(n9307) );
  OAI221_X1 U10569 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .C1(
        SI_12_), .C2(keyinput_f20), .A(n9307), .ZN(n9314) );
  AOI22_X1 U10570 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_f59), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n9308) );
  OAI221_X1 U10571 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_f59), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n9308), .ZN(n9313) );
  AOI22_X1 U10572 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_f39), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(keyinput_f56), .ZN(n9309) );
  OAI221_X1 U10573 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_f56), .A(n9309), .ZN(n9312) );
  AOI22_X1 U10574 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_f38), .B1(SI_2_), .B2(keyinput_f30), .ZN(n9310) );
  OAI221_X1 U10575 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .C1(
        SI_2_), .C2(keyinput_f30), .A(n9310), .ZN(n9311) );
  NOR4_X1 U10576 ( .A1(n9314), .A2(n9313), .A3(n9312), .A4(n9311), .ZN(n9341)
         );
  XOR2_X1 U10577 ( .A(SI_20_), .B(keyinput_f12), .Z(n9321) );
  AOI22_X1 U10578 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_f34), .B1(SI_9_), 
        .B2(keyinput_f23), .ZN(n9315) );
  OAI221_X1 U10579 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .C1(SI_9_), 
        .C2(keyinput_f23), .A(n9315), .ZN(n9320) );
  AOI22_X1 U10580 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_f49), .B1(SI_6_), 
        .B2(keyinput_f26), .ZN(n9316) );
  OAI221_X1 U10581 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_f49), .C1(SI_6_), .C2(keyinput_f26), .A(n9316), .ZN(n9319) );
  AOI22_X1 U10582 ( .A1(SI_30_), .A2(keyinput_f2), .B1(SI_27_), .B2(
        keyinput_f5), .ZN(n9317) );
  OAI221_X1 U10583 ( .B1(SI_30_), .B2(keyinput_f2), .C1(SI_27_), .C2(
        keyinput_f5), .A(n9317), .ZN(n9318) );
  NOR4_X1 U10584 ( .A1(n9321), .A2(n9320), .A3(n9319), .A4(n9318), .ZN(n9340)
         );
  AOI22_X1 U10585 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_f62), .B1(
        SI_23_), .B2(keyinput_f9), .ZN(n9322) );
  OAI221_X1 U10586 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .C1(
        SI_23_), .C2(keyinput_f9), .A(n9322), .ZN(n9329) );
  AOI22_X1 U10587 ( .A1(SI_31_), .A2(keyinput_f1), .B1(SI_19_), .B2(
        keyinput_f13), .ZN(n9323) );
  OAI221_X1 U10588 ( .B1(SI_31_), .B2(keyinput_f1), .C1(SI_19_), .C2(
        keyinput_f13), .A(n9323), .ZN(n9328) );
  AOI22_X1 U10589 ( .A1(n9422), .A2(keyinput_f54), .B1(n9425), .B2(
        keyinput_f52), .ZN(n9324) );
  OAI221_X1 U10590 ( .B1(n9422), .B2(keyinput_f54), .C1(n9425), .C2(
        keyinput_f52), .A(n9324), .ZN(n9327) );
  AOI22_X1 U10591 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_f43), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput_f37), .ZN(n9325) );
  OAI221_X1 U10592 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_f37), .A(n9325), .ZN(n9326) );
  NOR4_X1 U10593 ( .A1(n9329), .A2(n9328), .A3(n9327), .A4(n9326), .ZN(n9339)
         );
  AOI22_X1 U10594 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_f42), .B1(
        SI_17_), .B2(keyinput_f15), .ZN(n9330) );
  OAI221_X1 U10595 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .C1(
        SI_17_), .C2(keyinput_f15), .A(n9330), .ZN(n9337) );
  AOI22_X1 U10596 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(SI_26_), .B2(keyinput_f6), .ZN(n9331) );
  OAI221_X1 U10597 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        SI_26_), .C2(keyinput_f6), .A(n9331), .ZN(n9336) );
  AOI22_X1 U10598 ( .A1(SI_28_), .A2(keyinput_f4), .B1(SI_5_), .B2(
        keyinput_f27), .ZN(n9332) );
  OAI221_X1 U10599 ( .B1(SI_28_), .B2(keyinput_f4), .C1(SI_5_), .C2(
        keyinput_f27), .A(n9332), .ZN(n9335) );
  AOI22_X1 U10600 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_f57), .B1(
        P2_RD_REG_SCAN_IN), .B2(keyinput_f33), .ZN(n9333) );
  OAI221_X1 U10601 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput_f33), .A(n9333), .ZN(n9334) );
  NOR4_X1 U10602 ( .A1(n9337), .A2(n9336), .A3(n9335), .A4(n9334), .ZN(n9338)
         );
  NAND4_X1 U10603 ( .A1(n9341), .A2(n9340), .A3(n9339), .A4(n9338), .ZN(n9389)
         );
  INV_X1 U10604 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9419) );
  AOI22_X1 U10605 ( .A1(n9419), .A2(keyinput_f0), .B1(n9410), .B2(keyinput_f35), .ZN(n9342) );
  OAI221_X1 U10606 ( .B1(n9419), .B2(keyinput_f0), .C1(n9410), .C2(
        keyinput_f35), .A(n9342), .ZN(n9350) );
  AOI22_X1 U10607 ( .A1(n9428), .A2(keyinput_f17), .B1(n9395), .B2(
        keyinput_f16), .ZN(n9343) );
  OAI221_X1 U10608 ( .B1(n9428), .B2(keyinput_f17), .C1(n9395), .C2(
        keyinput_f16), .A(n9343), .ZN(n9349) );
  AOI22_X1 U10609 ( .A1(n9468), .A2(keyinput_f10), .B1(keyinput_f48), .B2(
        n7422), .ZN(n9344) );
  OAI221_X1 U10610 ( .B1(n9468), .B2(keyinput_f10), .C1(n7422), .C2(
        keyinput_f48), .A(n9344), .ZN(n9348) );
  AOI22_X1 U10611 ( .A1(n9408), .A2(keyinput_f45), .B1(n9346), .B2(
        keyinput_f51), .ZN(n9345) );
  OAI221_X1 U10612 ( .B1(n9408), .B2(keyinput_f45), .C1(n9346), .C2(
        keyinput_f51), .A(n9345), .ZN(n9347) );
  NOR4_X1 U10613 ( .A1(n9350), .A2(n9349), .A3(n9348), .A4(n9347), .ZN(n9387)
         );
  INV_X1 U10614 ( .A(SI_4_), .ZN(n9472) );
  AOI22_X1 U10615 ( .A1(n5231), .A2(keyinput_f58), .B1(n9472), .B2(
        keyinput_f28), .ZN(n9351) );
  OAI221_X1 U10616 ( .B1(n5231), .B2(keyinput_f58), .C1(n9472), .C2(
        keyinput_f28), .A(n9351), .ZN(n9359) );
  INV_X1 U10617 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9475) );
  AOI22_X1 U10618 ( .A1(n9475), .A2(keyinput_f61), .B1(n5445), .B2(keyinput_f8), .ZN(n9352) );
  OAI221_X1 U10619 ( .B1(n9475), .B2(keyinput_f61), .C1(n5445), .C2(
        keyinput_f8), .A(n9352), .ZN(n9358) );
  AOI22_X1 U10620 ( .A1(n9354), .A2(keyinput_f22), .B1(keyinput_f41), .B2(
        n5357), .ZN(n9353) );
  OAI221_X1 U10621 ( .B1(n9354), .B2(keyinput_f22), .C1(n5357), .C2(
        keyinput_f41), .A(n9353), .ZN(n9357) );
  AOI22_X1 U10622 ( .A1(n5005), .A2(keyinput_f21), .B1(keyinput_f47), .B2(
        n8207), .ZN(n9355) );
  OAI221_X1 U10623 ( .B1(n5005), .B2(keyinput_f21), .C1(n8207), .C2(
        keyinput_f47), .A(n9355), .ZN(n9356) );
  NOR4_X1 U10624 ( .A1(n9359), .A2(n9358), .A3(n9357), .A4(n9356), .ZN(n9386)
         );
  AOI22_X1 U10625 ( .A1(n9362), .A2(keyinput_f3), .B1(n9361), .B2(keyinput_f19), .ZN(n9360) );
  OAI221_X1 U10626 ( .B1(n9362), .B2(keyinput_f3), .C1(n9361), .C2(
        keyinput_f19), .A(n9360), .ZN(n9372) );
  AOI22_X1 U10627 ( .A1(n5020), .A2(keyinput_f18), .B1(keyinput_f24), .B2(
        n9364), .ZN(n9363) );
  OAI221_X1 U10628 ( .B1(n5020), .B2(keyinput_f18), .C1(n9364), .C2(
        keyinput_f24), .A(n9363), .ZN(n9371) );
  INV_X1 U10629 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9366) );
  AOI22_X1 U10630 ( .A1(n9366), .A2(keyinput_f53), .B1(n9437), .B2(
        keyinput_f31), .ZN(n9365) );
  OAI221_X1 U10631 ( .B1(n9366), .B2(keyinput_f53), .C1(n9437), .C2(
        keyinput_f31), .A(n9365), .ZN(n9370) );
  AOI22_X1 U10632 ( .A1(n9393), .A2(keyinput_f7), .B1(keyinput_f40), .B2(n9368), .ZN(n9367) );
  OAI221_X1 U10633 ( .B1(n9393), .B2(keyinput_f7), .C1(n9368), .C2(
        keyinput_f40), .A(n9367), .ZN(n9369) );
  NOR4_X1 U10634 ( .A1(n9372), .A2(n9371), .A3(n9370), .A4(n9369), .ZN(n9385)
         );
  AOI22_X1 U10635 ( .A1(n9374), .A2(keyinput_f46), .B1(n9435), .B2(
        keyinput_f50), .ZN(n9373) );
  OAI221_X1 U10636 ( .B1(n9374), .B2(keyinput_f46), .C1(n9435), .C2(
        keyinput_f50), .A(n9373), .ZN(n9383) );
  INV_X1 U10637 ( .A(SI_7_), .ZN(n9399) );
  AOI22_X1 U10638 ( .A1(n9399), .A2(keyinput_f25), .B1(keyinput_f60), .B2(
        n9473), .ZN(n9375) );
  OAI221_X1 U10639 ( .B1(n9399), .B2(keyinput_f25), .C1(n9473), .C2(
        keyinput_f60), .A(n9375), .ZN(n9382) );
  INV_X1 U10640 ( .A(SI_3_), .ZN(n9407) );
  INV_X1 U10641 ( .A(SI_18_), .ZN(n9377) );
  AOI22_X1 U10642 ( .A1(n9407), .A2(keyinput_f29), .B1(n9377), .B2(
        keyinput_f14), .ZN(n9376) );
  OAI221_X1 U10643 ( .B1(n9407), .B2(keyinput_f29), .C1(n9377), .C2(
        keyinput_f14), .A(n9376), .ZN(n9381) );
  XNOR2_X1 U10644 ( .A(SI_0_), .B(keyinput_f32), .ZN(n9379) );
  XNOR2_X1 U10645 ( .A(SI_21_), .B(keyinput_f11), .ZN(n9378) );
  NAND2_X1 U10646 ( .A1(n9379), .A2(n9378), .ZN(n9380) );
  NOR4_X1 U10647 ( .A1(n9383), .A2(n9382), .A3(n9381), .A4(n9380), .ZN(n9384)
         );
  NAND4_X1 U10648 ( .A1(n9387), .A2(n9386), .A3(n9385), .A4(n9384), .ZN(n9388)
         );
  OAI22_X1 U10649 ( .A1(n9389), .A2(n9388), .B1(keyinput_f63), .B2(
        P2_REG3_REG_15__SCAN_IN), .ZN(n9390) );
  AOI21_X1 U10650 ( .B1(keyinput_f63), .B2(P2_REG3_REG_15__SCAN_IN), .A(n9390), 
        .ZN(n9496) );
  AOI22_X1 U10651 ( .A1(n9393), .A2(keyinput_g7), .B1(keyinput_g57), .B2(n9392), .ZN(n9391) );
  OAI221_X1 U10652 ( .B1(n9393), .B2(keyinput_g7), .C1(n9392), .C2(
        keyinput_g57), .A(n9391), .ZN(n9403) );
  AOI22_X1 U10653 ( .A1(n9395), .A2(keyinput_g16), .B1(n5445), .B2(keyinput_g8), .ZN(n9394) );
  OAI221_X1 U10654 ( .B1(n9395), .B2(keyinput_g16), .C1(n5445), .C2(
        keyinput_g8), .A(n9394), .ZN(n9402) );
  AOI22_X1 U10655 ( .A1(n5034), .A2(keyinput_g15), .B1(keyinput_g59), .B2(
        n5075), .ZN(n9396) );
  OAI221_X1 U10656 ( .B1(n5034), .B2(keyinput_g15), .C1(n5075), .C2(
        keyinput_g59), .A(n9396), .ZN(n9401) );
  AOI22_X1 U10657 ( .A1(n9399), .A2(keyinput_g25), .B1(keyinput_g44), .B2(
        n9398), .ZN(n9397) );
  OAI221_X1 U10658 ( .B1(n9399), .B2(keyinput_g25), .C1(n9398), .C2(
        keyinput_g44), .A(n9397), .ZN(n9400) );
  NOR4_X1 U10659 ( .A1(n9403), .A2(n9402), .A3(n9401), .A4(n9400), .ZN(n9451)
         );
  AOI22_X1 U10660 ( .A1(n7590), .A2(keyinput_g1), .B1(n9405), .B2(keyinput_g55), .ZN(n9404) );
  OAI221_X1 U10661 ( .B1(n7590), .B2(keyinput_g1), .C1(n9405), .C2(
        keyinput_g55), .A(n9404), .ZN(n9417) );
  AOI22_X1 U10662 ( .A1(n9408), .A2(keyinput_g45), .B1(n9407), .B2(
        keyinput_g29), .ZN(n9406) );
  OAI221_X1 U10663 ( .B1(n9408), .B2(keyinput_g45), .C1(n9407), .C2(
        keyinput_g29), .A(n9406), .ZN(n9416) );
  AOI22_X1 U10664 ( .A1(n9410), .A2(keyinput_g35), .B1(n5588), .B2(
        keyinput_g42), .ZN(n9409) );
  OAI221_X1 U10665 ( .B1(n9410), .B2(keyinput_g35), .C1(n5588), .C2(
        keyinput_g42), .A(n9409), .ZN(n9415) );
  AOI22_X1 U10666 ( .A1(P2_U3152), .A2(keyinput_g34), .B1(n9412), .B2(
        keyinput_g6), .ZN(n9411) );
  OAI221_X1 U10667 ( .B1(P2_U3152), .B2(keyinput_g34), .C1(n9412), .C2(
        keyinput_g6), .A(n9411), .ZN(n9414) );
  NOR4_X1 U10668 ( .A1(n9417), .A2(n9416), .A3(n9415), .A4(n9414), .ZN(n9450)
         );
  AOI22_X1 U10669 ( .A1(n9420), .A2(keyinput_g5), .B1(keyinput_g0), .B2(n9419), 
        .ZN(n9418) );
  OAI221_X1 U10670 ( .B1(n9420), .B2(keyinput_g5), .C1(n9419), .C2(keyinput_g0), .A(n9418), .ZN(n9432) );
  AOI22_X1 U10671 ( .A1(n9423), .A2(keyinput_g9), .B1(keyinput_g54), .B2(n9422), .ZN(n9421) );
  OAI221_X1 U10672 ( .B1(n9423), .B2(keyinput_g9), .C1(n9422), .C2(
        keyinput_g54), .A(n9421), .ZN(n9431) );
  AOI22_X1 U10673 ( .A1(n9425), .A2(keyinput_g52), .B1(n5005), .B2(
        keyinput_g21), .ZN(n9424) );
  OAI221_X1 U10674 ( .B1(n9425), .B2(keyinput_g52), .C1(n5005), .C2(
        keyinput_g21), .A(n9424), .ZN(n9430) );
  AOI22_X1 U10675 ( .A1(n9428), .A2(keyinput_g17), .B1(keyinput_g30), .B2(
        n9427), .ZN(n9426) );
  OAI221_X1 U10676 ( .B1(n9428), .B2(keyinput_g17), .C1(n9427), .C2(
        keyinput_g30), .A(n9426), .ZN(n9429) );
  NOR4_X1 U10677 ( .A1(n9432), .A2(n9431), .A3(n9430), .A4(n9429), .ZN(n9449)
         );
  AOI22_X1 U10678 ( .A1(n9435), .A2(keyinput_g50), .B1(n9434), .B2(
        keyinput_g13), .ZN(n9433) );
  OAI221_X1 U10679 ( .B1(n9435), .B2(keyinput_g50), .C1(n9434), .C2(
        keyinput_g13), .A(n9433), .ZN(n9447) );
  AOI22_X1 U10680 ( .A1(n9438), .A2(keyinput_g26), .B1(keyinput_g31), .B2(
        n9437), .ZN(n9436) );
  OAI221_X1 U10681 ( .B1(n9438), .B2(keyinput_g26), .C1(n9437), .C2(
        keyinput_g31), .A(n9436), .ZN(n9446) );
  AOI22_X1 U10682 ( .A1(n9441), .A2(keyinput_g4), .B1(n9440), .B2(keyinput_g23), .ZN(n9439) );
  OAI221_X1 U10683 ( .B1(n9441), .B2(keyinput_g4), .C1(n9440), .C2(
        keyinput_g23), .A(n9439), .ZN(n9445) );
  XNOR2_X1 U10684 ( .A(SI_0_), .B(keyinput_g32), .ZN(n9443) );
  XNOR2_X1 U10685 ( .A(SI_30_), .B(keyinput_g2), .ZN(n9442) );
  NAND2_X1 U10686 ( .A1(n9443), .A2(n9442), .ZN(n9444) );
  NOR4_X1 U10687 ( .A1(n9447), .A2(n9446), .A3(n9445), .A4(n9444), .ZN(n9448)
         );
  NAND4_X1 U10688 ( .A1(n9451), .A2(n9450), .A3(n9449), .A4(n9448), .ZN(n9494)
         );
  AOI22_X1 U10689 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_g58), .B1(
        SI_21_), .B2(keyinput_g11), .ZN(n9452) );
  OAI221_X1 U10690 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .C1(
        SI_21_), .C2(keyinput_g11), .A(n9452), .ZN(n9459) );
  AOI22_X1 U10691 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_g51), .B1(
        SI_13_), .B2(keyinput_g19), .ZN(n9453) );
  OAI221_X1 U10692 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .C1(
        SI_13_), .C2(keyinput_g19), .A(n9453), .ZN(n9458) );
  AOI22_X1 U10693 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_g47), .B1(
        SI_14_), .B2(keyinput_g18), .ZN(n9454) );
  OAI221_X1 U10694 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .C1(
        SI_14_), .C2(keyinput_g18), .A(n9454), .ZN(n9457) );
  AOI22_X1 U10695 ( .A1(SI_5_), .A2(keyinput_g27), .B1(SI_8_), .B2(
        keyinput_g24), .ZN(n9455) );
  OAI221_X1 U10696 ( .B1(SI_5_), .B2(keyinput_g27), .C1(SI_8_), .C2(
        keyinput_g24), .A(n9455), .ZN(n9456) );
  NOR4_X1 U10697 ( .A1(n9459), .A2(n9458), .A3(n9457), .A4(n9456), .ZN(n9492)
         );
  XOR2_X1 U10698 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_g48), .Z(n9466) );
  AOI22_X1 U10699 ( .A1(SI_10_), .A2(keyinput_g22), .B1(SI_20_), .B2(
        keyinput_g12), .ZN(n9460) );
  OAI221_X1 U10700 ( .B1(SI_10_), .B2(keyinput_g22), .C1(SI_20_), .C2(
        keyinput_g12), .A(n9460), .ZN(n9465) );
  AOI22_X1 U10701 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_g56), .B1(
        P2_RD_REG_SCAN_IN), .B2(keyinput_g33), .ZN(n9461) );
  OAI221_X1 U10702 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput_g33), .A(n9461), .ZN(n9464) );
  AOI22_X1 U10703 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_g53), .B1(SI_12_), .B2(keyinput_g20), .ZN(n9462) );
  OAI221_X1 U10704 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_g53), .C1(
        SI_12_), .C2(keyinput_g20), .A(n9462), .ZN(n9463) );
  NOR4_X1 U10705 ( .A1(n9466), .A2(n9465), .A3(n9464), .A4(n9463), .ZN(n9491)
         );
  AOI22_X1 U10706 ( .A1(n9469), .A2(keyinput_g36), .B1(n9468), .B2(
        keyinput_g10), .ZN(n9467) );
  OAI221_X1 U10707 ( .B1(n9469), .B2(keyinput_g36), .C1(n9468), .C2(
        keyinput_g10), .A(n9467), .ZN(n9480) );
  AOI22_X1 U10708 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_g39), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .ZN(n9470) );
  OAI221_X1 U10709 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_g37), .A(n9470), .ZN(n9479) );
  AOI22_X1 U10710 ( .A1(n9473), .A2(keyinput_g60), .B1(n9472), .B2(
        keyinput_g28), .ZN(n9471) );
  OAI221_X1 U10711 ( .B1(n9473), .B2(keyinput_g60), .C1(n9472), .C2(
        keyinput_g28), .A(n9471), .ZN(n9478) );
  AOI22_X1 U10712 ( .A1(n9476), .A2(keyinput_g62), .B1(keyinput_g61), .B2(
        n9475), .ZN(n9474) );
  OAI221_X1 U10713 ( .B1(n9476), .B2(keyinput_g62), .C1(n9475), .C2(
        keyinput_g61), .A(n9474), .ZN(n9477) );
  NOR4_X1 U10714 ( .A1(n9480), .A2(n9479), .A3(n9478), .A4(n9477), .ZN(n9490)
         );
  AOI22_X1 U10715 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_g40), .B1(SI_18_), .B2(keyinput_g14), .ZN(n9481) );
  OAI221_X1 U10716 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .C1(
        SI_18_), .C2(keyinput_g14), .A(n9481), .ZN(n9488) );
  AOI22_X1 U10717 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_g49), .B1(
        P2_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .ZN(n9482) );
  OAI221_X1 U10718 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_g38), .A(n9482), .ZN(n9487) );
  AOI22_X1 U10719 ( .A1(SI_29_), .A2(keyinput_g3), .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .ZN(n9483) );
  OAI221_X1 U10720 ( .B1(SI_29_), .B2(keyinput_g3), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n9483), .ZN(n9486) );
  AOI22_X1 U10721 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_g43), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n9484) );
  OAI221_X1 U10722 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_g43), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_g41), .A(n9484), .ZN(n9485) );
  NOR4_X1 U10723 ( .A1(n9488), .A2(n9487), .A3(n9486), .A4(n9485), .ZN(n9489)
         );
  NAND4_X1 U10724 ( .A1(n9492), .A2(n9491), .A3(n9490), .A4(n9489), .ZN(n9493)
         );
  OAI22_X1 U10725 ( .A1(keyinput_g63), .A2(n9497), .B1(n9494), .B2(n9493), 
        .ZN(n9495) );
  AOI211_X1 U10726 ( .C1(keyinput_g63), .C2(n9497), .A(n9496), .B(n9495), .ZN(
        n9498) );
  XNOR2_X1 U10727 ( .A(n9499), .B(n9498), .ZN(n9503) );
  NOR2_X1 U10728 ( .A1(n9501), .A2(n9500), .ZN(n9502) );
  XOR2_X1 U10729 ( .A(n9503), .B(n9502), .Z(ADD_1071_U4) );
  AOI22_X1 U10730 ( .A1(n9926), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9519) );
  INV_X1 U10731 ( .A(n9504), .ZN(n9506) );
  AND2_X1 U10732 ( .A1(n9506), .A2(n9505), .ZN(n9507) );
  OR3_X1 U10733 ( .A1(n9929), .A2(n9508), .A3(n9507), .ZN(n9515) );
  INV_X1 U10734 ( .A(n9509), .ZN(n9513) );
  INV_X1 U10735 ( .A(n9510), .ZN(n9512) );
  OAI211_X1 U10736 ( .C1(n9513), .C2(n9512), .A(n9924), .B(n9511), .ZN(n9514)
         );
  OAI211_X1 U10737 ( .C1(n9927), .C2(n9516), .A(n9515), .B(n9514), .ZN(n9517)
         );
  INV_X1 U10738 ( .A(n9517), .ZN(n9518) );
  NAND2_X1 U10739 ( .A1(n9519), .A2(n9518), .ZN(P2_U3247) );
  INV_X1 U10740 ( .A(n9524), .ZN(n9526) );
  AOI211_X1 U10741 ( .C1(n9563), .C2(n9522), .A(n9521), .B(n9520), .ZN(n9523)
         );
  OAI21_X1 U10742 ( .B1(n9524), .B2(n9658), .A(n9523), .ZN(n9525) );
  AOI21_X1 U10743 ( .B1(n9646), .B2(n9526), .A(n9525), .ZN(n9528) );
  INV_X1 U10744 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9527) );
  AOI22_X1 U10745 ( .A1(n9879), .A2(n9528), .B1(n9527), .B2(n9877), .ZN(
        P1_U3484) );
  AOI22_X1 U10746 ( .A1(n9888), .A2(n9528), .B1(n6584), .B2(n9886), .ZN(
        P1_U3533) );
  INV_X1 U10747 ( .A(n9529), .ZN(n9530) );
  AOI21_X1 U10748 ( .B1(n9892), .B2(n9531), .A(n9530), .ZN(n9538) );
  NAND2_X1 U10749 ( .A1(n9533), .A2(n9532), .ZN(n9534) );
  AOI21_X1 U10750 ( .B1(n4387), .B2(n9534), .A(n9909), .ZN(n9535) );
  AOI21_X1 U10751 ( .B1(n9902), .B2(n9536), .A(n9535), .ZN(n9537) );
  OAI211_X1 U10752 ( .C1(n9923), .C2(n9539), .A(n9538), .B(n9537), .ZN(
        P2_U3217) );
  INV_X1 U10753 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9543) );
  AOI22_X1 U10754 ( .A1(n10077), .A2(n9558), .B1(n9543), .B2(n10075), .ZN(
        P2_U3551) );
  INV_X1 U10755 ( .A(n9544), .ZN(n9549) );
  OAI22_X1 U10756 ( .A1(n9546), .A2(n10049), .B1(n9545), .B2(n10048), .ZN(
        n9547) );
  AOI211_X1 U10757 ( .C1(n9549), .C2(n10054), .A(n9548), .B(n9547), .ZN(n9560)
         );
  AOI22_X1 U10758 ( .A1(n10077), .A2(n9560), .B1(n9550), .B2(n10075), .ZN(
        P2_U3534) );
  INV_X1 U10759 ( .A(n9551), .ZN(n10040) );
  OAI22_X1 U10760 ( .A1(n9552), .A2(n10049), .B1(n4706), .B2(n10048), .ZN(
        n9554) );
  AOI211_X1 U10761 ( .C1(n10040), .C2(n9555), .A(n9554), .B(n9553), .ZN(n9562)
         );
  AOI22_X1 U10762 ( .A1(n10077), .A2(n9562), .B1(n9556), .B2(n10075), .ZN(
        P2_U3533) );
  INV_X1 U10763 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9557) );
  AOI22_X1 U10764 ( .A1(n10057), .A2(n9558), .B1(n9557), .B2(n10055), .ZN(
        P2_U3519) );
  INV_X1 U10765 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9559) );
  AOI22_X1 U10766 ( .A1(n10057), .A2(n9560), .B1(n9559), .B2(n10055), .ZN(
        P2_U3493) );
  INV_X1 U10767 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9561) );
  AOI22_X1 U10768 ( .A1(n10057), .A2(n9562), .B1(n9561), .B2(n10055), .ZN(
        P2_U3490) );
  NAND2_X1 U10769 ( .A1(n9595), .A2(n9563), .ZN(n9659) );
  INV_X1 U10770 ( .A(n9659), .ZN(n9571) );
  NAND2_X1 U10771 ( .A1(n9564), .A2(n9616), .ZN(n9567) );
  INV_X1 U10772 ( .A(n9565), .ZN(n9566) );
  OAI211_X1 U10773 ( .C1(n9584), .C2(n9568), .A(n9567), .B(n9566), .ZN(n9569)
         );
  AOI21_X1 U10774 ( .B1(n9571), .B2(n9570), .A(n9569), .ZN(n9579) );
  NAND2_X1 U10775 ( .A1(n9573), .A2(n9572), .ZN(n9575) );
  XNOR2_X1 U10776 ( .A(n9575), .B(n9574), .ZN(n9577) );
  NAND2_X1 U10777 ( .A1(n9577), .A2(n9576), .ZN(n9578) );
  OAI211_X1 U10778 ( .C1(n9580), .C2(n9592), .A(n9579), .B(n9578), .ZN(
        P1_U3239) );
  OAI21_X1 U10779 ( .B1(n9582), .B2(n9588), .A(n9581), .ZN(n9591) );
  OAI22_X1 U10780 ( .A1(n9586), .A2(n9585), .B1(n9584), .B2(n9583), .ZN(n9590)
         );
  XOR2_X1 U10781 ( .A(n9588), .B(n9587), .Z(n9596) );
  NOR2_X1 U10782 ( .A1(n9596), .A2(n9864), .ZN(n9589) );
  AOI211_X1 U10783 ( .C1(n9613), .C2(n9591), .A(n9590), .B(n9589), .ZN(n9661)
         );
  INV_X1 U10784 ( .A(n9592), .ZN(n9594) );
  AOI222_X1 U10785 ( .A1(n9595), .A2(n9651), .B1(n9594), .B2(n9593), .C1(
        P1_REG2_REG_15__SCAN_IN), .C2(n9647), .ZN(n9602) );
  INV_X1 U10786 ( .A(n9596), .ZN(n9664) );
  OAI21_X1 U10787 ( .B1(n9599), .B2(n9598), .A(n9597), .ZN(n9660) );
  INV_X1 U10788 ( .A(n9660), .ZN(n9600) );
  AOI22_X1 U10789 ( .A1(n9664), .A2(n9632), .B1(n9631), .B2(n9600), .ZN(n9601)
         );
  OAI211_X1 U10790 ( .C1(n9149), .C2(n9661), .A(n9602), .B(n9601), .ZN(
        P1_U3276) );
  INV_X1 U10791 ( .A(n9611), .ZN(n9603) );
  XNOR2_X1 U10792 ( .A(n9604), .B(n9603), .ZN(n9668) );
  AND2_X1 U10793 ( .A1(n9605), .A2(n9622), .ZN(n9607) );
  OR2_X1 U10794 ( .A1(n9607), .A2(n9606), .ZN(n9666) );
  INV_X1 U10795 ( .A(n9666), .ZN(n9608) );
  AOI22_X1 U10796 ( .A1(n9668), .A2(n9632), .B1(n9631), .B2(n9608), .ZN(n9624)
         );
  OAI22_X1 U10797 ( .A1(n9128), .A2(n9610), .B1(n9609), .B2(n9633), .ZN(n9621)
         );
  NOR2_X1 U10798 ( .A1(n9612), .A2(n9611), .ZN(n9615) );
  OAI21_X1 U10799 ( .B1(n9615), .B2(n9614), .A(n9613), .ZN(n9618) );
  AOI22_X1 U10800 ( .A1(n9641), .A2(n9639), .B1(n9616), .B2(n9638), .ZN(n9617)
         );
  NAND2_X1 U10801 ( .A1(n9618), .A2(n9617), .ZN(n9619) );
  AOI21_X1 U10802 ( .B1(n9668), .B2(n9646), .A(n9619), .ZN(n9670) );
  NOR2_X1 U10803 ( .A1(n9670), .A2(n9647), .ZN(n9620) );
  AOI211_X1 U10804 ( .C1(n9651), .C2(n9622), .A(n9621), .B(n9620), .ZN(n9623)
         );
  NAND2_X1 U10805 ( .A1(n9624), .A2(n9623), .ZN(P1_U3278) );
  INV_X1 U10806 ( .A(n9625), .ZN(n9636) );
  XNOR2_X1 U10807 ( .A(n9626), .B(n9636), .ZN(n9674) );
  OR2_X1 U10808 ( .A1(n9627), .A2(n9671), .ZN(n9628) );
  NAND2_X1 U10809 ( .A1(n9629), .A2(n9628), .ZN(n9672) );
  INV_X1 U10810 ( .A(n9672), .ZN(n9630) );
  AOI22_X1 U10811 ( .A1(n9674), .A2(n9632), .B1(n9631), .B2(n9630), .ZN(n9653)
         );
  OAI22_X1 U10812 ( .A1(n9128), .A2(n9635), .B1(n9634), .B2(n9633), .ZN(n9649)
         );
  XNOR2_X1 U10813 ( .A(n9637), .B(n9636), .ZN(n9644) );
  AOI22_X1 U10814 ( .A1(n9641), .A2(n9640), .B1(n9639), .B2(n9638), .ZN(n9642)
         );
  OAI21_X1 U10815 ( .B1(n9644), .B2(n9643), .A(n9642), .ZN(n9645) );
  AOI21_X1 U10816 ( .B1(n9674), .B2(n9646), .A(n9645), .ZN(n9676) );
  NOR2_X1 U10817 ( .A1(n9676), .A2(n9647), .ZN(n9648) );
  AOI211_X1 U10818 ( .C1(n9651), .C2(n9650), .A(n9649), .B(n9648), .ZN(n9652)
         );
  NAND2_X1 U10819 ( .A1(n9653), .A2(n9652), .ZN(P1_U3280) );
  OAI21_X1 U10820 ( .B1(n9655), .B2(n9854), .A(n9654), .ZN(n9656) );
  AOI21_X1 U10821 ( .B1(n9657), .B2(n9860), .A(n9656), .ZN(n9678) );
  AOI22_X1 U10822 ( .A1(n9888), .A2(n9678), .B1(n6367), .B2(n9886), .ZN(
        P1_U3553) );
  INV_X1 U10823 ( .A(n9658), .ZN(n9868) );
  OAI21_X1 U10824 ( .B1(n9660), .B2(n9873), .A(n9659), .ZN(n9663) );
  INV_X1 U10825 ( .A(n9661), .ZN(n9662) );
  AOI211_X1 U10826 ( .C1(n9868), .C2(n9664), .A(n9663), .B(n9662), .ZN(n9680)
         );
  AOI22_X1 U10827 ( .A1(n9888), .A2(n9680), .B1(n5948), .B2(n9886), .ZN(
        P1_U3538) );
  OAI22_X1 U10828 ( .A1(n9666), .A2(n9873), .B1(n9665), .B2(n9854), .ZN(n9667)
         );
  AOI21_X1 U10829 ( .B1(n9668), .B2(n9868), .A(n9667), .ZN(n9669) );
  AOI22_X1 U10830 ( .A1(n9888), .A2(n9682), .B1(n5908), .B2(n9886), .ZN(
        P1_U3536) );
  OAI22_X1 U10831 ( .A1(n9672), .A2(n9873), .B1(n9671), .B2(n9854), .ZN(n9673)
         );
  AOI21_X1 U10832 ( .B1(n9674), .B2(n9868), .A(n9673), .ZN(n9675) );
  AND2_X1 U10833 ( .A1(n9676), .A2(n9675), .ZN(n9684) );
  AOI22_X1 U10834 ( .A1(n9888), .A2(n9684), .B1(n6738), .B2(n9886), .ZN(
        P1_U3534) );
  INV_X1 U10835 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9677) );
  AOI22_X1 U10836 ( .A1(n9879), .A2(n9678), .B1(n9677), .B2(n9877), .ZN(
        P1_U3521) );
  INV_X1 U10837 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9679) );
  AOI22_X1 U10838 ( .A1(n9879), .A2(n9680), .B1(n9679), .B2(n9877), .ZN(
        P1_U3499) );
  INV_X1 U10839 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9681) );
  AOI22_X1 U10840 ( .A1(n9879), .A2(n9682), .B1(n9681), .B2(n9877), .ZN(
        P1_U3493) );
  INV_X1 U10841 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9683) );
  AOI22_X1 U10842 ( .A1(n9879), .A2(n9684), .B1(n9683), .B2(n9877), .ZN(
        P1_U3487) );
  XNOR2_X1 U10843 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U10844 ( .A(n9685), .ZN(n9694) );
  AND2_X1 U10845 ( .A1(n9689), .A2(n5647), .ZN(n9687) );
  OAI21_X1 U10846 ( .B1(n9688), .B2(n9687), .A(n9686), .ZN(n9709) );
  INV_X1 U10847 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9695) );
  OAI21_X1 U10848 ( .B1(n5647), .B2(n9695), .A(n9689), .ZN(n9690) );
  OAI211_X1 U10849 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9692), .A(n9691), .B(
        n9690), .ZN(n9693) );
  AND3_X1 U10850 ( .A1(n9694), .A2(n9709), .A3(n9693), .ZN(n9697) );
  NOR3_X1 U10851 ( .A1(n9736), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n9695), .ZN(
        n9696) );
  AOI211_X1 U10852 ( .C1(P1_ADDR_REG_0__SCAN_IN), .C2(n9783), .A(n9697), .B(
        n9696), .ZN(n9698) );
  OAI21_X1 U10853 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n5644), .A(n9698), .ZN(
        P1_U3241) );
  INV_X1 U10854 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9718) );
  OAI211_X1 U10855 ( .C1(n9701), .C2(n9700), .A(n9797), .B(n9699), .ZN(n9702)
         );
  INV_X1 U10856 ( .A(n9702), .ZN(n9703) );
  AOI21_X1 U10857 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(P1_U3084), .A(n9703), 
        .ZN(n9717) );
  AOI211_X1 U10858 ( .C1(n9706), .C2(n9705), .A(n9704), .B(n9775), .ZN(n9714)
         );
  MUX2_X1 U10859 ( .A(n9708), .B(n9707), .S(n6355), .Z(n9712) );
  OAI211_X1 U10860 ( .C1(n9712), .C2(n9711), .A(n9710), .B(n9709), .ZN(n9713)
         );
  INV_X1 U10861 ( .A(n9713), .ZN(n9732) );
  AOI211_X1 U10862 ( .C1(n9789), .C2(n9715), .A(n9714), .B(n9732), .ZN(n9716)
         );
  OAI211_X1 U10863 ( .C1(n9802), .C2(n9718), .A(n9717), .B(n9716), .ZN(
        P1_U3243) );
  INV_X1 U10864 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9735) );
  OAI21_X1 U10865 ( .B1(n9721), .B2(n9720), .A(n9719), .ZN(n9723) );
  AOI22_X1 U10866 ( .A1(n9798), .A2(n9723), .B1(n9789), .B2(n9722), .ZN(n9734)
         );
  INV_X1 U10867 ( .A(n9724), .ZN(n9726) );
  OAI21_X1 U10868 ( .B1(n9727), .B2(n9726), .A(n9725), .ZN(n9728) );
  AOI21_X1 U10869 ( .B1(n9729), .B2(n9728), .A(n9736), .ZN(n9730) );
  NOR3_X1 U10870 ( .A1(n9732), .A2(n9731), .A3(n9730), .ZN(n9733) );
  OAI211_X1 U10871 ( .C1(n9802), .C2(n9735), .A(n9734), .B(n9733), .ZN(
        P1_U3245) );
  AOI211_X1 U10872 ( .C1(n9739), .C2(n9738), .A(n9737), .B(n9736), .ZN(n9740)
         );
  AOI211_X1 U10873 ( .C1(n9789), .C2(n9742), .A(n9741), .B(n9740), .ZN(n9748)
         );
  OAI21_X1 U10874 ( .B1(n9745), .B2(n9744), .A(n9743), .ZN(n9746) );
  NAND2_X1 U10875 ( .A1(n9798), .A2(n9746), .ZN(n9747) );
  OAI211_X1 U10876 ( .C1(n10123), .C2(n9802), .A(n9748), .B(n9747), .ZN(
        P1_U3246) );
  AOI22_X1 U10877 ( .A1(n9783), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n9749), .B2(
        n9789), .ZN(n9759) );
  XNOR2_X1 U10878 ( .A(n9751), .B(n9750), .ZN(n9757) );
  AOI211_X1 U10879 ( .C1(n9754), .C2(n9753), .A(n9752), .B(n9775), .ZN(n9755)
         );
  AOI211_X1 U10880 ( .C1(n9797), .C2(n9757), .A(n9756), .B(n9755), .ZN(n9758)
         );
  NAND2_X1 U10881 ( .A1(n9759), .A2(n9758), .ZN(P1_U3247) );
  OAI21_X1 U10882 ( .B1(n9762), .B2(n9761), .A(n9760), .ZN(n9768) );
  AOI211_X1 U10883 ( .C1(n9765), .C2(n9764), .A(n9763), .B(n9775), .ZN(n9766)
         );
  AOI211_X1 U10884 ( .C1(n9797), .C2(n9768), .A(n9767), .B(n9766), .ZN(n9771)
         );
  AOI22_X1 U10885 ( .A1(n9783), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(n9769), .B2(
        n9789), .ZN(n9770) );
  NAND2_X1 U10886 ( .A1(n9771), .A2(n9770), .ZN(P1_U3250) );
  OAI21_X1 U10887 ( .B1(n9774), .B2(n9773), .A(n9772), .ZN(n9781) );
  AOI211_X1 U10888 ( .C1(n9778), .C2(n9777), .A(n9776), .B(n9775), .ZN(n9779)
         );
  AOI211_X1 U10889 ( .C1(n9797), .C2(n9781), .A(n9780), .B(n9779), .ZN(n9785)
         );
  AOI22_X1 U10890 ( .A1(n9783), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(n9782), .B2(
        n9789), .ZN(n9784) );
  NAND2_X1 U10891 ( .A1(n9785), .A2(n9784), .ZN(P1_U3251) );
  INV_X1 U10892 ( .A(n9786), .ZN(n9787) );
  AOI21_X1 U10893 ( .B1(n9789), .B2(n9788), .A(n9787), .ZN(n9801) );
  AOI21_X1 U10894 ( .B1(n9792), .B2(n9791), .A(n9790), .ZN(n9799) );
  OAI21_X1 U10895 ( .B1(n9795), .B2(n9794), .A(n9793), .ZN(n9796) );
  AOI22_X1 U10896 ( .A1(n9799), .A2(n9798), .B1(n9797), .B2(n9796), .ZN(n9800)
         );
  OAI211_X1 U10897 ( .C1(n9802), .C2(n10115), .A(n9801), .B(n9800), .ZN(
        P1_U3259) );
  INV_X1 U10898 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n9803) );
  NOR2_X1 U10899 ( .A1(n9834), .A2(n9803), .ZN(P1_U3292) );
  INV_X1 U10900 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n9804) );
  NOR2_X1 U10901 ( .A1(n9834), .A2(n9804), .ZN(P1_U3293) );
  INV_X1 U10902 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n9805) );
  NOR2_X1 U10903 ( .A1(n9834), .A2(n9805), .ZN(P1_U3294) );
  INV_X1 U10904 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9806) );
  NOR2_X1 U10905 ( .A1(n9816), .A2(n9806), .ZN(P1_U3295) );
  INV_X1 U10906 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9807) );
  NOR2_X1 U10907 ( .A1(n9816), .A2(n9807), .ZN(P1_U3296) );
  INV_X1 U10908 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9808) );
  NOR2_X1 U10909 ( .A1(n9816), .A2(n9808), .ZN(P1_U3297) );
  INV_X1 U10910 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n9809) );
  NOR2_X1 U10911 ( .A1(n9816), .A2(n9809), .ZN(P1_U3298) );
  INV_X1 U10912 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9810) );
  NOR2_X1 U10913 ( .A1(n9816), .A2(n9810), .ZN(P1_U3299) );
  INV_X1 U10914 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9811) );
  NOR2_X1 U10915 ( .A1(n9816), .A2(n9811), .ZN(P1_U3300) );
  INV_X1 U10916 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9812) );
  NOR2_X1 U10917 ( .A1(n9816), .A2(n9812), .ZN(P1_U3301) );
  INV_X1 U10918 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9813) );
  NOR2_X1 U10919 ( .A1(n9816), .A2(n9813), .ZN(P1_U3302) );
  INV_X1 U10920 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9814) );
  NOR2_X1 U10921 ( .A1(n9816), .A2(n9814), .ZN(P1_U3303) );
  INV_X1 U10922 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9815) );
  NOR2_X1 U10923 ( .A1(n9816), .A2(n9815), .ZN(P1_U3304) );
  INV_X1 U10924 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n9817) );
  NOR2_X1 U10925 ( .A1(n9834), .A2(n9817), .ZN(P1_U3305) );
  INV_X1 U10926 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9818) );
  NOR2_X1 U10927 ( .A1(n9834), .A2(n9818), .ZN(P1_U3306) );
  INV_X1 U10928 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9819) );
  NOR2_X1 U10929 ( .A1(n9834), .A2(n9819), .ZN(P1_U3307) );
  INV_X1 U10930 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n9820) );
  NOR2_X1 U10931 ( .A1(n9834), .A2(n9820), .ZN(P1_U3308) );
  INV_X1 U10932 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9821) );
  NOR2_X1 U10933 ( .A1(n9834), .A2(n9821), .ZN(P1_U3309) );
  INV_X1 U10934 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9822) );
  NOR2_X1 U10935 ( .A1(n9834), .A2(n9822), .ZN(P1_U3310) );
  INV_X1 U10936 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9823) );
  NOR2_X1 U10937 ( .A1(n9834), .A2(n9823), .ZN(P1_U3311) );
  INV_X1 U10938 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9824) );
  NOR2_X1 U10939 ( .A1(n9834), .A2(n9824), .ZN(P1_U3312) );
  INV_X1 U10940 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n9825) );
  NOR2_X1 U10941 ( .A1(n9834), .A2(n9825), .ZN(P1_U3313) );
  INV_X1 U10942 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9826) );
  NOR2_X1 U10943 ( .A1(n9834), .A2(n9826), .ZN(P1_U3314) );
  INV_X1 U10944 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9827) );
  NOR2_X1 U10945 ( .A1(n9834), .A2(n9827), .ZN(P1_U3315) );
  INV_X1 U10946 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n9828) );
  NOR2_X1 U10947 ( .A1(n9834), .A2(n9828), .ZN(P1_U3316) );
  INV_X1 U10948 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9829) );
  NOR2_X1 U10949 ( .A1(n9834), .A2(n9829), .ZN(P1_U3317) );
  INV_X1 U10950 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9830) );
  NOR2_X1 U10951 ( .A1(n9834), .A2(n9830), .ZN(P1_U3318) );
  INV_X1 U10952 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9831) );
  NOR2_X1 U10953 ( .A1(n9834), .A2(n9831), .ZN(P1_U3319) );
  INV_X1 U10954 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9832) );
  NOR2_X1 U10955 ( .A1(n9834), .A2(n9832), .ZN(P1_U3320) );
  INV_X1 U10956 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n9833) );
  NOR2_X1 U10957 ( .A1(n9834), .A2(n9833), .ZN(P1_U3321) );
  OAI22_X1 U10958 ( .A1(n9836), .A2(n9873), .B1(n9835), .B2(n9854), .ZN(n9838)
         );
  AOI211_X1 U10959 ( .C1(n9868), .C2(n9839), .A(n9838), .B(n9837), .ZN(n9880)
         );
  INV_X1 U10960 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9840) );
  AOI22_X1 U10961 ( .A1(n9879), .A2(n9880), .B1(n9840), .B2(n9877), .ZN(
        P1_U3463) );
  OAI21_X1 U10962 ( .B1(n9842), .B2(n9854), .A(n9841), .ZN(n9844) );
  AOI211_X1 U10963 ( .C1(n9845), .C2(n9875), .A(n9844), .B(n9843), .ZN(n9881)
         );
  AOI22_X1 U10964 ( .A1(n9879), .A2(n9881), .B1(n5745), .B2(n9877), .ZN(
        P1_U3469) );
  OAI22_X1 U10965 ( .A1(n9847), .A2(n9873), .B1(n9846), .B2(n9854), .ZN(n9849)
         );
  AOI211_X1 U10966 ( .C1(n9868), .C2(n9850), .A(n9849), .B(n9848), .ZN(n9882)
         );
  INV_X1 U10967 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9851) );
  AOI22_X1 U10968 ( .A1(n9879), .A2(n9882), .B1(n9851), .B2(n9877), .ZN(
        P1_U3472) );
  OAI211_X1 U10969 ( .C1(n9855), .C2(n9854), .A(n9853), .B(n9852), .ZN(n9856)
         );
  AOI21_X1 U10970 ( .B1(n9875), .B2(n9857), .A(n9856), .ZN(n9883) );
  INV_X1 U10971 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9858) );
  AOI22_X1 U10972 ( .A1(n9879), .A2(n9883), .B1(n9858), .B2(n9877), .ZN(
        P1_U3475) );
  AOI21_X1 U10973 ( .B1(n9861), .B2(n9860), .A(n9859), .ZN(n9862) );
  OAI211_X1 U10974 ( .C1(n9865), .C2(n9864), .A(n9863), .B(n9862), .ZN(n9866)
         );
  AOI21_X1 U10975 ( .B1(n9868), .B2(n9867), .A(n9866), .ZN(n9885) );
  AOI22_X1 U10976 ( .A1(n9879), .A2(n9885), .B1(n5799), .B2(n9877), .ZN(
        P1_U3478) );
  INV_X1 U10977 ( .A(n9869), .ZN(n9870) );
  OAI211_X1 U10978 ( .C1(n9873), .C2(n9872), .A(n9871), .B(n9870), .ZN(n9874)
         );
  AOI21_X1 U10979 ( .B1(n9876), .B2(n9875), .A(n9874), .ZN(n9887) );
  INV_X1 U10980 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9878) );
  AOI22_X1 U10981 ( .A1(n9879), .A2(n9887), .B1(n9878), .B2(n9877), .ZN(
        P1_U3481) );
  AOI22_X1 U10982 ( .A1(n9888), .A2(n9880), .B1(n6382), .B2(n9886), .ZN(
        P1_U3526) );
  AOI22_X1 U10983 ( .A1(n9888), .A2(n9881), .B1(n5744), .B2(n9886), .ZN(
        P1_U3528) );
  AOI22_X1 U10984 ( .A1(n9888), .A2(n9882), .B1(n6411), .B2(n9886), .ZN(
        P1_U3529) );
  AOI22_X1 U10985 ( .A1(n9888), .A2(n9883), .B1(n5782), .B2(n9886), .ZN(
        P1_U3530) );
  AOI22_X1 U10986 ( .A1(n9888), .A2(n9885), .B1(n9884), .B2(n9886), .ZN(
        P1_U3531) );
  AOI22_X1 U10987 ( .A1(n9888), .A2(n9887), .B1(n5829), .B2(n9886), .ZN(
        P1_U3532) );
  INV_X1 U10988 ( .A(n9889), .ZN(n9890) );
  AOI21_X1 U10989 ( .B1(n9892), .B2(n9891), .A(n9890), .ZN(n9906) );
  INV_X1 U10990 ( .A(n7058), .ZN(n9895) );
  OAI21_X1 U10991 ( .B1(n9895), .B2(n9894), .A(n9893), .ZN(n9900) );
  NAND3_X1 U10992 ( .A1(n9898), .A2(n9897), .A3(n9896), .ZN(n9899) );
  NAND2_X1 U10993 ( .A1(n9900), .A2(n9899), .ZN(n9904) );
  AOI22_X1 U10994 ( .A1(n9904), .A2(n9903), .B1(n9902), .B2(n9901), .ZN(n9905)
         );
  OAI211_X1 U10995 ( .C1(n9923), .C2(n9907), .A(n9906), .B(n9905), .ZN(
        P2_U3226) );
  AOI211_X1 U10996 ( .C1(n9911), .C2(n9910), .A(n9909), .B(n9908), .ZN(n9920)
         );
  OAI22_X1 U10997 ( .A1(n9913), .A2(n9912), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5119), .ZN(n9919) );
  OAI22_X1 U10998 ( .A1(n9917), .A2(n9916), .B1(n9915), .B2(n9914), .ZN(n9918)
         );
  NOR3_X1 U10999 ( .A1(n9920), .A2(n9919), .A3(n9918), .ZN(n9921) );
  OAI21_X1 U11000 ( .B1(n9923), .B2(n9922), .A(n9921), .ZN(P2_U3229) );
  AOI22_X1 U11001 ( .A1(n9925), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9924), .ZN(n9934) );
  AOI22_X1 U11002 ( .A1(n9926), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9933) );
  OAI21_X1 U11003 ( .B1(n9928), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9927), .ZN(
        n9931) );
  NOR2_X1 U11004 ( .A1(n9929), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9930) );
  OAI21_X1 U11005 ( .B1(n9931), .B2(n9930), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9932) );
  OAI211_X1 U11006 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9934), .A(n9933), .B(
        n9932), .ZN(P2_U3245) );
  XNOR2_X1 U11007 ( .A(n9935), .B(n7307), .ZN(n10039) );
  INV_X1 U11008 ( .A(n9937), .ZN(n9938) );
  AOI211_X1 U11009 ( .C1(n9936), .C2(n7307), .A(n9939), .B(n9938), .ZN(n9940)
         );
  AOI211_X1 U11010 ( .C1(n9942), .C2(n10039), .A(n9941), .B(n9940), .ZN(n10036) );
  AOI222_X1 U11011 ( .A1(n9946), .A2(n9945), .B1(P2_REG2_REG_10__SCAN_IN), 
        .B2(n9944), .C1(n9960), .C2(n9943), .ZN(n9954) );
  INV_X1 U11012 ( .A(n9947), .ZN(n9948) );
  OAI21_X1 U11013 ( .B1(n10034), .B2(n9949), .A(n9948), .ZN(n10035) );
  INV_X1 U11014 ( .A(n10035), .ZN(n9950) );
  AOI22_X1 U11015 ( .A1(n10039), .A2(n9952), .B1(n9951), .B2(n9950), .ZN(n9953) );
  OAI211_X1 U11016 ( .C1(n9944), .C2(n10036), .A(n9954), .B(n9953), .ZN(
        P2_U3286) );
  INV_X1 U11017 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9970) );
  INV_X1 U11018 ( .A(n9955), .ZN(n9966) );
  INV_X1 U11019 ( .A(n9956), .ZN(n9963) );
  AOI22_X1 U11020 ( .A1(n9960), .A2(n9959), .B1(n9958), .B2(n9957), .ZN(n9961)
         );
  OAI21_X1 U11021 ( .B1(n9963), .B2(n9962), .A(n9961), .ZN(n9965) );
  AOI211_X1 U11022 ( .C1(n9967), .C2(n9966), .A(n9965), .B(n9964), .ZN(n9969)
         );
  AOI22_X1 U11023 ( .A1(n9944), .A2(n9970), .B1(n9969), .B2(n9968), .ZN(
        P2_U3291) );
  INV_X1 U11024 ( .A(n9971), .ZN(n9973) );
  NAND2_X1 U11025 ( .A1(n9973), .A2(n9972), .ZN(n9976) );
  AND2_X1 U11026 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9976), .ZN(P2_U3297) );
  AND2_X1 U11027 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9976), .ZN(P2_U3298) );
  AND2_X1 U11028 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9976), .ZN(P2_U3299) );
  AND2_X1 U11029 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9976), .ZN(P2_U3300) );
  AND2_X1 U11030 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9976), .ZN(P2_U3301) );
  AND2_X1 U11031 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9976), .ZN(P2_U3302) );
  AND2_X1 U11032 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9976), .ZN(P2_U3303) );
  AND2_X1 U11033 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9976), .ZN(P2_U3304) );
  AND2_X1 U11034 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9976), .ZN(P2_U3305) );
  AND2_X1 U11035 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9976), .ZN(P2_U3306) );
  AND2_X1 U11036 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9976), .ZN(P2_U3307) );
  AND2_X1 U11037 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9976), .ZN(P2_U3308) );
  AND2_X1 U11038 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9976), .ZN(P2_U3309) );
  AND2_X1 U11039 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9976), .ZN(P2_U3310) );
  AND2_X1 U11040 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9976), .ZN(P2_U3311) );
  AND2_X1 U11041 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9976), .ZN(P2_U3312) );
  AND2_X1 U11042 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9976), .ZN(P2_U3313) );
  AND2_X1 U11043 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9976), .ZN(P2_U3314) );
  AND2_X1 U11044 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9976), .ZN(P2_U3315) );
  AND2_X1 U11045 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9976), .ZN(P2_U3316) );
  AND2_X1 U11046 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9976), .ZN(P2_U3317) );
  AND2_X1 U11047 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9976), .ZN(P2_U3318) );
  AND2_X1 U11048 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9976), .ZN(P2_U3319) );
  AND2_X1 U11049 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9976), .ZN(P2_U3320) );
  AND2_X1 U11050 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9976), .ZN(P2_U3321) );
  AND2_X1 U11051 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9976), .ZN(P2_U3322) );
  AND2_X1 U11052 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9976), .ZN(P2_U3323) );
  AND2_X1 U11053 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9976), .ZN(P2_U3324) );
  AND2_X1 U11054 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9976), .ZN(P2_U3325) );
  AND2_X1 U11055 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9976), .ZN(P2_U3326) );
  AOI22_X1 U11056 ( .A1(n9975), .A2(n9976), .B1(n9979), .B2(n9974), .ZN(
        P2_U3437) );
  AOI22_X1 U11057 ( .A1(n9979), .A2(n9978), .B1(n9977), .B2(n9976), .ZN(
        P2_U3438) );
  INV_X1 U11058 ( .A(n9980), .ZN(n9986) );
  OAI22_X1 U11059 ( .A1(n9984), .A2(n9983), .B1(n9982), .B2(n9981), .ZN(n9985)
         );
  NOR2_X1 U11060 ( .A1(n9986), .A2(n9985), .ZN(n10059) );
  INV_X1 U11061 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9987) );
  AOI22_X1 U11062 ( .A1(n10057), .A2(n10059), .B1(n9987), .B2(n10055), .ZN(
        P2_U3451) );
  OAI22_X1 U11063 ( .A1(n9989), .A2(n10049), .B1(n9988), .B2(n10048), .ZN(
        n9991) );
  AOI211_X1 U11064 ( .C1(n10054), .C2(n9992), .A(n9991), .B(n9990), .ZN(n10061) );
  INV_X1 U11065 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9993) );
  AOI22_X1 U11066 ( .A1(n10057), .A2(n10061), .B1(n9993), .B2(n10055), .ZN(
        P2_U3454) );
  OAI22_X1 U11067 ( .A1(n9994), .A2(n10049), .B1(n6634), .B2(n10048), .ZN(
        n9996) );
  AOI211_X1 U11068 ( .C1(n10054), .C2(n9997), .A(n9996), .B(n9995), .ZN(n10063) );
  INV_X1 U11069 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9998) );
  AOI22_X1 U11070 ( .A1(n10057), .A2(n10063), .B1(n9998), .B2(n10055), .ZN(
        P2_U3457) );
  OAI22_X1 U11071 ( .A1(n10000), .A2(n10049), .B1(n9999), .B2(n10048), .ZN(
        n10002) );
  AOI211_X1 U11072 ( .C1(n10054), .C2(n10003), .A(n10002), .B(n10001), .ZN(
        n10065) );
  INV_X1 U11073 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10004) );
  AOI22_X1 U11074 ( .A1(n10057), .A2(n10065), .B1(n10004), .B2(n10055), .ZN(
        P2_U3463) );
  OAI22_X1 U11075 ( .A1(n10006), .A2(n10049), .B1(n10005), .B2(n10048), .ZN(
        n10008) );
  AOI211_X1 U11076 ( .C1(n10054), .C2(n10009), .A(n10008), .B(n10007), .ZN(
        n10066) );
  INV_X1 U11077 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10010) );
  AOI22_X1 U11078 ( .A1(n10057), .A2(n10066), .B1(n10010), .B2(n10055), .ZN(
        P2_U3469) );
  OAI22_X1 U11079 ( .A1(n10012), .A2(n10049), .B1(n10011), .B2(n10048), .ZN(
        n10014) );
  AOI211_X1 U11080 ( .C1(n10054), .C2(n10015), .A(n10014), .B(n10013), .ZN(
        n10068) );
  INV_X1 U11081 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10016) );
  AOI22_X1 U11082 ( .A1(n10057), .A2(n10068), .B1(n10016), .B2(n10055), .ZN(
        P2_U3472) );
  AOI22_X1 U11083 ( .A1(n10020), .A2(n10019), .B1(n10018), .B2(n10017), .ZN(
        n10024) );
  NAND3_X1 U11084 ( .A1(n10022), .A2(n10021), .A3(n10054), .ZN(n10023) );
  AND3_X1 U11085 ( .A1(n10025), .A2(n10024), .A3(n10023), .ZN(n10070) );
  INV_X1 U11086 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10026) );
  AOI22_X1 U11087 ( .A1(n10057), .A2(n10070), .B1(n10026), .B2(n10055), .ZN(
        P2_U3475) );
  INV_X1 U11088 ( .A(n10027), .ZN(n10028) );
  OAI22_X1 U11089 ( .A1(n10029), .A2(n10049), .B1(n10028), .B2(n10048), .ZN(
        n10031) );
  AOI211_X1 U11090 ( .C1(n10040), .C2(n10032), .A(n10031), .B(n10030), .ZN(
        n10072) );
  INV_X1 U11091 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10033) );
  AOI22_X1 U11092 ( .A1(n10057), .A2(n10072), .B1(n10033), .B2(n10055), .ZN(
        P2_U3478) );
  OAI22_X1 U11093 ( .A1(n10035), .A2(n10049), .B1(n10034), .B2(n10048), .ZN(
        n10038) );
  INV_X1 U11094 ( .A(n10036), .ZN(n10037) );
  AOI211_X1 U11095 ( .C1(n10040), .C2(n10039), .A(n10038), .B(n10037), .ZN(
        n10073) );
  INV_X1 U11096 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10041) );
  AOI22_X1 U11097 ( .A1(n10057), .A2(n10073), .B1(n10041), .B2(n10055), .ZN(
        P2_U3481) );
  OAI22_X1 U11098 ( .A1(n10043), .A2(n10049), .B1(n10042), .B2(n10048), .ZN(
        n10045) );
  AOI211_X1 U11099 ( .C1(n10046), .C2(n10054), .A(n10045), .B(n10044), .ZN(
        n10074) );
  INV_X1 U11100 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10047) );
  AOI22_X1 U11101 ( .A1(n10057), .A2(n10074), .B1(n10047), .B2(n10055), .ZN(
        P2_U3484) );
  OAI22_X1 U11102 ( .A1(n10050), .A2(n10049), .B1(n4707), .B2(n10048), .ZN(
        n10052) );
  AOI211_X1 U11103 ( .C1(n10054), .C2(n10053), .A(n10052), .B(n10051), .ZN(
        n10076) );
  INV_X1 U11104 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10056) );
  AOI22_X1 U11105 ( .A1(n10057), .A2(n10076), .B1(n10056), .B2(n10055), .ZN(
        P2_U3487) );
  INV_X1 U11106 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10058) );
  AOI22_X1 U11107 ( .A1(n10077), .A2(n10059), .B1(n10058), .B2(n10075), .ZN(
        P2_U3520) );
  INV_X1 U11108 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10060) );
  AOI22_X1 U11109 ( .A1(n10077), .A2(n10061), .B1(n10060), .B2(n10075), .ZN(
        P2_U3521) );
  INV_X1 U11110 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10062) );
  AOI22_X1 U11111 ( .A1(n10077), .A2(n10063), .B1(n10062), .B2(n10075), .ZN(
        P2_U3522) );
  INV_X1 U11112 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10064) );
  AOI22_X1 U11113 ( .A1(n10077), .A2(n10065), .B1(n10064), .B2(n10075), .ZN(
        P2_U3524) );
  AOI22_X1 U11114 ( .A1(n10077), .A2(n10066), .B1(n6462), .B2(n10075), .ZN(
        P2_U3526) );
  AOI22_X1 U11115 ( .A1(n10077), .A2(n10068), .B1(n10067), .B2(n10075), .ZN(
        P2_U3527) );
  AOI22_X1 U11116 ( .A1(n10077), .A2(n10070), .B1(n10069), .B2(n10075), .ZN(
        P2_U3528) );
  AOI22_X1 U11117 ( .A1(n10077), .A2(n10072), .B1(n10071), .B2(n10075), .ZN(
        P2_U3529) );
  AOI22_X1 U11118 ( .A1(n10077), .A2(n10073), .B1(n6599), .B2(n10075), .ZN(
        P2_U3530) );
  AOI22_X1 U11119 ( .A1(n10077), .A2(n10074), .B1(n6669), .B2(n10075), .ZN(
        P2_U3531) );
  AOI22_X1 U11120 ( .A1(n10077), .A2(n10076), .B1(n6852), .B2(n10075), .ZN(
        P2_U3532) );
  INV_X1 U11121 ( .A(n10078), .ZN(n10079) );
  NAND2_X1 U11122 ( .A1(n10080), .A2(n10079), .ZN(n10081) );
  XNOR2_X1 U11123 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10081), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11124 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11125 ( .B1(n10084), .B2(n10083), .A(n10082), .ZN(ADD_1071_U56) );
  OAI21_X1 U11126 ( .B1(n10087), .B2(n10086), .A(n10085), .ZN(ADD_1071_U57) );
  OAI21_X1 U11127 ( .B1(n10090), .B2(n10089), .A(n10088), .ZN(ADD_1071_U58) );
  OAI21_X1 U11128 ( .B1(n10093), .B2(n10092), .A(n10091), .ZN(ADD_1071_U59) );
  OAI21_X1 U11129 ( .B1(n10096), .B2(n10095), .A(n10094), .ZN(ADD_1071_U60) );
  OAI21_X1 U11130 ( .B1(n10099), .B2(n10098), .A(n10097), .ZN(ADD_1071_U61) );
  AOI21_X1 U11131 ( .B1(n10102), .B2(n10101), .A(n10100), .ZN(ADD_1071_U62) );
  AOI21_X1 U11132 ( .B1(n10105), .B2(n10104), .A(n10103), .ZN(ADD_1071_U63) );
  AOI21_X1 U11133 ( .B1(n10108), .B2(n10107), .A(n10106), .ZN(ADD_1071_U47) );
  XOR2_X1 U11134 ( .A(n10110), .B(n10109), .Z(ADD_1071_U54) );
  XNOR2_X1 U11135 ( .A(n10112), .B(n10111), .ZN(ADD_1071_U48) );
  OAI21_X1 U11136 ( .B1(n10115), .B2(n10114), .A(n10113), .ZN(n10116) );
  XNOR2_X1 U11137 ( .A(n10116), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XNOR2_X1 U11138 ( .A(n10118), .B(n10117), .ZN(ADD_1071_U49) );
  XNOR2_X1 U11139 ( .A(n10120), .B(n10119), .ZN(ADD_1071_U50) );
  AOI21_X1 U11140 ( .B1(n10122), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n10121), .ZN(
        n10124) );
  XNOR2_X1 U11141 ( .A(n10124), .B(n10123), .ZN(ADD_1071_U51) );
  XOR2_X1 U11142 ( .A(n10126), .B(n10125), .Z(ADD_1071_U53) );
  XNOR2_X1 U11143 ( .A(n10128), .B(n10127), .ZN(ADD_1071_U52) );
  XNOR2_X1 U4961 ( .A(n5458), .B(n5448), .ZN(n8213) );
  INV_X1 U4826 ( .A(n4313), .ZN(n4314) );
  CLKBUF_X1 U4829 ( .A(n5356), .Z(n5249) );
  CLKBUF_X2 U4860 ( .A(n8091), .Z(n4320) );
endmodule

