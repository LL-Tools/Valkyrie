

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput63,
         keyinput62, keyinput61, keyinput60, keyinput59, keyinput58,
         keyinput57, keyinput56, keyinput55, keyinput54, keyinput53,
         keyinput52, keyinput51, keyinput50, keyinput49, keyinput48,
         keyinput47, keyinput46, keyinput45, keyinput44, keyinput43,
         keyinput42, keyinput41, keyinput40, keyinput39, keyinput38,
         keyinput37, keyinput36, keyinput35, keyinput34, keyinput33,
         keyinput32, keyinput31, keyinput30, keyinput29, keyinput28,
         keyinput27, keyinput26, keyinput25, keyinput24, keyinput23,
         keyinput22, keyinput21, keyinput20, keyinput19, keyinput18,
         keyinput17, keyinput16, keyinput15, keyinput14, keyinput13,
         keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7,
         keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1,
         keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008;

  INV_X4 U7166 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X4 U7167 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  OAI21_X1 U7168 ( .B1(n8037), .B2(n8036), .A(n8039), .ZN(n8060) );
  AND2_X1 U7169 ( .A1(n11966), .A2(n7206), .ZN(n7205) );
  CLKBUF_X2 U7170 ( .A(n10179), .Z(n12365) );
  CLKBUF_X2 U7171 ( .A(n12921), .Z(n12948) );
  INV_X1 U7172 ( .A(n11940), .ZN(n12364) );
  OR2_X1 U7173 ( .A1(n9747), .A2(n9748), .ZN(n11941) );
  INV_X1 U7175 ( .A(n10161), .ZN(n13595) );
  INV_X1 U7176 ( .A(n8079), .ZN(n7580) );
  INV_X2 U7177 ( .A(n7484), .ZN(n7534) );
  NAND4_X1 U7178 ( .A1(n7590), .A2(n7150), .A3(n7214), .A4(n7213), .ZN(n7410)
         );
  NOR2_X1 U7179 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7374) );
  CLKBUF_X1 U7180 ( .A(n13002), .Z(n6418) );
  OAI21_X1 U7181 ( .B1(n10016), .B2(n10573), .A(n13245), .ZN(n13002) );
  OR2_X1 U7182 ( .A1(n14633), .A2(n14632), .ZN(n14630) );
  NOR2_X1 U7183 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n7377) );
  INV_X1 U7184 ( .A(n8327), .ZN(n8305) );
  INV_X1 U7185 ( .A(n12288), .ZN(n12294) );
  AND3_X1 U7186 ( .A1(n8357), .A2(n8356), .A3(n8355), .ZN(n10056) );
  CLKBUF_X3 U7187 ( .A(n7760), .Z(n6455) );
  NOR2_X1 U7188 ( .A1(n13120), .A2(n7138), .ZN(n7135) );
  INV_X1 U7189 ( .A(n7434), .ZN(n7859) );
  INV_X1 U7190 ( .A(n12161), .ZN(n12310) );
  CLKBUF_X2 U7191 ( .A(n12096), .Z(n9361) );
  AND3_X1 U7192 ( .A1(n8304), .A2(n8303), .A3(n8302), .ZN(n14815) );
  AND3_X1 U7193 ( .A1(n7308), .A2(n8326), .A3(n7307), .ZN(n10200) );
  INV_X1 U7194 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8723) );
  OR2_X1 U7195 ( .A1(n11965), .A2(n6498), .ZN(n11966) );
  INV_X2 U7197 ( .A(n7534), .ZN(n7798) );
  INV_X1 U7198 ( .A(n10995), .ZN(n10010) );
  OR2_X1 U7199 ( .A1(n9529), .A2(n9270), .ZN(n6494) );
  XNOR2_X1 U7201 ( .A(n11186), .B(n11185), .ZN(n11297) );
  NAND2_X1 U7202 ( .A1(n7410), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7412) );
  AND4_X1 U7203 ( .A1(n8892), .A2(n7281), .A3(n8891), .A4(n8890), .ZN(n10161)
         );
  INV_X1 U7204 ( .A(n6953), .ZN(n9454) );
  INV_X2 U7206 ( .A(n13257), .ZN(n13304) );
  XNOR2_X1 U7207 ( .A(n9454), .B(n9453), .ZN(n14043) );
  AND2_X2 U7208 ( .A1(n9978), .A2(n9977), .ZN(n6419) );
  NAND2_X2 U7209 ( .A1(n13900), .A2(n11848), .ZN(n13869) );
  NAND2_X2 U7210 ( .A1(n7361), .A2(n7297), .ZN(n13900) );
  AND2_X1 U7211 ( .A1(n9978), .A2(n9977), .ZN(n6420) );
  NAND2_X1 U7212 ( .A1(n10022), .A2(n10021), .ZN(n12921) );
  NAND2_X1 U7213 ( .A1(n13598), .A2(n10098), .ZN(n9926) );
  NAND2_X2 U7214 ( .A1(n14580), .A2(n9860), .ZN(n8107) );
  OAI21_X2 U7215 ( .B1(n13167), .B2(n13051), .A(n13160), .ZN(n13144) );
  NAND4_X2 U7216 ( .A1(n8826), .A2(n8825), .A3(n8824), .A4(n8823), .ZN(n13594)
         );
  OAI21_X2 U7217 ( .B1(n8015), .B2(n6899), .A(n6894), .ZN(n8037) );
  NAND2_X2 U7218 ( .A1(n12418), .A2(n12417), .ZN(n12443) );
  BUF_X2 U7219 ( .A(n8888), .Z(n6425) );
  NAND2_X2 U7220 ( .A1(n11701), .A2(n11700), .ZN(n11967) );
  NOR2_X2 U7221 ( .A1(n9387), .A2(n9386), .ZN(n9388) );
  NAND2_X2 U7222 ( .A1(n8701), .A2(n12257), .ZN(n12775) );
  NAND2_X2 U7223 ( .A1(n10115), .A2(n10114), .ZN(n10149) );
  XNOR2_X2 U7224 ( .A(n13952), .B(n13827), .ZN(n13813) );
  AOI21_X2 U7225 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n10636), .A(n14712), .ZN(
        n10590) );
  AND4_X4 U7226 ( .A1(n8349), .A2(n8348), .A3(n8347), .A4(n8346), .ZN(n8358)
         );
  XNOR2_X2 U7227 ( .A(n8060), .B(n8059), .ZN(n14008) );
  NAND4_X4 U7228 ( .A1(n8834), .A2(n8833), .A3(n8832), .A4(n8831), .ZN(n13597)
         );
  NOR2_X2 U7230 ( .A1(n12959), .A2(n12958), .ZN(n13007) );
  OR2_X2 U7231 ( .A1(n12868), .A2(n8723), .ZN(n8242) );
  BUF_X4 U7232 ( .A(n8345), .Z(n12087) );
  OAI21_X2 U7233 ( .B1(n12514), .B2(n12392), .A(n12435), .ZN(n12496) );
  XNOR2_X2 U7234 ( .A(n8070), .B(n8069), .ZN(n13427) );
  AOI21_X2 U7235 ( .B1(n11031), .B2(n11032), .A(n8414), .ZN(n11289) );
  AND2_X1 U7236 ( .A1(n14005), .A2(n14003), .ZN(n6421) );
  AND2_X2 U7237 ( .A1(n14005), .A2(n14003), .ZN(n8889) );
  NOR2_X1 U7238 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n7280) );
  XNOR2_X2 U7239 ( .A(n8773), .B(P1_IR_REG_30__SCAN_IN), .ZN(n8783) );
  XNOR2_X2 U7240 ( .A(n12398), .B(n12399), .ZN(n12501) );
  XOR2_X2 U7241 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), .Z(
        n9422) );
  AOI22_X2 U7242 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P3_ADDR_REG_2__SCAN_IN), 
        .B1(n14923), .B2(n14930), .ZN(n9420) );
  XNOR2_X1 U7243 ( .A(n8234), .B(n8233), .ZN(n6422) );
  INV_X1 U7244 ( .A(n12073), .ZN(n6423) );
  OAI21_X2 U7245 ( .B1(n10092), .B2(n10091), .A(n9927), .ZN(n10110) );
  XNOR2_X2 U7246 ( .A(n8354), .B(P3_IR_REG_2__SCAN_IN), .ZN(n10334) );
  OR2_X2 U7247 ( .A1(n10322), .A2(n8723), .ZN(n8354) );
  NAND2_X1 U7248 ( .A1(n11850), .A2(n11849), .ZN(n13858) );
  OAI22_X1 U7249 ( .A1(n13199), .A2(n6990), .B1(n6992), .B2(n6497), .ZN(n13162) );
  NAND2_X1 U7250 ( .A1(n11250), .A2(n7042), .ZN(n7044) );
  INV_X2 U7251 ( .A(n14346), .ZN(n10887) );
  AND2_X1 U7252 ( .A1(n10054), .A2(n9983), .ZN(n9990) );
  AND2_X1 U7253 ( .A1(n8142), .A2(n10290), .ZN(n10562) );
  NAND2_X1 U7254 ( .A1(n12916), .A2(n13071), .ZN(n10253) );
  INV_X1 U7255 ( .A(n14305), .ZN(n14328) );
  INV_X1 U7256 ( .A(n13594), .ZN(n10164) );
  INV_X2 U7257 ( .A(n13597), .ZN(n6611) );
  CLKBUF_X2 U7258 ( .A(n8107), .Z(n6467) );
  INV_X2 U7259 ( .A(n8107), .ZN(n8123) );
  INV_X1 U7260 ( .A(n8676), .ZN(n6424) );
  CLKBUF_X2 U7261 ( .A(n9235), .Z(n9262) );
  INV_X1 U7262 ( .A(n10455), .ZN(n8757) );
  NAND2_X1 U7263 ( .A1(n9754), .A2(n9747), .ZN(n11942) );
  NAND2_X1 U7264 ( .A1(n8669), .A2(n8668), .ZN(n10455) );
  INV_X1 U7265 ( .A(n8863), .ZN(n10098) );
  XNOR2_X1 U7266 ( .A(n6453), .B(n8816), .ZN(n11020) );
  BUF_X2 U7267 ( .A(n7485), .Z(n8096) );
  NOR2_X1 U7268 ( .A1(n10579), .A2(n6519), .ZN(n10580) );
  NAND2_X1 U7269 ( .A1(n7433), .A2(n8840), .ZN(n7455) );
  NAND2_X1 U7270 ( .A1(n7414), .A2(n6724), .ZN(n7457) );
  INV_X2 U7271 ( .A(n9501), .ZN(n9504) );
  INV_X2 U7272 ( .A(n7416), .ZN(n9501) );
  BUF_X1 U7273 ( .A(n8257), .Z(n10322) );
  OR2_X1 U7274 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n8808) );
  INV_X1 U7275 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6613) );
  NAND2_X1 U7276 ( .A1(n7093), .A2(n7094), .ZN(n9260) );
  MUX2_X1 U7277 ( .A(n12051), .B(n12050), .S(n12049), .Z(n12057) );
  AOI22_X1 U7278 ( .A1(n12045), .A2(n12049), .B1(n13560), .B2(n13930), .ZN(
        n13747) );
  OAI21_X1 U7279 ( .B1(n13034), .B2(n13033), .A(n13032), .ZN(n13036) );
  AND2_X1 U7280 ( .A1(n6710), .A2(n6506), .ZN(n13034) );
  NAND2_X1 U7281 ( .A1(n6436), .A2(n6435), .ZN(n13447) );
  AOI21_X1 U7282 ( .B1(n6438), .B2(n6440), .A(n12356), .ZN(n6435) );
  NAND2_X1 U7283 ( .A1(n13489), .A2(n6438), .ZN(n6436) );
  NAND2_X1 U7284 ( .A1(n6437), .A2(n12349), .ZN(n13555) );
  NAND2_X1 U7285 ( .A1(n8705), .A2(n12273), .ZN(n12688) );
  NAND2_X1 U7286 ( .A1(n6610), .A2(n6502), .ZN(n11857) );
  NAND2_X1 U7287 ( .A1(n6716), .A2(n6717), .ZN(n12983) );
  NAND2_X1 U7288 ( .A1(n13489), .A2(n13490), .ZN(n6437) );
  AND2_X1 U7289 ( .A1(n6439), .A2(n13556), .ZN(n6438) );
  NOR2_X1 U7290 ( .A1(n7347), .A2(n6718), .ZN(n6717) );
  OR2_X1 U7291 ( .A1(n13490), .A2(n6440), .ZN(n6439) );
  AND2_X1 U7292 ( .A1(n12355), .A2(n12354), .ZN(n12356) );
  INV_X1 U7293 ( .A(n12349), .ZN(n6440) );
  NAND2_X1 U7294 ( .A1(n13526), .A2(n7034), .ZN(n7032) );
  OR2_X1 U7295 ( .A1(n12743), .A2(n12738), .ZN(n8703) );
  NAND2_X1 U7296 ( .A1(n13480), .A2(n12321), .ZN(n13526) );
  INV_X1 U7297 ( .A(n13118), .ZN(n13315) );
  NAND2_X1 U7298 ( .A1(n12317), .A2(n7037), .ZN(n13480) );
  NAND2_X1 U7299 ( .A1(n9253), .A2(n9252), .ZN(n13927) );
  AND2_X1 U7300 ( .A1(n13870), .A2(n11871), .ZN(n13855) );
  NAND2_X1 U7301 ( .A1(n11946), .A2(n11945), .ZN(n12317) );
  NAND2_X1 U7302 ( .A1(n13872), .A2(n13871), .ZN(n13870) );
  NAND2_X1 U7303 ( .A1(n13466), .A2(n11927), .ZN(n11946) );
  NAND2_X1 U7304 ( .A1(n13497), .A2(n11915), .ZN(n13466) );
  AND2_X1 U7305 ( .A1(n11869), .A2(n11868), .ZN(n13872) );
  NAND2_X1 U7306 ( .A1(n7030), .A2(n13566), .ZN(n13497) );
  NAND2_X1 U7307 ( .A1(n13568), .A2(n13567), .ZN(n13566) );
  AND2_X1 U7308 ( .A1(n7344), .A2(n7031), .ZN(n7030) );
  OAI21_X1 U7309 ( .B1(n12727), .B2(n12110), .A(n12111), .ZN(n12717) );
  XNOR2_X1 U7310 ( .A(n11911), .B(n11909), .ZN(n13568) );
  OR2_X1 U7311 ( .A1(n11911), .A2(n11910), .ZN(n7344) );
  NAND2_X1 U7312 ( .A1(n14122), .A2(n11903), .ZN(n11911) );
  XNOR2_X1 U7313 ( .A(n7980), .B(SI_24_), .ZN(n7977) );
  NAND2_X1 U7314 ( .A1(n9151), .A2(n9150), .ZN(n13965) );
  NAND2_X1 U7315 ( .A1(n14121), .A2(n11899), .ZN(n14122) );
  NAND2_X1 U7316 ( .A1(n6618), .A2(n6916), .ZN(n7980) );
  NAND2_X1 U7317 ( .A1(n6430), .A2(n6429), .ZN(n11828) );
  AOI21_X1 U7318 ( .B1(n6431), .B2(n6434), .A(n7039), .ZN(n6429) );
  OAI21_X1 U7319 ( .B1(n11571), .B2(n6434), .A(n6431), .ZN(n14136) );
  NAND2_X1 U7320 ( .A1(n11576), .A2(n11575), .ZN(n14135) );
  NAND2_X1 U7321 ( .A1(n11571), .A2(n6431), .ZN(n6430) );
  XNOR2_X1 U7322 ( .A(n7899), .B(SI_20_), .ZN(n7898) );
  NAND2_X1 U7323 ( .A1(n11571), .A2(n6625), .ZN(n11576) );
  AND2_X1 U7324 ( .A1(n11783), .A2(n6432), .ZN(n6431) );
  OR2_X1 U7325 ( .A1(n11789), .A2(n7040), .ZN(n7039) );
  NAND2_X1 U7326 ( .A1(n9456), .A2(n9457), .ZN(n6967) );
  NAND2_X1 U7327 ( .A1(n7044), .A2(n6509), .ZN(n11571) );
  NAND2_X1 U7328 ( .A1(n11575), .A2(n6433), .ZN(n6432) );
  INV_X1 U7329 ( .A(n11575), .ZN(n6434) );
  NAND2_X1 U7330 ( .A1(n11047), .A2(n11046), .ZN(n11250) );
  INV_X1 U7331 ( .A(n6625), .ZN(n6433) );
  NAND2_X1 U7332 ( .A1(n11041), .A2(n7348), .ZN(n11047) );
  NAND2_X1 U7333 ( .A1(n10469), .A2(n10470), .ZN(n10823) );
  NAND2_X1 U7334 ( .A1(n10881), .A2(n10880), .ZN(n11041) );
  NAND2_X1 U7335 ( .A1(n10757), .A2(n10756), .ZN(n10785) );
  AOI21_X1 U7336 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n9404), .A(n9403), .ZN(
        n9458) );
  NAND2_X1 U7337 ( .A1(n9004), .A2(n9003), .ZN(n14172) );
  NAND2_X1 U7338 ( .A1(n7639), .A2(n7638), .ZN(n11146) );
  OAI21_X1 U7339 ( .B1(n10876), .B2(n10875), .A(n10874), .ZN(n10881) );
  NAND2_X1 U7340 ( .A1(n7666), .A2(n7665), .ZN(n11174) );
  NAND2_X1 U7341 ( .A1(n10357), .A2(n10356), .ZN(n10755) );
  AND2_X1 U7342 ( .A1(n8972), .A2(n8971), .ZN(n11426) );
  XNOR2_X1 U7343 ( .A(n7029), .B(n10536), .ZN(n10538) );
  NAND2_X1 U7344 ( .A1(n6911), .A2(n6913), .ZN(n7680) );
  NAND2_X1 U7345 ( .A1(n6442), .A2(n6441), .ZN(n7029) );
  AND2_X1 U7346 ( .A1(n13536), .A2(n7027), .ZN(n7026) );
  NAND2_X1 U7347 ( .A1(n9990), .A2(n9986), .ZN(n10055) );
  OAI21_X1 U7348 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n9400), .A(n9399), .ZN(
        n9414) );
  XNOR2_X1 U7349 ( .A(n6720), .B(n7610), .ZN(n9570) );
  INV_X2 U7350 ( .A(n14597), .ZN(n10992) );
  INV_X2 U7351 ( .A(n14603), .ZN(n10988) );
  AND2_X1 U7352 ( .A1(n12197), .A2(n12196), .ZN(n12113) );
  NOR2_X1 U7353 ( .A1(n9397), .A2(n9396), .ZN(n9417) );
  AND2_X1 U7354 ( .A1(n10459), .A2(n10458), .ZN(n6477) );
  INV_X8 U7355 ( .A(n6419), .ZN(n12444) );
  AND4_X1 U7356 ( .A1(n8296), .A2(n8295), .A3(n8294), .A4(n8293), .ZN(n12207)
         );
  NAND4_X1 U7357 ( .A1(n8283), .A2(n8282), .A3(n8281), .A4(n8280), .ZN(n12553)
         );
  NAND4_X1 U7358 ( .A1(n8381), .A2(n8380), .A3(n8379), .A4(n8378), .ZN(n12181)
         );
  AND4_X1 U7359 ( .A1(n8269), .A2(n8268), .A3(n8267), .A4(n8266), .ZN(n10818)
         );
  NAND2_X1 U7360 ( .A1(n6424), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8335) );
  AND4_X1 U7361 ( .A1(n8333), .A2(n8332), .A3(n8331), .A4(n8330), .ZN(n8342)
         );
  INV_X2 U7362 ( .A(n12921), .ZN(n12917) );
  AND2_X1 U7363 ( .A1(n9750), .A2(n6452), .ZN(n9755) );
  BUF_X4 U7364 ( .A(n8123), .Z(n6460) );
  BUF_X4 U7365 ( .A(n8123), .Z(n6461) );
  CLKBUF_X3 U7366 ( .A(n8344), .Z(n8484) );
  NAND2_X2 U7367 ( .A1(n12069), .A2(n8245), .ZN(n8676) );
  INV_X2 U7368 ( .A(n10541), .ZN(n12366) );
  NAND2_X1 U7369 ( .A1(n7481), .A2(n7480), .ZN(n10772) );
  AND2_X2 U7370 ( .A1(n12310), .A2(n10207), .ZN(n12288) );
  INV_X2 U7371 ( .A(n8327), .ZN(n12083) );
  INV_X8 U7372 ( .A(n9238), .ZN(n9192) );
  CLKBUF_X2 U7373 ( .A(n6466), .Z(n9265) );
  INV_X1 U7374 ( .A(n8246), .ZN(n12069) );
  OR2_X2 U7375 ( .A1(n11942), .A2(n6445), .ZN(n11940) );
  NAND4_X1 U7376 ( .A1(n7490), .A2(n7489), .A3(n7488), .A4(n7487), .ZN(n13071)
         );
  OR2_X2 U7377 ( .A1(n8246), .A2(n8245), .ZN(n8327) );
  NAND2_X1 U7378 ( .A1(n10995), .A2(n9860), .ZN(n10021) );
  CLKBUF_X1 U7379 ( .A(n9860), .Z(n11143) );
  NAND4_X1 U7380 ( .A1(n7448), .A2(n7447), .A3(n7446), .A4(n7445), .ZN(n8146)
         );
  CLKBUF_X2 U7381 ( .A(n9274), .Z(n6466) );
  INV_X1 U7382 ( .A(n14182), .ZN(n6445) );
  CLKBUF_X3 U7383 ( .A(n9247), .Z(n6462) );
  AND2_X2 U7384 ( .A1(n8165), .A2(n7400), .ZN(n9860) );
  CLKBUF_X3 U7385 ( .A(n9247), .Z(n6463) );
  NAND2_X1 U7386 ( .A1(n8888), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8844) );
  NAND2_X2 U7387 ( .A1(n9756), .A2(n11020), .ZN(n14182) );
  NAND2_X1 U7388 ( .A1(n9343), .A2(n11534), .ZN(n9754) );
  NOR2_X1 U7389 ( .A1(n9389), .A2(n9390), .ZN(n9391) );
  XNOR2_X1 U7390 ( .A(n8244), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8245) );
  MUX2_X1 U7391 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7399), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n7400) );
  XNOR2_X1 U7392 ( .A(n6454), .B(P1_IR_REG_24__SCAN_IN), .ZN(n11534) );
  INV_X1 U7393 ( .A(n12380), .ZN(n8812) );
  CLKBUF_X1 U7394 ( .A(n8680), .Z(n6630) );
  AND2_X1 U7395 ( .A1(n12380), .A2(n9908), .ZN(n9756) );
  OR2_X1 U7396 ( .A1(n7426), .A2(n7428), .ZN(n7430) );
  AND2_X1 U7397 ( .A1(n7387), .A2(n7386), .ZN(n7717) );
  INV_X2 U7398 ( .A(n8104), .ZN(n7960) );
  NAND2_X1 U7399 ( .A1(n8811), .A2(n6446), .ZN(n12380) );
  NAND2_X1 U7400 ( .A1(n8815), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6453) );
  OR2_X1 U7401 ( .A1(n7401), .A2(n14924), .ZN(n7426) );
  NAND2_X1 U7402 ( .A1(n8792), .A2(n8793), .ZN(n8846) );
  AND2_X1 U7403 ( .A1(n12042), .A2(n7386), .ZN(n7484) );
  OAI21_X1 U7404 ( .B1(n9334), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6454) );
  NAND2_X1 U7405 ( .A1(n8165), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8108) );
  NAND2_X1 U7406 ( .A1(n7288), .A2(n7287), .ZN(n8792) );
  NAND2_X1 U7407 ( .A1(n9335), .A2(n9337), .ZN(n14015) );
  XNOR2_X1 U7408 ( .A(n8234), .B(n8233), .ZN(n8681) );
  MUX2_X1 U7409 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8774), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n8775) );
  NAND2_X1 U7410 ( .A1(n8807), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8814) );
  OAI21_X1 U7411 ( .B1(n8807), .B2(n8808), .A(n6447), .ZN(n6446) );
  AND2_X1 U7412 ( .A1(n8810), .A2(n8809), .ZN(n8811) );
  NOR2_X1 U7413 ( .A1(n7023), .A2(n7022), .ZN(n7021) );
  INV_X1 U7414 ( .A(n9341), .ZN(n8790) );
  NAND2_X1 U7415 ( .A1(n8793), .A2(n6612), .ZN(n7024) );
  INV_X1 U7416 ( .A(n10334), .ZN(n10641) );
  AND3_X2 U7417 ( .A1(n9338), .A2(n6470), .A3(n7279), .ZN(n8776) );
  AOI21_X1 U7418 ( .B1(n6963), .B2(n6962), .A(n9383), .ZN(n9385) );
  AND3_X2 U7419 ( .A1(n6534), .A2(n8916), .A3(n6474), .ZN(n9338) );
  OAI21_X1 U7420 ( .B1(n9423), .B2(n9422), .A(n6542), .ZN(n6963) );
  AOI21_X1 U7421 ( .B1(n7289), .B2(n6613), .A(n6545), .ZN(n7287) );
  AND4_X1 U7422 ( .A1(n8769), .A2(n8768), .A3(n8767), .A4(n8798), .ZN(n6474)
         );
  NOR2_X2 U7423 ( .A1(n8877), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n8916) );
  AND2_X1 U7424 ( .A1(n7353), .A2(n8721), .ZN(n6952) );
  NOR2_X1 U7425 ( .A1(n8772), .A2(n6613), .ZN(n6612) );
  AND3_X1 U7426 ( .A1(n8804), .A2(n7025), .A3(n8797), .ZN(n8769) );
  NOR2_X1 U7427 ( .A1(n6613), .A2(n6448), .ZN(n6447) );
  AND4_X1 U7428 ( .A1(n8257), .A2(n8220), .A3(n8221), .A4(n8315), .ZN(n6815)
         );
  NAND2_X1 U7429 ( .A1(n8827), .A2(n7280), .ZN(n8877) );
  AND4_X1 U7430 ( .A1(n8225), .A2(n8224), .A3(n8223), .A4(n8425), .ZN(n8226)
         );
  NAND4_X1 U7431 ( .A1(n6922), .A2(n6921), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7262) );
  INV_X1 U7432 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7265) );
  INV_X1 U7433 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13096) );
  INV_X1 U7434 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7264) );
  INV_X1 U7435 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14613) );
  INV_X1 U7436 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n6922) );
  INV_X1 U7437 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n7404) );
  INV_X1 U7438 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6448) );
  INV_X1 U7439 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8666) );
  NOR2_X1 U7440 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n8798) );
  NOR2_X1 U7441 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n8257) );
  NOR2_X1 U7442 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6428) );
  NOR2_X1 U7443 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n6427) );
  NOR2_X1 U7444 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n6426) );
  INV_X1 U7445 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6451) );
  INV_X1 U7446 ( .A(P2_RD_REG_SCAN_IN), .ZN(n6921) );
  INV_X1 U7447 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8915) );
  INV_X1 U7448 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8921) );
  INV_X1 U7449 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8923) );
  NOR2_X2 U7450 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n8827) );
  INV_X4 U7451 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7452 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n8982) );
  INV_X1 U7453 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8425) );
  INV_X1 U7454 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7524) );
  NOR2_X1 U7455 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n8224) );
  NOR2_X1 U7456 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n8225) );
  INV_X1 U7457 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6450) );
  INV_X1 U7458 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7398) );
  INV_X1 U7459 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8369) );
  INV_X1 U7460 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8259) );
  NOR2_X1 U7461 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n7393) );
  NAND4_X1 U7462 ( .A1(n6428), .A2(n6427), .A3(n6426), .A4(n6451), .ZN(n9049)
         );
  NAND2_X1 U7463 ( .A1(n11834), .A2(n11833), .ZN(n14121) );
  AOI21_X1 U7464 ( .B1(n7027), .B2(n6444), .A(n6477), .ZN(n6441) );
  NAND2_X1 U7465 ( .A1(n6443), .A2(n7027), .ZN(n6442) );
  INV_X1 U7466 ( .A(n13537), .ZN(n6443) );
  INV_X1 U7467 ( .A(n13538), .ZN(n6444) );
  NAND2_X1 U7468 ( .A1(n13537), .A2(n13538), .ZN(n13536) );
  NAND2_X1 U7469 ( .A1(n12364), .A2(n13598), .ZN(n6452) );
  NOR2_X2 U7470 ( .A1(n9049), .A2(n6449), .ZN(n6534) );
  NAND4_X1 U7471 ( .A1(n8921), .A2(n8923), .A3(n8915), .A4(n6450), .ZN(n6449)
         );
  NAND2_X1 U7473 ( .A1(n11828), .A2(n11827), .ZN(n11834) );
  XNOR2_X1 U7474 ( .A(n7853), .B(SI_18_), .ZN(n7852) );
  XNOR2_X1 U7475 ( .A(n14071), .B(n12610), .ZN(n14081) );
  NAND2_X1 U7476 ( .A1(n8687), .A2(n8686), .ZN(n10714) );
  NAND2_X2 U7477 ( .A1(n8692), .A2(n12220), .ZN(n11345) );
  INV_X1 U7478 ( .A(n9870), .ZN(n13093) );
  NAND2_X1 U7479 ( .A1(n13745), .A2(n7350), .ZN(n11862) );
  NAND2_X1 U7480 ( .A1(n13747), .A2(n13746), .ZN(n13745) );
  NAND2_X1 U7481 ( .A1(n7434), .A2(n9504), .ZN(n7760) );
  AND2_X2 U7482 ( .A1(n8509), .A2(n6952), .ZN(n8716) );
  INV_X1 U7483 ( .A(n10552), .ZN(n6883) );
  NAND2_X2 U7484 ( .A1(n8822), .A2(n8821), .ZN(n10552) );
  NAND2_X1 U7485 ( .A1(n9559), .A2(n9501), .ZN(n6456) );
  NAND2_X1 U7486 ( .A1(n9559), .A2(n9501), .ZN(n6457) );
  NAND2_X1 U7487 ( .A1(n9559), .A2(n9501), .ZN(n8895) );
  NAND2_X1 U7488 ( .A1(n7304), .A2(n7302), .ZN(n13788) );
  NOR2_X2 U7489 ( .A1(n10079), .A2(n13540), .ZN(n14312) );
  AOI21_X2 U7491 ( .B1(n12662), .B2(n12141), .A(n12286), .ZN(n9376) );
  AOI21_X2 U7492 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n14033), .A(n11184), .ZN(
        n11186) );
  NAND2_X2 U7493 ( .A1(n11227), .A2(n11226), .ZN(n14170) );
  NAND2_X2 U7494 ( .A1(n8920), .A2(n8919), .ZN(n14346) );
  NAND2_X1 U7495 ( .A1(n10022), .A2(n10021), .ZN(n6459) );
  XNOR2_X2 U7496 ( .A(n11862), .B(n11861), .ZN(n13923) );
  NAND2_X1 U7497 ( .A1(n9338), .A2(n8788), .ZN(n9341) );
  XNOR2_X2 U7498 ( .A(n7456), .B(n7455), .ZN(n9506) );
  NAND2_X1 U7499 ( .A1(n13788), .A2(n11859), .ZN(n13761) );
  CLKBUF_X1 U7500 ( .A(n9274), .Z(n6465) );
  NOR2_X2 U7501 ( .A1(n8243), .A2(P3_IR_REG_29__SCAN_IN), .ZN(n12868) );
  INV_X2 U7502 ( .A(n8676), .ZN(n12082) );
  NAND4_X4 U7503 ( .A1(n8337), .A2(n8336), .A3(n8335), .A4(n8334), .ZN(n9718)
         );
  NOR2_X2 U7504 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7449) );
  OAI21_X2 U7505 ( .B1(n11158), .B2(n6713), .A(n7201), .ZN(n11520) );
  NAND3_X2 U7506 ( .A1(n6608), .A2(n7407), .A3(n9870), .ZN(n13341) );
  INV_X1 U7507 ( .A(n8783), .ZN(n14003) );
  AND2_X1 U7508 ( .A1(n8783), .A2(n8782), .ZN(n9247) );
  INV_X2 U7509 ( .A(n10080), .ZN(n9761) );
  AND4_X4 U7510 ( .A1(n8843), .A2(n8842), .A3(n8845), .A4(n8844), .ZN(n10080)
         );
  AND2_X1 U7511 ( .A1(n14005), .A2(n8783), .ZN(n9274) );
  AND2_X2 U7512 ( .A1(n8782), .A2(n14003), .ZN(n8888) );
  AOI21_X2 U7513 ( .B1(n13761), .B2(n13760), .A(n11860), .ZN(n12045) );
  OR2_X1 U7514 ( .A1(n13150), .A2(n12968), .ZN(n12012) );
  NOR2_X1 U7515 ( .A1(n6986), .A2(n6988), .ZN(n6985) );
  INV_X1 U7516 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7367) );
  NOR2_X1 U7517 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n7368) );
  INV_X1 U7518 ( .A(n13919), .ZN(n11880) );
  NAND2_X1 U7519 ( .A1(n14091), .A2(n12534), .ZN(n12296) );
  NAND2_X1 U7520 ( .A1(n7434), .A2(n9501), .ZN(n8104) );
  INV_X1 U7521 ( .A(n12031), .ZN(n7007) );
  NAND2_X1 U7522 ( .A1(n6745), .A2(n6747), .ZN(n6744) );
  INV_X1 U7523 ( .A(n6748), .ZN(n6747) );
  OR2_X1 U7524 ( .A1(n13805), .A2(n13779), .ZN(n11858) );
  NAND2_X1 U7525 ( .A1(n11857), .A2(n7305), .ZN(n7304) );
  NOR2_X1 U7526 ( .A1(n13793), .A2(n7306), .ZN(n7305) );
  INV_X1 U7527 ( .A(n11856), .ZN(n7306) );
  NAND2_X1 U7528 ( .A1(n7482), .A2(n7253), .ZN(n7252) );
  AND2_X1 U7529 ( .A1(n9066), .A2(n11341), .ZN(n7052) );
  AND2_X1 U7530 ( .A1(n9281), .A2(n13589), .ZN(n9065) );
  INV_X1 U7531 ( .A(n9096), .ZN(n7074) );
  NAND2_X1 U7532 ( .A1(n7814), .A2(n7815), .ZN(n7243) );
  INV_X1 U7533 ( .A(n7917), .ZN(n7249) );
  OAI21_X1 U7534 ( .B1(n7876), .B2(n7875), .A(n7877), .ZN(n7899) );
  NAND2_X1 U7535 ( .A1(n14616), .A2(n10646), .ZN(n14636) );
  NAND2_X1 U7536 ( .A1(n14636), .A2(n14635), .ZN(n14634) );
  OR2_X1 U7537 ( .A1(n12570), .A2(n12569), .ZN(n12571) );
  OR2_X1 U7538 ( .A1(n12529), .A2(n12415), .ZN(n12281) );
  INV_X1 U7539 ( .A(n12232), .ZN(n6831) );
  NAND2_X1 U7540 ( .A1(n6686), .A2(n6685), .ZN(n8604) );
  NAND2_X1 U7541 ( .A1(n6599), .A2(n8591), .ZN(n6685) );
  NAND2_X1 U7542 ( .A1(n14499), .A2(n6753), .ZN(n11730) );
  OR2_X1 U7543 ( .A1(n14510), .A2(n11455), .ZN(n6753) );
  NOR2_X1 U7544 ( .A1(n13222), .A2(n13246), .ZN(n7146) );
  NAND2_X1 U7545 ( .A1(n6529), .A2(n6469), .ZN(n7144) );
  INV_X1 U7546 ( .A(n7148), .ZN(n7145) );
  NOR2_X1 U7547 ( .A1(n7144), .A2(n13213), .ZN(n7142) );
  INV_X1 U7548 ( .A(n11427), .ZN(n6646) );
  OAI21_X1 U7549 ( .B1(n7410), .B2(P2_IR_REG_27__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7409) );
  AND2_X1 U7550 ( .A1(n7393), .A2(n7370), .ZN(n7371) );
  INV_X1 U7551 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n7370) );
  INV_X1 U7552 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7373) );
  INV_X1 U7553 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7372) );
  INV_X1 U7554 ( .A(n13590), .ZN(n11577) );
  NAND2_X1 U7555 ( .A1(n12058), .A2(n11879), .ZN(n13754) );
  OAI21_X1 U7556 ( .B1(n8060), .B2(n8059), .A(n8058), .ZN(n8085) );
  NOR2_X1 U7557 ( .A1(n6900), .A2(n6901), .ZN(n6899) );
  AND2_X1 U7558 ( .A1(n6897), .A2(n6895), .ZN(n6894) );
  NAND2_X1 U7559 ( .A1(n6900), .A2(n6898), .ZN(n6897) );
  AND2_X1 U7560 ( .A1(n7804), .A2(n7790), .ZN(n7802) );
  AND2_X1 U7561 ( .A1(n7785), .A2(n7784), .ZN(n7786) );
  NAND2_X1 U7562 ( .A1(n7222), .A2(n7221), .ZN(n7633) );
  AOI21_X1 U7563 ( .B1(n7224), .B2(n7226), .A(n6539), .ZN(n7221) );
  NOR2_X1 U7564 ( .A1(n9443), .A2(n9444), .ZN(n9396) );
  NAND2_X1 U7565 ( .A1(n11314), .A2(n7318), .ZN(n7317) );
  NOR2_X1 U7566 ( .A1(n7319), .A2(n11557), .ZN(n7318) );
  INV_X1 U7567 ( .A(n7320), .ZN(n7319) );
  INV_X1 U7568 ( .A(n10200), .ZN(n9982) );
  AND2_X1 U7569 ( .A1(n11812), .A2(n12247), .ZN(n11813) );
  AND2_X1 U7570 ( .A1(n14089), .A2(n12101), .ZN(n12102) );
  NOR2_X1 U7571 ( .A1(n14652), .A2(n10720), .ZN(n14651) );
  NAND2_X1 U7572 ( .A1(n6939), .A2(n6943), .ZN(n6938) );
  INV_X1 U7573 ( .A(n6941), .ZN(n6939) );
  AOI21_X1 U7574 ( .B1(n14732), .B2(n14733), .A(n6942), .ZN(n6941) );
  INV_X1 U7575 ( .A(n10634), .ZN(n6942) );
  INV_X1 U7576 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8223) );
  AOI21_X1 U7577 ( .B1(n14072), .B2(n12598), .A(n12599), .ZN(n12622) );
  AND2_X1 U7578 ( .A1(n12281), .A2(n12283), .ZN(n12669) );
  XNOR2_X1 U7579 ( .A(n12491), .B(n12538), .ZN(n12695) );
  AOI21_X1 U7580 ( .B1(n11799), .B2(n12126), .A(n8521), .ZN(n12762) );
  AND2_X1 U7581 ( .A1(n12385), .A2(n12764), .ZN(n8521) );
  AND4_X1 U7582 ( .A1(n8536), .A2(n8535), .A3(n8534), .A4(n8533), .ZN(n12478)
         );
  NAND2_X1 U7583 ( .A1(n8690), .A2(n6805), .ZN(n6804) );
  AND2_X1 U7584 ( .A1(n12213), .A2(n8689), .ZN(n6805) );
  NAND2_X1 U7585 ( .A1(n8496), .A2(n8495), .ZN(n12254) );
  XNOR2_X1 U7586 ( .A(n6816), .B(n8240), .ZN(n8680) );
  NAND2_X1 U7587 ( .A1(n8239), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6816) );
  NAND2_X1 U7588 ( .A1(n8232), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8234) );
  NAND2_X1 U7589 ( .A1(n6675), .A2(n6673), .ZN(n8648) );
  NAND2_X1 U7590 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n6674), .ZN(n6673) );
  OR2_X1 U7591 ( .A1(n8634), .A2(n8635), .ZN(n6675) );
  NAND2_X1 U7592 ( .A1(n8214), .A2(n8213), .ZN(n8539) );
  NAND2_X1 U7593 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n10457), .ZN(n8213) );
  OAI21_X1 U7594 ( .B1(n7163), .B2(n6492), .A(n6682), .ZN(n8204) );
  INV_X1 U7595 ( .A(n6683), .ZN(n6682) );
  NAND2_X1 U7596 ( .A1(n8201), .A2(n8200), .ZN(n8299) );
  NAND2_X1 U7597 ( .A1(n7163), .A2(n6468), .ZN(n8201) );
  AOI21_X1 U7598 ( .B1(n6709), .B2(n6707), .A(n12920), .ZN(n6706) );
  INV_X1 U7599 ( .A(n12965), .ZN(n6707) );
  NOR2_X1 U7600 ( .A1(n13120), .A2(n13131), .ZN(n6637) );
  AND4_X1 U7601 ( .A1(n7998), .A2(n7997), .A3(n7996), .A4(n7995), .ZN(n12968)
         );
  XNOR2_X1 U7602 ( .A(n11734), .B(n11744), .ZN(n14513) );
  NAND2_X1 U7603 ( .A1(n6981), .A2(n6979), .ZN(n13119) );
  AOI21_X1 U7604 ( .B1(n6982), .B2(n6984), .A(n6980), .ZN(n6979) );
  INV_X1 U7605 ( .A(n13120), .ZN(n6980) );
  AND2_X1 U7606 ( .A1(n12037), .A2(n8136), .ZN(n13120) );
  OR2_X1 U7607 ( .A1(n13315), .A2(n13048), .ZN(n8136) );
  NAND2_X1 U7608 ( .A1(n13189), .A2(n6662), .ZN(n6656) );
  XNOR2_X1 U7609 ( .A(n13349), .B(n12928), .ZN(n13213) );
  AOI21_X1 U7610 ( .B1(n7005), .B2(n7004), .A(n6524), .ZN(n7003) );
  INV_X1 U7611 ( .A(n12030), .ZN(n7004) );
  AND2_X1 U7612 ( .A1(n13359), .A2(n12007), .ZN(n7148) );
  NAND2_X1 U7613 ( .A1(n6667), .A2(n6665), .ZN(n13236) );
  INV_X1 U7614 ( .A(n6666), .ZN(n6665) );
  OAI22_X1 U7615 ( .A1(n13254), .A2(n6671), .B1(n13056), .B2(n13262), .ZN(
        n6666) );
  OAI21_X1 U7616 ( .B1(n11210), .B2(n7011), .A(n6540), .ZN(n11711) );
  INV_X1 U7617 ( .A(n7012), .ZN(n7011) );
  INV_X1 U7618 ( .A(n7019), .ZN(n7016) );
  NAND2_X1 U7619 ( .A1(n10847), .A2(n10846), .ZN(n10850) );
  NAND2_X1 U7620 ( .A1(n10511), .A2(n10510), .ZN(n10947) );
  NAND2_X1 U7621 ( .A1(n6973), .A2(n10285), .ZN(n10506) );
  NAND2_X1 U7622 ( .A1(n9872), .A2(n9871), .ZN(n13284) );
  OR2_X1 U7623 ( .A1(n7426), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n6608) );
  XNOR2_X1 U7624 ( .A(n7385), .B(P2_IR_REG_29__SCAN_IN), .ZN(n7386) );
  NOR2_X1 U7625 ( .A1(n11252), .A2(n7043), .ZN(n7042) );
  INV_X1 U7626 ( .A(n7343), .ZN(n7043) );
  NAND2_X1 U7627 ( .A1(n9559), .A2(n9504), .ZN(n9270) );
  OR2_X1 U7628 ( .A1(n11902), .A2(n11901), .ZN(n11903) );
  NAND2_X1 U7629 ( .A1(n9301), .A2(n9308), .ZN(n9328) );
  NAND2_X1 U7630 ( .A1(n13927), .A2(n13452), .ZN(n6752) );
  AOI21_X1 U7631 ( .B1(n6748), .B2(n6746), .A(n6543), .ZN(n6745) );
  INV_X1 U7632 ( .A(n6499), .ZN(n6746) );
  OR2_X1 U7633 ( .A1(n13784), .A2(n13799), .ZN(n7352) );
  NOR2_X1 U7634 ( .A1(n13785), .A2(n7303), .ZN(n7302) );
  INV_X1 U7635 ( .A(n11858), .ZN(n7303) );
  NOR2_X1 U7636 ( .A1(n13897), .A2(n7298), .ZN(n7297) );
  INV_X1 U7637 ( .A(n11846), .ZN(n7298) );
  AND2_X1 U7638 ( .A1(n11547), .A2(n11545), .ZN(n7296) );
  INV_X1 U7639 ( .A(n8895), .ZN(n9271) );
  AND2_X1 U7640 ( .A1(n11231), .A2(n11229), .ZN(n7278) );
  XNOR2_X1 U7641 ( .A(n7953), .B(n8235), .ZN(n9161) );
  INV_X1 U7642 ( .A(n12536), .ZN(n12671) );
  NAND2_X2 U7643 ( .A1(n7941), .A2(n7940), .ZN(n13344) );
  OAI21_X1 U7644 ( .B1(n13091), .B2(n14536), .A(n6769), .ZN(n6768) );
  NAND2_X1 U7645 ( .A1(n13092), .A2(n14542), .ZN(n6769) );
  OAI21_X1 U7646 ( .B1(n9261), .B2(n9260), .A(n9259), .ZN(n9355) );
  NAND2_X1 U7647 ( .A1(n7531), .A2(n7533), .ZN(n7250) );
  NAND2_X1 U7648 ( .A1(n8958), .A2(n8957), .ZN(n7059) );
  AND2_X1 U7649 ( .A1(n8960), .A2(n7062), .ZN(n7058) );
  NAND2_X1 U7650 ( .A1(n7089), .A2(n8907), .ZN(n7088) );
  NOR2_X1 U7651 ( .A1(n7060), .A2(n7057), .ZN(n7056) );
  NOR2_X1 U7652 ( .A1(n8973), .A2(n8974), .ZN(n7060) );
  INV_X1 U7653 ( .A(n8957), .ZN(n7057) );
  AOI21_X1 U7654 ( .B1(n7052), .B2(n7051), .A(n6531), .ZN(n7050) );
  INV_X1 U7655 ( .A(n9064), .ZN(n7051) );
  OR2_X1 U7656 ( .A1(n9063), .A2(n7049), .ZN(n7048) );
  INV_X1 U7657 ( .A(n9281), .ZN(n7049) );
  NAND2_X1 U7658 ( .A1(n7075), .A2(n7073), .ZN(n9108) );
  AOI21_X1 U7659 ( .B1(n7076), .B2(n7079), .A(n7074), .ZN(n7073) );
  AND2_X1 U7660 ( .A1(n9083), .A2(n7080), .ZN(n7079) );
  NOR2_X1 U7661 ( .A1(n9182), .A2(n9179), .ZN(n7086) );
  NAND2_X1 U7662 ( .A1(n9182), .A2(n9179), .ZN(n7085) );
  MUX2_X1 U7663 ( .A(n13049), .B(n8135), .S(n6460), .Z(n8050) );
  INV_X1 U7664 ( .A(n7219), .ZN(n7218) );
  OAI21_X1 U7665 ( .B1(n7703), .B2(n7220), .A(n7725), .ZN(n7219) );
  AND2_X1 U7666 ( .A1(n7218), .A2(n6740), .ZN(n6739) );
  NAND2_X1 U7667 ( .A1(n7679), .A2(n7678), .ZN(n6740) );
  OAI21_X1 U7668 ( .B1(n7900), .B2(n7248), .A(n7244), .ZN(n6619) );
  AOI21_X1 U7669 ( .B1(n7247), .B2(n7249), .A(n7245), .ZN(n7244) );
  INV_X1 U7670 ( .A(n7959), .ZN(n7245) );
  INV_X1 U7671 ( .A(n6909), .ZN(n6908) );
  OAI21_X1 U7672 ( .B1(n7802), .B2(n6910), .A(n7826), .ZN(n6909) );
  INV_X1 U7673 ( .A(n7804), .ZN(n6910) );
  AND2_X1 U7674 ( .A1(n6736), .A2(n7215), .ZN(n6735) );
  AOI21_X1 U7675 ( .B1(n7218), .B2(n7220), .A(n7216), .ZN(n7215) );
  NAND2_X1 U7676 ( .A1(n6739), .A2(n6737), .ZN(n6736) );
  INV_X1 U7677 ( .A(n7727), .ZN(n7216) );
  INV_X1 U7678 ( .A(n6739), .ZN(n6738) );
  OAI211_X1 U7679 ( .C1(n6810), .C2(n12274), .A(n7179), .B(n12687), .ZN(n7177)
         );
  NAND2_X1 U7680 ( .A1(n12276), .A2(n12695), .ZN(n7179) );
  NAND2_X1 U7681 ( .A1(n6627), .A2(n6512), .ZN(n12276) );
  INV_X1 U7682 ( .A(n7160), .ZN(n7159) );
  OAI21_X1 U7683 ( .B1(n8646), .B2(n12283), .A(n12288), .ZN(n7160) );
  AND2_X1 U7684 ( .A1(n12280), .A2(n12294), .ZN(n7162) );
  INV_X1 U7685 ( .A(n8202), .ZN(n7190) );
  NOR2_X1 U7686 ( .A1(n7071), .A2(n9225), .ZN(n7072) );
  NAND2_X1 U7687 ( .A1(n7071), .A2(n9225), .ZN(n7070) );
  NAND2_X1 U7688 ( .A1(n7072), .A2(n7070), .ZN(n7068) );
  OAI21_X1 U7689 ( .B1(n7680), .B2(n6738), .A(n6735), .ZN(n7781) );
  NOR2_X1 U7690 ( .A1(n7656), .A2(n7631), .ZN(n6912) );
  INV_X1 U7691 ( .A(n7635), .ZN(n6914) );
  NAND2_X1 U7692 ( .A1(n14634), .A2(n10647), .ZN(n10649) );
  NAND2_X1 U7693 ( .A1(n14671), .A2(n10651), .ZN(n10652) );
  NAND2_X1 U7694 ( .A1(n14715), .A2(n10654), .ZN(n10655) );
  NAND2_X1 U7695 ( .A1(n11197), .A2(n6596), .ZN(n11199) );
  NAND2_X1 U7696 ( .A1(n11470), .A2(n11471), .ZN(n11630) );
  OAI21_X1 U7697 ( .B1(n12682), .B2(n6822), .A(n8633), .ZN(n6821) );
  NAND2_X1 U7698 ( .A1(n12831), .A2(n12415), .ZN(n8633) );
  INV_X1 U7699 ( .A(n6845), .ZN(n6844) );
  AOI21_X1 U7700 ( .B1(n6845), .B2(n8577), .A(n8602), .ZN(n6843) );
  NOR2_X1 U7701 ( .A1(n6846), .A2(n12142), .ZN(n6845) );
  INV_X1 U7702 ( .A(n6848), .ZN(n6846) );
  OR2_X1 U7703 ( .A1(n12505), .A2(n12500), .ZN(n12143) );
  AND2_X1 U7704 ( .A1(n12505), .A2(n12500), .ZN(n12144) );
  INV_X1 U7705 ( .A(n6839), .ZN(n6838) );
  OAI21_X1 U7706 ( .B1(n6840), .B2(n11599), .A(n8503), .ZN(n6839) );
  OR2_X1 U7707 ( .A1(n12254), .A2(n12544), .ZN(n8503) );
  INV_X1 U7708 ( .A(n7363), .ZN(n6840) );
  INV_X1 U7709 ( .A(n12251), .ZN(n6790) );
  OAI21_X1 U7710 ( .B1(n12244), .B2(n6790), .A(n12127), .ZN(n6789) );
  INV_X1 U7711 ( .A(n6490), .ZN(n6828) );
  NAND2_X1 U7712 ( .A1(n12556), .A2(n14782), .ZN(n12179) );
  AND2_X1 U7713 ( .A1(n8728), .A2(n8740), .ZN(n8742) );
  AND2_X1 U7714 ( .A1(n7334), .A2(n8233), .ZN(n7333) );
  INV_X1 U7715 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8658) );
  NOR2_X1 U7716 ( .A1(n7176), .A2(n9828), .ZN(n7174) );
  INV_X1 U7717 ( .A(n8207), .ZN(n7172) );
  NAND2_X1 U7718 ( .A1(n6681), .A2(n6679), .ZN(n8206) );
  NAND2_X1 U7719 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n6680), .ZN(n6679) );
  NAND2_X1 U7720 ( .A1(n8443), .A2(n8441), .ZN(n6681) );
  INV_X1 U7721 ( .A(n7184), .ZN(n7183) );
  OAI21_X1 U7722 ( .B1(n8407), .B2(n7185), .A(n8422), .ZN(n7184) );
  INV_X1 U7723 ( .A(n8205), .ZN(n7185) );
  OAI21_X1 U7724 ( .B1(n6468), .B2(n6492), .A(n7188), .ZN(n6683) );
  INV_X1 U7725 ( .A(n7189), .ZN(n7188) );
  OAI21_X1 U7726 ( .B1(n8297), .B2(n7190), .A(n8312), .ZN(n7189) );
  INV_X1 U7727 ( .A(n9680), .ZN(n6764) );
  NAND2_X1 U7728 ( .A1(n6764), .A2(n6762), .ZN(n6761) );
  INV_X1 U7729 ( .A(n9642), .ZN(n6762) );
  NAND2_X1 U7730 ( .A1(n7134), .A2(n6986), .ZN(n7136) );
  OAI21_X1 U7731 ( .B1(n12034), .B2(n6994), .A(n13174), .ZN(n6993) );
  INV_X1 U7732 ( .A(n12035), .ZN(n6994) );
  AND2_X1 U7733 ( .A1(n6664), .A2(n6663), .ZN(n6662) );
  INV_X1 U7734 ( .A(n13174), .ZN(n6663) );
  INV_X1 U7735 ( .A(n6660), .ZN(n6659) );
  AOI21_X1 U7736 ( .B1(n6660), .B2(n6658), .A(n13161), .ZN(n6657) );
  INV_X1 U7737 ( .A(n6662), .ZN(n6658) );
  INV_X1 U7738 ( .A(n7003), .ZN(n6999) );
  OAI21_X1 U7739 ( .B1(n11213), .B2(n6646), .A(n11722), .ZN(n6645) );
  NAND2_X1 U7740 ( .A1(n6651), .A2(n6653), .ZN(n6650) );
  INV_X1 U7741 ( .A(n10980), .ZN(n6653) );
  AND2_X1 U7742 ( .A1(n10982), .A2(n6652), .ZN(n6651) );
  OR2_X1 U7743 ( .A1(n10849), .A2(n6653), .ZN(n6652) );
  NAND2_X1 U7744 ( .A1(n7411), .A2(n7408), .ZN(n7259) );
  AND2_X1 U7745 ( .A1(n13458), .A2(n7035), .ZN(n7034) );
  OR2_X1 U7746 ( .A1(n13527), .A2(n7036), .ZN(n7035) );
  INV_X1 U7747 ( .A(n12328), .ZN(n7036) );
  NAND2_X1 U7748 ( .A1(n9305), .A2(n9302), .ZN(n9311) );
  AND2_X1 U7749 ( .A1(n8817), .A2(n9747), .ZN(n7045) );
  INV_X1 U7750 ( .A(n12049), .ZN(n6751) );
  AND2_X1 U7751 ( .A1(n13562), .A2(n13778), .ZN(n11860) );
  OR2_X1 U7752 ( .A1(n12049), .A2(n12044), .ZN(n6750) );
  AOI21_X1 U7753 ( .B1(n6728), .B2(n11876), .A(n6727), .ZN(n6871) );
  INV_X1 U7754 ( .A(n6873), .ZN(n6728) );
  INV_X1 U7755 ( .A(n13813), .ZN(n6727) );
  NOR2_X1 U7756 ( .A1(n13960), .A2(n6886), .ZN(n6885) );
  INV_X1 U7757 ( .A(n6887), .ZN(n6886) );
  AOI21_X1 U7758 ( .B1(n7271), .B2(n6878), .A(n6877), .ZN(n6876) );
  INV_X1 U7759 ( .A(n11866), .ZN(n6877) );
  INV_X1 U7760 ( .A(n7276), .ZN(n7275) );
  OAI21_X1 U7761 ( .B1(n11654), .B2(n7277), .A(n11863), .ZN(n7276) );
  NOR2_X1 U7762 ( .A1(n7277), .A2(n6880), .ZN(n6879) );
  INV_X1 U7763 ( .A(n11540), .ZN(n6880) );
  OR2_X1 U7764 ( .A1(n14171), .A2(n7295), .ZN(n7294) );
  INV_X1 U7765 ( .A(n11228), .ZN(n7295) );
  INV_X1 U7766 ( .A(n10150), .ZN(n7285) );
  INV_X1 U7767 ( .A(n13596), .ZN(n10175) );
  NAND2_X1 U7768 ( .A1(n6732), .A2(SI_20_), .ZN(n7900) );
  AND2_X1 U7769 ( .A1(n6562), .A2(n8797), .ZN(n7081) );
  NAND2_X1 U7770 ( .A1(n6725), .A2(n7855), .ZN(n7876) );
  NAND2_X1 U7771 ( .A1(n7854), .A2(SI_18_), .ZN(n7855) );
  NAND2_X1 U7772 ( .A1(n7852), .A2(n7851), .ZN(n6725) );
  OAI21_X1 U7773 ( .B1(n7680), .B2(n7679), .A(n7678), .ZN(n7704) );
  NOR2_X1 U7774 ( .A1(n8980), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n8983) );
  NAND2_X1 U7775 ( .A1(n6694), .A2(n7492), .ZN(n6695) );
  INV_X1 U7776 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14930) );
  XNOR2_X1 U7777 ( .A(n9391), .B(n14668), .ZN(n9433) );
  OAI22_X1 U7778 ( .A1(n9440), .A2(n9394), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n14687), .ZN(n9395) );
  INV_X1 U7779 ( .A(n11557), .ZN(n7316) );
  NAND2_X1 U7780 ( .A1(n10823), .A2(n10822), .ZN(n7332) );
  NOR2_X1 U7781 ( .A1(n6522), .A2(n7321), .ZN(n7320) );
  INV_X1 U7782 ( .A(n11313), .ZN(n7321) );
  INV_X1 U7783 ( .A(n11374), .ZN(n11358) );
  AOI21_X1 U7784 ( .B1(n7325), .B2(n7323), .A(n6549), .ZN(n7322) );
  INV_X1 U7785 ( .A(n7325), .ZN(n7324) );
  OR2_X1 U7786 ( .A1(n11673), .A2(n11674), .ZN(n7313) );
  NAND2_X1 U7787 ( .A1(n12295), .A2(n7157), .ZN(n12293) );
  AND2_X1 U7788 ( .A1(n12090), .A2(n12089), .ZN(n12640) );
  AND4_X1 U7789 ( .A1(n8520), .A2(n8519), .A3(n8518), .A4(n8517), .ZN(n12386)
         );
  NOR2_X1 U7790 ( .A1(n10481), .A2(n8329), .ZN(n10480) );
  OR2_X1 U7791 ( .A1(n10480), .A2(n7101), .ZN(n7100) );
  AND2_X1 U7792 ( .A1(n10322), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7101) );
  AND2_X1 U7793 ( .A1(n7102), .A2(n7100), .ZN(n10579) );
  INV_X1 U7794 ( .A(n10324), .ZN(n7102) );
  XNOR2_X1 U7795 ( .A(n10649), .B(n14661), .ZN(n14659) );
  NAND2_X1 U7796 ( .A1(n14673), .A2(n14672), .ZN(n14671) );
  XNOR2_X1 U7797 ( .A(n10652), .B(n10613), .ZN(n14701) );
  OAI21_X1 U7798 ( .B1(n14651), .B2(n7120), .A(n7122), .ZN(n10587) );
  NAND2_X1 U7799 ( .A1(n14669), .A2(n10586), .ZN(n7122) );
  NAND2_X1 U7800 ( .A1(n7121), .A2(n10586), .ZN(n7120) );
  NAND2_X1 U7801 ( .A1(n14716), .A2(n14717), .ZN(n14715) );
  XNOR2_X1 U7802 ( .A(n10655), .B(n10625), .ZN(n14745) );
  NAND2_X1 U7803 ( .A1(n10660), .A2(n10659), .ZN(n11197) );
  NAND2_X1 U7804 ( .A1(n14734), .A2(n6577), .ZN(n6937) );
  XNOR2_X1 U7805 ( .A(n11199), .B(n11185), .ZN(n11299) );
  NAND2_X1 U7806 ( .A1(n6933), .A2(n6932), .ZN(n11303) );
  NAND2_X1 U7807 ( .A1(n6936), .A2(n6934), .ZN(n6932) );
  NAND2_X1 U7808 ( .A1(n11201), .A2(n11202), .ZN(n11470) );
  AOI21_X1 U7809 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n11469), .A(n11467), .ZN(
        n11625) );
  XNOR2_X1 U7810 ( .A(n11630), .B(n11626), .ZN(n11472) );
  OR2_X1 U7811 ( .A1(n11468), .A2(n8452), .ZN(n7115) );
  NOR2_X1 U7812 ( .A1(n11643), .A2(n6584), .ZN(n12570) );
  NAND3_X1 U7813 ( .A1(n6815), .A2(n7328), .A3(n8226), .ZN(n8507) );
  AND2_X1 U7814 ( .A1(n8222), .A2(n8227), .ZN(n7328) );
  NAND2_X1 U7815 ( .A1(n6948), .A2(n6947), .ZN(n6946) );
  NAND2_X1 U7816 ( .A1(n12587), .A2(n14025), .ZN(n6947) );
  INV_X1 U7817 ( .A(n14074), .ZN(n6948) );
  OR2_X1 U7818 ( .A1(n12588), .A2(n12589), .ZN(n6945) );
  AOI21_X1 U7819 ( .B1(n6799), .B2(n6801), .A(n6797), .ZN(n6796) );
  INV_X1 U7820 ( .A(n12283), .ZN(n6797) );
  NAND2_X1 U7821 ( .A1(n12688), .A2(n12687), .ZN(n12686) );
  NOR2_X1 U7822 ( .A1(n6809), .A2(n6808), .ZN(n6807) );
  INV_X1 U7823 ( .A(n12150), .ZN(n6808) );
  NAND2_X1 U7824 ( .A1(n12761), .A2(n8537), .ZN(n12749) );
  OR2_X1 U7825 ( .A1(n12774), .A2(n12478), .ZN(n12150) );
  INV_X1 U7826 ( .A(n11599), .ZN(n12244) );
  NAND2_X1 U7827 ( .A1(n6834), .A2(n6473), .ZN(n6833) );
  NAND2_X1 U7828 ( .A1(n11289), .A2(n6490), .ZN(n6832) );
  AND4_X1 U7829 ( .A1(n8437), .A2(n8436), .A3(n8435), .A4(n8434), .ZN(n11503)
         );
  AOI21_X1 U7830 ( .B1(n6793), .B2(n6795), .A(n6517), .ZN(n6792) );
  NAND2_X1 U7831 ( .A1(n9567), .A2(n9964), .ZN(n12308) );
  OR2_X1 U7832 ( .A1(n12096), .A2(n9502), .ZN(n7308) );
  OR2_X1 U7833 ( .A1(n12303), .A2(n12294), .ZN(n10129) );
  NAND2_X1 U7834 ( .A1(n12098), .A2(n12097), .ZN(n14089) );
  NAND2_X1 U7835 ( .A1(n12867), .A2(n8353), .ZN(n12098) );
  NAND2_X1 U7836 ( .A1(n8514), .A2(n8513), .ZN(n12385) );
  AND3_X1 U7837 ( .A1(n8429), .A2(n8428), .A3(n8427), .ZN(n14105) );
  NAND2_X1 U7838 ( .A1(n8682), .A2(n12288), .ZN(n14760) );
  NAND2_X1 U7839 ( .A1(n8243), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8244) );
  AOI21_X1 U7840 ( .B1(n8620), .B2(n8619), .A(n8618), .ZN(n8634) );
  AND2_X1 U7841 ( .A1(n11616), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8618) );
  NOR2_X2 U7842 ( .A1(n8507), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n8509) );
  NAND2_X1 U7843 ( .A1(n6598), .A2(n7194), .ZN(n7191) );
  INV_X1 U7844 ( .A(n7195), .ZN(n7192) );
  NAND2_X1 U7845 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n12382), .ZN(n7195) );
  OR2_X1 U7846 ( .A1(n8668), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n8713) );
  NAND2_X1 U7847 ( .A1(n8219), .A2(n8218), .ZN(n8566) );
  AND2_X1 U7848 ( .A1(n8659), .A2(n8658), .ZN(n8664) );
  NAND2_X1 U7849 ( .A1(n8664), .A2(n8666), .ZN(n8668) );
  XNOR2_X1 U7850 ( .A(n8217), .B(n10994), .ZN(n8553) );
  OAI21_X1 U7851 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(n10097), .A(n8212), .ZN(
        n8524) );
  OAI21_X1 U7852 ( .B1(P2_DATAO_REG_15__SCAN_IN), .B2(n10142), .A(n8209), .ZN(
        n8491) );
  NAND2_X1 U7853 ( .A1(n8206), .A2(n9886), .ZN(n8207) );
  XNOR2_X1 U7854 ( .A(n8206), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8446) );
  XNOR2_X1 U7855 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8297) );
  AND2_X1 U7856 ( .A1(n7167), .A2(n8199), .ZN(n7166) );
  NAND2_X1 U7857 ( .A1(n7168), .A2(n8198), .ZN(n7167) );
  INV_X1 U7858 ( .A(n8197), .ZN(n7168) );
  NOR2_X1 U7859 ( .A1(n7169), .A2(n7165), .ZN(n7164) );
  INV_X1 U7860 ( .A(n8198), .ZN(n7169) );
  AND2_X1 U7861 ( .A1(n8385), .A2(n8259), .ZN(n8387) );
  INV_X1 U7862 ( .A(n8149), .ZN(n10282) );
  NAND2_X1 U7863 ( .A1(n10899), .A2(n10898), .ZN(n6723) );
  NAND2_X1 U7864 ( .A1(n10735), .A2(n10734), .ZN(n10740) );
  NOR2_X1 U7865 ( .A1(n7200), .A2(n7199), .ZN(n7198) );
  INV_X1 U7866 ( .A(n6723), .ZN(n7199) );
  INV_X1 U7867 ( .A(n10866), .ZN(n7200) );
  NAND2_X1 U7868 ( .A1(n10752), .A2(n10744), .ZN(n6721) );
  XNOR2_X1 U7869 ( .A(n6459), .B(n10026), .ZN(n11956) );
  OR4_X1 U7870 ( .A1(n13198), .A2(n13213), .A3(n13222), .A4(n8159), .ZN(n8160)
         );
  OR4_X1 U7871 ( .A1(n13246), .A2(n13254), .A3(n12027), .A4(n8158), .ZN(n8159)
         );
  AND2_X1 U7872 ( .A1(n12042), .A2(n13435), .ZN(n7485) );
  AND2_X1 U7873 ( .A1(n7387), .A2(n13435), .ZN(n7486) );
  XNOR2_X1 U7874 ( .A(n9647), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n14401) );
  NOR2_X1 U7875 ( .A1(n14415), .A2(n6774), .ZN(n14429) );
  AND2_X1 U7876 ( .A1(n14411), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6774) );
  OR2_X1 U7877 ( .A1(n14429), .A2(n14428), .ZN(n6773) );
  NOR2_X1 U7878 ( .A1(n9793), .A2(n9792), .ZN(n9791) );
  NOR2_X1 U7879 ( .A1(n6757), .A2(n6763), .ZN(n6756) );
  AND2_X1 U7880 ( .A1(n9947), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6763) );
  INV_X1 U7881 ( .A(n6759), .ZN(n6757) );
  OR2_X1 U7882 ( .A1(n14472), .A2(n14473), .ZN(n6779) );
  NAND2_X1 U7883 ( .A1(n11732), .A2(n11733), .ZN(n11734) );
  NAND2_X1 U7884 ( .A1(n14513), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n14512) );
  INV_X1 U7885 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7392) );
  NAND2_X1 U7886 ( .A1(n8072), .A2(n8071), .ZN(n13103) );
  NAND2_X1 U7887 ( .A1(n8106), .A2(n8105), .ZN(n13097) );
  NAND2_X1 U7888 ( .A1(n6550), .A2(n7132), .ZN(n7129) );
  AND2_X1 U7889 ( .A1(n7132), .A2(n12012), .ZN(n7130) );
  NAND2_X1 U7890 ( .A1(n13130), .A2(n13118), .ZN(n13113) );
  INV_X1 U7891 ( .A(n8135), .ZN(n13128) );
  NAND2_X1 U7892 ( .A1(n7131), .A2(n12010), .ZN(n7134) );
  NAND2_X1 U7893 ( .A1(n13140), .A2(n12012), .ZN(n7131) );
  AOI21_X1 U7894 ( .B1(n6493), .B2(n6662), .A(n6661), .ZN(n6660) );
  NOR2_X1 U7895 ( .A1(n13184), .A2(n13052), .ZN(n6661) );
  OR2_X1 U7896 ( .A1(n13344), .A2(n12986), .ZN(n6664) );
  INV_X1 U7897 ( .A(n7147), .ZN(n7140) );
  NAND2_X1 U7898 ( .A1(n13236), .A2(n7146), .ZN(n7143) );
  INV_X1 U7899 ( .A(n7144), .ZN(n7141) );
  AND2_X1 U7900 ( .A1(n7125), .A2(n7126), .ZN(n6670) );
  NAND2_X1 U7901 ( .A1(n13274), .A2(n13057), .ZN(n7125) );
  NAND2_X1 U7902 ( .A1(n12028), .A2(n12027), .ZN(n13275) );
  NAND2_X1 U7903 ( .A1(n13282), .A2(n7362), .ZN(n7127) );
  NAND2_X1 U7904 ( .A1(n13295), .A2(n13058), .ZN(n7126) );
  OAI21_X1 U7905 ( .B1(n6486), .B2(n6997), .A(n6995), .ZN(n13296) );
  INV_X1 U7906 ( .A(n6996), .ZN(n6995) );
  OAI21_X1 U7907 ( .B1(n6998), .B2(n6997), .A(n13297), .ZN(n6996) );
  INV_X1 U7908 ( .A(n12024), .ZN(n6997) );
  NAND2_X1 U7909 ( .A1(n13286), .A2(n13295), .ZN(n13287) );
  AND2_X1 U7910 ( .A1(n11763), .A2(n11770), .ZN(n6998) );
  AOI21_X1 U7911 ( .B1(n7015), .B2(n7013), .A(n6507), .ZN(n7012) );
  INV_X1 U7912 ( .A(n6544), .ZN(n7013) );
  OR2_X1 U7913 ( .A1(n13398), .A2(n11990), .ZN(n11427) );
  NAND2_X1 U7914 ( .A1(n11136), .A2(n6931), .ZN(n11432) );
  NAND2_X1 U7915 ( .A1(n7020), .A2(n8138), .ZN(n7019) );
  XNOR2_X1 U7916 ( .A(n13398), .B(n13062), .ZN(n11213) );
  NOR2_X2 U7917 ( .A1(n11137), .A2(n13403), .ZN(n11136) );
  OAI21_X1 U7918 ( .B1(n10850), .B2(n6653), .A(n6651), .ZN(n11067) );
  NAND2_X1 U7919 ( .A1(n10850), .A2(n10849), .ZN(n10981) );
  NAND2_X1 U7920 ( .A1(n6978), .A2(n6518), .ZN(n10975) );
  NAND2_X1 U7921 ( .A1(n6972), .A2(n10508), .ZN(n10668) );
  NAND2_X1 U7922 ( .A1(n7124), .A2(n8146), .ZN(n8147) );
  OAI21_X1 U7923 ( .B1(n9891), .B2(n9888), .A(n9887), .ZN(n10280) );
  INV_X1 U7924 ( .A(n13284), .ZN(n13268) );
  CLKBUF_X1 U7925 ( .A(n10022), .Z(n9868) );
  INV_X1 U7926 ( .A(n12023), .ZN(n13310) );
  NAND2_X1 U7927 ( .A1(n7902), .A2(n7901), .ZN(n13354) );
  NAND2_X1 U7928 ( .A1(n7831), .A2(n7830), .ZN(n13369) );
  NAND2_X1 U7929 ( .A1(n6719), .A2(n7592), .ZN(n10890) );
  NAND2_X1 U7930 ( .A1(n9570), .A2(n7960), .ZN(n6719) );
  NAND2_X1 U7931 ( .A1(n7501), .A2(n7500), .ZN(n14566) );
  OR2_X1 U7932 ( .A1(n8104), .A2(n9529), .ZN(n7461) );
  INV_X1 U7933 ( .A(n14592), .ZN(n14567) );
  NAND2_X1 U7934 ( .A1(n9864), .A2(n9863), .ZN(n10007) );
  INV_X1 U7935 ( .A(n7259), .ZN(n7258) );
  INV_X1 U7936 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7257) );
  AND2_X1 U7937 ( .A1(n7371), .A2(n7381), .ZN(n7150) );
  INV_X1 U7938 ( .A(n7791), .ZN(n7213) );
  OR2_X1 U7939 ( .A1(n7636), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8174) );
  OAI21_X1 U7940 ( .B1(n8165), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8170) );
  INV_X1 U7941 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8169) );
  OR2_X1 U7942 ( .A1(n7402), .A2(n14924), .ZN(n7403) );
  OR2_X1 U7943 ( .A1(n7709), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n7728) );
  NOR2_X1 U7944 ( .A1(n13483), .A2(n7038), .ZN(n7037) );
  INV_X1 U7945 ( .A(n12316), .ZN(n7038) );
  INV_X1 U7946 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8961) );
  OR2_X1 U7947 ( .A1(n9113), .A2(n9112), .ZN(n9127) );
  AND2_X1 U7948 ( .A1(n9754), .A2(n9549), .ZN(n9763) );
  XNOR2_X1 U7949 ( .A(n9328), .B(n9320), .ZN(n7269) );
  NAND2_X1 U7950 ( .A1(n7095), .A2(n9255), .ZN(n7094) );
  NAND2_X1 U7951 ( .A1(n11592), .A2(n11593), .ZN(n13701) );
  NAND2_X1 U7952 ( .A1(n9273), .A2(n9272), .ZN(n13738) );
  OR2_X1 U7953 ( .A1(n14004), .A2(n9270), .ZN(n9273) );
  INV_X1 U7954 ( .A(n12058), .ZN(n13753) );
  NOR2_X1 U7955 ( .A1(n13837), .A2(n6874), .ZN(n6873) );
  INV_X1 U7956 ( .A(n11873), .ZN(n6874) );
  NAND2_X1 U7957 ( .A1(n6868), .A2(n6871), .ZN(n13812) );
  OR2_X1 U7958 ( .A1(n11874), .A2(n6872), .ZN(n6868) );
  XNOR2_X1 U7959 ( .A(n13835), .B(n13583), .ZN(n13837) );
  INV_X1 U7960 ( .A(n11853), .ZN(n7301) );
  NAND2_X1 U7961 ( .A1(n11852), .A2(n11851), .ZN(n13856) );
  INV_X1 U7962 ( .A(n13858), .ZN(n11852) );
  NAND2_X1 U7963 ( .A1(n7273), .A2(n7275), .ZN(n14148) );
  NAND2_X1 U7964 ( .A1(n11541), .A2(n6879), .ZN(n7273) );
  NAND2_X1 U7965 ( .A1(n11340), .A2(n11339), .ZN(n11342) );
  INV_X1 U7966 ( .A(n11222), .ZN(n10791) );
  NAND2_X1 U7967 ( .A1(n13593), .A2(n10887), .ZN(n6867) );
  NAND2_X1 U7968 ( .A1(n10229), .A2(n10887), .ZN(n10358) );
  OAI21_X1 U7969 ( .B1(n13929), .B2(n14349), .A(n6890), .ZN(n6889) );
  AOI21_X1 U7970 ( .B1(n13927), .B2(n14345), .A(n13926), .ZN(n6890) );
  INV_X1 U7971 ( .A(n13562), .ZN(n13936) );
  NAND2_X1 U7972 ( .A1(n12366), .A2(n9911), .ZN(n14349) );
  OR2_X1 U7973 ( .A1(n9757), .A2(n9914), .ZN(n14371) );
  OR2_X1 U7974 ( .A1(n8101), .A2(n8100), .ZN(n8103) );
  OAI21_X1 U7975 ( .B1(n8015), .B2(n8014), .A(n7986), .ZN(n8001) );
  NAND2_X1 U7976 ( .A1(n7246), .A2(n7917), .ZN(n7953) );
  AOI22_X1 U7977 ( .A1(n7898), .A2(n6730), .B1(n6732), .B2(n6729), .ZN(n7246)
         );
  NOR2_X1 U7978 ( .A1(n7913), .A2(n7896), .ZN(n6730) );
  NOR2_X1 U7979 ( .A1(n7913), .A2(n10453), .ZN(n6729) );
  INV_X1 U7980 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8813) );
  NAND2_X1 U7981 ( .A1(n6907), .A2(n7804), .ZN(n7827) );
  NAND2_X1 U7982 ( .A1(n7803), .A2(n7802), .ZN(n6907) );
  XNOR2_X1 U7983 ( .A(n7726), .B(n7725), .ZN(n9827) );
  NAND2_X1 U7984 ( .A1(n7217), .A2(n7705), .ZN(n7726) );
  NAND2_X1 U7985 ( .A1(n7704), .A2(n7703), .ZN(n7217) );
  INV_X1 U7986 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8770) );
  CLKBUF_X1 U7987 ( .A(n8827), .Z(n8828) );
  NAND2_X1 U7988 ( .A1(n14035), .A2(n14034), .ZN(n6970) );
  OAI21_X1 U7989 ( .B1(n14036), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6505), .ZN(
        n6953) );
  NOR2_X1 U7990 ( .A1(n9412), .A2(n9411), .ZN(n9403) );
  NOR2_X1 U7991 ( .A1(n14050), .A2(n14051), .ZN(n9480) );
  AND4_X1 U7992 ( .A1(n8421), .A2(n8420), .A3(n8419), .A4(n8418), .ZN(n11315)
         );
  OR2_X1 U7993 ( .A1(n12389), .A2(n12478), .ZN(n12390) );
  AOI21_X1 U7994 ( .B1(n7312), .B2(n11674), .A(n6533), .ZN(n7309) );
  AND3_X1 U7995 ( .A1(n8319), .A2(n8318), .A3(n8317), .ZN(n10838) );
  INV_X1 U7996 ( .A(n12531), .ZN(n12509) );
  AND2_X1 U7997 ( .A1(n12304), .A2(n12303), .ZN(n12305) );
  XNOR2_X1 U7998 ( .A(n12138), .B(n12623), .ZN(n12140) );
  INV_X1 U7999 ( .A(n12307), .ZN(n7155) );
  INV_X1 U8000 ( .A(n11315), .ZN(n12548) );
  XNOR2_X1 U8001 ( .A(n11625), .B(n11626), .ZN(n11468) );
  NAND2_X1 U8002 ( .A1(n7103), .A2(n7104), .ZN(n14066) );
  INV_X1 U8003 ( .A(n14079), .ZN(n14083) );
  NOR2_X1 U8004 ( .A1(n12622), .A2(n6606), .ZN(n6783) );
  NAND2_X1 U8005 ( .A1(n6503), .A2(n6781), .ZN(n6780) );
  INV_X1 U8006 ( .A(n12634), .ZN(n6781) );
  NAND2_X1 U8007 ( .A1(n12681), .A2(n7364), .ZN(n12667) );
  NAND2_X1 U8008 ( .A1(n10455), .A2(n12623), .ZN(n12302) );
  AND2_X1 U8009 ( .A1(n9374), .A2(n9373), .ZN(n12078) );
  NOR2_X1 U8010 ( .A1(n6489), .A2(n9494), .ZN(n6852) );
  NOR2_X1 U8011 ( .A1(n6489), .A2(n14832), .ZN(n6853) );
  AND2_X1 U8012 ( .A1(n8582), .A2(n8581), .ZN(n12842) );
  NAND2_X1 U8013 ( .A1(n8465), .A2(n8464), .ZN(n11624) );
  INV_X1 U8014 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10321) );
  NAND2_X1 U8015 ( .A1(n6705), .A2(n6706), .ZN(n12946) );
  AOI21_X1 U8016 ( .B1(n6471), .B2(n6708), .A(n6548), .ZN(n6703) );
  INV_X1 U8017 ( .A(n7203), .ZN(n6713) );
  AOI21_X1 U8018 ( .B1(n7203), .B2(n7204), .A(n7202), .ZN(n7201) );
  AOI21_X1 U8019 ( .B1(n11172), .B2(n11159), .A(n6536), .ZN(n7203) );
  NAND2_X1 U8020 ( .A1(n7616), .A2(n7615), .ZN(n11090) );
  NAND2_X1 U8021 ( .A1(n7879), .A2(n7878), .ZN(n13359) );
  NAND2_X1 U8022 ( .A1(n7919), .A2(n7918), .ZN(n13349) );
  NAND2_X1 U8023 ( .A1(n6710), .A2(n6709), .ZN(n13032) );
  INV_X1 U8024 ( .A(n13023), .ZN(n13035) );
  NAND2_X1 U8025 ( .A1(n7763), .A2(n7762), .ZN(n13387) );
  OAI21_X1 U8026 ( .B1(n13211), .B2(n8077), .A(n7912), .ZN(n13012) );
  NOR2_X1 U8027 ( .A1(n14534), .A2(n13079), .ZN(n13080) );
  OAI21_X1 U8028 ( .B1(n13144), .B2(n6984), .A(n6982), .ZN(n13121) );
  AND2_X1 U8029 ( .A1(n6640), .A2(n6639), .ZN(n13317) );
  INV_X1 U8030 ( .A(n13111), .ZN(n6639) );
  NAND2_X1 U8031 ( .A1(n6642), .A2(n6641), .ZN(n6640) );
  NAND2_X1 U8032 ( .A1(n6643), .A2(n13120), .ZN(n6642) );
  NAND2_X1 U8033 ( .A1(n6991), .A2(n12035), .ZN(n13175) );
  NAND2_X1 U8034 ( .A1(n13199), .A2(n12034), .ZN(n6991) );
  INV_X1 U8035 ( .A(n8145), .ZN(n7124) );
  NAND2_X1 U8036 ( .A1(n14556), .A2(n10012), .ZN(n13245) );
  INV_X1 U8037 ( .A(n14556), .ZN(n14553) );
  AND2_X1 U8038 ( .A1(n10258), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14556) );
  NAND2_X1 U8039 ( .A1(n9237), .A2(n9236), .ZN(n13454) );
  NAND2_X1 U8040 ( .A1(n9033), .A2(n9032), .ZN(n14210) );
  NAND2_X1 U8041 ( .A1(n11570), .A2(n11569), .ZN(n6625) );
  INV_X1 U8042 ( .A(n7041), .ZN(n7040) );
  NAND2_X1 U8043 ( .A1(n14136), .A2(n7041), .ZN(n11788) );
  NAND2_X1 U8044 ( .A1(n9191), .A2(n9190), .ZN(n13805) );
  NAND2_X1 U8045 ( .A1(n9105), .A2(n9104), .ZN(n14180) );
  AND2_X1 U8046 ( .A1(n9328), .A2(n9327), .ZN(n9318) );
  NAND2_X1 U8047 ( .A1(n9264), .A2(n9263), .ZN(n13732) );
  AND2_X1 U8048 ( .A1(n8796), .A2(n8795), .ZN(n13919) );
  XNOR2_X1 U8049 ( .A(n6858), .B(n11878), .ZN(n13916) );
  OAI21_X1 U8050 ( .B1(n6743), .B2(n6742), .A(n6541), .ZN(n6858) );
  INV_X1 U8051 ( .A(n6745), .ZN(n6742) );
  NAND2_X1 U8052 ( .A1(n6961), .A2(n9455), .ZN(n14045) );
  NOR2_X1 U8053 ( .A1(n14046), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n6958) );
  NAND2_X1 U8054 ( .A1(n6959), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n6957) );
  NAND2_X1 U8055 ( .A1(n6956), .A2(n14046), .ZN(n6955) );
  NOR2_X1 U8056 ( .A1(n14245), .A2(n14244), .ZN(n14243) );
  XNOR2_X1 U8057 ( .A(n9486), .B(n9485), .ZN(n14020) );
  OR2_X1 U8058 ( .A1(n7505), .A2(n7504), .ZN(n7506) );
  INV_X1 U8059 ( .A(n7577), .ZN(n7261) );
  OAI21_X1 U8060 ( .B1(n9192), .B2(n10111), .A(n7066), .ZN(n7065) );
  INV_X1 U8061 ( .A(n8907), .ZN(n7090) );
  INV_X1 U8062 ( .A(n8938), .ZN(n7089) );
  NAND2_X1 U8063 ( .A1(n7624), .A2(n7623), .ZN(n7642) );
  AOI22_X1 U8064 ( .A1(n7061), .A2(n8973), .B1(n7054), .B2(n8974), .ZN(n7053)
         );
  NAND2_X1 U8065 ( .A1(n6496), .A2(n7056), .ZN(n7055) );
  NAND2_X1 U8066 ( .A1(n7059), .A2(n7058), .ZN(n7061) );
  NAND2_X1 U8067 ( .A1(n7237), .A2(n7236), .ZN(n7691) );
  NAND2_X1 U8068 ( .A1(n7667), .A2(n7669), .ZN(n7236) );
  NAND2_X1 U8069 ( .A1(n9008), .A2(n9005), .ZN(n7091) );
  NOR2_X1 U8070 ( .A1(n9005), .A2(n9008), .ZN(n7092) );
  NAND2_X1 U8071 ( .A1(n7234), .A2(n7233), .ZN(n7736) );
  NAND2_X1 U8072 ( .A1(n7714), .A2(n7716), .ZN(n7233) );
  INV_X1 U8073 ( .A(n9021), .ZN(n9024) );
  AOI21_X1 U8074 ( .B1(n12177), .B2(n12176), .A(n12175), .ZN(n12188) );
  OR2_X1 U8075 ( .A1(n12173), .A2(n12172), .ZN(n12177) );
  INV_X1 U8076 ( .A(n9081), .ZN(n7080) );
  AND2_X1 U8077 ( .A1(n7050), .A2(n7048), .ZN(n7046) );
  AND2_X1 U8078 ( .A1(n14155), .A2(n7077), .ZN(n7076) );
  NAND2_X1 U8079 ( .A1(n9081), .A2(n7078), .ZN(n7077) );
  NAND2_X1 U8080 ( .A1(n6622), .A2(n6621), .ZN(n9165) );
  NAND2_X1 U8081 ( .A1(n9152), .A2(n9154), .ZN(n6621) );
  AOI21_X1 U8082 ( .B1(n12250), .B2(n12249), .A(n6786), .ZN(n12256) );
  NAND2_X1 U8083 ( .A1(n7228), .A2(n7227), .ZN(n7882) );
  NAND2_X1 U8084 ( .A1(n7862), .A2(n7864), .ZN(n7227) );
  NAND2_X1 U8085 ( .A1(n7231), .A2(n7230), .ZN(n7922) );
  NAND2_X1 U8086 ( .A1(n7903), .A2(n7905), .ZN(n7230) );
  AOI21_X1 U8087 ( .B1(n7086), .B2(n7085), .A(n7084), .ZN(n7083) );
  INV_X1 U8088 ( .A(n9196), .ZN(n7084) );
  INV_X1 U8089 ( .A(n7678), .ZN(n6737) );
  INV_X1 U8090 ( .A(n7705), .ZN(n7220) );
  NAND2_X1 U8091 ( .A1(n6629), .A2(n6628), .ZN(n6627) );
  NOR2_X1 U8092 ( .A1(n12272), .A2(n12710), .ZN(n6628) );
  OR2_X1 U8093 ( .A1(n12270), .A2(n12271), .ZN(n6629) );
  OR2_X1 U8094 ( .A1(n12539), .A2(n12294), .ZN(n6626) );
  OR2_X1 U8095 ( .A1(n12114), .A2(n9987), .ZN(n12162) );
  NAND2_X1 U8096 ( .A1(n7942), .A2(n7944), .ZN(n7239) );
  AND2_X1 U8097 ( .A1(n8049), .A2(n8004), .ZN(n8021) );
  NOR2_X1 U8098 ( .A1(n13598), .A2(n8863), .ZN(n8861) );
  AND2_X1 U8099 ( .A1(n7986), .A2(SI_26_), .ZN(n6903) );
  INV_X1 U8100 ( .A(n8589), .ZN(n6688) );
  AND2_X1 U8101 ( .A1(n6594), .A2(n8591), .ZN(n6687) );
  OR2_X1 U8102 ( .A1(n7965), .A2(n7966), .ZN(n8020) );
  INV_X1 U8103 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7408) );
  INV_X1 U8104 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7478) );
  INV_X1 U8105 ( .A(n6879), .ZN(n6878) );
  NAND2_X1 U8106 ( .A1(n11653), .A2(n11656), .ZN(n7277) );
  AOI21_X1 U8107 ( .B1(n8014), .B2(n6903), .A(n6902), .ZN(n6901) );
  INV_X1 U8108 ( .A(n7999), .ZN(n6902) );
  AOI21_X1 U8109 ( .B1(n8014), .B2(n7986), .A(SI_26_), .ZN(n6900) );
  INV_X1 U8110 ( .A(n7986), .ZN(n6898) );
  NAND2_X1 U8111 ( .A1(n6901), .A2(n6896), .ZN(n6895) );
  INV_X1 U8112 ( .A(n6903), .ZN(n6896) );
  INV_X1 U8113 ( .A(n6619), .ZN(n6618) );
  NOR2_X1 U8114 ( .A1(n7248), .A2(n7896), .ZN(n6917) );
  NAND2_X1 U8115 ( .A1(n7856), .A2(n10044), .ZN(n7877) );
  AOI21_X1 U8116 ( .B1(n6908), .B2(n6910), .A(n6905), .ZN(n6904) );
  INV_X1 U8117 ( .A(n7828), .ZN(n6905) );
  NAND2_X1 U8118 ( .A1(n7805), .A2(n8511), .ZN(n7828) );
  AOI21_X1 U8119 ( .B1(n6735), .B2(n6738), .A(n6479), .ZN(n6734) );
  INV_X1 U8120 ( .A(n7783), .ZN(n6741) );
  INV_X1 U8121 ( .A(n7225), .ZN(n7224) );
  OAI21_X1 U8122 ( .B1(n7586), .B2(n7226), .A(n7611), .ZN(n7225) );
  INV_X1 U8123 ( .A(n7589), .ZN(n7226) );
  NAND2_X1 U8124 ( .A1(n7476), .A2(n7474), .ZN(n6698) );
  INV_X1 U8125 ( .A(n7476), .ZN(n6694) );
  INV_X1 U8126 ( .A(n7491), .ZN(n7492) );
  OAI21_X1 U8127 ( .B1(n7459), .B2(n9532), .A(n6617), .ZN(n7494) );
  NAND2_X1 U8128 ( .A1(n7459), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6617) );
  AND2_X1 U8129 ( .A1(n8743), .A2(n9563), .ZN(n9975) );
  INV_X1 U8130 ( .A(n12495), .ZN(n7323) );
  AND2_X1 U8131 ( .A1(n12290), .A2(n12291), .ZN(n7157) );
  OAI21_X1 U8132 ( .B1(n8646), .B2(n12281), .A(n7162), .ZN(n7161) );
  OAI21_X1 U8133 ( .B1(n12284), .B2(n12285), .A(n7159), .ZN(n7158) );
  INV_X1 U8134 ( .A(n12296), .ZN(n12101) );
  NAND2_X1 U8135 ( .A1(n7097), .A2(n8324), .ZN(n7342) );
  NOR2_X1 U8136 ( .A1(n10309), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n7097) );
  INV_X1 U8137 ( .A(n10633), .ZN(n6943) );
  INV_X1 U8138 ( .A(n11304), .ZN(n6934) );
  INV_X1 U8139 ( .A(n6800), .ZN(n6799) );
  OAI21_X1 U8140 ( .B1(n12687), .B2(n6801), .A(n12281), .ZN(n6800) );
  INV_X1 U8141 ( .A(n12277), .ZN(n6801) );
  NAND2_X1 U8142 ( .A1(n12834), .A2(n7178), .ZN(n12282) );
  OR2_X1 U8143 ( .A1(n8583), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8594) );
  INV_X1 U8144 ( .A(n7355), .ZN(n6809) );
  OR2_X1 U8145 ( .A1(n10911), .A2(n11108), .ZN(n11105) );
  INV_X1 U8146 ( .A(n6794), .ZN(n6793) );
  OAI21_X1 U8147 ( .B1(n12113), .B2(n6795), .A(n12199), .ZN(n6794) );
  INV_X1 U8148 ( .A(n12197), .ZN(n6795) );
  NAND2_X1 U8149 ( .A1(n10200), .A2(n12557), .ZN(n12166) );
  OR2_X1 U8150 ( .A1(n12652), .A2(n12419), .ZN(n12291) );
  OR2_X1 U8151 ( .A1(n9377), .A2(n12451), .ZN(n12297) );
  INV_X1 U8152 ( .A(SI_17_), .ZN(n8511) );
  INV_X1 U8153 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8240) );
  AND2_X1 U8154 ( .A1(n8230), .A2(n8231), .ZN(n7334) );
  NAND2_X1 U8155 ( .A1(n11391), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7194) );
  NAND2_X1 U8156 ( .A1(n8216), .A2(n8215), .ZN(n8217) );
  NAND2_X1 U8157 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n10557), .ZN(n8215) );
  NOR2_X1 U8158 ( .A1(n8540), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n8659) );
  INV_X1 U8159 ( .A(n8200), .ZN(n7186) );
  INV_X1 U8160 ( .A(n8284), .ZN(n6684) );
  AND2_X1 U8161 ( .A1(n7991), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n7969) );
  NOR2_X1 U8162 ( .A1(n7743), .A2(n7742), .ZN(n7772) );
  INV_X1 U8163 ( .A(n7135), .ZN(n7133) );
  AOI21_X1 U8164 ( .B1(n7135), .B2(n13131), .A(n12013), .ZN(n7132) );
  NOR2_X1 U8165 ( .A1(n13315), .A2(n12922), .ZN(n12013) );
  NAND2_X1 U8166 ( .A1(n6928), .A2(n13332), .ZN(n6927) );
  INV_X1 U8167 ( .A(n6929), .ZN(n6928) );
  OR2_X1 U8168 ( .A1(n13338), .A2(n13344), .ZN(n6929) );
  NAND2_X1 U8169 ( .A1(n12008), .A2(n13012), .ZN(n7147) );
  AND2_X1 U8170 ( .A1(n7840), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n7865) );
  NOR2_X1 U8171 ( .A1(n13258), .A2(n13359), .ZN(n13224) );
  NOR2_X1 U8172 ( .A1(n13254), .A2(n6669), .ZN(n6668) );
  INV_X1 U8173 ( .A(n6670), .ZN(n6669) );
  NAND2_X1 U8174 ( .A1(n7012), .A2(n7014), .ZN(n7010) );
  AND2_X1 U8175 ( .A1(n7648), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7670) );
  NAND2_X1 U8176 ( .A1(n6924), .A2(n6923), .ZN(n10525) );
  NAND2_X1 U8177 ( .A1(n10278), .A2(n10281), .ZN(n6975) );
  NAND2_X1 U8178 ( .A1(n8145), .A2(n7123), .ZN(n10286) );
  INV_X1 U8179 ( .A(n8146), .ZN(n7123) );
  AND2_X1 U8180 ( .A1(n7428), .A2(n7398), .ZN(n7211) );
  NOR2_X1 U8181 ( .A1(n9127), .A2(n11949), .ZN(n9128) );
  AND2_X1 U8182 ( .A1(n9295), .A2(n11878), .ZN(n9296) );
  AND2_X1 U8183 ( .A1(n7068), .A2(n9242), .ZN(n7067) );
  NOR2_X1 U8184 ( .A1(n13764), .A2(n13454), .ZN(n12058) );
  NOR2_X1 U8185 ( .A1(n13965), .A2(n9280), .ZN(n6887) );
  NAND2_X1 U8186 ( .A1(n11907), .A2(n11908), .ZN(n9281) );
  OR2_X1 U8187 ( .A1(n11907), .A2(n11908), .ZN(n11656) );
  INV_X1 U8188 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8950) );
  INV_X1 U8189 ( .A(n10109), .ZN(n10103) );
  NAND2_X1 U8190 ( .A1(n8859), .A2(n10080), .ZN(n9928) );
  NAND2_X1 U8191 ( .A1(n9338), .A2(n6470), .ZN(n8794) );
  INV_X1 U8192 ( .A(n7290), .ZN(n7289) );
  OAI21_X1 U8193 ( .B1(n8789), .B2(n6613), .A(P1_IR_REG_27__SCAN_IN), .ZN(
        n7290) );
  INV_X1 U8194 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8791) );
  INV_X1 U8195 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7025) );
  XNOR2_X1 U8196 ( .A(n9310), .B(P1_IR_REG_23__SCAN_IN), .ZN(n9743) );
  NAND2_X1 U8197 ( .A1(n8802), .A2(n8797), .ZN(n9084) );
  NAND2_X1 U8198 ( .A1(n7788), .A2(n9787), .ZN(n7804) );
  XNOR2_X1 U8199 ( .A(n7781), .B(SI_14_), .ZN(n7750) );
  AND2_X1 U8200 ( .A1(n7705), .A2(n7683), .ZN(n7703) );
  AOI21_X1 U8201 ( .B1(n7657), .B2(n6914), .A(n6538), .ZN(n6913) );
  AND2_X1 U8202 ( .A1(n14930), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n9383) );
  INV_X1 U8203 ( .A(n9420), .ZN(n6962) );
  AOI21_X1 U8204 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n14728), .A(n9398), .ZN(
        n9450) );
  NAND2_X1 U8205 ( .A1(n8432), .A2(n8431), .ZN(n8466) );
  NOR2_X1 U8206 ( .A1(n12457), .A2(n7326), .ZN(n7325) );
  INV_X1 U8207 ( .A(n12395), .ZN(n7326) );
  NAND2_X1 U8208 ( .A1(n11314), .A2(n11313), .ZN(n11376) );
  NOR2_X1 U8209 ( .A1(n7314), .A2(n11813), .ZN(n7312) );
  INV_X1 U8210 ( .A(n11815), .ZN(n7314) );
  AND2_X1 U8211 ( .A1(n8497), .A2(n11816), .ZN(n8515) );
  INV_X1 U8212 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n12477) );
  NOR2_X1 U8213 ( .A1(n8546), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8556) );
  AND2_X1 U8214 ( .A1(n8556), .A2(n14920), .ZN(n8569) );
  NAND2_X1 U8215 ( .A1(n8569), .A2(n12458), .ZN(n8571) );
  NAND2_X1 U8216 ( .A1(n12165), .A2(n12444), .ZN(n9980) );
  NAND2_X1 U8217 ( .A1(n8515), .A2(n12477), .ZN(n8531) );
  NOR2_X1 U8218 ( .A1(n8482), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8497) );
  AND4_X1 U8219 ( .A1(n8254), .A2(n8253), .A3(n8252), .A4(n8251), .ZN(n10926)
         );
  OR2_X1 U8220 ( .A1(n8345), .A2(n8329), .ZN(n8330) );
  NAND2_X1 U8221 ( .A1(n10312), .A2(n10313), .ZN(n10642) );
  NAND2_X1 U8222 ( .A1(n14658), .A2(n10650), .ZN(n14673) );
  NAND2_X1 U8223 ( .A1(n14700), .A2(n10653), .ZN(n14716) );
  NOR2_X1 U8224 ( .A1(n10588), .A2(n14688), .ZN(n14714) );
  INV_X1 U8225 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n10836) );
  NAND2_X1 U8226 ( .A1(n6940), .A2(n14732), .ZN(n14731) );
  OR2_X1 U8227 ( .A1(n14734), .A2(n14733), .ZN(n6940) );
  NAND2_X1 U8228 ( .A1(n14744), .A2(n10656), .ZN(n10660) );
  NAND2_X1 U8229 ( .A1(n11298), .A2(n11200), .ZN(n11201) );
  NAND2_X1 U8230 ( .A1(n11631), .A2(n11632), .ZN(n11633) );
  NAND2_X1 U8231 ( .A1(n11633), .A2(n11637), .ZN(n12562) );
  NOR2_X1 U8232 ( .A1(n11480), .A2(n6949), .ZN(n11643) );
  NAND2_X1 U8233 ( .A1(n6951), .A2(n6950), .ZN(n6949) );
  INV_X1 U8234 ( .A(n11479), .ZN(n6950) );
  INV_X1 U8235 ( .A(n11478), .ZN(n6951) );
  NAND2_X1 U8236 ( .A1(n12562), .A2(n12566), .ZN(n12592) );
  INV_X1 U8237 ( .A(n12571), .ZN(n12584) );
  NAND2_X1 U8238 ( .A1(n7106), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7105) );
  NAND2_X1 U8239 ( .A1(n12607), .A2(n7106), .ZN(n7103) );
  OR2_X1 U8240 ( .A1(n12559), .A2(n12560), .ZN(n7108) );
  AND2_X1 U8241 ( .A1(n6945), .A2(n6944), .ZN(n12632) );
  OR2_X1 U8242 ( .A1(n6946), .A2(n14041), .ZN(n6944) );
  OR2_X1 U8243 ( .A1(n12640), .A2(n12639), .ZN(n14088) );
  AND2_X1 U8244 ( .A1(n12291), .A2(n12289), .ZN(n12445) );
  OAI22_X1 U8245 ( .A1(n12683), .A2(n6819), .B1(n8632), .B2(n6820), .ZN(n12656) );
  NAND2_X1 U8246 ( .A1(n7364), .A2(n6823), .ZN(n6819) );
  INV_X1 U8247 ( .A(n6821), .ZN(n6820) );
  INV_X1 U8248 ( .A(n12141), .ZN(n8646) );
  NAND2_X1 U8249 ( .A1(n12683), .A2(n12682), .ZN(n12681) );
  NAND2_X1 U8250 ( .A1(n6842), .A2(n6513), .ZN(n12696) );
  NAND2_X1 U8251 ( .A1(n6843), .A2(n6844), .ZN(n6841) );
  NAND2_X1 U8252 ( .A1(n12845), .A2(n12500), .ZN(n6848) );
  NAND2_X1 U8253 ( .A1(n12717), .A2(n8578), .ZN(n6847) );
  AND2_X1 U8254 ( .A1(n6847), .A2(n6845), .ZN(n12708) );
  AND2_X1 U8255 ( .A1(n12106), .A2(n12143), .ZN(n12721) );
  AOI21_X1 U8256 ( .B1(n6838), .B2(n6840), .A(n6525), .ZN(n6837) );
  AOI21_X1 U8257 ( .B1(n6788), .B2(n6790), .A(n6786), .ZN(n6785) );
  INV_X1 U8258 ( .A(n6789), .ZN(n6788) );
  NAND2_X1 U8259 ( .A1(n11600), .A2(n11599), .ZN(n11598) );
  NAND2_X1 U8260 ( .A1(n6826), .A2(n6824), .ZN(n11490) );
  AOI21_X1 U8261 ( .B1(n6827), .B2(n6830), .A(n6825), .ZN(n6824) );
  AOI21_X1 U8262 ( .B1(n6829), .B2(n6828), .A(n11488), .ZN(n6827) );
  OR2_X1 U8263 ( .A1(n8695), .A2(n8694), .ZN(n11493) );
  NOR2_X1 U8264 ( .A1(n8415), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8432) );
  AND2_X1 U8265 ( .A1(n12220), .A2(n12227), .ZN(n12226) );
  INV_X1 U8266 ( .A(n14815), .ZN(n12208) );
  NAND2_X1 U8267 ( .A1(n10923), .A2(n12113), .ZN(n10925) );
  OR2_X1 U8268 ( .A1(n8264), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8278) );
  AND2_X1 U8269 ( .A1(n12190), .A2(n12189), .ZN(n12186) );
  AND2_X1 U8270 ( .A1(n10726), .A2(n8391), .ZN(n10717) );
  NAND2_X1 U8271 ( .A1(n10727), .A2(n12121), .ZN(n10726) );
  AND3_X1 U8272 ( .A1(n8374), .A2(n8373), .A3(n8372), .ZN(n10057) );
  NAND2_X1 U8273 ( .A1(n6817), .A2(n8360), .ZN(n10445) );
  NOR2_X1 U8274 ( .A1(n12118), .A2(n6818), .ZN(n6817) );
  INV_X1 U8275 ( .A(n8359), .ZN(n6818) );
  NAND2_X1 U8276 ( .A1(n12165), .A2(n12166), .ZN(n9987) );
  INV_X1 U8277 ( .A(n14760), .ZN(n12765) );
  INV_X1 U8278 ( .A(n14088), .ZN(n14092) );
  OR2_X1 U8279 ( .A1(n9356), .A2(n12419), .ZN(n7366) );
  OAI21_X1 U8280 ( .B1(n12649), .B2(n14828), .A(n12654), .ZN(n8764) );
  NAND2_X1 U8281 ( .A1(n14879), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6691) );
  AOI21_X1 U8282 ( .B1(n8648), .B2(n8649), .A(n6672), .ZN(n9358) );
  AND2_X1 U8283 ( .A1(n11842), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6672) );
  XNOR2_X1 U8284 ( .A(n8724), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8740) );
  OR2_X1 U8285 ( .A1(n8718), .A2(n8723), .ZN(n8724) );
  NAND2_X1 U8286 ( .A1(n8606), .A2(n8605), .ZN(n8620) );
  XNOR2_X1 U8287 ( .A(n8715), .B(n8714), .ZN(n10305) );
  INV_X1 U8288 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8714) );
  OAI21_X1 U8289 ( .B1(n8713), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8715) );
  INV_X1 U8290 ( .A(n8509), .ZN(n8540) );
  NAND2_X1 U8291 ( .A1(n8211), .A2(n8210), .ZN(n8506) );
  NAND2_X1 U8292 ( .A1(n8491), .A2(n8489), .ZN(n8211) );
  NAND3_X1 U8293 ( .A1(n7173), .A2(n8208), .A3(n7171), .ZN(n8476) );
  NAND2_X1 U8294 ( .A1(n7172), .A2(n8457), .ZN(n7171) );
  NAND2_X1 U8295 ( .A1(n7181), .A2(n7180), .ZN(n8443) );
  AOI21_X1 U8296 ( .B1(n7183), .B2(n7185), .A(n6587), .ZN(n7180) );
  INV_X1 U8297 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8424) );
  OR2_X1 U8298 ( .A1(n8274), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8300) );
  INV_X2 U8299 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8272) );
  XNOR2_X1 U8300 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8382) );
  XNOR2_X1 U8301 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8366) );
  AND2_X1 U8302 ( .A1(n8188), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8338) );
  INV_X1 U8303 ( .A(n12944), .ZN(n6712) );
  INV_X1 U8304 ( .A(n12943), .ZN(n6711) );
  INV_X1 U8305 ( .A(n12945), .ZN(n6704) );
  INV_X1 U8306 ( .A(n6709), .ZN(n6708) );
  AOI21_X1 U8307 ( .B1(n12917), .B2(n10025), .A(n7349), .ZN(n10028) );
  INV_X1 U8308 ( .A(n11283), .ZN(n7202) );
  INV_X1 U8309 ( .A(n11172), .ZN(n7204) );
  NOR2_X1 U8310 ( .A1(n12994), .A2(n7208), .ZN(n7207) );
  INV_X1 U8311 ( .A(n12934), .ZN(n7208) );
  AND2_X1 U8312 ( .A1(n11182), .A2(n11171), .ZN(n11172) );
  NAND2_X1 U8313 ( .A1(n11157), .A2(n11156), .ZN(n11173) );
  INV_X1 U8314 ( .A(n11158), .ZN(n11157) );
  AND2_X1 U8315 ( .A1(n9866), .A2(n11143), .ZN(n10017) );
  INV_X1 U8316 ( .A(n12995), .ZN(n13038) );
  AND2_X1 U8317 ( .A1(n13033), .A2(n6506), .ZN(n6709) );
  NAND2_X1 U8318 ( .A1(n10995), .A2(n13093), .ZN(n10013) );
  INV_X1 U8319 ( .A(n8096), .ZN(n8076) );
  AND2_X1 U8320 ( .A1(n14401), .A2(n6590), .ZN(n14403) );
  NOR2_X1 U8321 ( .A1(n6770), .A2(n14403), .ZN(n14417) );
  NOR2_X1 U8322 ( .A1(n9647), .A2(n6771), .ZN(n6770) );
  AND2_X1 U8323 ( .A1(n6773), .A2(n6772), .ZN(n9793) );
  NAND2_X1 U8324 ( .A1(n9656), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6772) );
  OR2_X1 U8325 ( .A1(n9643), .A2(n9642), .ZN(n9682) );
  NAND2_X1 U8326 ( .A1(n6764), .A2(n6760), .ZN(n6759) );
  INV_X1 U8327 ( .A(n9681), .ZN(n6760) );
  INV_X1 U8328 ( .A(n6755), .ZN(n6754) );
  AOI21_X1 U8329 ( .B1(n6756), .B2(n6761), .A(n14443), .ZN(n6755) );
  OR2_X1 U8330 ( .A1(n9643), .A2(n6761), .ZN(n6758) );
  NOR2_X1 U8331 ( .A1(n8174), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n7685) );
  NAND2_X1 U8332 ( .A1(n10427), .A2(n6775), .ZN(n14489) );
  NOR2_X1 U8333 ( .A1(n6777), .A2(n6776), .ZN(n6775) );
  NOR2_X1 U8334 ( .A1(n10441), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6776) );
  INV_X1 U8335 ( .A(n10426), .ZN(n6777) );
  AOI21_X1 U8336 ( .B1(n14489), .B2(n14487), .A(n14488), .ZN(n14486) );
  NAND2_X1 U8337 ( .A1(n14501), .A2(n14500), .ZN(n14499) );
  XNOR2_X1 U8338 ( .A(n11730), .B(n11742), .ZN(n11457) );
  XNOR2_X1 U8339 ( .A(n13078), .B(n13087), .ZN(n14535) );
  NAND2_X1 U8340 ( .A1(n14525), .A2(n13077), .ZN(n13078) );
  NOR2_X1 U8341 ( .A1(n14535), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n14534) );
  AND2_X1 U8342 ( .A1(n8087), .A2(n8086), .ZN(n12023) );
  AOI21_X1 U8343 ( .B1(n6985), .B2(n6983), .A(n6526), .ZN(n6982) );
  INV_X1 U8344 ( .A(n12036), .ZN(n6983) );
  INV_X1 U8345 ( .A(n6985), .ZN(n6984) );
  NAND2_X1 U8346 ( .A1(n7136), .A2(n7137), .ZN(n6643) );
  AOI21_X1 U8347 ( .B1(n7136), .B2(n7135), .A(n13268), .ZN(n6641) );
  NAND2_X1 U8348 ( .A1(n6655), .A2(n6654), .ZN(n13140) );
  NAND2_X1 U8349 ( .A1(n13189), .A2(n6657), .ZN(n6655) );
  AOI21_X1 U8350 ( .B1(n6657), .B2(n6659), .A(n6530), .ZN(n6654) );
  NOR2_X1 U8351 ( .A1(n13207), .A2(n6927), .ZN(n13164) );
  OR2_X1 U8352 ( .A1(n6994), .A2(n6497), .ZN(n6990) );
  INV_X1 U8353 ( .A(n6993), .ZN(n6992) );
  NOR2_X1 U8354 ( .A1(n13207), .A2(n6929), .ZN(n13179) );
  NOR2_X1 U8355 ( .A1(n13207), .A2(n13344), .ZN(n13194) );
  NAND2_X1 U8356 ( .A1(n13222), .A2(n6999), .ZN(n7001) );
  OR2_X1 U8357 ( .A1(n7888), .A2(n12960), .ZN(n7906) );
  NAND2_X1 U8358 ( .A1(n7865), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7888) );
  NAND2_X1 U8359 ( .A1(n6930), .A2(n13262), .ZN(n13258) );
  AND2_X1 U8360 ( .A1(n6647), .A2(n6589), .ZN(n11724) );
  OAI21_X1 U8361 ( .B1(n11214), .B2(n6646), .A(n6644), .ZN(n6647) );
  INV_X1 U8362 ( .A(n6645), .ZN(n6644) );
  INV_X1 U8363 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11525) );
  OR2_X1 U8364 ( .A1(n7697), .A2(n11525), .ZN(n7719) );
  NAND2_X1 U8365 ( .A1(n11067), .A2(n11066), .ZN(n11070) );
  AND2_X1 U8366 ( .A1(n7152), .A2(n6650), .ZN(n6649) );
  NAND2_X1 U8367 ( .A1(n10850), .A2(n6651), .ZN(n6648) );
  AND2_X1 U8368 ( .A1(n11068), .A2(n11066), .ZN(n7152) );
  AND2_X1 U8369 ( .A1(n10522), .A2(n10520), .ZN(n7149) );
  NAND2_X1 U8370 ( .A1(n10669), .A2(n10518), .ZN(n10943) );
  AND2_X1 U8371 ( .A1(n8140), .A2(n10515), .ZN(n10504) );
  NAND2_X1 U8372 ( .A1(n13071), .A2(n8141), .ZN(n8142) );
  NAND2_X1 U8373 ( .A1(n10282), .A2(n10772), .ZN(n10565) );
  NAND2_X1 U8374 ( .A1(n10287), .A2(n10286), .ZN(n10778) );
  NAND2_X1 U8375 ( .A1(n9869), .A2(n10025), .ZN(n8144) );
  INV_X1 U8376 ( .A(n9876), .ZN(n10023) );
  OR2_X1 U8377 ( .A1(n14555), .A2(n10006), .ZN(n10191) );
  AND2_X1 U8378 ( .A1(n6987), .A2(n6989), .ZN(n13132) );
  NAND2_X1 U8379 ( .A1(n6987), .A2(n6985), .ZN(n13319) );
  AND2_X1 U8380 ( .A1(n9633), .A2(n9634), .ZN(n10258) );
  CLKBUF_X1 U8381 ( .A(n8180), .Z(n8181) );
  INV_X1 U8382 ( .A(n7956), .ZN(n7954) );
  OR2_X1 U8383 ( .A1(n7523), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n7526) );
  INV_X1 U8384 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7369) );
  NAND2_X1 U8385 ( .A1(n9144), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9172) );
  INV_X1 U8386 ( .A(n9184), .ZN(n9171) );
  INV_X1 U8387 ( .A(n9156), .ZN(n9144) );
  AND2_X1 U8388 ( .A1(n9070), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9091) );
  INV_X1 U8389 ( .A(n13500), .ZN(n7031) );
  AOI21_X1 U8390 ( .B1(n7034), .B2(n7036), .A(n6520), .ZN(n7033) );
  AOI21_X1 U8391 ( .B1(n10179), .B2(n10098), .A(n9749), .ZN(n9750) );
  OAI211_X1 U8392 ( .C1(n9754), .C2(n9753), .A(n9752), .B(n9751), .ZN(n9836)
         );
  INV_X1 U8393 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n11949) );
  NAND2_X1 U8394 ( .A1(n13526), .A2(n13527), .ZN(n13525) );
  INV_X1 U8395 ( .A(n9172), .ZN(n9155) );
  NAND2_X1 U8396 ( .A1(n10178), .A2(n10177), .ZN(n13537) );
  INV_X1 U8397 ( .A(n10183), .ZN(n6631) );
  AND2_X1 U8398 ( .A1(n9091), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9097) );
  OR3_X1 U8399 ( .A1(n9041), .A2(n9035), .A3(n9034), .ZN(n9056) );
  INV_X1 U8400 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n14977) );
  INV_X1 U8401 ( .A(n6463), .ZN(n9130) );
  NAND2_X1 U8402 ( .A1(n8889), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n7281) );
  OR2_X1 U8403 ( .A1(n9806), .A2(n9805), .ZN(n9807) );
  OR2_X1 U8404 ( .A1(n9015), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9016) );
  NAND2_X1 U8405 ( .A1(n11589), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6624) );
  INV_X1 U8406 ( .A(n13763), .ZN(n6743) );
  AND2_X1 U8407 ( .A1(n6750), .A2(n6561), .ZN(n6748) );
  NAND2_X1 U8408 ( .A1(n6749), .A2(n6750), .ZN(n12052) );
  AND2_X1 U8409 ( .A1(n9229), .A2(n9218), .ZN(n13768) );
  INV_X1 U8410 ( .A(n9199), .ZN(n9183) );
  NAND2_X1 U8411 ( .A1(n11857), .A2(n11856), .ZN(n13792) );
  NAND2_X1 U8412 ( .A1(n6869), .A2(n6726), .ZN(n13798) );
  AOI21_X1 U8413 ( .B1(n6871), .B2(n6872), .A(n6547), .ZN(n6726) );
  NAND2_X1 U8414 ( .A1(n13812), .A2(n11877), .ZN(n13796) );
  NAND2_X1 U8415 ( .A1(n13873), .A2(n6476), .ZN(n13816) );
  AOI21_X1 U8416 ( .B1(n7300), .B2(n13859), .A(n6523), .ZN(n7299) );
  NAND2_X1 U8417 ( .A1(n13873), .A2(n6885), .ZN(n13831) );
  NAND2_X1 U8418 ( .A1(n13873), .A2(n13971), .ZN(n13860) );
  NAND2_X1 U8419 ( .A1(n9111), .A2(n9110), .ZN(n13874) );
  OR2_X1 U8420 ( .A1(n14158), .A2(n14180), .ZN(n13902) );
  AND2_X1 U8421 ( .A1(n9121), .A2(n9120), .ZN(n13893) );
  NAND2_X1 U8422 ( .A1(n7274), .A2(n11656), .ZN(n11865) );
  NAND2_X1 U8423 ( .A1(n11655), .A2(n11654), .ZN(n7274) );
  NAND2_X1 U8424 ( .A1(n6892), .A2(n6891), .ZN(n11660) );
  AOI21_X1 U8425 ( .B1(n6472), .B2(n7295), .A(n6521), .ZN(n7291) );
  NAND2_X1 U8426 ( .A1(n14170), .A2(n14171), .ZN(n7293) );
  NOR2_X1 U8427 ( .A1(n14174), .A2(n11787), .ZN(n11327) );
  AND2_X1 U8428 ( .A1(n8996), .A2(n8778), .ZN(n9009) );
  NAND2_X1 U8429 ( .A1(n14282), .A2(n11232), .ZN(n14164) );
  OR2_X1 U8430 ( .A1(n14290), .A2(n14287), .ZN(n14173) );
  OR2_X1 U8431 ( .A1(n14172), .A2(n14173), .ZN(n14174) );
  OR2_X1 U8432 ( .A1(n9911), .A2(n9760), .ZN(n13892) );
  NOR2_X1 U8433 ( .A1(n10765), .A2(n6866), .ZN(n6859) );
  INV_X1 U8434 ( .A(n6867), .ZN(n6866) );
  INV_X1 U8435 ( .A(n6864), .ZN(n6862) );
  OAI21_X1 U8436 ( .B1(n10765), .B2(n6865), .A(n10764), .ZN(n6864) );
  NAND2_X1 U8437 ( .A1(n10351), .A2(n6867), .ZN(n6865) );
  NOR2_X1 U8438 ( .A1(n10759), .A2(n11258), .ZN(n10800) );
  NAND2_X1 U8439 ( .A1(n6882), .A2(n6881), .ZN(n10759) );
  INV_X1 U8440 ( .A(n10358), .ZN(n6882) );
  INV_X1 U8441 ( .A(n7283), .ZN(n7282) );
  NAND2_X1 U8442 ( .A1(n10149), .A2(n10148), .ZN(n7284) );
  AND2_X1 U8443 ( .A1(n6482), .A2(n14309), .ZN(n10229) );
  NAND2_X1 U8444 ( .A1(n14309), .A2(n10121), .ZN(n10228) );
  NAND2_X1 U8445 ( .A1(n10108), .A2(n10107), .ZN(n10160) );
  AND2_X1 U8446 ( .A1(n14312), .A2(n14328), .ZN(n14309) );
  INV_X1 U8447 ( .A(n14182), .ZN(n14310) );
  INV_X1 U8448 ( .A(n14371), .ZN(n14345) );
  NAND2_X1 U8449 ( .A1(n9345), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9546) );
  INV_X1 U8450 ( .A(n9743), .ZN(n9345) );
  NAND2_X1 U8451 ( .A1(n8103), .A2(n8067), .ZN(n8070) );
  INV_X1 U8452 ( .A(n8794), .ZN(n7023) );
  NOR2_X1 U8453 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7022) );
  NAND2_X1 U8454 ( .A1(n9338), .A2(n8771), .ZN(n8793) );
  INV_X1 U8455 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8789) );
  INV_X1 U8456 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8788) );
  NAND2_X1 U8457 ( .A1(n8805), .A2(n8804), .ZN(n9334) );
  INV_X1 U8458 ( .A(n8810), .ZN(n8805) );
  NAND2_X1 U8459 ( .A1(n6731), .A2(n7900), .ZN(n7915) );
  NAND2_X1 U8460 ( .A1(n7898), .A2(n7897), .ZN(n6731) );
  INV_X1 U8461 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9101) );
  CLKBUF_X1 U8462 ( .A(n9049), .Z(n9050) );
  XNOR2_X1 U8463 ( .A(n7750), .B(n7782), .ZN(n10050) );
  NAND2_X1 U8464 ( .A1(n6915), .A2(n7635), .ZN(n7658) );
  NAND2_X1 U8465 ( .A1(n7633), .A2(n7632), .ZN(n6915) );
  OR2_X1 U8466 ( .A1(n9051), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n8980) );
  OR2_X1 U8467 ( .A1(n8945), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9051) );
  NAND2_X1 U8468 ( .A1(n7223), .A2(n7589), .ZN(n6720) );
  CLKBUF_X1 U8469 ( .A(n7519), .Z(n7496) );
  NOR2_X1 U8470 ( .A1(n14613), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n9424) );
  XNOR2_X1 U8471 ( .A(n9385), .B(n9384), .ZN(n9430) );
  NOR2_X1 U8472 ( .A1(n9436), .A2(n9437), .ZN(n9438) );
  NOR2_X1 U8473 ( .A1(n9393), .A2(n9392), .ZN(n9440) );
  NAND2_X1 U8474 ( .A1(n9447), .A2(n9446), .ZN(n9448) );
  INV_X1 U8475 ( .A(n9455), .ZN(n6956) );
  INV_X1 U8476 ( .A(n14046), .ZN(n6960) );
  OAI21_X1 U8477 ( .B1(n9402), .B2(n10662), .A(n9401), .ZN(n9412) );
  OAI21_X1 U8478 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n9406), .A(n9405), .ZN(
        n9410) );
  NOR2_X1 U8479 ( .A1(n9470), .A2(n14260), .ZN(n9475) );
  NOR2_X1 U8480 ( .A1(n9484), .A2(n9483), .ZN(n9488) );
  AND2_X1 U8481 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n9482), .ZN(n9483) );
  NAND2_X1 U8482 ( .A1(n7317), .A2(n7315), .ZN(n11559) );
  OAI21_X1 U8483 ( .B1(n6478), .B2(n11560), .A(n7316), .ZN(n7315) );
  AND3_X1 U8484 ( .A1(n8413), .A2(n8412), .A3(n8411), .ZN(n10967) );
  AND4_X1 U8485 ( .A1(n8311), .A2(n8310), .A3(n8309), .A4(n8308), .ZN(n11057)
         );
  NAND2_X1 U8486 ( .A1(n12494), .A2(n12395), .ZN(n12456) );
  NAND2_X1 U8487 ( .A1(n8568), .A2(n8567), .ZN(n12460) );
  INV_X1 U8488 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n11816) );
  INV_X1 U8489 ( .A(n11813), .ZN(n7311) );
  NAND2_X1 U8490 ( .A1(n7313), .A2(n7312), .ZN(n12384) );
  INV_X1 U8491 ( .A(n12544), .ZN(n12476) );
  CLKBUF_X1 U8492 ( .A(n12484), .Z(n12485) );
  NAND2_X1 U8493 ( .A1(n8593), .A2(n8592), .ZN(n12491) );
  NAND2_X1 U8494 ( .A1(n10396), .A2(n10395), .ZN(n10402) );
  NAND2_X1 U8495 ( .A1(n10831), .A2(n7332), .ZN(n10834) );
  OAI21_X1 U8496 ( .B1(n10307), .B2(n10321), .A(n7098), .ZN(n12157) );
  NAND2_X1 U8497 ( .A1(n10307), .A2(n9498), .ZN(n7098) );
  NAND2_X1 U8498 ( .A1(n12496), .A2(n12495), .ZN(n12494) );
  AND4_X1 U8499 ( .A1(n8406), .A2(n8405), .A3(n8404), .A4(n8403), .ZN(n11317)
         );
  AND4_X1 U8500 ( .A1(n8552), .A2(n8551), .A3(n8550), .A4(n8549), .ZN(n12514)
         );
  OR2_X1 U8501 ( .A1(n12387), .A2(n12386), .ZN(n12388) );
  CLKBUF_X1 U8502 ( .A(n12519), .Z(n12520) );
  NAND2_X1 U8503 ( .A1(n8623), .A2(n8622), .ZN(n12529) );
  OR2_X1 U8504 ( .A1(n12096), .A2(n11691), .ZN(n8622) );
  NAND2_X1 U8505 ( .A1(n9995), .A2(n9994), .ZN(n12531) );
  INV_X1 U8506 ( .A(n7313), .ZN(n11814) );
  INV_X1 U8507 ( .A(n12450), .ZN(n12523) );
  NAND2_X1 U8508 ( .A1(n8645), .A2(n8644), .ZN(n12536) );
  INV_X1 U8509 ( .A(n12514), .ZN(n12766) );
  INV_X1 U8510 ( .A(n12478), .ZN(n12543) );
  INV_X1 U8511 ( .A(n12386), .ZN(n12764) );
  INV_X1 U8512 ( .A(n11503), .ZN(n12547) );
  INV_X1 U8513 ( .A(n11317), .ZN(n12549) );
  INV_X1 U8514 ( .A(n12207), .ZN(n12551) );
  NAND2_X1 U8515 ( .A1(n12082), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8280) );
  INV_X1 U8516 ( .A(P3_U3897), .ZN(n12552) );
  AND2_X1 U8517 ( .A1(P3_U3151), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7099) );
  INV_X1 U8518 ( .A(n7100), .ZN(n10325) );
  INV_X1 U8519 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n9384) );
  NOR2_X1 U8520 ( .A1(n8388), .A2(n8387), .ZN(n14647) );
  INV_X1 U8521 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14687) );
  NOR2_X1 U8522 ( .A1(n14651), .A2(n10585), .ZN(n14670) );
  XNOR2_X1 U8523 ( .A(n10587), .B(n10613), .ZN(n14689) );
  OAI21_X1 U8524 ( .B1(n14730), .B2(n7110), .A(n7109), .ZN(n11184) );
  NAND2_X1 U8525 ( .A1(n7111), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7110) );
  NAND2_X1 U8526 ( .A1(n10591), .A2(n7111), .ZN(n7109) );
  NOR2_X1 U8527 ( .A1(n11297), .A2(n8417), .ZN(n11296) );
  AND2_X1 U8528 ( .A1(n6937), .A2(n6935), .ZN(n11305) );
  OAI21_X1 U8529 ( .B1(n11297), .B2(n7118), .A(n7117), .ZN(n11467) );
  NAND2_X1 U8530 ( .A1(n7119), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7118) );
  NAND2_X1 U8531 ( .A1(n11187), .A2(n7119), .ZN(n7117) );
  INV_X1 U8532 ( .A(n11189), .ZN(n7119) );
  INV_X1 U8533 ( .A(n7115), .ZN(n11627) );
  OAI21_X1 U8534 ( .B1(n11468), .B2(n7113), .A(n7112), .ZN(n12558) );
  NAND2_X1 U8535 ( .A1(n7116), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7113) );
  INV_X1 U8536 ( .A(n11639), .ZN(n7116) );
  INV_X1 U8537 ( .A(n11628), .ZN(n7114) );
  XNOR2_X1 U8538 ( .A(n12592), .B(n12605), .ZN(n12563) );
  NOR2_X1 U8539 ( .A1(n7330), .A2(n7329), .ZN(n8492) );
  INV_X1 U8540 ( .A(n8226), .ZN(n7329) );
  AND2_X1 U8541 ( .A1(n10319), .A2(n10318), .ZN(n14080) );
  XNOR2_X1 U8542 ( .A(n6946), .B(n14041), .ZN(n12588) );
  INV_X1 U8543 ( .A(n6945), .ZN(n12627) );
  AND2_X1 U8544 ( .A1(n12081), .A2(n12080), .ZN(n14091) );
  NAND2_X1 U8545 ( .A1(n8638), .A2(n8637), .ZN(n12781) );
  OR2_X1 U8546 ( .A1(n12096), .A2(n12071), .ZN(n8637) );
  NAND2_X1 U8547 ( .A1(n12686), .A2(n12277), .ZN(n12668) );
  NAND2_X1 U8548 ( .A1(n6811), .A2(n12275), .ZN(n12700) );
  NAND2_X1 U8549 ( .A1(n12775), .A2(n12150), .ZN(n12753) );
  NAND2_X1 U8550 ( .A1(n8530), .A2(n8529), .ZN(n12774) );
  NAND2_X1 U8551 ( .A1(n11602), .A2(n12244), .ZN(n6787) );
  NAND2_X1 U8552 ( .A1(n6832), .A2(n6833), .ZN(n11502) );
  NAND2_X1 U8553 ( .A1(n11289), .A2(n8430), .ZN(n6835) );
  AND2_X1 U8554 ( .A1(n14770), .A2(n10713), .ZN(n12778) );
  NAND2_X1 U8555 ( .A1(n6804), .A2(n12214), .ZN(n11030) );
  AND3_X1 U8556 ( .A1(n8263), .A2(n8262), .A3(n8261), .ZN(n10722) );
  INV_X1 U8557 ( .A(n12757), .ZN(n12773) );
  INV_X1 U8558 ( .A(n12778), .ZN(n12663) );
  OR2_X1 U8559 ( .A1(n12308), .A2(n10132), .ZN(n14755) );
  INV_X1 U8560 ( .A(n14755), .ZN(n12755) );
  NAND2_X1 U8561 ( .A1(n10136), .A2(n14755), .ZN(n14770) );
  OR2_X1 U8562 ( .A1(n10136), .A2(n10131), .ZN(n12757) );
  AND2_X2 U8563 ( .A1(n10130), .A2(n8751), .ZN(n14846) );
  NAND2_X1 U8564 ( .A1(n8764), .A2(n14833), .ZN(n6814) );
  OR2_X1 U8565 ( .A1(n14833), .A2(n6813), .ZN(n6812) );
  INV_X1 U8566 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n6813) );
  INV_X1 U8567 ( .A(n12529), .ZN(n12831) );
  INV_X1 U8568 ( .A(n12460), .ZN(n12849) );
  AND2_X1 U8569 ( .A1(n8555), .A2(n8554), .ZN(n12853) );
  NAND2_X1 U8570 ( .A1(n8545), .A2(n8544), .ZN(n12857) );
  INV_X1 U8571 ( .A(n12385), .ZN(n12866) );
  INV_X1 U8572 ( .A(n12246), .ZN(n11759) );
  INV_X1 U8573 ( .A(n12157), .ZN(n10274) );
  NAND2_X1 U8574 ( .A1(n14833), .A2(n14812), .ZN(n12865) );
  NAND2_X1 U8575 ( .A1(n9567), .A2(n9562), .ZN(n14965) );
  XNOR2_X1 U8576 ( .A(n6690), .B(n12095), .ZN(n12867) );
  OAI21_X1 U8577 ( .B1(n12092), .B2(n12091), .A(n6691), .ZN(n6690) );
  INV_X1 U8578 ( .A(n8245), .ZN(n12877) );
  INV_X1 U8579 ( .A(n8740), .ZN(n11693) );
  NAND2_X1 U8580 ( .A1(n8719), .A2(n6632), .ZN(n11610) );
  AOI21_X1 U8581 ( .B1(n8717), .B2(P3_IR_REG_25__SCAN_IN), .A(n6546), .ZN(
        n6632) );
  XNOR2_X1 U8582 ( .A(n8722), .B(n8721), .ZN(n11463) );
  INV_X1 U8583 ( .A(SI_23_), .ZN(n11103) );
  NAND2_X1 U8584 ( .A1(n6689), .A2(n7191), .ZN(n8590) );
  NAND2_X1 U8585 ( .A1(n8566), .A2(n6594), .ZN(n6689) );
  NAND2_X1 U8586 ( .A1(n7193), .A2(n7195), .ZN(n8580) );
  NAND2_X1 U8587 ( .A1(n8566), .A2(n8564), .ZN(n7193) );
  XNOR2_X1 U8588 ( .A(n8661), .B(n8660), .ZN(n12161) );
  INV_X1 U8589 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8660) );
  INV_X1 U8590 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8662) );
  INV_X1 U8591 ( .A(SI_19_), .ZN(n10044) );
  INV_X1 U8592 ( .A(n14071), .ZN(n14025) );
  INV_X1 U8593 ( .A(SI_16_), .ZN(n9787) );
  INV_X1 U8594 ( .A(SI_15_), .ZN(n9631) );
  NAND2_X1 U8595 ( .A1(n7175), .A2(n8207), .ZN(n8458) );
  NAND2_X1 U8596 ( .A1(n8446), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7175) );
  INV_X1 U8597 ( .A(SI_12_), .ZN(n14938) );
  INV_X1 U8598 ( .A(n11476), .ZN(n11469) );
  INV_X1 U8599 ( .A(SI_11_), .ZN(n9538) );
  NAND2_X1 U8600 ( .A1(n7182), .A2(n8205), .ZN(n8423) );
  NAND2_X1 U8601 ( .A1(n8408), .A2(n8407), .ZN(n7182) );
  NAND2_X1 U8602 ( .A1(n7187), .A2(n8202), .ZN(n8313) );
  NAND2_X1 U8603 ( .A1(n8299), .A2(n8297), .ZN(n7187) );
  INV_X1 U8604 ( .A(n14719), .ZN(n10636) );
  NAND2_X1 U8605 ( .A1(n7163), .A2(n7166), .ZN(n8285) );
  NAND2_X1 U8606 ( .A1(n7170), .A2(n8197), .ZN(n8271) );
  NAND2_X1 U8607 ( .A1(n8256), .A2(n8255), .ZN(n7170) );
  NAND2_X1 U8608 ( .A1(n8324), .A2(n7096), .ZN(n8370) );
  NOR2_X1 U8609 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7096) );
  NAND2_X1 U8610 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8325) );
  AND2_X1 U8611 ( .A1(n11994), .A2(n11694), .ZN(n7196) );
  INV_X1 U8612 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n14937) );
  NAND2_X1 U8613 ( .A1(n11964), .A2(n10245), .ZN(n10346) );
  OR2_X1 U8614 ( .A1(n7434), .A2(n9647), .ZN(n7420) );
  OR2_X1 U8615 ( .A1(n8104), .A2(n9506), .ZN(n7422) );
  NAND2_X1 U8616 ( .A1(n11967), .A2(n11966), .ZN(n12974) );
  INV_X1 U8617 ( .A(n12975), .ZN(n7206) );
  INV_X1 U8618 ( .A(n12984), .ZN(n6718) );
  INV_X1 U8619 ( .A(n7347), .ZN(n6715) );
  NAND2_X1 U8620 ( .A1(n6721), .A2(n6723), .ZN(n6722) );
  INV_X1 U8621 ( .A(n6721), .ZN(n10745) );
  NAND2_X1 U8622 ( .A1(n10212), .A2(n8143), .ZN(n10215) );
  NAND2_X1 U8623 ( .A1(n7209), .A2(n12934), .ZN(n12993) );
  NAND2_X1 U8624 ( .A1(n12885), .A2(n12884), .ZN(n13025) );
  OAI211_X1 U8625 ( .C1(n11999), .C2(n6498), .A(n6701), .B(n6699), .ZN(n11701)
         );
  OR2_X1 U8626 ( .A1(n6498), .A2(n11699), .ZN(n6701) );
  NAND2_X1 U8627 ( .A1(n11999), .A2(n6700), .ZN(n6699) );
  AND2_X1 U8628 ( .A1(n6498), .A2(n11699), .ZN(n6700) );
  INV_X1 U8629 ( .A(n11989), .ZN(n13013) );
  AOI211_X1 U8630 ( .C1(n8164), .C2(n10195), .A(n11143), .B(n8163), .ZN(n8167)
         );
  NAND4_X1 U8631 ( .A1(n7541), .A2(n7540), .A3(n7539), .A4(n7538), .ZN(n13069)
         );
  NAND4_X1 U8632 ( .A1(n7516), .A2(n7515), .A3(n7514), .A4(n7513), .ZN(n13070)
         );
  OR2_X1 U8633 ( .A1(n7508), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7473) );
  NAND2_X1 U8634 ( .A1(n7485), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7389) );
  INV_X1 U8635 ( .A(n6773), .ZN(n14427) );
  NAND2_X1 U8636 ( .A1(n6758), .A2(n6759), .ZN(n9941) );
  INV_X1 U8637 ( .A(n6779), .ZN(n14471) );
  AND2_X1 U8638 ( .A1(n6779), .A2(n6778), .ZN(n10427) );
  NAND2_X1 U8639 ( .A1(n10434), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U8640 ( .A1(n14512), .A2(n11735), .ZN(n11739) );
  INV_X1 U8641 ( .A(n14483), .ZN(n14542) );
  OAI21_X1 U8642 ( .B1(n14497), .B2(n13096), .A(n13095), .ZN(n6766) );
  NAND2_X1 U8643 ( .A1(n13099), .A2(n13379), .ZN(n13305) );
  XNOR2_X1 U8644 ( .A(n13106), .B(n13098), .ZN(n13099) );
  INV_X1 U8645 ( .A(n13097), .ZN(n13308) );
  XNOR2_X1 U8646 ( .A(n12039), .B(n12014), .ZN(n13312) );
  NAND2_X1 U8647 ( .A1(n13119), .A2(n12037), .ZN(n12039) );
  NAND2_X1 U8648 ( .A1(n7989), .A2(n7988), .ZN(n8135) );
  NAND2_X1 U8649 ( .A1(n6656), .A2(n6660), .ZN(n13157) );
  OAI21_X1 U8650 ( .B1(n13189), .B2(n6493), .A(n6664), .ZN(n13173) );
  NAND2_X1 U8651 ( .A1(n7143), .A2(n7141), .ZN(n13203) );
  OAI21_X1 U8652 ( .B1(n13275), .B2(n7006), .A(n7003), .ZN(n13223) );
  AOI21_X1 U8653 ( .B1(n13236), .B2(n13235), .A(n7148), .ZN(n13218) );
  NAND2_X1 U8654 ( .A1(n7008), .A2(n12031), .ZN(n13247) );
  NAND2_X1 U8655 ( .A1(n13275), .A2(n12030), .ZN(n7008) );
  AOI21_X1 U8656 ( .B1(n7127), .B2(n6670), .A(n12006), .ZN(n13253) );
  NAND2_X1 U8657 ( .A1(n7127), .A2(n7126), .ZN(n13266) );
  NAND2_X1 U8658 ( .A1(n13382), .A2(n12024), .ZN(n13298) );
  NAND2_X1 U8659 ( .A1(n6486), .A2(n6998), .ZN(n13382) );
  NAND2_X1 U8660 ( .A1(n6486), .A2(n11770), .ZN(n11772) );
  NAND2_X1 U8661 ( .A1(n7794), .A2(n7793), .ZN(n13378) );
  NAND2_X1 U8662 ( .A1(n7009), .A2(n7012), .ZN(n11709) );
  NAND2_X1 U8663 ( .A1(n11210), .A2(n7015), .ZN(n7009) );
  NAND2_X1 U8664 ( .A1(n11428), .A2(n11427), .ZN(n11723) );
  INV_X1 U8665 ( .A(n11136), .ZN(n11217) );
  NAND2_X1 U8666 ( .A1(n7017), .A2(n7019), .ZN(n11435) );
  NAND2_X1 U8667 ( .A1(n7018), .A2(n6544), .ZN(n7017) );
  INV_X1 U8668 ( .A(n11210), .ZN(n7018) );
  NAND2_X1 U8669 ( .A1(n10981), .A2(n10980), .ZN(n10983) );
  NAND2_X1 U8670 ( .A1(n6978), .A2(n10512), .ZN(n10513) );
  AND2_X1 U8671 ( .A1(n13257), .A2(n13093), .ZN(n13302) );
  NAND2_X1 U8672 ( .A1(n13317), .A2(n6638), .ZN(n13410) );
  AND2_X1 U8673 ( .A1(n13316), .A2(n6504), .ZN(n6638) );
  OR2_X1 U8674 ( .A1(n9921), .A2(n10190), .ZN(n14597) );
  OR2_X1 U8675 ( .A1(n10007), .A2(n14553), .ZN(n14551) );
  NOR2_X1 U8676 ( .A1(n7256), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n7255) );
  NAND2_X1 U8677 ( .A1(n7258), .A2(n7257), .ZN(n7256) );
  XNOR2_X1 U8678 ( .A(n7384), .B(n7383), .ZN(n12042) );
  INV_X1 U8679 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n7383) );
  OR2_X1 U8680 ( .A1(n13428), .A2(n14924), .ZN(n7384) );
  INV_X1 U8681 ( .A(n7386), .ZN(n13435) );
  INV_X1 U8682 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13439) );
  INV_X1 U8683 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11613) );
  NAND2_X1 U8684 ( .A1(n7213), .A2(n7214), .ZN(n8173) );
  XNOR2_X1 U8685 ( .A(n8172), .B(P2_IR_REG_24__SCAN_IN), .ZN(n11532) );
  INV_X1 U8686 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11391) );
  INV_X1 U8687 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10994) );
  INV_X1 U8688 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10097) );
  INV_X1 U8689 ( .A(n11737), .ZN(n13083) );
  INV_X1 U8690 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10142) );
  INV_X1 U8691 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10051) );
  XNOR2_X1 U8692 ( .A(n7710), .B(n7729), .ZN(n14510) );
  INV_X1 U8693 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9627) );
  INV_X1 U8694 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9554) );
  INV_X1 U8695 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9540) );
  INV_X1 U8696 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9536) );
  OR2_X1 U8697 ( .A1(n11040), .A2(n11039), .ZN(n7348) );
  AND2_X1 U8698 ( .A1(n14123), .A2(n14120), .ZN(n11899) );
  NAND2_X1 U8699 ( .A1(n13525), .A2(n12328), .ZN(n13457) );
  AOI22_X1 U8700 ( .A1(n13447), .A2(n13448), .B1(n12362), .B2(n12361), .ZN(
        n12371) );
  NAND2_X1 U8701 ( .A1(n11250), .A2(n7343), .ZN(n11251) );
  NAND2_X1 U8702 ( .A1(n12317), .A2(n12316), .ZN(n13482) );
  INV_X1 U8703 ( .A(n14291), .ZN(n11792) );
  NAND2_X1 U8704 ( .A1(n9207), .A2(n9206), .ZN(n13942) );
  NAND2_X1 U8705 ( .A1(n13566), .A2(n7344), .ZN(n13499) );
  NAND2_X1 U8706 ( .A1(n9080), .A2(n9079), .ZN(n14195) );
  AND2_X1 U8707 ( .A1(n7044), .A2(n6500), .ZN(n11419) );
  AND2_X1 U8708 ( .A1(n9759), .A2(n10034), .ZN(n14141) );
  AND2_X1 U8709 ( .A1(n14137), .A2(n14134), .ZN(n11783) );
  OR2_X1 U8710 ( .A1(n9765), .A2(n9758), .ZN(n13564) );
  NAND2_X1 U8711 ( .A1(n9224), .A2(n9223), .ZN(n13562) );
  INV_X1 U8712 ( .A(n13564), .ZN(n14139) );
  INV_X1 U8713 ( .A(n14146), .ZN(n13576) );
  XNOR2_X1 U8714 ( .A(n8829), .B(P1_IR_REG_2__SCAN_IN), .ZN(n13623) );
  XNOR2_X1 U8715 ( .A(n9031), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11392) );
  XNOR2_X1 U8716 ( .A(n13733), .B(n13732), .ZN(n13912) );
  INV_X1 U8717 ( .A(n13738), .ZN(n13915) );
  NAND2_X1 U8718 ( .A1(n14008), .A2(n9262), .ZN(n9253) );
  NAND2_X1 U8719 ( .A1(n7304), .A2(n11858), .ZN(n13786) );
  NAND2_X1 U8720 ( .A1(n6870), .A2(n11876), .ZN(n13814) );
  NAND2_X1 U8721 ( .A1(n11874), .A2(n6873), .ZN(n6870) );
  CLKBUF_X1 U8722 ( .A(n13810), .Z(n13811) );
  NAND2_X1 U8723 ( .A1(n11874), .A2(n11873), .ZN(n13826) );
  NAND2_X1 U8724 ( .A1(n13856), .A2(n11853), .ZN(n13849) );
  NAND2_X1 U8725 ( .A1(n7361), .A2(n11846), .ZN(n13898) );
  NAND2_X1 U8726 ( .A1(n9090), .A2(n9089), .ZN(n14154) );
  NAND2_X1 U8727 ( .A1(n7273), .A2(n7271), .ZN(n14151) );
  NAND2_X1 U8728 ( .A1(n11546), .A2(n11545), .ZN(n11548) );
  NAND2_X1 U8729 ( .A1(n9048), .A2(n6491), .ZN(n11832) );
  NAND2_X1 U8730 ( .A1(n11230), .A2(n11229), .ZN(n14280) );
  OR2_X1 U8731 ( .A1(n9905), .A2(n9766), .ZN(n14302) );
  NAND2_X1 U8732 ( .A1(n6863), .A2(n6867), .ZN(n10766) );
  OR2_X1 U8733 ( .A1(n10352), .A2(n10351), .ZN(n6863) );
  OR2_X1 U8734 ( .A1(n14318), .A2(n14349), .ZN(n13887) );
  NOR2_X1 U8735 ( .A1(n13880), .A2(n14357), .ZN(n13885) );
  NAND2_X1 U8736 ( .A1(n11885), .A2(n14302), .ZN(n14303) );
  INV_X1 U8737 ( .A(n14160), .ZN(n14314) );
  OR2_X1 U8738 ( .A1(n11885), .A2(n11272), .ZN(n14160) );
  INV_X1 U8739 ( .A(n14302), .ZN(n14285) );
  INV_X1 U8740 ( .A(n13883), .ZN(n14306) );
  NAND2_X1 U8741 ( .A1(n13916), .A2(n14353), .ZN(n13922) );
  NAND2_X1 U8742 ( .A1(n6634), .A2(n6511), .ZN(n13986) );
  INV_X1 U8743 ( .A(n6889), .ZN(n6634) );
  INV_X1 U8744 ( .A(n13925), .ZN(n6633) );
  AND2_X1 U8745 ( .A1(n13931), .A2(n7351), .ZN(n13932) );
  INV_X2 U8746 ( .A(n14376), .ZN(n14378) );
  OR2_X1 U8747 ( .A1(n11534), .A2(n9547), .ZN(n9741) );
  INV_X1 U8748 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7279) );
  NAND2_X1 U8749 ( .A1(n8103), .A2(n8102), .ZN(n14004) );
  INV_X1 U8750 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11616) );
  XNOR2_X1 U8751 ( .A(n7939), .B(n7938), .ZN(n11444) );
  INV_X1 U8752 ( .A(n9908), .ZN(n14017) );
  XNOR2_X1 U8753 ( .A(n9162), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14016) );
  INV_X1 U8754 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8816) );
  INV_X1 U8755 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10144) );
  INV_X1 U8756 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10070) );
  INV_X1 U8757 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9625) );
  INV_X1 U8758 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9592) );
  INV_X1 U8759 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9586) );
  INV_X1 U8760 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9573) );
  INV_X1 U8761 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9558) );
  INV_X1 U8762 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n14864) );
  NAND2_X1 U8763 ( .A1(n8878), .A2(n8877), .ZN(n9772) );
  NAND2_X1 U8764 ( .A1(n8828), .A2(n8770), .ZN(n8875) );
  NAND2_X1 U8765 ( .A1(n8855), .A2(n8854), .ZN(n13605) );
  INV_X1 U8766 ( .A(n6963), .ZN(n9421) );
  XNOR2_X1 U8767 ( .A(n9435), .B(n9434), .ZN(n14997) );
  XNOR2_X1 U8768 ( .A(n9438), .B(n6971), .ZN(n14035) );
  INV_X1 U8769 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6971) );
  XNOR2_X1 U8770 ( .A(n9445), .B(n6969), .ZN(n15000) );
  INV_X1 U8771 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6969) );
  XNOR2_X1 U8772 ( .A(n9448), .B(n9449), .ZN(n14036) );
  NAND2_X1 U8773 ( .A1(n14248), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6965) );
  OR2_X1 U8774 ( .A1(n14248), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6966) );
  AND2_X1 U8775 ( .A1(n9468), .A2(n9469), .ZN(n14259) );
  AND2_X1 U8776 ( .A1(n9475), .A2(n9474), .ZN(n14262) );
  AND2_X1 U8777 ( .A1(n9477), .A2(n9476), .ZN(n14050) );
  INV_X1 U8778 ( .A(n14263), .ZN(n9476) );
  OR2_X1 U8779 ( .A1(n14262), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n9477) );
  OR2_X1 U8780 ( .A1(n12312), .A2(n12311), .ZN(n7156) );
  NAND2_X1 U8781 ( .A1(n12140), .A2(n6602), .ZN(n7154) );
  OAI21_X1 U8782 ( .B1(n12306), .B2(n12305), .A(n9970), .ZN(n7153) );
  AOI21_X1 U8783 ( .B1(n14718), .B2(P3_IR_REG_0__SCAN_IN), .A(n7099), .ZN(
        n14611) );
  NOR2_X1 U8784 ( .A1(n14606), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14609) );
  AOI21_X1 U8785 ( .B1(n6782), .B2(n14746), .A(n6780), .ZN(n12635) );
  XNOR2_X1 U8786 ( .A(n6783), .B(n12624), .ZN(n6782) );
  NOR2_X1 U8787 ( .A1(n6852), .A2(n6853), .ZN(n6850) );
  NOR2_X1 U8788 ( .A1(n6852), .A2(n14828), .ZN(n6851) );
  OAI22_X1 U8789 ( .A1(n13040), .A2(n11955), .B1(n13045), .B2(n7124), .ZN(
        n11961) );
  AND2_X1 U8790 ( .A1(n13044), .A2(n6485), .ZN(n6615) );
  OAI211_X1 U8791 ( .C1(n13094), .C2(n13093), .A(n6767), .B(n6765), .ZN(
        P2_U3233) );
  INV_X1 U8792 ( .A(n6766), .ZN(n6765) );
  NAND2_X1 U8793 ( .A1(n6768), .A2(n13093), .ZN(n6767) );
  OAI21_X1 U8794 ( .B1(n13313), .B2(n13304), .A(n6918), .ZN(P2_U3236) );
  AND2_X1 U8795 ( .A1(n6920), .A2(n6919), .ZN(n6918) );
  AOI21_X1 U8796 ( .B1(n13309), .B2(n13302), .A(n12040), .ZN(n6919) );
  OR2_X1 U8797 ( .A1(n13312), .A2(n13299), .ZN(n6920) );
  OAI22_X1 U8798 ( .A1(n13170), .A2(n10997), .B1(n13294), .B2(n7124), .ZN(
        n10998) );
  NAND2_X1 U8799 ( .A1(n6926), .A2(n6925), .ZN(P2_U3496) );
  OR2_X1 U8800 ( .A1(n10992), .A2(n8075), .ZN(n6925) );
  NAND2_X1 U8801 ( .A1(n13409), .A2(n10992), .ZN(n6926) );
  AND2_X1 U8802 ( .A1(n9351), .A2(n7359), .ZN(n9352) );
  AOI21_X1 U8803 ( .B1(n6537), .B2(n9319), .A(n9318), .ZN(n9354) );
  NAND2_X1 U8804 ( .A1(n14045), .A2(n14046), .ZN(n14044) );
  OAI21_X1 U8805 ( .B1(n14020), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6508), .ZN(
        n6954) );
  INV_X1 U8806 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14924) );
  INV_X1 U8807 ( .A(n7486), .ZN(n8079) );
  INV_X1 U8808 ( .A(n9834), .ZN(n10541) );
  AND2_X1 U8809 ( .A1(n7166), .A2(n6684), .ZN(n6468) );
  NAND2_X1 U8810 ( .A1(n6714), .A2(n6583), .ZN(n6716) );
  OR2_X1 U8811 ( .A1(n13222), .A2(n7145), .ZN(n6469) );
  AND2_X1 U8812 ( .A1(n8771), .A2(n8772), .ZN(n6470) );
  AND2_X1 U8813 ( .A1(n6706), .A2(n6704), .ZN(n6471) );
  AND2_X1 U8814 ( .A1(n11262), .A2(n7294), .ZN(n6472) );
  INV_X1 U8815 ( .A(n13859), .ZN(n11851) );
  NAND2_X1 U8816 ( .A1(n12547), .A2(n11385), .ZN(n6473) );
  NAND2_X1 U8817 ( .A1(n12277), .A2(n12282), .ZN(n12682) );
  INV_X1 U8818 ( .A(n9290), .ZN(n11341) );
  MUX2_X1 U8819 ( .A(n14397), .B(n13445), .S(n7434), .Z(n10025) );
  AND4_X1 U8820 ( .A1(n7368), .A2(n7367), .A3(n7478), .A4(n7524), .ZN(n6475)
         );
  AND2_X1 U8821 ( .A1(n6885), .A2(n6884), .ZN(n6476) );
  INV_X1 U8822 ( .A(n12500), .ZN(n12540) );
  AND3_X1 U8823 ( .A1(n8249), .A2(n8248), .A3(n8247), .ZN(n12500) );
  NAND2_X1 U8824 ( .A1(n13873), .A2(n6887), .ZN(n6888) );
  NAND2_X1 U8825 ( .A1(n6495), .A2(n11358), .ZN(n6478) );
  NAND2_X1 U8826 ( .A1(n8609), .A2(n8608), .ZN(n12469) );
  INV_X1 U8827 ( .A(n12469), .ZN(n12834) );
  OR2_X1 U8828 ( .A1(n6553), .A2(n6741), .ZN(n6479) );
  OR2_X1 U8829 ( .A1(n12025), .A2(n7816), .ZN(n6480) );
  AND2_X1 U8830 ( .A1(n10903), .A2(n6722), .ZN(n6481) );
  AND2_X1 U8831 ( .A1(n10121), .A2(n6883), .ZN(n6482) );
  INV_X1 U8832 ( .A(n7717), .ZN(n7508) );
  AND2_X1 U8833 ( .A1(n6480), .A2(n6582), .ZN(n6483) );
  AND2_X1 U8834 ( .A1(n6532), .A2(n9281), .ZN(n6484) );
  AND2_X1 U8835 ( .A1(n13369), .A2(n12005), .ZN(n12006) );
  INV_X1 U8836 ( .A(n12234), .ZN(n6825) );
  OR2_X1 U8837 ( .A1(n13326), .A2(n13045), .ZN(n6485) );
  INV_X1 U8838 ( .A(n10522), .ZN(n6977) );
  INV_X1 U8839 ( .A(n14526), .ZN(n14536) );
  INV_X1 U8840 ( .A(n10507), .ZN(n6923) );
  INV_X1 U8841 ( .A(n14065), .ZN(n7106) );
  OR2_X1 U8842 ( .A1(n11769), .A2(n11768), .ZN(n6486) );
  OR2_X1 U8843 ( .A1(n13816), .A2(n13805), .ZN(n6487) );
  NAND2_X1 U8844 ( .A1(n11315), .A2(n11324), .ZN(n6488) );
  NOR2_X1 U8845 ( .A1(n12075), .A2(n12865), .ZN(n6489) );
  XNOR2_X1 U8846 ( .A(n8135), .B(n13049), .ZN(n6986) );
  AND2_X1 U8847 ( .A1(n6473), .A2(n8430), .ZN(n6490) );
  AOI21_X1 U8848 ( .B1(n12019), .B2(n13284), .A(n12018), .ZN(n13313) );
  AND2_X1 U8849 ( .A1(n6857), .A2(n6856), .ZN(n6491) );
  AND2_X1 U8850 ( .A1(n9124), .A2(n11871), .ZN(n13871) );
  OR2_X1 U8851 ( .A1(n12032), .A2(n7007), .ZN(n7006) );
  OR2_X1 U8852 ( .A1(n7190), .A2(n7186), .ZN(n6492) );
  NOR2_X1 U8853 ( .A1(n12009), .A2(n13053), .ZN(n6493) );
  OR3_X1 U8854 ( .A1(n11373), .A2(n12548), .A3(n11375), .ZN(n6495) );
  OAI211_X2 U8855 ( .C1(n9521), .C2(n6457), .A(n6494), .B(n8830), .ZN(n13540)
         );
  AND3_X1 U8856 ( .A1(n7087), .A2(n7088), .A3(n8937), .ZN(n6496) );
  AND2_X1 U8857 ( .A1(n10286), .A2(n8147), .ZN(n10278) );
  AND2_X1 U8858 ( .A1(n8003), .A2(n8002), .ZN(n13326) );
  INV_X1 U8859 ( .A(n13326), .ZN(n13150) );
  INV_X1 U8860 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6680) );
  AND2_X1 U8861 ( .A1(n13338), .A2(n13052), .ZN(n6497) );
  XOR2_X1 U8862 ( .A(n13387), .B(n12948), .Z(n6498) );
  AND2_X1 U8863 ( .A1(n6751), .A2(n13762), .ZN(n6499) );
  INV_X1 U8864 ( .A(n11941), .ZN(n10179) );
  NAND2_X1 U8865 ( .A1(n11415), .A2(n11414), .ZN(n6500) );
  AND4_X1 U8866 ( .A1(n7976), .A2(n7975), .A3(n7974), .A4(n7973), .ZN(n12952)
         );
  INV_X1 U8867 ( .A(n12952), .ZN(n13049) );
  XOR2_X1 U8868 ( .A(n13344), .B(n12948), .Z(n6501) );
  OR2_X1 U8869 ( .A1(n13952), .A2(n13827), .ZN(n6502) );
  AND2_X1 U8870 ( .A1(n9138), .A2(n9137), .ZN(n13971) );
  OR2_X1 U8871 ( .A1(n12633), .A2(n14709), .ZN(n6503) );
  OR2_X1 U8872 ( .A1(n13318), .A2(n14571), .ZN(n6504) );
  NAND2_X1 U8873 ( .A1(n14016), .A2(n9559), .ZN(n13835) );
  INV_X1 U8874 ( .A(n13835), .ZN(n13960) );
  XNOR2_X1 U8875 ( .A(n14978), .B(n7419), .ZN(n9647) );
  OR2_X1 U8876 ( .A1(n9449), .A2(n9448), .ZN(n6505) );
  NAND2_X1 U8877 ( .A1(n12914), .A2(n12915), .ZN(n6506) );
  AND2_X1 U8878 ( .A1(n12695), .A2(n12275), .ZN(n6810) );
  AND2_X1 U8879 ( .A1(n13398), .A2(n13062), .ZN(n6507) );
  INV_X1 U8880 ( .A(n7483), .ZN(n7253) );
  OR2_X1 U8881 ( .A1(n9486), .A2(n9485), .ZN(n6508) );
  INV_X1 U8882 ( .A(n11876), .ZN(n6872) );
  AND2_X1 U8883 ( .A1(n6500), .A2(n11418), .ZN(n6509) );
  NOR2_X1 U8884 ( .A1(n12845), .A2(n12500), .ZN(n8577) );
  XNOR2_X1 U8885 ( .A(n13046), .B(n13097), .ZN(n6510) );
  AND2_X1 U8886 ( .A1(n13928), .A2(n6633), .ZN(n6511) );
  INV_X1 U8887 ( .A(n6986), .ZN(n13131) );
  OR2_X1 U8888 ( .A1(n12842), .A2(n6626), .ZN(n6512) );
  INV_X1 U8889 ( .A(n6830), .ZN(n6829) );
  NAND2_X1 U8890 ( .A1(n6833), .A2(n6831), .ZN(n6830) );
  AND2_X1 U8891 ( .A1(n12701), .A2(n6841), .ZN(n6513) );
  INV_X1 U8892 ( .A(n9254), .ZN(n7095) );
  AND2_X1 U8893 ( .A1(n7143), .A2(n7142), .ZN(n6514) );
  INV_X1 U8894 ( .A(n9227), .ZN(n7071) );
  AND2_X1 U8895 ( .A1(n6847), .A2(n6848), .ZN(n6515) );
  AND2_X1 U8896 ( .A1(n13856), .A2(n7300), .ZN(n6516) );
  INV_X1 U8897 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7428) );
  AND2_X1 U8898 ( .A1(n11058), .A2(n14811), .ZN(n6517) );
  AND2_X1 U8899 ( .A1(n6977), .A2(n10512), .ZN(n6518) );
  INV_X1 U8900 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7396) );
  AND2_X1 U8901 ( .A1(n8017), .A2(n8016), .ZN(n13332) );
  INV_X1 U8902 ( .A(n13332), .ZN(n13167) );
  AND2_X1 U8903 ( .A1(n10641), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n6519) );
  AND2_X1 U8904 ( .A1(n12334), .A2(n12333), .ZN(n6520) );
  INV_X1 U8905 ( .A(n11653), .ZN(n11864) );
  INV_X1 U8906 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9085) );
  NOR2_X1 U8907 ( .A1(n11787), .A2(n14129), .ZN(n6521) );
  NAND2_X1 U8908 ( .A1(n11355), .A2(n11354), .ZN(n6522) );
  NOR2_X1 U8909 ( .A1(n13965), .A2(n13828), .ZN(n6523) );
  NOR2_X1 U8910 ( .A1(n13359), .A2(n13055), .ZN(n6524) );
  NOR2_X1 U8911 ( .A1(n11822), .A2(n12476), .ZN(n6525) );
  NOR2_X1 U8912 ( .A1(n13128), .A2(n12952), .ZN(n6526) );
  OR2_X1 U8913 ( .A1(n7052), .A2(n6484), .ZN(n6527) );
  XOR2_X1 U8914 ( .A(n9493), .B(n7360), .Z(n6528) );
  INV_X1 U8915 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7210) );
  OR2_X1 U8916 ( .A1(n13230), .A2(n13054), .ZN(n6529) );
  AND2_X1 U8917 ( .A1(n13167), .A2(n12985), .ZN(n6530) );
  AND2_X1 U8918 ( .A1(n9067), .A2(n9238), .ZN(n6531) );
  NOR2_X1 U8919 ( .A1(n9290), .A2(n9064), .ZN(n6532) );
  NOR2_X1 U8920 ( .A1(n12383), .A2(n12476), .ZN(n6533) );
  INV_X1 U8921 ( .A(n8974), .ZN(n7062) );
  INV_X1 U8922 ( .A(n7138), .ZN(n7137) );
  NOR2_X1 U8923 ( .A1(n13128), .A2(n13049), .ZN(n7138) );
  AND2_X1 U8924 ( .A1(n6814), .A2(n6812), .ZN(n6535) );
  INV_X1 U8925 ( .A(n12006), .ZN(n6671) );
  AND2_X1 U8926 ( .A1(n11277), .A2(n11276), .ZN(n6536) );
  AND2_X1 U8927 ( .A1(n7267), .A2(n7266), .ZN(n6537) );
  AND2_X1 U8928 ( .A1(n7659), .A2(SI_10_), .ZN(n6538) );
  AND2_X1 U8929 ( .A1(n7612), .A2(SI_8_), .ZN(n6539) );
  INV_X1 U8930 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7381) );
  AND2_X1 U8931 ( .A1(n7010), .A2(n11708), .ZN(n6540) );
  AND2_X1 U8932 ( .A1(n6744), .A2(n6752), .ZN(n6541) );
  NAND2_X1 U8933 ( .A1(n13600), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n6542) );
  NOR2_X1 U8934 ( .A1(n13927), .A2(n13452), .ZN(n6543) );
  NAND2_X1 U8935 ( .A1(n13403), .A2(n13063), .ZN(n6544) );
  INV_X1 U8936 ( .A(n12845), .ZN(n12505) );
  AND2_X1 U8937 ( .A1(n8237), .A2(n8236), .ZN(n12845) );
  AND2_X1 U8938 ( .A1(n8791), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6545) );
  AND2_X1 U8939 ( .A1(n8723), .A2(n8230), .ZN(n6546) );
  NAND2_X1 U8940 ( .A1(n13793), .A2(n11877), .ZN(n6547) );
  AND2_X1 U8941 ( .A1(n6712), .A2(n6711), .ZN(n6548) );
  AND2_X1 U8942 ( .A1(n12397), .A2(n12396), .ZN(n6549) );
  INV_X1 U8943 ( .A(n7364), .ZN(n6822) );
  OR2_X1 U8944 ( .A1(n12834), .A2(n12670), .ZN(n7364) );
  INV_X1 U8945 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7411) );
  NAND2_X1 U8946 ( .A1(n11346), .A2(n6488), .ZN(n6834) );
  OR2_X1 U8947 ( .A1(n7133), .A2(n12011), .ZN(n6550) );
  AND3_X1 U8948 ( .A1(n12278), .A2(n12277), .A3(n7177), .ZN(n6551) );
  NAND2_X1 U8949 ( .A1(n7962), .A2(n7961), .ZN(n13338) );
  OR2_X1 U8950 ( .A1(n8161), .A2(n6636), .ZN(n6552) );
  AND2_X1 U8951 ( .A1(n7780), .A2(SI_14_), .ZN(n6553) );
  NOR2_X1 U8952 ( .A1(n13850), .A2(n7301), .ZN(n7300) );
  AND2_X1 U8953 ( .A1(n7147), .A2(n7146), .ZN(n6554) );
  AND2_X1 U8954 ( .A1(n6716), .A2(n6715), .ZN(n6555) );
  AND2_X1 U8955 ( .A1(n10400), .A2(n10395), .ZN(n6556) );
  AND2_X1 U8956 ( .A1(n12886), .A2(n12884), .ZN(n6557) );
  INV_X1 U8957 ( .A(n9083), .ZN(n7078) );
  OR2_X1 U8958 ( .A1(n7095), .A2(n9255), .ZN(n6558) );
  OR2_X1 U8959 ( .A1(n7533), .A2(n7531), .ZN(n6559) );
  OR2_X1 U8960 ( .A1(n9154), .A2(n9152), .ZN(n6560) );
  NAND2_X1 U8961 ( .A1(n13454), .A2(n13560), .ZN(n6561) );
  AND2_X1 U8962 ( .A1(n9101), .A2(n9085), .ZN(n6562) );
  INV_X1 U8963 ( .A(n10758), .ZN(n10789) );
  OR2_X1 U8964 ( .A1(n7261), .A2(n7578), .ZN(n6563) );
  OR2_X1 U8965 ( .A1(n7577), .A2(n7579), .ZN(n6564) );
  AND2_X1 U8966 ( .A1(n7108), .A2(n7107), .ZN(n6565) );
  AND2_X1 U8967 ( .A1(n7211), .A2(n7210), .ZN(n6566) );
  INV_X1 U8968 ( .A(n6989), .ZN(n6988) );
  NAND2_X1 U8969 ( .A1(n13326), .A2(n12968), .ZN(n6989) );
  INV_X1 U8970 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8233) );
  NAND2_X1 U8971 ( .A1(n7715), .A2(n7235), .ZN(n6567) );
  NAND2_X1 U8972 ( .A1(n7668), .A2(n7238), .ZN(n6568) );
  NAND2_X1 U8973 ( .A1(n7943), .A2(n7241), .ZN(n6569) );
  INV_X1 U8974 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8721) );
  AND2_X1 U8975 ( .A1(n6952), .A2(n7334), .ZN(n6570) );
  NAND2_X1 U8976 ( .A1(n7090), .A2(n8938), .ZN(n6571) );
  OR2_X1 U8977 ( .A1(n7410), .A2(n7259), .ZN(n6572) );
  INV_X1 U8978 ( .A(n7006), .ZN(n7005) );
  OR2_X1 U8979 ( .A1(n13354), .A2(n13054), .ZN(n6573) );
  NAND2_X1 U8980 ( .A1(n7863), .A2(n7229), .ZN(n6574) );
  NAND2_X1 U8981 ( .A1(n7904), .A2(n7232), .ZN(n6575) );
  INV_X1 U8982 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8804) );
  INV_X1 U8983 ( .A(n7272), .ZN(n7271) );
  NAND2_X1 U8984 ( .A1(n7275), .A2(n14155), .ZN(n7272) );
  INV_X1 U8985 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8772) );
  INV_X1 U8986 ( .A(n7248), .ZN(n7247) );
  OAI21_X1 U8987 ( .B1(n7914), .B2(n7249), .A(n7952), .ZN(n7248) );
  NAND2_X1 U8988 ( .A1(n9055), .A2(n9054), .ZN(n11907) );
  INV_X1 U8989 ( .A(n11907), .ZN(n6891) );
  AND2_X1 U8990 ( .A1(n8617), .A2(n8616), .ZN(n12670) );
  INV_X1 U8991 ( .A(n12670), .ZN(n7178) );
  AND2_X1 U8992 ( .A1(n11173), .A2(n11172), .ZN(n6576) );
  NAND2_X1 U8993 ( .A1(n6649), .A2(n6648), .ZN(n11131) );
  OR2_X1 U8994 ( .A1(n11521), .A2(n11522), .ZN(n11695) );
  NAND2_X1 U8995 ( .A1(n8652), .A2(n8651), .ZN(n12652) );
  AND2_X1 U8996 ( .A1(n6943), .A2(n14732), .ZN(n6577) );
  INV_X1 U8997 ( .A(n12252), .ZN(n6786) );
  INV_X1 U8998 ( .A(n8457), .ZN(n7176) );
  NAND2_X1 U8999 ( .A1(n11598), .A2(n7363), .ZN(n11682) );
  NAND2_X1 U9000 ( .A1(n11541), .A2(n11540), .ZN(n11655) );
  NAND2_X1 U9001 ( .A1(n6787), .A2(n12251), .ZN(n11685) );
  NAND2_X1 U9002 ( .A1(n7293), .A2(n11228), .ZN(n11263) );
  XNOR2_X1 U9003 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8255) );
  INV_X1 U9004 ( .A(n8255), .ZN(n7165) );
  INV_X1 U9005 ( .A(n6464), .ZN(n9117) );
  INV_X1 U9006 ( .A(n13952), .ZN(n6884) );
  NAND2_X1 U9007 ( .A1(n7861), .A2(n7860), .ZN(n13365) );
  OR2_X1 U9008 ( .A1(n9084), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n6578) );
  NAND2_X1 U9009 ( .A1(n11724), .A2(n11768), .ZN(n11762) );
  INV_X1 U9010 ( .A(n12225), .ZN(n6806) );
  NOR2_X1 U9011 ( .A1(n11296), .A2(n11187), .ZN(n6579) );
  INV_X1 U9012 ( .A(n6892), .ZN(n11550) );
  NOR2_X1 U9013 ( .A1(n11328), .A2(n14210), .ZN(n6892) );
  OR2_X1 U9014 ( .A1(n12912), .A2(n12911), .ZN(n6580) );
  AND2_X1 U9015 ( .A1(n12494), .A2(n7325), .ZN(n6581) );
  OR2_X1 U9016 ( .A1(n7814), .A2(n7815), .ZN(n6582) );
  NAND2_X1 U9017 ( .A1(n13053), .A2(n10256), .ZN(n6583) );
  OR2_X1 U9018 ( .A1(n11642), .A2(n11645), .ZN(n6584) );
  INV_X1 U9019 ( .A(n6930), .ZN(n13271) );
  NOR2_X2 U9020 ( .A1(n13287), .A2(n13369), .ZN(n6930) );
  AND2_X1 U9021 ( .A1(n7115), .A2(n7114), .ZN(n6585) );
  AND2_X1 U9022 ( .A1(n7313), .A2(n7311), .ZN(n6586) );
  INV_X1 U9023 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9828) );
  INV_X1 U9024 ( .A(n13295), .ZN(n13374) );
  AND2_X1 U9025 ( .A1(n7813), .A2(n7812), .ZN(n13295) );
  AND2_X1 U9026 ( .A1(n9625), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6587) );
  AND2_X1 U9027 ( .A1(n6832), .A2(n6829), .ZN(n6588) );
  INV_X1 U9028 ( .A(n6936), .ZN(n6935) );
  NAND2_X1 U9029 ( .A1(n6938), .A2(n11190), .ZN(n6936) );
  INV_X1 U9030 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9783) );
  OR2_X1 U9031 ( .A1(n13392), .A2(n11720), .ZN(n6589) );
  AND2_X1 U9032 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n6590) );
  AND2_X1 U9033 ( .A1(n6577), .A2(n6934), .ZN(n6591) );
  AND2_X1 U9034 ( .A1(n6967), .A2(n6968), .ZN(n6592) );
  INV_X2 U9035 ( .A(n14388), .ZN(n14391) );
  NAND2_X1 U9036 ( .A1(n13257), .A2(n10574), .ZN(n13294) );
  NAND2_X1 U9037 ( .A1(n7713), .A2(n7712), .ZN(n13398) );
  INV_X1 U9038 ( .A(n13398), .ZN(n6931) );
  AND2_X1 U9039 ( .A1(n10746), .A2(n10745), .ZN(n6593) );
  AND2_X1 U9040 ( .A1(n8564), .A2(n7194), .ZN(n6594) );
  INV_X1 U9041 ( .A(n12605), .ZN(n12593) );
  INV_X1 U9042 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11145) );
  NAND2_X1 U9043 ( .A1(n10925), .A2(n12197), .ZN(n10908) );
  NAND2_X1 U9044 ( .A1(n6855), .A2(n10162), .ZN(n10222) );
  NAND2_X1 U9045 ( .A1(n7284), .A2(n10150), .ZN(n10221) );
  NAND2_X1 U9046 ( .A1(n10740), .A2(n10866), .ZN(n10746) );
  NAND2_X1 U9047 ( .A1(n10521), .A2(n10520), .ZN(n10523) );
  NOR2_X1 U9048 ( .A1(n14729), .A2(n10591), .ZN(n6595) );
  OR2_X1 U9049 ( .A1(n11198), .A2(n10657), .ZN(n6596) );
  INV_X1 U9050 ( .A(n7015), .ZN(n7014) );
  NOR2_X1 U9051 ( .A1(n7016), .A2(n11434), .ZN(n7015) );
  NOR2_X1 U9052 ( .A1(n14670), .A2(n14669), .ZN(n6597) );
  OR2_X1 U9053 ( .A1(n8579), .A2(n7192), .ZN(n6598) );
  INV_X1 U9054 ( .A(n7151), .ZN(n7382) );
  NAND2_X1 U9055 ( .A1(n7191), .A2(n6688), .ZN(n6599) );
  AND2_X1 U9056 ( .A1(n6835), .A2(n6488), .ZN(n6600) );
  INV_X1 U9057 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9886) );
  INV_X1 U9058 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n6674) );
  INV_X1 U9059 ( .A(n11045), .ZN(n6881) );
  NAND2_X1 U9060 ( .A1(n7688), .A2(n7687), .ZN(n13403) );
  INV_X1 U9061 ( .A(n13403), .ZN(n7020) );
  INV_X1 U9062 ( .A(n14054), .ZN(n12609) );
  NAND2_X1 U9063 ( .A1(n10776), .A2(n8141), .ZN(n10571) );
  INV_X1 U9064 ( .A(n10571), .ZN(n6924) );
  AND2_X1 U9065 ( .A1(n6758), .A2(n6756), .ZN(n6601) );
  AND2_X1 U9066 ( .A1(n9970), .A2(n9974), .ZN(n6602) );
  AND2_X1 U9067 ( .A1(n8360), .A2(n8359), .ZN(n6603) );
  INV_X1 U9068 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13442) );
  AND2_X1 U9069 ( .A1(n9970), .A2(n7155), .ZN(n6604) );
  INV_X1 U9070 ( .A(SI_26_), .ZN(n11691) );
  OR2_X1 U9071 ( .A1(n14054), .A2(n12585), .ZN(n6605) );
  INV_X1 U9072 ( .A(n10556), .ZN(n11272) );
  AND2_X1 U9073 ( .A1(n14041), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n6606) );
  AND2_X1 U9074 ( .A1(n7382), .A2(n7255), .ZN(n13428) );
  INV_X1 U9075 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6771) );
  OAI222_X1 U9076 ( .A1(P3_U3151), .A2(n6630), .B1(n12880), .B2(n12879), .C1(
        n14863), .C2(n12874), .ZN(P3_U3267) );
  AOI21_X1 U9077 ( .B1(n13628), .B2(n13627), .A(n13626), .ZN(n13625) );
  INV_X1 U9078 ( .A(n6607), .ZN(n13727) );
  XNOR2_X1 U9079 ( .A(n13715), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n6607) );
  NAND2_X1 U9080 ( .A1(n13701), .A2(n6624), .ZN(n13712) );
  NOR2_X1 U9081 ( .A1(n11404), .A2(n14265), .ZN(n11407) );
  NOR2_X1 U9082 ( .A1(n9816), .A2(n9815), .ZN(n10378) );
  NOR2_X1 U9083 ( .A1(n9708), .A2(n9707), .ZN(n9706) );
  AOI21_X1 U9084 ( .B1(n11372), .B2(n10381), .A(n13687), .ZN(n10384) );
  AOI21_X1 U9085 ( .B1(n11401), .B2(n14216), .A(n11400), .ZN(n11403) );
  OAI21_X1 U9086 ( .B1(n9697), .B2(n9695), .A(n9696), .ZN(n9814) );
  AOI21_X1 U9087 ( .B1(n13636), .B2(n13635), .A(n13634), .ZN(n13638) );
  NAND2_X1 U9088 ( .A1(n7251), .A2(n7250), .ZN(n7554) );
  NAND2_X1 U9089 ( .A1(n7240), .A2(n7239), .ZN(n7965) );
  NAND2_X1 U9090 ( .A1(n7820), .A2(n7819), .ZN(n7834) );
  NAND2_X1 U9091 ( .A1(n7254), .A2(n7252), .ZN(n7505) );
  OAI21_X1 U9092 ( .B1(n7354), .B2(n8090), .A(n8089), .ZN(n8119) );
  XNOR2_X2 U9093 ( .A(n7403), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9870) );
  NAND2_X1 U9094 ( .A1(n6534), .A2(n8916), .ZN(n9076) );
  INV_X1 U9095 ( .A(n13810), .ZN(n6610) );
  INV_X1 U9096 ( .A(n8782), .ZN(n14005) );
  INV_X1 U9097 ( .A(n11342), .ZN(n6609) );
  NAND2_X1 U9098 ( .A1(n13869), .A2(n11870), .ZN(n11850) );
  NAND2_X1 U9099 ( .A1(n13858), .A2(n7300), .ZN(n6614) );
  NAND2_X1 U9100 ( .A1(n10110), .A2(n10109), .ZN(n10113) );
  OAI21_X1 U9101 ( .B1(n10149), .B2(n7285), .A(n7282), .ZN(n7286) );
  NAND2_X2 U9102 ( .A1(n6609), .A2(n9290), .ZN(n11546) );
  NAND2_X1 U9103 ( .A1(n14307), .A2(n14308), .ZN(n10115) );
  NAND2_X1 U9104 ( .A1(n6614), .A2(n7299), .ZN(n13836) );
  XNOR2_X2 U9105 ( .A(n13540), .B(n6611), .ZN(n10109) );
  NAND2_X1 U9106 ( .A1(n11546), .A2(n7296), .ZN(n11652) );
  XNOR2_X2 U9107 ( .A(n10552), .B(n10164), .ZN(n10223) );
  NAND2_X1 U9108 ( .A1(n6616), .A2(n6615), .ZN(P2_U3212) );
  NAND2_X1 U9109 ( .A1(n13036), .A2(n13035), .ZN(n6616) );
  NAND2_X1 U9110 ( .A1(n11971), .A2(n11978), .ZN(n12885) );
  NAND2_X2 U9111 ( .A1(n12983), .A2(n6580), .ZN(n12966) );
  NAND2_X1 U9112 ( .A1(n6906), .A2(n6904), .ZN(n7853) );
  NAND2_X2 U9113 ( .A1(n7205), .A2(n11967), .ZN(n11977) );
  NAND2_X1 U9114 ( .A1(n7209), .A2(n7207), .ZN(n12991) );
  XNOR2_X1 U9115 ( .A(n12909), .B(n6501), .ZN(n12931) );
  NAND2_X1 U9116 ( .A1(n8688), .A2(n12190), .ZN(n10923) );
  OAI22_X2 U9117 ( .A1(n12731), .A2(n8704), .B1(n12849), .B2(n12541), .ZN(
        n12720) );
  AOI21_X2 U9118 ( .B1(n9376), .B2(n12289), .A(n9375), .ZN(n12100) );
  NAND2_X1 U9119 ( .A1(n12078), .A2(n6854), .ZN(n9495) );
  AND2_X2 U9120 ( .A1(n13146), .A2(n13128), .ZN(n13130) );
  NAND3_X1 U9121 ( .A1(n9245), .A2(n6620), .A3(n6558), .ZN(n7093) );
  NAND2_X1 U9122 ( .A1(n9244), .A2(n9243), .ZN(n6620) );
  NAND3_X1 U9123 ( .A1(n9143), .A2(n9142), .A3(n6560), .ZN(n6622) );
  OR2_X1 U9124 ( .A1(n9889), .A2(n8145), .ZN(n10773) );
  NAND2_X1 U9125 ( .A1(n11714), .A2(n11713), .ZN(n11760) );
  OR2_X2 U9126 ( .A1(n10855), .A2(n11090), .ZN(n10985) );
  NAND2_X1 U9127 ( .A1(n13224), .A2(n13230), .ZN(n13226) );
  NAND2_X1 U9128 ( .A1(n6692), .A2(n7572), .ZN(n7587) );
  OR2_X1 U9129 ( .A1(n9195), .A2(n9196), .ZN(n9197) );
  OAI21_X1 U9130 ( .B1(n9258), .B2(n9257), .A(n9256), .ZN(n9259) );
  OAI211_X1 U9131 ( .C1(n13312), .C2(n14571), .A(n13311), .B(n13313), .ZN(
        n13409) );
  NAND2_X4 U9132 ( .A1(n8846), .A2(n14009), .ZN(n9559) );
  NAND2_X2 U9133 ( .A1(n7024), .A2(n7021), .ZN(n14009) );
  NAND2_X1 U9134 ( .A1(n11327), .A2(n14219), .ZN(n11328) );
  NOR2_X4 U9135 ( .A1(n13874), .A2(n13902), .ZN(n13873) );
  NOR2_X2 U9136 ( .A1(n11660), .A2(n14195), .ZN(n14159) );
  NAND2_X1 U9137 ( .A1(n7292), .A2(n7291), .ZN(n11338) );
  XNOR2_X1 U9138 ( .A(n10237), .B(n11956), .ZN(n10027) );
  NAND2_X1 U9139 ( .A1(n12991), .A2(n12901), .ZN(n12959) );
  NAND2_X1 U9140 ( .A1(n12936), .A2(n12935), .ZN(n7209) );
  NAND2_X1 U9141 ( .A1(n10241), .A2(n11957), .ZN(n11964) );
  NAND2_X1 U9142 ( .A1(n11520), .A2(n11519), .ZN(n11521) );
  NOR2_X1 U9143 ( .A1(n9430), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n9387) );
  XNOR2_X1 U9144 ( .A(n9388), .B(n14650), .ZN(n9418) );
  NAND2_X1 U9145 ( .A1(n6623), .A2(n9432), .ZN(n9435) );
  NAND2_X1 U9146 ( .A1(n14996), .A2(n14995), .ZN(n6623) );
  NAND2_X1 U9147 ( .A1(n9455), .A2(n6960), .ZN(n6959) );
  NAND2_X2 U9148 ( .A1(n10961), .A2(n10960), .ZN(n11314) );
  NAND2_X1 U9149 ( .A1(n7310), .A2(n7309), .ZN(n12474) );
  INV_X1 U9150 ( .A(n7327), .ZN(n12398) );
  XNOR2_X1 U9151 ( .A(n6954), .B(n6528), .ZN(SUB_1596_U4) );
  NAND2_X1 U9152 ( .A1(n7464), .A2(n7465), .ZN(n7463) );
  NAND3_X1 U9153 ( .A1(n7444), .A2(n7442), .A3(n7443), .ZN(n7464) );
  NAND3_X1 U9154 ( .A1(n7507), .A2(n7506), .A3(n6559), .ZN(n7251) );
  OAI211_X1 U9155 ( .C1(n7253), .C2(n7482), .A(n7469), .B(n7468), .ZN(n7254)
         );
  NOR2_X1 U9156 ( .A1(n9833), .A2(n10176), .ZN(n9838) );
  OAI211_X1 U9157 ( .C1(n6551), .C2(n7161), .A(n12445), .B(n7158), .ZN(n12295)
         );
  NAND2_X1 U9158 ( .A1(n8802), .A2(n8801), .ZN(n8810) );
  XNOR2_X1 U9159 ( .A(n10182), .B(n6631), .ZN(n13538) );
  NAND2_X1 U9160 ( .A1(n10061), .A2(n10060), .ZN(n10396) );
  NAND2_X1 U9161 ( .A1(n12437), .A2(n12436), .ZN(n12435) );
  NAND2_X1 U9162 ( .A1(n9981), .A2(n9980), .ZN(n10054) );
  AOI21_X2 U9163 ( .B1(n11314), .B2(n7320), .A(n6478), .ZN(n11558) );
  INV_X1 U9164 ( .A(n14308), .ZN(n14298) );
  NAND2_X1 U9165 ( .A1(n10107), .A2(n8883), .ZN(n14308) );
  NAND2_X2 U9166 ( .A1(n6635), .A2(n7458), .ZN(n7475) );
  NAND2_X1 U9167 ( .A1(n7455), .A2(n7456), .ZN(n6635) );
  INV_X2 U9168 ( .A(n7417), .ZN(n7459) );
  NAND2_X1 U9169 ( .A1(n6693), .A2(n7546), .ZN(n7569) );
  NAND4_X1 U9170 ( .A1(n6510), .A2(n8162), .A3(n12038), .A4(n6637), .ZN(n6636)
         );
  NOR2_X2 U9171 ( .A1(n7379), .A2(n7380), .ZN(n7214) );
  AND2_X2 U9172 ( .A1(n6475), .A2(n7452), .ZN(n7590) );
  NAND2_X1 U9173 ( .A1(n11214), .A2(n11213), .ZN(n11428) );
  OAI21_X1 U9174 ( .B1(n13189), .B2(n6659), .A(n6657), .ZN(n13155) );
  NAND2_X1 U9175 ( .A1(n7127), .A2(n6668), .ZN(n6667) );
  NAND4_X1 U9176 ( .A1(n7154), .A2(n7153), .A3(n7156), .A4(n6676), .ZN(
        P3_U3296) );
  NAND2_X1 U9177 ( .A1(n6677), .A2(n6604), .ZN(n6676) );
  XNOR2_X1 U9178 ( .A(n6678), .B(n12623), .ZN(n6677) );
  OR2_X1 U9179 ( .A1(n12104), .A2(n12103), .ZN(n6678) );
  NAND2_X1 U9180 ( .A1(n8566), .A2(n6687), .ZN(n6686) );
  NAND2_X1 U9181 ( .A1(n7569), .A2(n7568), .ZN(n6692) );
  NAND2_X1 U9182 ( .A1(n7544), .A2(n7543), .ZN(n6693) );
  INV_X1 U9183 ( .A(n6893), .ZN(n6697) );
  NAND2_X1 U9184 ( .A1(n7519), .A2(n7518), .ZN(n7522) );
  NAND3_X1 U9185 ( .A1(n6696), .A2(n7495), .A3(n6695), .ZN(n7519) );
  NAND3_X1 U9186 ( .A1(n6697), .A2(n6698), .A3(n7492), .ZN(n6696) );
  OAI21_X1 U9187 ( .B1(n6893), .B2(n7474), .A(n7476), .ZN(n7493) );
  NAND2_X1 U9188 ( .A1(n11999), .A2(n11699), .ZN(n11965) );
  NAND2_X1 U9189 ( .A1(n12966), .A2(n6471), .ZN(n6702) );
  OR2_X1 U9190 ( .A1(n12966), .A2(n6708), .ZN(n6705) );
  NAND2_X1 U9191 ( .A1(n6702), .A2(n6703), .ZN(n12951) );
  NAND2_X1 U9192 ( .A1(n12966), .A2(n12965), .ZN(n6710) );
  INV_X1 U9193 ( .A(n12931), .ZN(n6714) );
  XNOR2_X1 U9194 ( .A(n10902), .B(n10898), .ZN(n10752) );
  NAND2_X2 U9195 ( .A1(n7263), .A2(n7262), .ZN(n7416) );
  NAND3_X1 U9196 ( .A1(n7263), .A2(n7262), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n6724) );
  INV_X1 U9197 ( .A(n7899), .ZN(n6732) );
  NAND2_X1 U9198 ( .A1(n6733), .A2(n6734), .ZN(n7787) );
  NAND2_X1 U9199 ( .A1(n7680), .A2(n6735), .ZN(n6733) );
  NAND2_X1 U9200 ( .A1(n13763), .A2(n6499), .ZN(n6749) );
  NAND2_X1 U9201 ( .A1(n13763), .A2(n13762), .ZN(n12043) );
  AND2_X1 U9202 ( .A1(n6749), .A2(n6748), .ZN(n13744) );
  AOI21_X1 U9203 ( .B1(n9643), .B2(n6756), .A(n6754), .ZN(n14442) );
  MUX2_X1 U9204 ( .A(n14835), .B(P3_REG1_REG_2__SCAN_IN), .S(n10334), .Z(
        n10313) );
  NAND2_X1 U9205 ( .A1(n12171), .A2(n12174), .ZN(n12116) );
  NAND2_X1 U9206 ( .A1(n10201), .A2(n14754), .ZN(n12171) );
  NAND2_X1 U9207 ( .A1(n11602), .A2(n6788), .ZN(n6784) );
  NAND2_X1 U9208 ( .A1(n6784), .A2(n6785), .ZN(n11801) );
  NAND2_X1 U9209 ( .A1(n6791), .A2(n6792), .ZN(n11012) );
  NAND2_X1 U9210 ( .A1(n10923), .A2(n6793), .ZN(n6791) );
  NAND2_X1 U9211 ( .A1(n8509), .A2(n7353), .ZN(n8720) );
  NAND2_X1 U9212 ( .A1(n6570), .A2(n8509), .ZN(n8232) );
  NAND2_X1 U9213 ( .A1(n12688), .A2(n6799), .ZN(n6798) );
  NAND2_X2 U9214 ( .A1(n6798), .A2(n6796), .ZN(n12662) );
  NAND2_X1 U9215 ( .A1(n6804), .A2(n6802), .ZN(n8691) );
  NOR2_X1 U9216 ( .A1(n6806), .A2(n6803), .ZN(n6802) );
  INV_X1 U9217 ( .A(n12214), .ZN(n6803) );
  NAND2_X1 U9218 ( .A1(n8690), .A2(n8689), .ZN(n11104) );
  NAND2_X1 U9219 ( .A1(n12775), .A2(n6807), .ZN(n8702) );
  NAND2_X1 U9220 ( .A1(n12711), .A2(n12142), .ZN(n6811) );
  NAND2_X1 U9221 ( .A1(n6811), .A2(n6810), .ZN(n8705) );
  XNOR2_X1 U9222 ( .A(n9376), .B(n12445), .ZN(n12649) );
  NAND2_X1 U9223 ( .A1(n6815), .A2(n8222), .ZN(n7330) );
  NAND2_X4 U9224 ( .A1(n10307), .A2(n9501), .ZN(n12096) );
  NAND2_X4 U9225 ( .A1(n8680), .A2(n6422), .ZN(n10307) );
  NAND2_X1 U9226 ( .A1(n10445), .A2(n8375), .ZN(n10727) );
  NAND2_X1 U9227 ( .A1(n12656), .A2(n8646), .ZN(n12655) );
  INV_X1 U9228 ( .A(n8632), .ZN(n6823) );
  NAND2_X1 U9229 ( .A1(n11289), .A2(n6827), .ZN(n6826) );
  NAND2_X1 U9230 ( .A1(n11600), .A2(n6838), .ZN(n6836) );
  NAND2_X1 U9231 ( .A1(n6836), .A2(n6837), .ZN(n11799) );
  NAND2_X1 U9232 ( .A1(n12717), .A2(n6843), .ZN(n6842) );
  NAND2_X1 U9233 ( .A1(n7365), .A2(n14106), .ZN(n6854) );
  OAI21_X1 U9234 ( .B1(n12078), .B2(n6852), .A(n6849), .ZN(P3_U3456) );
  AOI21_X1 U9235 ( .B1(n7365), .B2(n6851), .A(n6850), .ZN(n6849) );
  NAND2_X1 U9236 ( .A1(n10222), .A2(n10163), .ZN(n10166) );
  NAND2_X1 U9237 ( .A1(n10160), .A2(n10159), .ZN(n6855) );
  OAI22_X1 U9238 ( .A1(n8895), .A2(n9542), .B1(n9559), .B2(n9609), .ZN(n8820)
         );
  OAI22_X1 U9239 ( .A1(n8895), .A2(n14864), .B1(n9559), .B2(n9717), .ZN(n8918)
         );
  OAI22_X1 U9240 ( .A1(n8895), .A2(n9573), .B1(n9559), .B2(n9617), .ZN(n8947)
         );
  OAI22_X1 U9241 ( .A1(n8895), .A2(n9558), .B1(n9559), .B2(n9813), .ZN(n8925)
         );
  OAI22_X1 U9242 ( .A1(n8895), .A2(n9586), .B1(n9559), .B2(n9700), .ZN(n8970)
         );
  OAI22_X1 U9243 ( .A1(n8895), .A2(n10053), .B1(n9559), .B2(n11591), .ZN(n9078) );
  OAI22_X1 U9244 ( .A1(n6457), .A2(n10144), .B1(n9559), .B2(n13702), .ZN(n9088) );
  OAI22_X1 U9245 ( .A1(n8895), .A2(n10457), .B1(n9559), .B2(n13711), .ZN(n9103) );
  OAI22_X1 U9246 ( .A1(n8895), .A2(n10557), .B1(n9559), .B2(n10556), .ZN(n9109) );
  NAND2_X1 U9247 ( .A1(n9271), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n6856) );
  OR2_X1 U9248 ( .A1(n10415), .A2(n9559), .ZN(n6857) );
  NAND2_X1 U9249 ( .A1(n10352), .A2(n6859), .ZN(n6861) );
  NAND2_X1 U9250 ( .A1(n6860), .A2(n10788), .ZN(n10793) );
  NAND3_X1 U9251 ( .A1(n10758), .A2(n6861), .A3(n6862), .ZN(n6860) );
  INV_X1 U9252 ( .A(n10793), .ZN(n10792) );
  NAND2_X1 U9253 ( .A1(n6861), .A2(n6862), .ZN(n10790) );
  NAND2_X1 U9254 ( .A1(n6871), .A2(n11874), .ZN(n6869) );
  OR2_X1 U9255 ( .A1(n7272), .A2(n11541), .ZN(n6875) );
  NAND2_X1 U9256 ( .A1(n6875), .A2(n6876), .ZN(n13888) );
  INV_X1 U9257 ( .A(n6888), .ZN(n13830) );
  AND2_X1 U9258 ( .A1(n13755), .A2(n13754), .ZN(n13925) );
  XNOR2_X1 U9259 ( .A(n6893), .B(n7474), .ZN(n9529) );
  XNOR2_X2 U9260 ( .A(n7475), .B(SI_2_), .ZN(n6893) );
  XNOR2_X1 U9261 ( .A(n8037), .B(n7987), .ZN(n11841) );
  NAND2_X1 U9262 ( .A1(n7803), .A2(n6908), .ZN(n6906) );
  NAND2_X1 U9263 ( .A1(n7633), .A2(n6912), .ZN(n6911) );
  NAND2_X1 U9264 ( .A1(n7898), .A2(n6917), .ZN(n6916) );
  NOR2_X2 U9265 ( .A1(n10525), .A2(n10694), .ZN(n10950) );
  NOR2_X2 U9266 ( .A1(n10773), .A2(n10772), .ZN(n10776) );
  NOR3_X4 U9267 ( .A1(n6927), .A2(n13207), .A3(n13150), .ZN(n13146) );
  NOR2_X2 U9268 ( .A1(n11760), .A2(n13378), .ZN(n13286) );
  NOR2_X2 U9269 ( .A1(n11432), .A2(n13392), .ZN(n11714) );
  NAND2_X1 U9270 ( .A1(n14734), .A2(n6591), .ZN(n6933) );
  NAND2_X1 U9271 ( .A1(n6937), .A2(n6938), .ZN(n11191) );
  NOR2_X2 U9272 ( .A1(n10308), .A2(n6423), .ZN(n14746) );
  NAND2_X1 U9273 ( .A1(n14043), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n6961) );
  OAI211_X2 U9274 ( .C1(n6961), .C2(n6958), .A(n6957), .B(n6955), .ZN(n14244)
         );
  INV_X1 U9275 ( .A(n14243), .ZN(n6968) );
  OAI21_X2 U9276 ( .B1(n6964), .B2(n14243), .A(n6965), .ZN(n14252) );
  NAND2_X1 U9277 ( .A1(n6967), .A2(n6966), .ZN(n6964) );
  NAND3_X1 U9278 ( .A1(n6968), .A2(n6967), .A3(n14248), .ZN(n14247) );
  NAND2_X1 U9279 ( .A1(n14252), .A2(n14251), .ZN(n14250) );
  XNOR2_X1 U9280 ( .A(n9433), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n9434) );
  NAND2_X1 U9281 ( .A1(n6970), .A2(n9442), .ZN(n9445) );
  NAND2_X1 U9282 ( .A1(n10506), .A2(n10505), .ZN(n6972) );
  NAND2_X1 U9283 ( .A1(n10563), .A2(n10566), .ZN(n6973) );
  NAND2_X1 U9284 ( .A1(n6974), .A2(n10281), .ZN(n10771) );
  NAND2_X1 U9285 ( .A1(n10280), .A2(n10279), .ZN(n6974) );
  OAI211_X1 U9286 ( .C1(n10280), .C2(n6976), .A(n6975), .B(n10288), .ZN(n10284) );
  INV_X1 U9287 ( .A(n10281), .ZN(n6976) );
  NAND2_X1 U9288 ( .A1(n10947), .A2(n10946), .ZN(n6978) );
  NAND2_X1 U9289 ( .A1(n13144), .A2(n6982), .ZN(n6981) );
  NAND2_X1 U9290 ( .A1(n13144), .A2(n12036), .ZN(n6987) );
  NAND2_X1 U9291 ( .A1(n13162), .A2(n13161), .ZN(n13160) );
  INV_X1 U9292 ( .A(n7000), .ZN(n13214) );
  OAI211_X1 U9293 ( .C1(n13275), .C2(n7002), .A(n7001), .B(n6573), .ZN(n7000)
         );
  NAND2_X1 U9294 ( .A1(n7005), .A2(n13222), .ZN(n7002) );
  NAND2_X1 U9295 ( .A1(n13536), .A2(n10184), .ZN(n10185) );
  NOR2_X1 U9296 ( .A1(n10186), .A2(n7028), .ZN(n7027) );
  INV_X1 U9297 ( .A(n10184), .ZN(n7028) );
  NAND2_X1 U9298 ( .A1(n7032), .A2(n7033), .ZN(n13517) );
  OR2_X1 U9299 ( .A1(n11784), .A2(n11785), .ZN(n7041) );
  INV_X1 U9300 ( .A(n7044), .ZN(n11416) );
  AND2_X4 U9301 ( .A1(n7045), .A2(n9311), .ZN(n9238) );
  NAND2_X1 U9302 ( .A1(n9313), .A2(n7045), .ZN(n9314) );
  NAND2_X1 U9303 ( .A1(n7047), .A2(n7046), .ZN(n9069) );
  NAND3_X1 U9304 ( .A1(n9026), .A2(n9025), .A3(n6527), .ZN(n7047) );
  NAND2_X1 U9305 ( .A1(n7059), .A2(n8960), .ZN(n7054) );
  NAND2_X1 U9306 ( .A1(n7055), .A2(n7053), .ZN(n8990) );
  OAI21_X1 U9307 ( .B1(n8869), .B2(n7065), .A(n7063), .ZN(n8882) );
  NAND2_X1 U9308 ( .A1(n7064), .A2(n8868), .ZN(n7063) );
  NAND2_X1 U9309 ( .A1(n8869), .A2(n7065), .ZN(n7064) );
  NAND2_X1 U9310 ( .A1(n9192), .A2(n13597), .ZN(n7066) );
  NAND2_X1 U9311 ( .A1(n9165), .A2(n9166), .ZN(n9164) );
  OAI21_X1 U9312 ( .B1(n9226), .B2(n7072), .A(n7070), .ZN(n9241) );
  NAND2_X1 U9313 ( .A1(n7069), .A2(n7067), .ZN(n9240) );
  NAND2_X1 U9314 ( .A1(n9226), .A2(n7070), .ZN(n7069) );
  NAND2_X1 U9315 ( .A1(n9082), .A2(n7076), .ZN(n7075) );
  NAND2_X1 U9316 ( .A1(n8802), .A2(n7081), .ZN(n8807) );
  NAND2_X1 U9317 ( .A1(n9180), .A2(n7085), .ZN(n7082) );
  OAI21_X1 U9318 ( .B1(n9180), .B2(n7086), .A(n7085), .ZN(n9195) );
  NAND2_X1 U9319 ( .A1(n7082), .A2(n7083), .ZN(n9194) );
  NAND3_X1 U9320 ( .A1(n8906), .A2(n6571), .A3(n8905), .ZN(n7087) );
  OAI21_X1 U9321 ( .B1(n9006), .B2(n7092), .A(n7091), .ZN(n9021) );
  INV_X1 U9322 ( .A(n9260), .ZN(n9258) );
  AND3_X2 U9323 ( .A1(n7104), .A2(n7103), .A3(n6605), .ZN(n12610) );
  OR2_X2 U9324 ( .A1(n12559), .A2(n7105), .ZN(n7104) );
  INV_X1 U9325 ( .A(n7108), .ZN(n12606) );
  INV_X1 U9326 ( .A(n12607), .ZN(n7107) );
  NOR2_X1 U9327 ( .A1(n14730), .A2(n10624), .ZN(n14729) );
  INV_X1 U9328 ( .A(n10592), .ZN(n7111) );
  XNOR2_X1 U9329 ( .A(n10590), .B(n10625), .ZN(n14730) );
  NAND2_X1 U9330 ( .A1(n11628), .A2(n7116), .ZN(n7112) );
  INV_X1 U9331 ( .A(n10585), .ZN(n7121) );
  NAND2_X1 U9332 ( .A1(n7128), .A2(n7129), .ZN(n12015) );
  NAND2_X1 U9333 ( .A1(n13140), .A2(n7130), .ZN(n7128) );
  INV_X1 U9334 ( .A(n7134), .ZN(n13125) );
  NAND2_X1 U9335 ( .A1(n13236), .A2(n6554), .ZN(n7139) );
  OAI21_X1 U9336 ( .B1(n7140), .B2(n7142), .A(n7139), .ZN(n13189) );
  NAND2_X1 U9337 ( .A1(n7149), .A2(n10521), .ZN(n10847) );
  NAND4_X1 U9338 ( .A1(n7590), .A2(n7213), .A3(n7371), .A4(n7214), .ZN(n7151)
         );
  NAND2_X2 U9339 ( .A1(n8180), .A2(n8183), .ZN(n7434) );
  XNOR2_X2 U9340 ( .A(n7412), .B(n7411), .ZN(n8183) );
  XNOR2_X1 U9341 ( .A(n7409), .B(n7408), .ZN(n8180) );
  NAND2_X1 U9342 ( .A1(n8256), .A2(n7164), .ZN(n7163) );
  NAND2_X1 U9343 ( .A1(n8446), .A2(n7174), .ZN(n7173) );
  NAND2_X1 U9344 ( .A1(n8408), .A2(n7183), .ZN(n7181) );
  NAND2_X2 U9345 ( .A1(n11695), .A2(n7196), .ZN(n11999) );
  NAND2_X1 U9346 ( .A1(n9867), .A2(n13093), .ZN(n10022) );
  NAND2_X1 U9347 ( .A1(n10740), .A2(n7198), .ZN(n7197) );
  NAND2_X1 U9348 ( .A1(n7197), .A2(n6481), .ZN(n11155) );
  NAND2_X1 U9349 ( .A1(n12885), .A2(n6557), .ZN(n13026) );
  NAND3_X1 U9350 ( .A1(n11964), .A2(n10245), .A3(n10250), .ZN(n10492) );
  NAND2_X1 U9351 ( .A1(n10492), .A2(n10252), .ZN(n10266) );
  NAND2_X1 U9352 ( .A1(n7402), .A2(n7211), .ZN(n7427) );
  AND2_X1 U9353 ( .A1(n7402), .A2(n7398), .ZN(n7401) );
  NAND2_X1 U9354 ( .A1(n7402), .A2(n6566), .ZN(n8165) );
  NAND3_X1 U9355 ( .A1(n7212), .A2(n7339), .A3(n6461), .ZN(n7442) );
  INV_X1 U9356 ( .A(n8144), .ZN(n7212) );
  AND2_X2 U9357 ( .A1(n7449), .A2(n7369), .ZN(n7452) );
  NAND2_X1 U9358 ( .A1(n7587), .A2(n7224), .ZN(n7222) );
  NAND2_X1 U9359 ( .A1(n7587), .A2(n7586), .ZN(n7223) );
  NAND3_X1 U9360 ( .A1(n7839), .A2(n7838), .A3(n6574), .ZN(n7228) );
  INV_X1 U9361 ( .A(n7862), .ZN(n7229) );
  NAND3_X1 U9362 ( .A1(n7887), .A2(n7886), .A3(n6575), .ZN(n7231) );
  INV_X1 U9363 ( .A(n7903), .ZN(n7232) );
  NAND3_X1 U9364 ( .A1(n7696), .A2(n7695), .A3(n6567), .ZN(n7234) );
  INV_X1 U9365 ( .A(n7714), .ZN(n7235) );
  NAND3_X1 U9366 ( .A1(n7647), .A2(n7646), .A3(n6568), .ZN(n7237) );
  INV_X1 U9367 ( .A(n7667), .ZN(n7238) );
  NAND3_X1 U9368 ( .A1(n7927), .A2(n7926), .A3(n6569), .ZN(n7240) );
  INV_X1 U9369 ( .A(n7942), .ZN(n7241) );
  NAND3_X1 U9370 ( .A1(n7771), .A2(n7770), .A3(n7243), .ZN(n7242) );
  NAND2_X1 U9371 ( .A1(n7242), .A2(n6483), .ZN(n7820) );
  NAND2_X1 U9372 ( .A1(n7260), .A2(n6563), .ZN(n7595) );
  NAND3_X1 U9373 ( .A1(n7559), .A2(n6564), .A3(n7558), .ZN(n7260) );
  NAND4_X1 U9374 ( .A1(n13096), .A2(n7265), .A3(P3_ADDR_REG_19__SCAN_IN), .A4(
        n7264), .ZN(n7263) );
  NAND3_X1 U9375 ( .A1(n7267), .A2(n7266), .A3(n7268), .ZN(n9351) );
  NAND2_X1 U9376 ( .A1(n7270), .A2(n9299), .ZN(n7266) );
  NAND2_X1 U9377 ( .A1(n7269), .A2(n9762), .ZN(n7267) );
  INV_X1 U9378 ( .A(n9325), .ZN(n7268) );
  XNOR2_X1 U9379 ( .A(n9298), .B(n10556), .ZN(n7270) );
  NAND2_X1 U9380 ( .A1(n11230), .A2(n7278), .ZN(n14282) );
  NAND2_X1 U9381 ( .A1(n13855), .A2(n13859), .ZN(n13854) );
  XNOR2_X1 U9382 ( .A(n14335), .B(n10161), .ZN(n10148) );
  OAI21_X1 U9383 ( .B1(n7285), .B2(n10148), .A(n10223), .ZN(n7283) );
  NAND2_X1 U9384 ( .A1(n7286), .A2(n10151), .ZN(n10355) );
  NAND2_X1 U9385 ( .A1(n8790), .A2(n7289), .ZN(n7288) );
  NAND2_X1 U9386 ( .A1(n8790), .A2(n8789), .ZN(n9335) );
  NAND2_X1 U9387 ( .A1(n14170), .A2(n6472), .ZN(n7292) );
  OR2_X2 U9388 ( .A1(n14156), .A2(n14155), .ZN(n7361) );
  NAND2_X1 U9389 ( .A1(n8353), .A2(n9500), .ZN(n7307) );
  NAND2_X1 U9390 ( .A1(n8342), .A2(n10200), .ZN(n9979) );
  NAND2_X1 U9391 ( .A1(n11673), .A2(n7312), .ZN(n7310) );
  OAI21_X1 U9392 ( .B1(n12496), .B2(n7324), .A(n7322), .ZN(n7327) );
  NAND2_X1 U9393 ( .A1(n10396), .A2(n6556), .ZN(n10468) );
  NAND4_X1 U9394 ( .A1(n8222), .A2(n8221), .A3(n8220), .A4(n10322), .ZN(n8314)
         );
  INV_X1 U9395 ( .A(n7330), .ZN(n8409) );
  AND2_X1 U9396 ( .A1(n10831), .A2(n10832), .ZN(n7331) );
  NAND2_X1 U9397 ( .A1(n7332), .A2(n7331), .ZN(n10961) );
  NAND2_X1 U9398 ( .A1(n8716), .A2(n7333), .ZN(n8239) );
  AND2_X1 U9399 ( .A1(n8716), .A2(n8230), .ZN(n8718) );
  XNOR2_X1 U9400 ( .A(n8085), .B(n8084), .ZN(n13433) );
  NAND2_X1 U9401 ( .A1(n7486), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7470) );
  NAND2_X1 U9402 ( .A1(n7486), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7448) );
  NAND2_X1 U9403 ( .A1(n11131), .A2(n11130), .ZN(n11212) );
  NAND2_X1 U9404 ( .A1(n7486), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7436) );
  NAND2_X1 U9405 ( .A1(n14752), .A2(n12174), .ZN(n10444) );
  NAND2_X1 U9406 ( .A1(n7717), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7435) );
  INV_X1 U9407 ( .A(n9210), .ZN(n9213) );
  OAI21_X1 U9408 ( .B1(n9324), .B2(n9323), .A(n9561), .ZN(n9325) );
  NOR4_X1 U9409 ( .A1(n12299), .A2(n12135), .A3(n12285), .A4(n12134), .ZN(
        n12137) );
  OR2_X1 U9410 ( .A1(n12299), .A2(n12102), .ZN(n12103) );
  OAI22_X1 U9411 ( .A1(n13007), .A2(n12908), .B1(n12907), .B2(n12906), .ZN(
        n12909) );
  INV_X1 U9412 ( .A(n8358), .ZN(n10201) );
  XNOR2_X1 U9413 ( .A(n8148), .B(n10026), .ZN(n9891) );
  NAND2_X1 U9414 ( .A1(n8246), .A2(n12877), .ZN(n8345) );
  NAND2_X1 U9415 ( .A1(n9837), .A2(n9838), .ZN(n10178) );
  NAND2_X1 U9416 ( .A1(n9755), .A2(n9836), .ZN(n9835) );
  NAND2_X1 U9417 ( .A1(n11235), .A2(n11261), .ZN(n11266) );
  NAND2_X1 U9418 ( .A1(n11652), .A2(n11651), .ZN(n11843) );
  NAND2_X1 U9419 ( .A1(n12052), .A2(n14353), .ZN(n12055) );
  AND2_X1 U9420 ( .A1(n10179), .A2(n13540), .ZN(n10180) );
  INV_X2 U9421 ( .A(n6455), .ZN(n7497) );
  NAND2_X1 U9422 ( .A1(n8397), .A2(n8396), .ZN(n7335) );
  INV_X1 U9423 ( .A(n12652), .ZN(n9356) );
  AND2_X1 U9424 ( .A1(n7471), .A2(n7470), .ZN(n7336) );
  AND2_X1 U9425 ( .A1(n8836), .A2(n8835), .ZN(n7337) );
  NAND2_X1 U9426 ( .A1(n6462), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7338) );
  OR2_X1 U9427 ( .A1(n8148), .A2(n11003), .ZN(n7339) );
  OR2_X1 U9428 ( .A1(n12407), .A2(n12838), .ZN(n7340) );
  NOR2_X1 U9429 ( .A1(n8696), .A2(n11493), .ZN(n7341) );
  OR2_X1 U9430 ( .A1(n11249), .A2(n11248), .ZN(n7343) );
  OR2_X1 U9431 ( .A1(n12853), .A2(n12394), .ZN(n7345) );
  NOR2_X1 U9432 ( .A1(n10973), .A2(n10972), .ZN(n7346) );
  AND2_X1 U9433 ( .A1(n12909), .A2(n6501), .ZN(n7347) );
  NOR2_X1 U9434 ( .A1(n10024), .A2(n10023), .ZN(n7349) );
  OR2_X1 U9435 ( .A1(n11879), .A2(n13452), .ZN(n7350) );
  OR2_X1 U9436 ( .A1(n13930), .A2(n14371), .ZN(n7351) );
  AND4_X1 U9437 ( .A1(n8229), .A2(n8228), .A3(n8666), .A4(n8658), .ZN(n7353)
         );
  INV_X1 U9438 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n8908) );
  INV_X1 U9439 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n12458) );
  INV_X1 U9440 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10005) );
  INV_X1 U9441 ( .A(n13897), .ZN(n11847) );
  AND2_X1 U9442 ( .A1(n7964), .A2(n7963), .ZN(n7354) );
  INV_X1 U9443 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10559) );
  INV_X1 U9444 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7742) );
  INV_X1 U9445 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10557) );
  INV_X1 U9446 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10457) );
  INV_X1 U9447 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10053) );
  NAND2_X1 U9448 ( .A1(n12857), .A2(n12766), .ZN(n7355) );
  AND2_X2 U9449 ( .A1(n8763), .A2(n9994), .ZN(n14833) );
  INV_X1 U9450 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10390) );
  AND2_X1 U9451 ( .A1(n9297), .A2(n9296), .ZN(n7356) );
  NOR2_X1 U9452 ( .A1(n13921), .A2(n13920), .ZN(n7357) );
  NOR2_X1 U9453 ( .A1(n12831), .A2(n12415), .ZN(n8632) );
  INV_X1 U9454 ( .A(n12922), .ZN(n13048) );
  AND4_X1 U9455 ( .A1(n8034), .A2(n8033), .A3(n8032), .A4(n8031), .ZN(n12922)
         );
  INV_X1 U9456 ( .A(n12985), .ZN(n13051) );
  AND4_X1 U9457 ( .A1(n8013), .A2(n8012), .A3(n8011), .A4(n8010), .ZN(n12985)
         );
  INV_X1 U9458 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14650) );
  NAND4_X1 U9459 ( .A1(n8057), .A2(n8056), .A3(n8055), .A4(n8054), .ZN(n7358)
         );
  INV_X1 U9460 ( .A(n13927), .ZN(n11879) );
  INV_X1 U9461 ( .A(n13103), .ZN(n13098) );
  AND3_X1 U9462 ( .A1(n9350), .A2(n9349), .A3(n9348), .ZN(n7359) );
  XOR2_X1 U9463 ( .A(n9492), .B(P1_ADDR_REG_19__SCAN_IN), .Z(n7360) );
  INV_X4 U9464 ( .A(n9501), .ZN(n9505) );
  OR2_X1 U9465 ( .A1(n13295), .A2(n13058), .ZN(n7362) );
  NAND2_X2 U9466 ( .A1(n10192), .A2(n13245), .ZN(n13257) );
  AND2_X1 U9467 ( .A1(n14808), .A2(n14821), .ZN(n14828) );
  INV_X1 U9468 ( .A(n14767), .ZN(n12768) );
  INV_X1 U9469 ( .A(n12623), .ZN(n12105) );
  INV_X1 U9470 ( .A(n13387), .ZN(n11713) );
  INV_X1 U9471 ( .A(n12545), .ZN(n11672) );
  OR2_X1 U9472 ( .A1(n11759), .A2(n12247), .ZN(n7363) );
  INV_X1 U9473 ( .A(n12542), .ZN(n12394) );
  NAND2_X1 U9474 ( .A1(n8631), .A2(n8630), .ZN(n12537) );
  XOR2_X1 U9475 ( .A(n12100), .B(n12135), .Z(n7365) );
  INV_X1 U9476 ( .A(n7465), .ZN(n7466) );
  NAND2_X1 U9477 ( .A1(n8944), .A2(n8943), .ZN(n8958) );
  INV_X1 U9478 ( .A(n9211), .ZN(n9212) );
  INV_X1 U9479 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8227) );
  INV_X1 U9480 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8231) );
  INV_X1 U9481 ( .A(n7913), .ZN(n7914) );
  INV_X1 U9482 ( .A(n12241), .ZN(n8697) );
  OR2_X1 U9483 ( .A1(n12113), .A2(n12199), .ZN(n10911) );
  INV_X1 U9484 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8230) );
  OAI22_X1 U9485 ( .A1(n10080), .A2(n11941), .B1(n14322), .B2(n11942), .ZN(
        n9830) );
  NOR3_X1 U9486 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .A3(
        P1_IR_REG_26__SCAN_IN), .ZN(n8771) );
  INV_X1 U9487 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n8431) );
  OR2_X1 U9488 ( .A1(n12774), .A2(n12543), .ZN(n8537) );
  AND2_X1 U9489 ( .A1(n7968), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n7991) );
  XNOR2_X1 U9490 ( .A(n10021), .B(n9866), .ZN(n9867) );
  NOR2_X1 U9491 ( .A1(n7821), .A2(n14533), .ZN(n7840) );
  NOR2_X1 U9492 ( .A1(n7625), .A2(n14937), .ZN(n7648) );
  OR2_X1 U9493 ( .A1(n7796), .A2(n7795), .ZN(n7821) );
  INV_X1 U9494 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7535) );
  INV_X1 U9495 ( .A(n12038), .ZN(n12014) );
  AOI21_X1 U9496 ( .B1(n10975), .B2(n10974), .A(n7346), .ZN(n10977) );
  INV_X1 U9497 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7613) );
  NAND2_X1 U9498 ( .A1(n11913), .A2(n11914), .ZN(n11915) );
  INV_X1 U9499 ( .A(n9762), .ZN(n9299) );
  OR2_X1 U9500 ( .A1(n9911), .A2(n9757), .ZN(n9344) );
  NOR2_X1 U9501 ( .A1(n8800), .A2(n8799), .ZN(n8801) );
  NOR2_X1 U9502 ( .A1(n9417), .A2(n9416), .ZN(n9398) );
  INV_X1 U9503 ( .A(n12537), .ZN(n12415) );
  INV_X1 U9504 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n8290) );
  INV_X1 U9505 ( .A(n10401), .ZN(n10400) );
  OR2_X1 U9506 ( .A1(n8345), .A2(n14605), .ZN(n8336) );
  OR2_X1 U9507 ( .A1(n8624), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8639) );
  NOR2_X1 U9508 ( .A1(n8594), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8611) );
  NOR2_X1 U9509 ( .A1(n8639), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8653) );
  OAI21_X1 U9510 ( .B1(n12749), .B2(n12107), .A(n12108), .ZN(n12739) );
  INV_X1 U9511 ( .A(n10648), .ZN(n14661) );
  INV_X1 U9512 ( .A(n12163), .ZN(n10207) );
  NAND2_X2 U9513 ( .A1(n8342), .A2(n9982), .ZN(n12165) );
  NAND2_X1 U9514 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n10053), .ZN(n8210) );
  OR2_X1 U9515 ( .A1(n8438), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n8447) );
  INV_X1 U9516 ( .A(n7945), .ZN(n7946) );
  OR2_X1 U9517 ( .A1(n7719), .A2(n7718), .ZN(n7743) );
  OR2_X1 U9518 ( .A1(n7604), .A2(n7603), .ZN(n7625) );
  NOR2_X1 U9519 ( .A1(n7906), .A2(n13017), .ZN(n7928) );
  INV_X1 U9520 ( .A(n10504), .ZN(n10505) );
  INV_X1 U9521 ( .A(n13071), .ZN(n10262) );
  INV_X1 U9522 ( .A(n10011), .ZN(n10012) );
  OAI211_X1 U9523 ( .C1(n7434), .C2(n9653), .A(n7461), .B(n7460), .ZN(n8145)
         );
  AND2_X1 U9524 ( .A1(n14548), .A2(n9857), .ZN(n10006) );
  NAND2_X1 U9525 ( .A1(n10182), .A2(n10183), .ZN(n10184) );
  AOI21_X1 U9526 ( .B1(n12364), .B2(n13597), .A(n10180), .ZN(n10182) );
  NAND2_X1 U9527 ( .A1(n13427), .A2(n9262), .ZN(n9264) );
  OR2_X1 U9528 ( .A1(n12046), .A2(n14349), .ZN(n12047) );
  AND2_X1 U9529 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8887) );
  NAND2_X1 U9530 ( .A1(n7706), .A2(n9574), .ZN(n7727) );
  INV_X1 U9531 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n9400) );
  OAI21_X1 U9532 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n9466), .A(n9465), .ZN(
        n9471) );
  NOR2_X1 U9533 ( .A1(n8278), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8291) );
  OR3_X1 U9534 ( .A1(n8466), .A2(P3_REG3_REG_14__SCAN_IN), .A3(
        P3_REG3_REG_13__SCAN_IN), .ZN(n8482) );
  OR2_X1 U9535 ( .A1(n8401), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8415) );
  AND2_X1 U9536 ( .A1(n8291), .A2(n8290), .ZN(n8306) );
  INV_X1 U9537 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10472) );
  NAND2_X1 U9538 ( .A1(n8306), .A2(n10836), .ZN(n8401) );
  INV_X1 U9539 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n14920) );
  OR2_X1 U9540 ( .A1(n8571), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8583) );
  OR2_X1 U9541 ( .A1(n8531), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8546) );
  INV_X1 U9542 ( .A(n10474), .ZN(n12503) );
  OR2_X1 U9543 ( .A1(n12637), .A2(n8654), .ZN(n12448) );
  AND4_X1 U9544 ( .A1(n8488), .A2(n8487), .A3(n8486), .A4(n8485), .ZN(n12247)
         );
  INV_X1 U9545 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n14923) );
  INV_X1 U9546 ( .A(n14033), .ZN(n11198) );
  AND2_X1 U9547 ( .A1(n8653), .A2(n12449), .ZN(n12637) );
  INV_X1 U9548 ( .A(n12695), .ZN(n12701) );
  NAND2_X1 U9549 ( .A1(n8741), .A2(n9566), .ZN(n10127) );
  INV_X1 U9550 ( .A(SI_22_), .ZN(n8235) );
  INV_X1 U9551 ( .A(n14828), .ZN(n14106) );
  AND2_X1 U9552 ( .A1(n8758), .A2(n12307), .ZN(n14767) );
  OR2_X1 U9553 ( .A1(n8760), .A2(n8759), .ZN(n9998) );
  NAND2_X1 U9554 ( .A1(n8524), .A2(n8522), .ZN(n8214) );
  INV_X1 U9555 ( .A(n10345), .ZN(n10250) );
  OR2_X1 U9556 ( .A1(n14551), .A2(n10191), .ZN(n10016) );
  INV_X1 U9557 ( .A(n12999), .ZN(n13040) );
  NAND2_X1 U9558 ( .A1(n7717), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7447) );
  INV_X1 U9559 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n14533) );
  INV_X1 U9560 ( .A(n13224), .ZN(n13239) );
  INV_X1 U9561 ( .A(n12997), .ZN(n13037) );
  INV_X1 U9562 ( .A(n13068), .ZN(n10742) );
  INV_X1 U9563 ( .A(n13379), .ZN(n13289) );
  AND2_X1 U9564 ( .A1(n9870), .A2(n10995), .ZN(n10195) );
  INV_X1 U9565 ( .A(n12027), .ZN(n13278) );
  NAND2_X1 U9566 ( .A1(n10023), .A2(n10195), .ZN(n10011) );
  NAND2_X1 U9567 ( .A1(n8171), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8172) );
  INV_X1 U9568 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9034) );
  INV_X1 U9569 ( .A(n13778), .ZN(n13493) );
  NAND2_X1 U9570 ( .A1(n9009), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9041) );
  INV_X1 U9571 ( .A(n14141), .ZN(n13513) );
  INV_X1 U9572 ( .A(n13765), .ZN(n13560) );
  NOR2_X1 U9573 ( .A1(n9056), .A2(n14977), .ZN(n9070) );
  AND2_X1 U9574 ( .A1(n9246), .A2(n9230), .ZN(n13449) );
  NAND2_X1 U9575 ( .A1(n9097), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9113) );
  INV_X1 U9576 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n13600) );
  INV_X1 U9577 ( .A(n9614), .ZN(n9600) );
  NAND2_X1 U9578 ( .A1(n11855), .A2(n11854), .ZN(n13810) );
  NOR2_X1 U9579 ( .A1(n8962), .A2(n8961), .ZN(n8996) );
  INV_X1 U9580 ( .A(n13591), .ZN(n11246) );
  OR2_X1 U9581 ( .A1(n14318), .A2(n10037), .ZN(n13883) );
  NAND2_X1 U9582 ( .A1(n8812), .A2(n14017), .ZN(n9911) );
  NAND2_X1 U9583 ( .A1(n10166), .A2(n10165), .ZN(n10352) );
  NOR2_X1 U9584 ( .A1(n9744), .A2(n9546), .ZN(n10034) );
  INV_X1 U9585 ( .A(n14015), .ZN(n9547) );
  AND2_X1 U9586 ( .A1(n7828), .A2(n7807), .ZN(n7826) );
  AND2_X1 U9587 ( .A1(n7727), .A2(n7708), .ZN(n7725) );
  CLKBUF_X1 U9588 ( .A(n7569), .Z(n7548) );
  NOR2_X1 U9589 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9433), .ZN(n9392) );
  AOI22_X1 U9590 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n9408), .B1(n9410), .B2(
        n9407), .ZN(n9464) );
  INV_X1 U9591 ( .A(n12763), .ZN(n14762) );
  AND3_X1 U9592 ( .A1(n8587), .A2(n8586), .A3(n8585), .ZN(n12487) );
  INV_X1 U9593 ( .A(n10319), .ZN(n10308) );
  INV_X1 U9594 ( .A(n14709), .ZN(n14735) );
  INV_X1 U9595 ( .A(n14740), .ZN(n14718) );
  AND3_X1 U9596 ( .A1(n10307), .A2(n10317), .A3(n12288), .ZN(n12763) );
  AND2_X1 U9597 ( .A1(n12236), .A2(n12235), .ZN(n12232) );
  NOR2_X1 U9598 ( .A1(n14846), .A2(n8677), .ZN(n9379) );
  AND3_X1 U9599 ( .A1(n8746), .A2(n8756), .A3(n8760), .ZN(n10130) );
  OR2_X1 U9600 ( .A1(n14833), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9494) );
  INV_X1 U9601 ( .A(n14827), .ZN(n14812) );
  INV_X1 U9602 ( .A(n12308), .ZN(n9994) );
  INV_X1 U9603 ( .A(n8742), .ZN(n9562) );
  AND2_X1 U9604 ( .A1(n9504), .A2(P3_U3151), .ZN(n14038) );
  AND2_X1 U9605 ( .A1(n14592), .A2(n10018), .ZN(n10019) );
  AND3_X1 U9606 ( .A1(n7801), .A2(n7800), .A3(n7799), .ZN(n12004) );
  AND2_X1 U9607 ( .A1(n9664), .A2(n9638), .ZN(n14526) );
  NAND2_X1 U9608 ( .A1(n9637), .A2(n9636), .ZN(n9664) );
  INV_X1 U9609 ( .A(n13294), .ZN(n13241) );
  NAND2_X1 U9610 ( .A1(n10023), .A2(n10013), .ZN(n14592) );
  AND2_X1 U9611 ( .A1(n13341), .A2(n9868), .ZN(n14571) );
  INV_X1 U9612 ( .A(n14571), .ZN(n14589) );
  AND2_X1 U9613 ( .A1(n9846), .A2(n9862), .ZN(n14548) );
  INV_X1 U9614 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7729) );
  OR2_X1 U9615 ( .A1(n9763), .A2(n9561), .ZN(n9577) );
  AND2_X1 U9616 ( .A1(n14141), .A2(n14131), .ZN(n13557) );
  NAND2_X1 U9617 ( .A1(n9767), .A2(n14302), .ZN(n14142) );
  AND2_X1 U9618 ( .A1(n9136), .A2(n9135), .ZN(n13476) );
  INV_X1 U9619 ( .A(n14270), .ZN(n13725) );
  NOR2_X1 U9620 ( .A1(n9600), .A2(n9760), .ZN(n13723) );
  NAND2_X1 U9621 ( .A1(n12055), .A2(n12054), .ZN(n12056) );
  INV_X1 U9622 ( .A(n13887), .ZN(n14315) );
  INV_X1 U9623 ( .A(n9916), .ZN(n10032) );
  INV_X1 U9624 ( .A(n14353), .ZN(n14357) );
  NAND2_X1 U9625 ( .A1(n9910), .A2(n9909), .ZN(n14353) );
  INV_X1 U9626 ( .A(n14349), .ZN(n14375) );
  AND3_X1 U9627 ( .A1(n9545), .A2(n9544), .A3(n9547), .ZN(n9740) );
  AND2_X1 U9628 ( .A1(n10316), .A2(n10315), .ZN(n14743) );
  AND2_X1 U9629 ( .A1(n9973), .A2(n9972), .ZN(n12450) );
  INV_X1 U9630 ( .A(n12528), .ZN(n12518) );
  AND2_X1 U9631 ( .A1(n12090), .A2(n8679), .ZN(n12451) );
  INV_X1 U9632 ( .A(n12487), .ZN(n12539) );
  INV_X1 U9633 ( .A(n14743), .ZN(n14727) );
  INV_X1 U9634 ( .A(n14080), .ZN(n14750) );
  AND2_X1 U9635 ( .A1(n10925), .A2(n10924), .ZN(n14800) );
  INV_X2 U9636 ( .A(n14770), .ZN(n14772) );
  NAND2_X1 U9637 ( .A1(n14846), .A2(n14812), .ZN(n12826) );
  INV_X1 U9638 ( .A(n14846), .ZN(n14844) );
  INV_X1 U9639 ( .A(n12491), .ZN(n12838) );
  INV_X1 U9640 ( .A(n12254), .ZN(n11822) );
  INV_X1 U9641 ( .A(n14833), .ZN(n14832) );
  AND2_X1 U9642 ( .A1(n10305), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9567) );
  INV_X1 U9643 ( .A(SI_13_), .ZN(n9574) );
  INV_X1 U9644 ( .A(n14497), .ZN(n14540) );
  NAND2_X1 U9645 ( .A1(n10261), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13015) );
  NAND2_X1 U9646 ( .A1(n10020), .A2(n10019), .ZN(n13023) );
  INV_X1 U9647 ( .A(n12953), .ZN(n13047) );
  OR2_X1 U9648 ( .A1(n14392), .A2(P2_U3088), .ZN(n14547) );
  INV_X1 U9649 ( .A(n13302), .ZN(n13170) );
  NAND2_X1 U9650 ( .A1(n13257), .A2(n10561), .ZN(n13299) );
  OR3_X1 U9651 ( .A1(n9921), .A2(n14551), .A3(n9920), .ZN(n14603) );
  NOR2_X1 U9652 ( .A1(n14553), .A2(n14548), .ZN(n14549) );
  INV_X1 U9653 ( .A(n14549), .ZN(n14550) );
  INV_X1 U9654 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n14948) );
  INV_X1 U9655 ( .A(n13874), .ZN(n13977) );
  INV_X1 U9656 ( .A(n14154), .ZN(n14190) );
  NAND2_X1 U9657 ( .A1(n10171), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14146) );
  INV_X1 U9658 ( .A(n14142), .ZN(n13579) );
  INV_X1 U9659 ( .A(n13476), .ZN(n13876) );
  INV_X1 U9660 ( .A(n13726), .ZN(n14272) );
  INV_X1 U9661 ( .A(n13723), .ZN(n14274) );
  INV_X1 U9662 ( .A(n14303), .ZN(n13880) );
  INV_X1 U9663 ( .A(n14303), .ZN(n14284) );
  INV_X1 U9664 ( .A(n14303), .ZN(n14318) );
  NAND2_X1 U9665 ( .A1(n9917), .A2(n10032), .ZN(n14388) );
  NAND2_X1 U9666 ( .A1(n9917), .A2(n9916), .ZN(n14376) );
  INV_X1 U9667 ( .A(n9546), .ZN(n9549) );
  INV_X1 U9668 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14011) );
  INV_X1 U9669 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n14852) );
  INV_X1 U9670 ( .A(n11589), .ZN(n13702) );
  AND2_X2 U9671 ( .A1(n9567), .A2(n9496), .ZN(P3_U3897) );
  NOR2_X1 U9672 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7375) );
  NAND4_X1 U9673 ( .A1(n7375), .A2(n7374), .A3(n7373), .A4(n7372), .ZN(n7791)
         );
  INV_X1 U9674 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n7376) );
  NAND4_X1 U9675 ( .A1(n7377), .A2(n7404), .A3(n7210), .A4(n7376), .ZN(n7380)
         );
  INV_X1 U9676 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7378) );
  NAND4_X1 U9677 ( .A1(n7428), .A2(n7398), .A3(n7378), .A4(n7396), .ZN(n7379)
         );
  NAND2_X1 U9678 ( .A1(n6572), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7385) );
  NAND2_X1 U9679 ( .A1(n7484), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7391) );
  INV_X1 U9680 ( .A(n12042), .ZN(n7387) );
  NAND2_X1 U9681 ( .A1(n7486), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7390) );
  NAND2_X1 U9682 ( .A1(n7717), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7388) );
  NAND4_X2 U9683 ( .A1(n7391), .A2(n7390), .A3(n7389), .A4(n7388), .ZN(n8148)
         );
  NAND2_X1 U9684 ( .A1(n7393), .A2(n7392), .ZN(n7394) );
  NOR2_X1 U9685 ( .A1(n7791), .A2(n7394), .ZN(n7395) );
  NAND2_X1 U9686 ( .A1(n7395), .A2(n7590), .ZN(n7808) );
  INV_X1 U9687 ( .A(n7808), .ZN(n7397) );
  NAND2_X1 U9688 ( .A1(n7397), .A2(n7396), .ZN(n7810) );
  NOR2_X2 U9689 ( .A1(n7810), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n7402) );
  NAND2_X1 U9690 ( .A1(n7427), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7399) );
  NAND2_X1 U9691 ( .A1(n7404), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n7406) );
  NAND2_X1 U9692 ( .A1(n14924), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n7405) );
  AND2_X1 U9693 ( .A1(n7406), .A2(n7405), .ZN(n7407) );
  INV_X1 U9694 ( .A(n13341), .ZN(n14580) );
  NAND2_X1 U9695 ( .A1(n7416), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7414) );
  INV_X1 U9696 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7413) );
  INV_X1 U9697 ( .A(SI_1_), .ZN(n9502) );
  XNOR2_X2 U9698 ( .A(n7457), .B(n9502), .ZN(n7456) );
  AND2_X1 U9699 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7415) );
  NAND2_X1 U9700 ( .A1(n9501), .A2(n7415), .ZN(n7433) );
  INV_X1 U9701 ( .A(n7416), .ZN(n7417) );
  AND2_X1 U9702 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7418) );
  NAND2_X1 U9703 ( .A1(n7459), .A2(n7418), .ZN(n8840) );
  OR2_X1 U9704 ( .A1(n7760), .A2(n7413), .ZN(n7421) );
  NAND2_X1 U9705 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n14978) );
  INV_X1 U9706 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7419) );
  NAND3_X2 U9707 ( .A1(n7422), .A2(n7421), .A3(n7420), .ZN(n10026) );
  OAI21_X1 U9708 ( .B1(n8148), .B2(n6461), .A(n10026), .ZN(n7425) );
  NAND2_X1 U9709 ( .A1(n8148), .A2(n8123), .ZN(n7423) );
  INV_X1 U9710 ( .A(n10026), .ZN(n11003) );
  NAND2_X1 U9711 ( .A1(n7423), .A2(n11003), .ZN(n7424) );
  NAND2_X1 U9712 ( .A1(n7425), .A2(n7424), .ZN(n7444) );
  NAND2_X1 U9713 ( .A1(n8148), .A2(n11003), .ZN(n7441) );
  NAND2_X1 U9714 ( .A1(n14924), .A2(n7428), .ZN(n7429) );
  NAND3_X2 U9715 ( .A1(n7430), .A2(n7427), .A3(n7429), .ZN(n10995) );
  INV_X1 U9716 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n14397) );
  INV_X1 U9717 ( .A(SI_0_), .ZN(n7431) );
  INV_X1 U9718 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8188) );
  OAI21_X1 U9719 ( .B1(n9504), .B2(n7431), .A(n8188), .ZN(n7432) );
  NAND2_X1 U9720 ( .A1(n7433), .A2(n7432), .ZN(n13445) );
  NAND2_X1 U9721 ( .A1(n7484), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7438) );
  NAND2_X1 U9722 ( .A1(n7485), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7437) );
  NAND4_X1 U9723 ( .A1(n7438), .A2(n7437), .A3(n7436), .A4(n7435), .ZN(n9869)
         );
  OAI21_X1 U9724 ( .B1(n10021), .B2(n10025), .A(n9869), .ZN(n7440) );
  AOI21_X1 U9725 ( .B1(n10021), .B2(n10025), .A(n6461), .ZN(n7439) );
  NAND3_X1 U9726 ( .A1(n7441), .A2(n7440), .A3(n7439), .ZN(n7443) );
  NAND2_X1 U9727 ( .A1(n7485), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7446) );
  NAND2_X1 U9728 ( .A1(n7484), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7445) );
  NOR2_X1 U9729 ( .A1(n7449), .A2(n14924), .ZN(n7450) );
  MUX2_X1 U9730 ( .A(n14924), .B(n7450), .S(P2_IR_REG_2__SCAN_IN), .Z(n7451)
         );
  INV_X1 U9731 ( .A(n7451), .ZN(n7454) );
  INV_X1 U9732 ( .A(n7452), .ZN(n7453) );
  NAND2_X1 U9733 ( .A1(n7454), .A2(n7453), .ZN(n9653) );
  NAND2_X1 U9734 ( .A1(n7457), .A2(SI_1_), .ZN(n7458) );
  INV_X1 U9735 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9530) );
  INV_X1 U9736 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9521) );
  MUX2_X1 U9737 ( .A(n9530), .B(n9521), .S(n7459), .Z(n7474) );
  OR2_X1 U9738 ( .A1(n6455), .A2(n9530), .ZN(n7460) );
  MUX2_X1 U9739 ( .A(n8146), .B(n8145), .S(n8107), .Z(n7465) );
  MUX2_X1 U9740 ( .A(n8146), .B(n8145), .S(n6460), .Z(n7462) );
  NAND2_X1 U9741 ( .A1(n7463), .A2(n7462), .ZN(n7469) );
  INV_X1 U9742 ( .A(n7464), .ZN(n7467) );
  NAND2_X1 U9743 ( .A1(n7467), .A2(n7466), .ZN(n7468) );
  NAND2_X1 U9744 ( .A1(n7485), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7471) );
  NAND2_X1 U9745 ( .A1(n7484), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7472) );
  NAND3_X1 U9746 ( .A1(n7336), .A2(n7473), .A3(n7472), .ZN(n8149) );
  NAND2_X1 U9747 ( .A1(n7475), .A2(SI_2_), .ZN(n7476) );
  XNOR2_X1 U9748 ( .A(n7494), .B(SI_3_), .ZN(n7491) );
  XNOR2_X1 U9749 ( .A(n7493), .B(n7491), .ZN(n9527) );
  NAND2_X1 U9750 ( .A1(n9527), .A2(n7960), .ZN(n7481) );
  NOR2_X1 U9751 ( .A1(n7452), .A2(n14924), .ZN(n7477) );
  MUX2_X1 U9752 ( .A(n14924), .B(n7477), .S(P2_IR_REG_3__SCAN_IN), .Z(n7479)
         );
  AND2_X1 U9753 ( .A1(n7452), .A2(n7478), .ZN(n7498) );
  NOR2_X1 U9754 ( .A1(n7479), .A2(n7498), .ZN(n9656) );
  AOI22_X1 U9755 ( .A1(n7497), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n7859), .B2(
        n9656), .ZN(n7480) );
  MUX2_X1 U9756 ( .A(n8149), .B(n10772), .S(n6460), .Z(n7483) );
  MUX2_X1 U9757 ( .A(n8149), .B(n10772), .S(n8107), .Z(n7482) );
  NAND2_X1 U9758 ( .A1(n7798), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7490) );
  AND2_X1 U9759 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7509) );
  INV_X1 U9760 ( .A(n7509), .ZN(n7511) );
  OAI21_X1 U9761 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n7511), .ZN(n10575) );
  OR2_X1 U9762 ( .A1(n7508), .A2(n10575), .ZN(n7489) );
  NAND2_X1 U9763 ( .A1(n8096), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7488) );
  NAND2_X1 U9764 ( .A1(n7486), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7487) );
  NAND2_X1 U9765 ( .A1(n7494), .A2(SI_3_), .ZN(n7495) );
  MUX2_X1 U9766 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n9505), .Z(n7520) );
  XNOR2_X1 U9767 ( .A(n7520), .B(SI_4_), .ZN(n7517) );
  XNOR2_X1 U9768 ( .A(n7496), .B(n7517), .ZN(n9533) );
  NAND2_X1 U9769 ( .A1(n9533), .A2(n7960), .ZN(n7501) );
  INV_X1 U9770 ( .A(n7498), .ZN(n7523) );
  NAND2_X1 U9771 ( .A1(n7523), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7499) );
  XNOR2_X1 U9772 ( .A(n7499), .B(P2_IR_REG_4__SCAN_IN), .ZN(n9659) );
  AOI22_X1 U9773 ( .A1(n7497), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7859), .B2(
        n9659), .ZN(n7500) );
  MUX2_X1 U9774 ( .A(n13071), .B(n14566), .S(n8107), .Z(n7504) );
  NAND2_X1 U9775 ( .A1(n7505), .A2(n7504), .ZN(n7503) );
  MUX2_X1 U9776 ( .A(n14566), .B(n13071), .S(n8107), .Z(n7502) );
  NAND2_X1 U9777 ( .A1(n7503), .A2(n7502), .ZN(n7507) );
  NAND2_X1 U9778 ( .A1(n7486), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7516) );
  NAND2_X1 U9779 ( .A1(n7509), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7536) );
  INV_X1 U9780 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7510) );
  NAND2_X1 U9781 ( .A1(n7511), .A2(n7510), .ZN(n7512) );
  NAND2_X1 U9782 ( .A1(n7536), .A2(n7512), .ZN(n10684) );
  OR2_X1 U9783 ( .A1(n7508), .A2(n10684), .ZN(n7515) );
  NAND2_X1 U9784 ( .A1(n7798), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7514) );
  NAND2_X1 U9785 ( .A1(n8096), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7513) );
  INV_X1 U9786 ( .A(n7517), .ZN(n7518) );
  NAND2_X1 U9787 ( .A1(n7520), .A2(SI_4_), .ZN(n7521) );
  NAND2_X1 U9788 ( .A1(n7522), .A2(n7521), .ZN(n7544) );
  MUX2_X1 U9789 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n9505), .Z(n7545) );
  XNOR2_X1 U9790 ( .A(n7545), .B(SI_5_), .ZN(n7542) );
  XNOR2_X1 U9791 ( .A(n7544), .B(n7542), .ZN(n9539) );
  NAND2_X1 U9792 ( .A1(n9539), .A2(n7960), .ZN(n7530) );
  NAND2_X1 U9793 ( .A1(n7526), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7525) );
  MUX2_X1 U9794 ( .A(n7525), .B(P2_IR_REG_31__SCAN_IN), .S(n7524), .Z(n7528)
         );
  INV_X1 U9795 ( .A(n7526), .ZN(n7527) );
  NAND2_X1 U9796 ( .A1(n7527), .A2(n7524), .ZN(n7573) );
  NAND2_X1 U9797 ( .A1(n7528), .A2(n7573), .ZN(n9672) );
  INV_X1 U9798 ( .A(n9672), .ZN(n9679) );
  AOI22_X1 U9799 ( .A1(n7497), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7859), .B2(
        n9679), .ZN(n7529) );
  NAND2_X1 U9800 ( .A1(n7530), .A2(n7529), .ZN(n10507) );
  MUX2_X1 U9801 ( .A(n13070), .B(n10507), .S(n6461), .Z(n7532) );
  MUX2_X1 U9802 ( .A(n13070), .B(n10507), .S(n8107), .Z(n7531) );
  INV_X1 U9803 ( .A(n7532), .ZN(n7533) );
  NAND2_X1 U9804 ( .A1(n7798), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7541) );
  NOR2_X1 U9805 ( .A1(n7536), .A2(n7535), .ZN(n7560) );
  INV_X1 U9806 ( .A(n7560), .ZN(n7562) );
  NAND2_X1 U9807 ( .A1(n7536), .A2(n7535), .ZN(n7537) );
  NAND2_X1 U9808 ( .A1(n7562), .A2(n7537), .ZN(n10690) );
  OR2_X1 U9809 ( .A1(n7508), .A2(n10690), .ZN(n7540) );
  NAND2_X1 U9810 ( .A1(n7580), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7539) );
  NAND2_X1 U9811 ( .A1(n8096), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7538) );
  INV_X1 U9812 ( .A(n7542), .ZN(n7543) );
  NAND2_X1 U9813 ( .A1(n7545), .A2(SI_5_), .ZN(n7546) );
  MUX2_X1 U9814 ( .A(n9554), .B(n14864), .S(n9505), .Z(n7570) );
  XNOR2_X1 U9815 ( .A(n7570), .B(SI_6_), .ZN(n7568) );
  INV_X1 U9816 ( .A(n7568), .ZN(n7547) );
  XNOR2_X1 U9817 ( .A(n7548), .B(n7547), .ZN(n9552) );
  NAND2_X1 U9818 ( .A1(n9552), .A2(n7960), .ZN(n7551) );
  NAND2_X1 U9819 ( .A1(n7573), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7549) );
  XNOR2_X1 U9820 ( .A(n7549), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9947) );
  AOI22_X1 U9821 ( .A1(n7497), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7859), .B2(
        n9947), .ZN(n7550) );
  NAND2_X1 U9822 ( .A1(n7551), .A2(n7550), .ZN(n10694) );
  MUX2_X1 U9823 ( .A(n13069), .B(n10694), .S(n6467), .Z(n7555) );
  NAND2_X1 U9824 ( .A1(n7554), .A2(n7555), .ZN(n7553) );
  MUX2_X1 U9825 ( .A(n13069), .B(n10694), .S(n6461), .Z(n7552) );
  NAND2_X1 U9826 ( .A1(n7553), .A2(n7552), .ZN(n7559) );
  INV_X1 U9827 ( .A(n7554), .ZN(n7557) );
  INV_X1 U9828 ( .A(n7555), .ZN(n7556) );
  NAND2_X1 U9829 ( .A1(n7557), .A2(n7556), .ZN(n7558) );
  NAND2_X1 U9830 ( .A1(n7580), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7567) );
  NAND2_X1 U9831 ( .A1(n7560), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7604) );
  INV_X1 U9832 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7561) );
  NAND2_X1 U9833 ( .A1(n7562), .A2(n7561), .ZN(n7563) );
  NAND2_X1 U9834 ( .A1(n7604), .A2(n7563), .ZN(n10951) );
  OR2_X1 U9835 ( .A1(n8077), .A2(n10951), .ZN(n7566) );
  NAND2_X1 U9836 ( .A1(n7798), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7565) );
  NAND2_X1 U9837 ( .A1(n8096), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7564) );
  NAND4_X1 U9838 ( .A1(n7567), .A2(n7566), .A3(n7565), .A4(n7564), .ZN(n13068)
         );
  INV_X1 U9839 ( .A(n7570), .ZN(n7571) );
  NAND2_X1 U9840 ( .A1(n7571), .A2(SI_6_), .ZN(n7572) );
  MUX2_X1 U9841 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n9505), .Z(n7588) );
  XNOR2_X1 U9842 ( .A(n7588), .B(SI_7_), .ZN(n7585) );
  XNOR2_X1 U9843 ( .A(n7587), .B(n7585), .ZN(n9555) );
  NAND2_X1 U9844 ( .A1(n9555), .A2(n7960), .ZN(n7576) );
  OAI21_X1 U9845 ( .B1(n7573), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7574) );
  XNOR2_X1 U9846 ( .A(n7574), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9951) );
  AOI22_X1 U9847 ( .A1(n7497), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7859), .B2(
        n9951), .ZN(n7575) );
  NAND2_X1 U9848 ( .A1(n7576), .A2(n7575), .ZN(n10953) );
  MUX2_X1 U9849 ( .A(n13068), .B(n10953), .S(n6460), .Z(n7578) );
  MUX2_X1 U9850 ( .A(n13068), .B(n10953), .S(n6467), .Z(n7577) );
  INV_X1 U9851 ( .A(n7578), .ZN(n7579) );
  NAND2_X1 U9852 ( .A1(n7798), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7584) );
  INV_X1 U9853 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7602) );
  XNOR2_X1 U9854 ( .A(n7604), .B(n7602), .ZN(n10888) );
  OR2_X1 U9855 ( .A1(n8077), .A2(n10888), .ZN(n7583) );
  NAND2_X1 U9856 ( .A1(n8096), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7582) );
  NAND2_X1 U9857 ( .A1(n7580), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7581) );
  NAND4_X1 U9858 ( .A1(n7584), .A2(n7583), .A3(n7582), .A4(n7581), .ZN(n13067)
         );
  INV_X1 U9859 ( .A(n7585), .ZN(n7586) );
  NAND2_X1 U9860 ( .A1(n7588), .A2(SI_7_), .ZN(n7589) );
  MUX2_X1 U9861 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n9505), .Z(n7612) );
  XNOR2_X1 U9862 ( .A(n7612), .B(SI_8_), .ZN(n7610) );
  OR2_X1 U9863 ( .A1(n7590), .A2(n14924), .ZN(n7591) );
  XNOR2_X1 U9864 ( .A(n7591), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9954) );
  AOI22_X1 U9865 ( .A1(n7497), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7859), .B2(
        n9954), .ZN(n7592) );
  MUX2_X1 U9866 ( .A(n13067), .B(n10890), .S(n6467), .Z(n7596) );
  NAND2_X1 U9867 ( .A1(n7595), .A2(n7596), .ZN(n7594) );
  MUX2_X1 U9868 ( .A(n13067), .B(n10890), .S(n6460), .Z(n7593) );
  NAND2_X1 U9869 ( .A1(n7594), .A2(n7593), .ZN(n7600) );
  INV_X1 U9870 ( .A(n7595), .ZN(n7598) );
  INV_X1 U9871 ( .A(n7596), .ZN(n7597) );
  NAND2_X1 U9872 ( .A1(n7598), .A2(n7597), .ZN(n7599) );
  NAND2_X1 U9873 ( .A1(n7600), .A2(n7599), .ZN(n7619) );
  NAND2_X1 U9874 ( .A1(n7580), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7609) );
  INV_X1 U9875 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7601) );
  OAI21_X1 U9876 ( .B1(n7604), .B2(n7602), .A(n7601), .ZN(n7605) );
  NAND2_X1 U9877 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .ZN(n7603) );
  NAND2_X1 U9878 ( .A1(n7605), .A2(n7625), .ZN(n11091) );
  OR2_X1 U9879 ( .A1(n8077), .A2(n11091), .ZN(n7608) );
  NAND2_X1 U9880 ( .A1(n7798), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7607) );
  NAND2_X1 U9881 ( .A1(n8096), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7606) );
  NAND4_X1 U9882 ( .A1(n7609), .A2(n7608), .A3(n7607), .A4(n7606), .ZN(n13066)
         );
  INV_X1 U9883 ( .A(n7610), .ZN(n7611) );
  MUX2_X1 U9884 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n9505), .Z(n7634) );
  XNOR2_X1 U9885 ( .A(n7634), .B(SI_9_), .ZN(n7631) );
  XNOR2_X1 U9886 ( .A(n7633), .B(n7631), .ZN(n9583) );
  NAND2_X1 U9887 ( .A1(n9583), .A2(n7960), .ZN(n7616) );
  NAND2_X1 U9888 ( .A1(n7590), .A2(n7613), .ZN(n7636) );
  NAND2_X1 U9889 ( .A1(n7636), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7614) );
  XNOR2_X1 U9890 ( .A(n7614), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10424) );
  AOI22_X1 U9891 ( .A1(n7497), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7859), .B2(
        n10424), .ZN(n7615) );
  MUX2_X1 U9892 ( .A(n13066), .B(n11090), .S(n6461), .Z(n7620) );
  NAND2_X1 U9893 ( .A1(n7619), .A2(n7620), .ZN(n7618) );
  MUX2_X1 U9894 ( .A(n13066), .B(n11090), .S(n6467), .Z(n7617) );
  NAND2_X1 U9895 ( .A1(n7618), .A2(n7617), .ZN(n7624) );
  INV_X1 U9896 ( .A(n7619), .ZN(n7622) );
  INV_X1 U9897 ( .A(n7620), .ZN(n7621) );
  NAND2_X1 U9898 ( .A1(n7622), .A2(n7621), .ZN(n7623) );
  NAND2_X1 U9899 ( .A1(n7798), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7630) );
  INV_X1 U9900 ( .A(n7648), .ZN(n7650) );
  NAND2_X1 U9901 ( .A1(n7625), .A2(n14937), .ZN(n7626) );
  NAND2_X1 U9902 ( .A1(n7650), .A2(n7626), .ZN(n11082) );
  OR2_X1 U9903 ( .A1(n8077), .A2(n11082), .ZN(n7629) );
  NAND2_X1 U9904 ( .A1(n7580), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7628) );
  NAND2_X1 U9905 ( .A1(n8096), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7627) );
  NAND4_X1 U9906 ( .A1(n7630), .A2(n7629), .A3(n7628), .A4(n7627), .ZN(n13065)
         );
  INV_X1 U9907 ( .A(n7631), .ZN(n7632) );
  NAND2_X1 U9908 ( .A1(n7634), .A2(SI_9_), .ZN(n7635) );
  MUX2_X1 U9909 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n9505), .Z(n7659) );
  XNOR2_X1 U9910 ( .A(n7659), .B(SI_10_), .ZN(n7656) );
  XNOR2_X1 U9911 ( .A(n7658), .B(n7656), .ZN(n9589) );
  NAND2_X1 U9912 ( .A1(n9589), .A2(n7960), .ZN(n7639) );
  NAND2_X1 U9913 ( .A1(n8174), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7637) );
  XNOR2_X1 U9914 ( .A(n7637), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10434) );
  AOI22_X1 U9915 ( .A1(n7497), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7859), .B2(
        n10434), .ZN(n7638) );
  MUX2_X1 U9916 ( .A(n13065), .B(n11146), .S(n6467), .Z(n7643) );
  NAND2_X1 U9917 ( .A1(n7642), .A2(n7643), .ZN(n7641) );
  MUX2_X1 U9918 ( .A(n13065), .B(n11146), .S(n6460), .Z(n7640) );
  NAND2_X1 U9919 ( .A1(n7641), .A2(n7640), .ZN(n7647) );
  INV_X1 U9920 ( .A(n7642), .ZN(n7645) );
  INV_X1 U9921 ( .A(n7643), .ZN(n7644) );
  NAND2_X1 U9922 ( .A1(n7645), .A2(n7644), .ZN(n7646) );
  NAND2_X1 U9923 ( .A1(n7798), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7655) );
  INV_X1 U9924 ( .A(n7670), .ZN(n7672) );
  INV_X1 U9925 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7649) );
  NAND2_X1 U9926 ( .A1(n7650), .A2(n7649), .ZN(n7651) );
  NAND2_X1 U9927 ( .A1(n7672), .A2(n7651), .ZN(n11179) );
  OR2_X1 U9928 ( .A1(n8077), .A2(n11179), .ZN(n7654) );
  NAND2_X1 U9929 ( .A1(n7580), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7653) );
  NAND2_X1 U9930 ( .A1(n8096), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7652) );
  NAND4_X1 U9931 ( .A1(n7655), .A2(n7654), .A3(n7653), .A4(n7652), .ZN(n13064)
         );
  INV_X1 U9932 ( .A(n7656), .ZN(n7657) );
  MUX2_X1 U9933 ( .A(n9627), .B(n9625), .S(n9505), .Z(n7660) );
  NAND2_X1 U9934 ( .A1(n7660), .A2(n9538), .ZN(n7678) );
  INV_X1 U9935 ( .A(n7660), .ZN(n7661) );
  NAND2_X1 U9936 ( .A1(n7661), .A2(SI_11_), .ZN(n7662) );
  NAND2_X1 U9937 ( .A1(n7678), .A2(n7662), .ZN(n7679) );
  XNOR2_X1 U9938 ( .A(n7680), .B(n7679), .ZN(n9624) );
  NAND2_X1 U9939 ( .A1(n9624), .A2(n7960), .ZN(n7666) );
  INV_X1 U9940 ( .A(n7685), .ZN(n7663) );
  NAND2_X1 U9941 ( .A1(n7663), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7664) );
  XNOR2_X1 U9942 ( .A(n7664), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10441) );
  AOI22_X1 U9943 ( .A1(n7497), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7859), .B2(
        n10441), .ZN(n7665) );
  MUX2_X1 U9944 ( .A(n13064), .B(n11174), .S(n6460), .Z(n7668) );
  MUX2_X1 U9945 ( .A(n13064), .B(n11174), .S(n6467), .Z(n7667) );
  INV_X1 U9946 ( .A(n7668), .ZN(n7669) );
  INV_X1 U9947 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11453) );
  OR2_X1 U9948 ( .A1(n8079), .A2(n11453), .ZN(n7677) );
  NAND2_X1 U9949 ( .A1(n7670), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7697) );
  INV_X1 U9950 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7671) );
  NAND2_X1 U9951 ( .A1(n7672), .A2(n7671), .ZN(n7673) );
  NAND2_X1 U9952 ( .A1(n7697), .A2(n7673), .ZN(n11281) );
  OR2_X1 U9953 ( .A1(n8077), .A2(n11281), .ZN(n7676) );
  NAND2_X1 U9954 ( .A1(n7798), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7675) );
  NAND2_X1 U9955 ( .A1(n8096), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7674) );
  NAND4_X1 U9956 ( .A1(n7677), .A2(n7676), .A3(n7675), .A4(n7674), .ZN(n13063)
         );
  MUX2_X1 U9957 ( .A(n9783), .B(n6680), .S(n9505), .Z(n7681) );
  NAND2_X1 U9958 ( .A1(n7681), .A2(n14938), .ZN(n7705) );
  INV_X1 U9959 ( .A(n7681), .ZN(n7682) );
  NAND2_X1 U9960 ( .A1(n7682), .A2(SI_12_), .ZN(n7683) );
  XNOR2_X1 U9961 ( .A(n7704), .B(n7703), .ZN(n9782) );
  NAND2_X1 U9962 ( .A1(n9782), .A2(n7960), .ZN(n7688) );
  INV_X1 U9963 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n7684) );
  NAND2_X1 U9964 ( .A1(n7685), .A2(n7684), .ZN(n7709) );
  NAND2_X1 U9965 ( .A1(n7709), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7686) );
  XNOR2_X1 U9966 ( .A(n7686), .B(P2_IR_REG_12__SCAN_IN), .ZN(n14494) );
  AOI22_X1 U9967 ( .A1(n7497), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7859), .B2(
        n14494), .ZN(n7687) );
  MUX2_X1 U9968 ( .A(n13063), .B(n13403), .S(n6467), .Z(n7692) );
  NAND2_X1 U9969 ( .A1(n7691), .A2(n7692), .ZN(n7690) );
  MUX2_X1 U9970 ( .A(n13063), .B(n13403), .S(n6461), .Z(n7689) );
  NAND2_X1 U9971 ( .A1(n7690), .A2(n7689), .ZN(n7696) );
  INV_X1 U9972 ( .A(n7691), .ZN(n7694) );
  INV_X1 U9973 ( .A(n7692), .ZN(n7693) );
  NAND2_X1 U9974 ( .A1(n7694), .A2(n7693), .ZN(n7695) );
  NAND2_X1 U9975 ( .A1(n7580), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7702) );
  NAND2_X1 U9976 ( .A1(n7697), .A2(n11525), .ZN(n7698) );
  NAND2_X1 U9977 ( .A1(n7719), .A2(n7698), .ZN(n11524) );
  OR2_X1 U9978 ( .A1(n8077), .A2(n11524), .ZN(n7701) );
  NAND2_X1 U9979 ( .A1(n7798), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7700) );
  NAND2_X1 U9980 ( .A1(n8096), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7699) );
  NAND4_X1 U9981 ( .A1(n7702), .A2(n7701), .A3(n7700), .A4(n7699), .ZN(n13062)
         );
  MUX2_X1 U9982 ( .A(n9828), .B(n9886), .S(n9505), .Z(n7706) );
  INV_X1 U9983 ( .A(n7706), .ZN(n7707) );
  NAND2_X1 U9984 ( .A1(n7707), .A2(SI_13_), .ZN(n7708) );
  NAND2_X1 U9985 ( .A1(n9827), .A2(n7960), .ZN(n7713) );
  NAND2_X1 U9986 ( .A1(n7728), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7710) );
  INV_X1 U9987 ( .A(n14510), .ZN(n7711) );
  AOI22_X1 U9988 ( .A1(n7711), .A2(n7859), .B1(n7497), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n7712) );
  MUX2_X1 U9989 ( .A(n13062), .B(n13398), .S(n6460), .Z(n7715) );
  MUX2_X1 U9990 ( .A(n13062), .B(n13398), .S(n6467), .Z(n7714) );
  INV_X1 U9991 ( .A(n7715), .ZN(n7716) );
  INV_X1 U9992 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11741) );
  OR2_X1 U9993 ( .A1(n7534), .A2(n11741), .ZN(n7724) );
  INV_X1 U9994 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14935) );
  OR2_X1 U9995 ( .A1(n8076), .A2(n14935), .ZN(n7723) );
  NAND2_X1 U9996 ( .A1(n7580), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7722) );
  INV_X1 U9997 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7718) );
  NAND2_X1 U9998 ( .A1(n7719), .A2(n7718), .ZN(n7720) );
  AND2_X1 U9999 ( .A1(n7743), .A2(n7720), .ZN(n11984) );
  NAND2_X1 U10000 ( .A1(n7717), .A2(n11984), .ZN(n7721) );
  NAND4_X1 U10001 ( .A1(n7724), .A2(n7723), .A3(n7722), .A4(n7721), .ZN(n13061) );
  MUX2_X1 U10002 ( .A(n10051), .B(n10070), .S(n9505), .Z(n7782) );
  NAND2_X1 U10003 ( .A1(n10050), .A2(n7960), .ZN(n7733) );
  INV_X1 U10004 ( .A(n7728), .ZN(n7730) );
  NAND2_X1 U10005 ( .A1(n7730), .A2(n7729), .ZN(n7758) );
  NAND2_X1 U10006 ( .A1(n7758), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7731) );
  XNOR2_X1 U10007 ( .A(n7731), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U10008 ( .A1(n11731), .A2(n7859), .B1(n7497), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n7732) );
  NAND2_X2 U10009 ( .A1(n7733), .A2(n7732), .ZN(n13392) );
  MUX2_X1 U10010 ( .A(n13061), .B(n13392), .S(n6467), .Z(n7737) );
  NAND2_X1 U10011 ( .A1(n7736), .A2(n7737), .ZN(n7735) );
  MUX2_X1 U10012 ( .A(n13061), .B(n13392), .S(n6461), .Z(n7734) );
  NAND2_X1 U10013 ( .A1(n7735), .A2(n7734), .ZN(n7741) );
  INV_X1 U10014 ( .A(n7736), .ZN(n7739) );
  INV_X1 U10015 ( .A(n7737), .ZN(n7738) );
  NAND2_X1 U10016 ( .A1(n7739), .A2(n7738), .ZN(n7740) );
  NAND2_X1 U10017 ( .A1(n7741), .A2(n7740), .ZN(n7766) );
  INV_X1 U10018 ( .A(n7772), .ZN(n7773) );
  NAND2_X1 U10019 ( .A1(n7743), .A2(n7742), .ZN(n7744) );
  NAND2_X1 U10020 ( .A1(n7773), .A2(n7744), .ZN(n11716) );
  OR2_X1 U10021 ( .A1(n11716), .A2(n8077), .ZN(n7749) );
  INV_X1 U10022 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7745) );
  OR2_X1 U10023 ( .A1(n8079), .A2(n7745), .ZN(n7748) );
  NAND2_X1 U10024 ( .A1(n7798), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7747) );
  NAND2_X1 U10025 ( .A1(n8096), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7746) );
  NAND4_X1 U10026 ( .A1(n7749), .A2(n7748), .A3(n7747), .A4(n7746), .ZN(n13060) );
  INV_X1 U10027 ( .A(n7782), .ZN(n7780) );
  NAND2_X1 U10028 ( .A1(n7750), .A2(n7780), .ZN(n7753) );
  INV_X1 U10029 ( .A(n7781), .ZN(n7751) );
  NAND2_X1 U10030 ( .A1(n7751), .A2(SI_14_), .ZN(n7752) );
  NAND2_X1 U10031 ( .A1(n7753), .A2(n7752), .ZN(n7757) );
  MUX2_X1 U10032 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n9505), .Z(n7754) );
  NAND2_X1 U10033 ( .A1(n7754), .A2(SI_15_), .ZN(n7783) );
  INV_X1 U10034 ( .A(n7754), .ZN(n7755) );
  NAND2_X1 U10035 ( .A1(n7755), .A2(n9631), .ZN(n7784) );
  NAND2_X1 U10036 ( .A1(n7783), .A2(n7784), .ZN(n7756) );
  XNOR2_X1 U10037 ( .A(n7757), .B(n7756), .ZN(n10139) );
  NAND2_X1 U10038 ( .A1(n10139), .A2(n7960), .ZN(n7763) );
  OAI21_X1 U10039 ( .B1(n7758), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7759) );
  XNOR2_X1 U10040 ( .A(n7759), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14511) );
  NOR2_X1 U10041 ( .A1(n6455), .A2(n10142), .ZN(n7761) );
  AOI21_X1 U10042 ( .B1(n14511), .B2(n7859), .A(n7761), .ZN(n7762) );
  MUX2_X1 U10043 ( .A(n13060), .B(n13387), .S(n6460), .Z(n7767) );
  NAND2_X1 U10044 ( .A1(n7766), .A2(n7767), .ZN(n7765) );
  MUX2_X1 U10045 ( .A(n13060), .B(n13387), .S(n6467), .Z(n7764) );
  NAND2_X1 U10046 ( .A1(n7765), .A2(n7764), .ZN(n7771) );
  INV_X1 U10047 ( .A(n7766), .ZN(n7769) );
  INV_X1 U10048 ( .A(n7767), .ZN(n7768) );
  NAND2_X1 U10049 ( .A1(n7769), .A2(n7768), .ZN(n7770) );
  INV_X1 U10050 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n7779) );
  NAND2_X1 U10051 ( .A1(n7772), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7796) );
  INV_X1 U10052 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n14867) );
  NAND2_X1 U10053 ( .A1(n7773), .A2(n14867), .ZN(n7774) );
  NAND2_X1 U10054 ( .A1(n7796), .A2(n7774), .ZN(n12979) );
  OR2_X1 U10055 ( .A1(n12979), .A2(n8077), .ZN(n7778) );
  NAND2_X1 U10056 ( .A1(n7580), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7776) );
  NAND2_X1 U10057 ( .A1(n7798), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7775) );
  AND2_X1 U10058 ( .A1(n7776), .A2(n7775), .ZN(n7777) );
  OAI211_X1 U10059 ( .C1(n8076), .C2(n7779), .A(n7778), .B(n7777), .ZN(n13059)
         );
  INV_X1 U10060 ( .A(SI_14_), .ZN(n9588) );
  NAND3_X1 U10061 ( .A1(n7783), .A2(n7782), .A3(n9588), .ZN(n7785) );
  NAND2_X1 U10062 ( .A1(n7787), .A2(n7786), .ZN(n7803) );
  MUX2_X1 U10063 ( .A(n10005), .B(n10053), .S(n9505), .Z(n7788) );
  INV_X1 U10064 ( .A(n7788), .ZN(n7789) );
  NAND2_X1 U10065 ( .A1(n7789), .A2(SI_16_), .ZN(n7790) );
  XNOR2_X1 U10066 ( .A(n7803), .B(n7802), .ZN(n10004) );
  NAND2_X1 U10067 ( .A1(n10004), .A2(n7960), .ZN(n7794) );
  OAI21_X1 U10068 ( .B1(n8174), .B2(n7791), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n7792) );
  XNOR2_X1 U10069 ( .A(n7792), .B(P2_IR_REG_16__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U10070 ( .A1(n7497), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7859), 
        .B2(n11737), .ZN(n7793) );
  MUX2_X1 U10071 ( .A(n13059), .B(n13378), .S(n6467), .Z(n7815) );
  INV_X1 U10072 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7795) );
  NAND2_X1 U10073 ( .A1(n7796), .A2(n7795), .ZN(n7797) );
  AND2_X1 U10074 ( .A1(n7821), .A2(n7797), .ZN(n13292) );
  NAND2_X1 U10075 ( .A1(n13292), .A2(n7717), .ZN(n7801) );
  AOI22_X1 U10076 ( .A1(n7798), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n7580), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n7800) );
  INV_X1 U10077 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14912) );
  OR2_X1 U10078 ( .A1(n8076), .A2(n14912), .ZN(n7799) );
  MUX2_X1 U10079 ( .A(n10097), .B(n10144), .S(n9504), .Z(n7805) );
  INV_X1 U10080 ( .A(n7805), .ZN(n7806) );
  NAND2_X1 U10081 ( .A1(n7806), .A2(SI_17_), .ZN(n7807) );
  XNOR2_X1 U10082 ( .A(n7827), .B(n7826), .ZN(n10096) );
  NAND2_X1 U10083 ( .A1(n10096), .A2(n7960), .ZN(n7813) );
  NAND2_X1 U10084 ( .A1(n7808), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7809) );
  MUX2_X1 U10085 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7809), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n7811) );
  AND2_X1 U10086 ( .A1(n7811), .A2(n7810), .ZN(n14520) );
  AOI22_X1 U10087 ( .A1(n7497), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7859), 
        .B2(n14520), .ZN(n7812) );
  MUX2_X1 U10088 ( .A(n12004), .B(n13295), .S(n6461), .Z(n7816) );
  INV_X1 U10089 ( .A(n12004), .ZN(n13058) );
  AND2_X1 U10090 ( .A1(n13374), .A2(n13058), .ZN(n12025) );
  INV_X1 U10091 ( .A(n13059), .ZN(n12001) );
  INV_X1 U10092 ( .A(n13378), .ZN(n12000) );
  MUX2_X1 U10093 ( .A(n12001), .B(n12000), .S(n6461), .Z(n7814) );
  INV_X1 U10094 ( .A(n7816), .ZN(n7818) );
  NOR2_X1 U10095 ( .A1(n13374), .A2(n13058), .ZN(n7817) );
  OR2_X1 U10096 ( .A1(n7818), .A2(n7817), .ZN(n7819) );
  INV_X1 U10097 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n7825) );
  INV_X1 U10098 ( .A(n7840), .ZN(n7842) );
  NAND2_X1 U10099 ( .A1(n7821), .A2(n14533), .ZN(n7822) );
  NAND2_X1 U10100 ( .A1(n7842), .A2(n7822), .ZN(n13028) );
  OR2_X1 U10101 ( .A1(n13028), .A2(n8077), .ZN(n7824) );
  AOI22_X1 U10102 ( .A1(n7798), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n7580), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n7823) );
  OAI211_X1 U10103 ( .C1(n8076), .C2(n7825), .A(n7824), .B(n7823), .ZN(n13057)
         );
  MUX2_X1 U10104 ( .A(n10390), .B(n10457), .S(n9504), .Z(n7850) );
  XNOR2_X1 U10105 ( .A(n7852), .B(n7850), .ZN(n10389) );
  NAND2_X1 U10106 ( .A1(n10389), .A2(n7960), .ZN(n7831) );
  NAND2_X1 U10107 ( .A1(n7810), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7829) );
  XNOR2_X1 U10108 ( .A(n7829), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13087) );
  AOI22_X1 U10109 ( .A1(n7497), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7859), 
        .B2(n13087), .ZN(n7830) );
  MUX2_X1 U10110 ( .A(n13057), .B(n13369), .S(n6467), .Z(n7835) );
  NAND2_X1 U10111 ( .A1(n7834), .A2(n7835), .ZN(n7833) );
  MUX2_X1 U10112 ( .A(n13057), .B(n13369), .S(n6461), .Z(n7832) );
  NAND2_X1 U10113 ( .A1(n7833), .A2(n7832), .ZN(n7839) );
  INV_X1 U10114 ( .A(n7834), .ZN(n7837) );
  INV_X1 U10115 ( .A(n7835), .ZN(n7836) );
  NAND2_X1 U10116 ( .A1(n7837), .A2(n7836), .ZN(n7838) );
  INV_X1 U10117 ( .A(n7865), .ZN(n7867) );
  INV_X1 U10118 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7841) );
  NAND2_X1 U10119 ( .A1(n7842), .A2(n7841), .ZN(n7843) );
  AND2_X1 U10120 ( .A1(n7867), .A2(n7843), .ZN(n13260) );
  NAND2_X1 U10121 ( .A1(n13260), .A2(n7717), .ZN(n7849) );
  INV_X1 U10122 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n7846) );
  NAND2_X1 U10123 ( .A1(n7580), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n7845) );
  NAND2_X1 U10124 ( .A1(n8096), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n7844) );
  OAI211_X1 U10125 ( .C1(n7534), .C2(n7846), .A(n7845), .B(n7844), .ZN(n7847)
         );
  INV_X1 U10126 ( .A(n7847), .ZN(n7848) );
  NAND2_X1 U10127 ( .A1(n7849), .A2(n7848), .ZN(n13056) );
  INV_X1 U10128 ( .A(n7850), .ZN(n7851) );
  INV_X1 U10129 ( .A(n7853), .ZN(n7854) );
  MUX2_X1 U10130 ( .A(n10559), .B(n10557), .S(n9504), .Z(n7856) );
  INV_X1 U10131 ( .A(n7856), .ZN(n7857) );
  NAND2_X1 U10132 ( .A1(n7857), .A2(SI_19_), .ZN(n7858) );
  NAND2_X1 U10133 ( .A1(n7877), .A2(n7858), .ZN(n7875) );
  XNOR2_X1 U10134 ( .A(n7876), .B(n7875), .ZN(n10555) );
  NAND2_X1 U10135 ( .A1(n10555), .A2(n7960), .ZN(n7861) );
  AOI22_X1 U10136 ( .A1(n7497), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9870), 
        .B2(n7859), .ZN(n7860) );
  MUX2_X1 U10137 ( .A(n13056), .B(n13365), .S(n6460), .Z(n7863) );
  MUX2_X1 U10138 ( .A(n13056), .B(n13365), .S(n6467), .Z(n7862) );
  INV_X1 U10139 ( .A(n7863), .ZN(n7864) );
  INV_X1 U10140 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7866) );
  NAND2_X1 U10141 ( .A1(n7867), .A2(n7866), .ZN(n7868) );
  NAND2_X1 U10142 ( .A1(n7888), .A2(n7868), .ZN(n13244) );
  OR2_X1 U10143 ( .A1(n13244), .A2(n8077), .ZN(n7874) );
  INV_X1 U10144 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n7871) );
  NAND2_X1 U10145 ( .A1(n7580), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n7870) );
  NAND2_X1 U10146 ( .A1(n8096), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n7869) );
  OAI211_X1 U10147 ( .C1(n7534), .C2(n7871), .A(n7870), .B(n7869), .ZN(n7872)
         );
  INV_X1 U10148 ( .A(n7872), .ZN(n7873) );
  NAND2_X1 U10149 ( .A1(n7874), .A2(n7873), .ZN(n13055) );
  INV_X1 U10150 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11022) );
  MUX2_X1 U10151 ( .A(n10994), .B(n11022), .S(n9504), .Z(n7896) );
  XNOR2_X1 U10152 ( .A(n7898), .B(n7896), .ZN(n10993) );
  NAND2_X1 U10153 ( .A1(n10993), .A2(n7960), .ZN(n7879) );
  OR2_X1 U10154 ( .A1(n6455), .A2(n10994), .ZN(n7878) );
  MUX2_X1 U10155 ( .A(n13055), .B(n13359), .S(n6467), .Z(n7883) );
  NAND2_X1 U10156 ( .A1(n7882), .A2(n7883), .ZN(n7881) );
  MUX2_X1 U10157 ( .A(n13055), .B(n13359), .S(n6461), .Z(n7880) );
  NAND2_X1 U10158 ( .A1(n7881), .A2(n7880), .ZN(n7887) );
  INV_X1 U10159 ( .A(n7882), .ZN(n7885) );
  INV_X1 U10160 ( .A(n7883), .ZN(n7884) );
  NAND2_X1 U10161 ( .A1(n7885), .A2(n7884), .ZN(n7886) );
  INV_X1 U10162 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12960) );
  NAND2_X1 U10163 ( .A1(n7888), .A2(n12960), .ZN(n7889) );
  AND2_X1 U10164 ( .A1(n7906), .A2(n7889), .ZN(n13227) );
  NAND2_X1 U10165 ( .A1(n13227), .A2(n7717), .ZN(n7895) );
  INV_X1 U10166 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n7892) );
  NAND2_X1 U10167 ( .A1(n7580), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7891) );
  NAND2_X1 U10168 ( .A1(n8096), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7890) );
  OAI211_X1 U10169 ( .C1(n7534), .C2(n7892), .A(n7891), .B(n7890), .ZN(n7893)
         );
  INV_X1 U10170 ( .A(n7893), .ZN(n7894) );
  NAND2_X1 U10171 ( .A1(n7895), .A2(n7894), .ZN(n13054) );
  INV_X1 U10172 ( .A(n7896), .ZN(n7897) );
  INV_X1 U10173 ( .A(SI_20_), .ZN(n10453) );
  MUX2_X1 U10174 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n9504), .Z(n7916) );
  XNOR2_X1 U10175 ( .A(n7916), .B(SI_21_), .ZN(n7913) );
  XNOR2_X1 U10176 ( .A(n7915), .B(n7913), .ZN(n11142) );
  NAND2_X1 U10177 ( .A1(n11142), .A2(n7960), .ZN(n7902) );
  OR2_X1 U10178 ( .A1(n6455), .A2(n11145), .ZN(n7901) );
  MUX2_X1 U10179 ( .A(n13054), .B(n13354), .S(n6460), .Z(n7904) );
  MUX2_X1 U10180 ( .A(n13054), .B(n13354), .S(n6467), .Z(n7903) );
  INV_X1 U10181 ( .A(n7904), .ZN(n7905) );
  INV_X1 U10182 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13017) );
  AND2_X1 U10183 ( .A1(n7906), .A2(n13017), .ZN(n7907) );
  OR2_X1 U10184 ( .A1(n7907), .A2(n7928), .ZN(n13211) );
  INV_X1 U10185 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n7910) );
  NAND2_X1 U10186 ( .A1(n7580), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n7909) );
  NAND2_X1 U10187 ( .A1(n8096), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n7908) );
  OAI211_X1 U10188 ( .C1(n7534), .C2(n7910), .A(n7909), .B(n7908), .ZN(n7911)
         );
  INV_X1 U10189 ( .A(n7911), .ZN(n7912) );
  NAND2_X1 U10190 ( .A1(n7916), .A2(SI_21_), .ZN(n7917) );
  MUX2_X1 U10191 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n9504), .Z(n7956) );
  XNOR2_X1 U10192 ( .A(n9161), .B(n7954), .ZN(n11388) );
  NAND2_X1 U10193 ( .A1(n11388), .A2(n7960), .ZN(n7919) );
  OR2_X1 U10194 ( .A1(n6455), .A2(n11391), .ZN(n7918) );
  MUX2_X1 U10195 ( .A(n13012), .B(n13349), .S(n6467), .Z(n7923) );
  NAND2_X1 U10196 ( .A1(n7922), .A2(n7923), .ZN(n7921) );
  MUX2_X1 U10197 ( .A(n13012), .B(n13349), .S(n6460), .Z(n7920) );
  NAND2_X1 U10198 ( .A1(n7921), .A2(n7920), .ZN(n7927) );
  INV_X1 U10199 ( .A(n7922), .ZN(n7925) );
  INV_X1 U10200 ( .A(n7923), .ZN(n7924) );
  NAND2_X1 U10201 ( .A1(n7925), .A2(n7924), .ZN(n7926) );
  OR2_X1 U10202 ( .A1(n7928), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n7929) );
  NAND2_X1 U10203 ( .A1(n7928), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n7945) );
  NAND2_X1 U10204 ( .A1(n7929), .A2(n7945), .ZN(n13197) );
  OR2_X1 U10205 ( .A1(n13197), .A2(n8077), .ZN(n7935) );
  INV_X1 U10206 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n7932) );
  NAND2_X1 U10207 ( .A1(n7580), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n7931) );
  NAND2_X1 U10208 ( .A1(n8096), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n7930) );
  OAI211_X1 U10209 ( .C1(n7534), .C2(n7932), .A(n7931), .B(n7930), .ZN(n7933)
         );
  INV_X1 U10210 ( .A(n7933), .ZN(n7934) );
  NAND2_X1 U10211 ( .A1(n7935), .A2(n7934), .ZN(n13053) );
  NAND2_X1 U10212 ( .A1(n9161), .A2(n7956), .ZN(n7937) );
  NAND2_X1 U10213 ( .A1(n7953), .A2(SI_22_), .ZN(n7936) );
  NAND2_X1 U10214 ( .A1(n7937), .A2(n7936), .ZN(n7939) );
  MUX2_X1 U10215 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n9504), .Z(n7957) );
  XNOR2_X1 U10216 ( .A(n7957), .B(SI_23_), .ZN(n7938) );
  NAND2_X1 U10217 ( .A1(n11444), .A2(n7960), .ZN(n7941) );
  INV_X1 U10218 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11442) );
  OR2_X1 U10219 ( .A1(n6455), .A2(n11442), .ZN(n7940) );
  MUX2_X1 U10220 ( .A(n13053), .B(n13344), .S(n6461), .Z(n7943) );
  MUX2_X1 U10221 ( .A(n13053), .B(n13344), .S(n6467), .Z(n7942) );
  INV_X1 U10222 ( .A(n7943), .ZN(n7944) );
  NAND2_X1 U10223 ( .A1(n7580), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n7950) );
  NAND2_X1 U10224 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n7946), .ZN(n8006) );
  OAI21_X1 U10225 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n7946), .A(n8006), .ZN(
        n13181) );
  OR2_X1 U10226 ( .A1(n8077), .A2(n13181), .ZN(n7949) );
  NAND2_X1 U10227 ( .A1(n7798), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n7948) );
  NAND2_X1 U10228 ( .A1(n8096), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n7947) );
  NAND4_X1 U10229 ( .A1(n7950), .A2(n7949), .A3(n7948), .A4(n7947), .ZN(n13052) );
  INV_X1 U10230 ( .A(n7957), .ZN(n7951) );
  AOI22_X1 U10231 ( .A1(n8235), .A2(n7954), .B1(n7951), .B2(n11103), .ZN(n7952) );
  OAI21_X1 U10232 ( .B1(n7954), .B2(n8235), .A(n11103), .ZN(n7958) );
  AND2_X1 U10233 ( .A1(SI_22_), .A2(SI_23_), .ZN(n7955) );
  AOI22_X1 U10234 ( .A1(n7958), .A2(n7957), .B1(n7956), .B2(n7955), .ZN(n7959)
         );
  MUX2_X1 U10235 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n9504), .Z(n7978) );
  XNOR2_X1 U10236 ( .A(n7977), .B(n7978), .ZN(n11531) );
  NAND2_X1 U10237 ( .A1(n11531), .A2(n7960), .ZN(n7962) );
  OR2_X1 U10238 ( .A1(n6455), .A2(n14948), .ZN(n7961) );
  MUX2_X1 U10239 ( .A(n13052), .B(n13338), .S(n8107), .Z(n7966) );
  NAND2_X1 U10240 ( .A1(n7965), .A2(n7966), .ZN(n7964) );
  MUX2_X1 U10241 ( .A(n13052), .B(n13338), .S(n6461), .Z(n7963) );
  NAND2_X1 U10242 ( .A1(n7580), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n7976) );
  INV_X1 U10243 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n7967) );
  OR2_X1 U10244 ( .A1(n7534), .A2(n7967), .ZN(n7975) );
  INV_X1 U10245 ( .A(n8006), .ZN(n7968) );
  NAND2_X1 U10246 ( .A1(n7969), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8028) );
  INV_X1 U10247 ( .A(n7969), .ZN(n7993) );
  INV_X1 U10248 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7970) );
  NAND2_X1 U10249 ( .A1(n7993), .A2(n7970), .ZN(n7971) );
  NAND2_X1 U10250 ( .A1(n8028), .A2(n7971), .ZN(n13133) );
  OR2_X1 U10251 ( .A1(n8077), .A2(n13133), .ZN(n7974) );
  INV_X1 U10252 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n7972) );
  OR2_X1 U10253 ( .A1(n8076), .A2(n7972), .ZN(n7973) );
  INV_X1 U10254 ( .A(n7977), .ZN(n7979) );
  NAND2_X1 U10255 ( .A1(n7979), .A2(n7978), .ZN(n7982) );
  NAND2_X1 U10256 ( .A1(n7980), .A2(SI_24_), .ZN(n7981) );
  NAND2_X1 U10257 ( .A1(n7982), .A2(n7981), .ZN(n8015) );
  MUX2_X1 U10258 ( .A(n11613), .B(n11616), .S(n9505), .Z(n7983) );
  INV_X1 U10259 ( .A(SI_25_), .ZN(n11608) );
  NAND2_X1 U10260 ( .A1(n7983), .A2(n11608), .ZN(n7986) );
  INV_X1 U10261 ( .A(n7983), .ZN(n7984) );
  NAND2_X1 U10262 ( .A1(n7984), .A2(SI_25_), .ZN(n7985) );
  NAND2_X1 U10263 ( .A1(n7986), .A2(n7985), .ZN(n8014) );
  MUX2_X1 U10264 ( .A(n13442), .B(n6674), .S(n9504), .Z(n7999) );
  INV_X1 U10265 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14882) );
  INV_X1 U10266 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n11842) );
  MUX2_X1 U10267 ( .A(n14882), .B(n11842), .S(n9504), .Z(n8035) );
  XNOR2_X1 U10268 ( .A(n8035), .B(SI_27_), .ZN(n7987) );
  NAND2_X1 U10269 ( .A1(n11841), .A2(n7960), .ZN(n7989) );
  OR2_X1 U10270 ( .A1(n6455), .A2(n14882), .ZN(n7988) );
  MUX2_X1 U10271 ( .A(n12952), .B(n13128), .S(n6467), .Z(n8051) );
  NAND2_X1 U10272 ( .A1(n8051), .A2(n8050), .ZN(n8049) );
  NAND2_X1 U10273 ( .A1(n7580), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n7998) );
  INV_X1 U10274 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n7990) );
  OR2_X1 U10275 ( .A1(n7534), .A2(n7990), .ZN(n7997) );
  INV_X1 U10276 ( .A(n7991), .ZN(n8008) );
  INV_X1 U10277 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13039) );
  NAND2_X1 U10278 ( .A1(n8008), .A2(n13039), .ZN(n7992) );
  NAND2_X1 U10279 ( .A1(n7993), .A2(n7992), .ZN(n13147) );
  OR2_X1 U10280 ( .A1(n8077), .A2(n13147), .ZN(n7996) );
  INV_X1 U10281 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n7994) );
  OR2_X1 U10282 ( .A1(n8076), .A2(n7994), .ZN(n7995) );
  XNOR2_X1 U10283 ( .A(n7999), .B(SI_26_), .ZN(n8000) );
  XNOR2_X1 U10284 ( .A(n8001), .B(n8000), .ZN(n13441) );
  NAND2_X1 U10285 ( .A1(n13441), .A2(n7960), .ZN(n8003) );
  OR2_X1 U10286 ( .A1(n6455), .A2(n13442), .ZN(n8002) );
  MUX2_X1 U10287 ( .A(n12968), .B(n13326), .S(n6467), .Z(n8046) );
  INV_X1 U10288 ( .A(n12968), .ZN(n13050) );
  MUX2_X1 U10289 ( .A(n13050), .B(n13150), .S(n6461), .Z(n8045) );
  NAND2_X1 U10290 ( .A1(n8046), .A2(n8045), .ZN(n8004) );
  NAND2_X1 U10291 ( .A1(n7580), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8013) );
  INV_X1 U10292 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14854) );
  OR2_X1 U10293 ( .A1(n7534), .A2(n14854), .ZN(n8012) );
  INV_X1 U10294 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8005) );
  NAND2_X1 U10295 ( .A1(n8006), .A2(n8005), .ZN(n8007) );
  NAND2_X1 U10296 ( .A1(n8008), .A2(n8007), .ZN(n13165) );
  OR2_X1 U10297 ( .A1(n8077), .A2(n13165), .ZN(n8011) );
  INV_X1 U10298 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8009) );
  OR2_X1 U10299 ( .A1(n8076), .A2(n8009), .ZN(n8010) );
  XNOR2_X1 U10300 ( .A(n8015), .B(n8014), .ZN(n11611) );
  NAND2_X1 U10301 ( .A1(n11611), .A2(n7960), .ZN(n8017) );
  OR2_X1 U10302 ( .A1(n6455), .A2(n11613), .ZN(n8016) );
  MUX2_X1 U10303 ( .A(n12985), .B(n13332), .S(n6467), .Z(n8023) );
  MUX2_X1 U10304 ( .A(n13051), .B(n13167), .S(n6460), .Z(n8022) );
  NAND2_X1 U10305 ( .A1(n8023), .A2(n8022), .ZN(n8018) );
  AND2_X1 U10306 ( .A1(n8021), .A2(n8018), .ZN(n8019) );
  NAND2_X1 U10307 ( .A1(n8020), .A2(n8019), .ZN(n8090) );
  INV_X1 U10308 ( .A(n8021), .ZN(n8024) );
  OR3_X1 U10309 ( .A1(n8024), .A2(n8023), .A3(n8022), .ZN(n8057) );
  NAND2_X1 U10310 ( .A1(n7580), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8034) );
  INV_X1 U10311 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8025) );
  OR2_X1 U10312 ( .A1(n7534), .A2(n8025), .ZN(n8033) );
  INV_X1 U10313 ( .A(n8028), .ZN(n8026) );
  NAND2_X1 U10314 ( .A1(n8026), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n12020) );
  INV_X1 U10315 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8027) );
  NAND2_X1 U10316 ( .A1(n8028), .A2(n8027), .ZN(n8029) );
  NAND2_X1 U10317 ( .A1(n12020), .A2(n8029), .ZN(n13114) );
  OR2_X1 U10318 ( .A1(n8077), .A2(n13114), .ZN(n8032) );
  INV_X1 U10319 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8030) );
  OR2_X1 U10320 ( .A1(n8076), .A2(n8030), .ZN(n8031) );
  INV_X1 U10321 ( .A(n8035), .ZN(n8038) );
  NOR2_X1 U10322 ( .A1(n8038), .A2(SI_27_), .ZN(n8036) );
  NAND2_X1 U10323 ( .A1(n8038), .A2(SI_27_), .ZN(n8039) );
  MUX2_X1 U10324 ( .A(n13439), .B(n14011), .S(n9504), .Z(n8040) );
  NAND2_X1 U10325 ( .A1(n8040), .A2(n14863), .ZN(n8058) );
  INV_X1 U10326 ( .A(n8040), .ZN(n8041) );
  NAND2_X1 U10327 ( .A1(n8041), .A2(SI_28_), .ZN(n8042) );
  NAND2_X1 U10328 ( .A1(n8058), .A2(n8042), .ZN(n8059) );
  NAND2_X1 U10329 ( .A1(n14008), .A2(n7960), .ZN(n8044) );
  OR2_X1 U10330 ( .A1(n6455), .A2(n13439), .ZN(n8043) );
  AND2_X2 U10331 ( .A1(n8044), .A2(n8043), .ZN(n13118) );
  MUX2_X1 U10332 ( .A(n12922), .B(n13118), .S(n6460), .Z(n8092) );
  MUX2_X1 U10333 ( .A(n13048), .B(n13315), .S(n8107), .Z(n8091) );
  NAND2_X1 U10334 ( .A1(n8092), .A2(n8091), .ZN(n8056) );
  INV_X1 U10335 ( .A(n8045), .ZN(n8048) );
  INV_X1 U10336 ( .A(n8046), .ZN(n8047) );
  NAND3_X1 U10337 ( .A1(n8049), .A2(n8048), .A3(n8047), .ZN(n8055) );
  INV_X1 U10338 ( .A(n8050), .ZN(n8053) );
  INV_X1 U10339 ( .A(n8051), .ZN(n8052) );
  NAND2_X1 U10340 ( .A1(n8053), .A2(n8052), .ZN(n8054) );
  INV_X1 U10341 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13434) );
  INV_X1 U10342 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14007) );
  MUX2_X1 U10343 ( .A(n13434), .B(n14007), .S(n9504), .Z(n8061) );
  XNOR2_X1 U10344 ( .A(n8061), .B(SI_29_), .ZN(n8084) );
  NAND2_X1 U10345 ( .A1(n8085), .A2(n8084), .ZN(n8063) );
  INV_X1 U10346 ( .A(SI_29_), .ZN(n12875) );
  NAND2_X1 U10347 ( .A1(n8061), .A2(n12875), .ZN(n8062) );
  NAND2_X1 U10348 ( .A1(n8063), .A2(n8062), .ZN(n8101) );
  MUX2_X1 U10349 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n9504), .Z(n8064) );
  NAND2_X1 U10350 ( .A1(n8064), .A2(SI_30_), .ZN(n8067) );
  INV_X1 U10351 ( .A(n8064), .ZN(n8065) );
  INV_X1 U10352 ( .A(SI_30_), .ZN(n14880) );
  NAND2_X1 U10353 ( .A1(n8065), .A2(n14880), .ZN(n8066) );
  NAND2_X1 U10354 ( .A1(n8067), .A2(n8066), .ZN(n8100) );
  MUX2_X1 U10355 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n9504), .Z(n8068) );
  XNOR2_X1 U10356 ( .A(n8068), .B(SI_31_), .ZN(n8069) );
  NAND2_X1 U10357 ( .A1(n13427), .A2(n7960), .ZN(n8072) );
  INV_X1 U10358 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12094) );
  OR2_X1 U10359 ( .A1(n6455), .A2(n12094), .ZN(n8071) );
  INV_X1 U10360 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n14883) );
  NAND2_X1 U10361 ( .A1(n7580), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8074) );
  NAND2_X1 U10362 ( .A1(n8096), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8073) );
  OAI211_X1 U10363 ( .C1(n7534), .C2(n14883), .A(n8074), .B(n8073), .ZN(n13101) );
  XNOR2_X1 U10364 ( .A(n13103), .B(n13101), .ZN(n8162) );
  NAND2_X1 U10365 ( .A1(n7484), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8083) );
  INV_X1 U10366 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8075) );
  OR2_X1 U10367 ( .A1(n8076), .A2(n8075), .ZN(n8082) );
  OR2_X1 U10368 ( .A1(n8077), .A2(n12020), .ZN(n8081) );
  INV_X1 U10369 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8078) );
  OR2_X1 U10370 ( .A1(n8079), .A2(n8078), .ZN(n8080) );
  AND4_X1 U10371 ( .A1(n8083), .A2(n8082), .A3(n8081), .A4(n8080), .ZN(n12953)
         );
  NAND2_X1 U10372 ( .A1(n13433), .A2(n7960), .ZN(n8087) );
  OR2_X1 U10373 ( .A1(n6455), .A2(n13434), .ZN(n8086) );
  MUX2_X1 U10374 ( .A(n12953), .B(n12023), .S(n6461), .Z(n8113) );
  MUX2_X1 U10375 ( .A(n13047), .B(n13310), .S(n8107), .Z(n8112) );
  NAND2_X1 U10376 ( .A1(n8113), .A2(n8112), .ZN(n8094) );
  NAND2_X1 U10377 ( .A1(n8162), .A2(n8094), .ZN(n8088) );
  NOR2_X1 U10378 ( .A1(n7358), .A2(n8088), .ZN(n8089) );
  INV_X1 U10379 ( .A(n8091), .ZN(n8095) );
  INV_X1 U10380 ( .A(n8092), .ZN(n8093) );
  NAND4_X1 U10381 ( .A1(n8162), .A2(n8095), .A3(n8094), .A4(n8093), .ZN(n8118)
         );
  INV_X1 U10382 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8099) );
  NAND2_X1 U10383 ( .A1(n7580), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8098) );
  NAND2_X1 U10384 ( .A1(n8096), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8097) );
  OAI211_X1 U10385 ( .C1(n7534), .C2(n8099), .A(n8098), .B(n8097), .ZN(n13046)
         );
  NAND2_X1 U10386 ( .A1(n8101), .A2(n8100), .ZN(n8102) );
  OR2_X1 U10387 ( .A1(n14004), .A2(n8104), .ZN(n8106) );
  INV_X1 U10388 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12066) );
  OR2_X1 U10389 ( .A1(n6455), .A2(n12066), .ZN(n8105) );
  MUX2_X1 U10390 ( .A(n13046), .B(n13097), .S(n8107), .Z(n8121) );
  NAND2_X1 U10391 ( .A1(n13101), .A2(n6467), .ZN(n8109) );
  XNOR2_X2 U10392 ( .A(n8108), .B(P2_IR_REG_22__SCAN_IN), .ZN(n9866) );
  NAND2_X1 U10393 ( .A1(n10195), .A2(n9866), .ZN(n8129) );
  NAND4_X1 U10394 ( .A1(n8109), .A2(n11143), .A3(n8129), .A4(n10013), .ZN(
        n8110) );
  AND2_X1 U10395 ( .A1(n8110), .A2(n13046), .ZN(n8111) );
  AOI21_X1 U10396 ( .B1(n13097), .B2(n6461), .A(n8111), .ZN(n8120) );
  OAI22_X1 U10397 ( .A1(n8121), .A2(n8120), .B1(n8113), .B2(n8112), .ZN(n8116)
         );
  OR2_X1 U10398 ( .A1(n13103), .A2(n13101), .ZN(n8122) );
  NAND2_X1 U10399 ( .A1(n13103), .A2(n13101), .ZN(n8114) );
  NAND2_X1 U10400 ( .A1(n8122), .A2(n8114), .ZN(n8115) );
  NAND2_X1 U10401 ( .A1(n8116), .A2(n8115), .ZN(n8117) );
  NAND3_X1 U10402 ( .A1(n8119), .A2(n8118), .A3(n8117), .ZN(n8128) );
  NAND2_X1 U10403 ( .A1(n8121), .A2(n8120), .ZN(n8127) );
  INV_X1 U10404 ( .A(n8122), .ZN(n8125) );
  MUX2_X1 U10405 ( .A(n13101), .B(n13103), .S(n6460), .Z(n8124) );
  NOR2_X1 U10406 ( .A1(n8125), .A2(n8124), .ZN(n8126) );
  AOI21_X2 U10407 ( .B1(n8128), .B2(n8127), .A(n8126), .ZN(n8164) );
  NAND2_X1 U10408 ( .A1(n10010), .A2(n11143), .ZN(n9872) );
  OAI21_X1 U10409 ( .B1(n9872), .B2(n13093), .A(n8129), .ZN(n8130) );
  INV_X1 U10410 ( .A(n8130), .ZN(n8134) );
  NAND2_X1 U10411 ( .A1(n11143), .A2(n13093), .ZN(n8131) );
  OAI211_X1 U10412 ( .C1(n10021), .C2(n9866), .A(n8131), .B(n10013), .ZN(n8132) );
  NAND2_X1 U10413 ( .A1(n8164), .A2(n8132), .ZN(n8133) );
  OAI21_X1 U10414 ( .B1(n8164), .B2(n8134), .A(n8133), .ZN(n8168) );
  NAND2_X1 U10415 ( .A1(n13315), .A2(n13048), .ZN(n12037) );
  NAND2_X1 U10416 ( .A1(n13150), .A2(n12968), .ZN(n12010) );
  NAND2_X1 U10417 ( .A1(n12012), .A2(n12010), .ZN(n13143) );
  XNOR2_X1 U10418 ( .A(n13167), .B(n12985), .ZN(n13161) );
  INV_X1 U10419 ( .A(n13052), .ZN(n12927) );
  XNOR2_X1 U10420 ( .A(n13338), .B(n12927), .ZN(n13174) );
  INV_X1 U10421 ( .A(n13053), .ZN(n12986) );
  XNOR2_X1 U10422 ( .A(n13344), .B(n12986), .ZN(n13198) );
  INV_X1 U10423 ( .A(n13012), .ZN(n12928) );
  INV_X1 U10424 ( .A(n13054), .ZN(n12998) );
  XNOR2_X1 U10425 ( .A(n13354), .B(n12998), .ZN(n13222) );
  INV_X1 U10426 ( .A(n13055), .ZN(n12007) );
  XNOR2_X1 U10427 ( .A(n13359), .B(n12007), .ZN(n13246) );
  INV_X1 U10428 ( .A(n13056), .ZN(n12996) );
  XNOR2_X1 U10429 ( .A(n13365), .B(n12996), .ZN(n13254) );
  INV_X1 U10430 ( .A(n13057), .ZN(n12005) );
  XNOR2_X1 U10431 ( .A(n13369), .B(n12005), .ZN(n12027) );
  XNOR2_X1 U10432 ( .A(n13374), .B(n12004), .ZN(n13297) );
  XNOR2_X1 U10433 ( .A(n13378), .B(n12001), .ZN(n11763) );
  INV_X1 U10434 ( .A(n13060), .ZN(n11764) );
  NAND2_X1 U10435 ( .A1(n13387), .A2(n11764), .ZN(n11761) );
  OR2_X1 U10436 ( .A1(n13387), .A2(n11764), .ZN(n8137) );
  NAND2_X1 U10437 ( .A1(n11761), .A2(n8137), .ZN(n11719) );
  OR2_X1 U10438 ( .A1(n13392), .A2(n13061), .ZN(n11708) );
  NAND2_X1 U10439 ( .A1(n13392), .A2(n13061), .ZN(n11710) );
  NAND2_X1 U10440 ( .A1(n11708), .A2(n11710), .ZN(n11436) );
  INV_X1 U10441 ( .A(n13063), .ZN(n8138) );
  OR2_X1 U10442 ( .A1(n13403), .A2(n8138), .ZN(n11211) );
  NAND2_X1 U10443 ( .A1(n13403), .A2(n8138), .ZN(n8139) );
  NAND2_X1 U10444 ( .A1(n11211), .A2(n8139), .ZN(n11128) );
  XNOR2_X1 U10445 ( .A(n11146), .B(n13065), .ZN(n10982) );
  XNOR2_X1 U10446 ( .A(n10953), .B(n10742), .ZN(n10946) );
  XNOR2_X1 U10447 ( .A(n10694), .B(n13069), .ZN(n10670) );
  INV_X1 U10448 ( .A(n13070), .ZN(n10672) );
  OR2_X1 U10449 ( .A1(n10507), .A2(n10672), .ZN(n8140) );
  NAND2_X1 U10450 ( .A1(n10507), .A2(n10672), .ZN(n10515) );
  INV_X1 U10451 ( .A(n14566), .ZN(n8141) );
  NAND2_X1 U10452 ( .A1(n14566), .A2(n10262), .ZN(n10290) );
  INV_X1 U10453 ( .A(n9869), .ZN(n8143) );
  AND2_X1 U10454 ( .A1(n10215), .A2(n8144), .ZN(n10199) );
  NAND4_X1 U10455 ( .A1(n10199), .A2(n10278), .A3(n10010), .A4(n9891), .ZN(
        n8151) );
  INV_X1 U10456 ( .A(n10772), .ZN(n14561) );
  NAND2_X1 U10457 ( .A1(n14561), .A2(n8149), .ZN(n8150) );
  NAND2_X1 U10458 ( .A1(n8150), .A2(n10565), .ZN(n10288) );
  NOR2_X1 U10459 ( .A1(n8151), .A2(n10288), .ZN(n8152) );
  NAND4_X1 U10460 ( .A1(n10670), .A2(n10504), .A3(n10562), .A4(n8152), .ZN(
        n8153) );
  NOR2_X1 U10461 ( .A1(n10946), .A2(n8153), .ZN(n8154) );
  XNOR2_X1 U10462 ( .A(n11090), .B(n13066), .ZN(n10849) );
  XNOR2_X1 U10463 ( .A(n10890), .B(n13067), .ZN(n10522) );
  NAND4_X1 U10464 ( .A1(n10982), .A2(n8154), .A3(n10849), .A4(n10522), .ZN(
        n8155) );
  NOR2_X1 U10465 ( .A1(n11128), .A2(n8155), .ZN(n8156) );
  XNOR2_X1 U10466 ( .A(n11174), .B(n13064), .ZN(n11068) );
  NAND4_X1 U10467 ( .A1(n11436), .A2(n8156), .A3(n11213), .A4(n11068), .ZN(
        n8157) );
  OR4_X1 U10468 ( .A1(n13297), .A2(n11763), .A3(n11719), .A4(n8157), .ZN(n8158) );
  OR4_X1 U10469 ( .A1(n13143), .A2(n13161), .A3(n13174), .A4(n8160), .ZN(n8161) );
  XNOR2_X1 U10470 ( .A(n13310), .B(n13047), .ZN(n12038) );
  XNOR2_X1 U10471 ( .A(n6552), .B(n13093), .ZN(n8163) );
  XNOR2_X1 U10472 ( .A(n8170), .B(n8169), .ZN(n9634) );
  OR2_X1 U10473 ( .A1(n9634), .A2(P2_U3088), .ZN(n11440) );
  INV_X1 U10474 ( .A(n11440), .ZN(n8166) );
  OAI21_X1 U10475 ( .B1(n8168), .B2(n8167), .A(n8166), .ZN(n8187) );
  NAND2_X1 U10476 ( .A1(n8170), .A2(n8169), .ZN(n8171) );
  OAI21_X1 U10477 ( .B1(n8174), .B2(n8173), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8175) );
  MUX2_X1 U10478 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8175), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8176) );
  NAND2_X1 U10479 ( .A1(n8176), .A2(n7151), .ZN(n11612) );
  NAND2_X1 U10480 ( .A1(n7151), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8177) );
  MUX2_X1 U10481 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8177), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8178) );
  NAND2_X1 U10482 ( .A1(n8178), .A2(n7410), .ZN(n13443) );
  NOR2_X1 U10483 ( .A1(n11612), .A2(n13443), .ZN(n8179) );
  NAND2_X1 U10484 ( .A1(n11532), .A2(n8179), .ZN(n9633) );
  INV_X1 U10485 ( .A(n8181), .ZN(n8182) );
  NAND2_X1 U10486 ( .A1(n10017), .A2(n8182), .ZN(n12995) );
  NOR4_X1 U10487 ( .A1(n14553), .A2(n12995), .A3(n8183), .A4(n10013), .ZN(
        n8185) );
  OAI21_X1 U10488 ( .B1(n11440), .B2(n9866), .A(P2_B_REG_SCAN_IN), .ZN(n8184)
         );
  OR2_X1 U10489 ( .A1(n8185), .A2(n8184), .ZN(n8186) );
  NAND2_X1 U10490 ( .A1(n8187), .A2(n8186), .ZN(P2_U3328) );
  AOI22_X1 U10491 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n10559), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n10557), .ZN(n8538) );
  XNOR2_X1 U10492 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n8441) );
  XNOR2_X1 U10493 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8323) );
  NAND2_X1 U10494 ( .A1(n8323), .A2(n8338), .ZN(n8190) );
  NAND2_X1 U10495 ( .A1(n7413), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8189) );
  NAND2_X1 U10496 ( .A1(n8190), .A2(n8189), .ZN(n8352) );
  XNOR2_X1 U10497 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8350) );
  NAND2_X1 U10498 ( .A1(n8352), .A2(n8350), .ZN(n8192) );
  NAND2_X1 U10499 ( .A1(n9530), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8191) );
  NAND2_X1 U10500 ( .A1(n8192), .A2(n8191), .ZN(n8368) );
  NAND2_X1 U10501 ( .A1(n8368), .A2(n8366), .ZN(n8194) );
  INV_X1 U10502 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9532) );
  NAND2_X1 U10503 ( .A1(n9532), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8193) );
  NAND2_X1 U10504 ( .A1(n8194), .A2(n8193), .ZN(n8384) );
  NAND2_X1 U10505 ( .A1(n8384), .A2(n8382), .ZN(n8196) );
  NAND2_X1 U10506 ( .A1(n9536), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8195) );
  NAND2_X1 U10507 ( .A1(n8196), .A2(n8195), .ZN(n8256) );
  NAND2_X1 U10508 ( .A1(n9540), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U10509 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n14864), .ZN(n8198) );
  NAND2_X1 U10510 ( .A1(n9554), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8199) );
  XNOR2_X1 U10511 ( .A(n9558), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n8284) );
  NAND2_X1 U10512 ( .A1(n9558), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U10513 ( .A1(n9573), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8202) );
  XNOR2_X1 U10514 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n8312) );
  NAND2_X1 U10515 ( .A1(n9586), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8203) );
  NAND2_X1 U10516 ( .A1(n8204), .A2(n8203), .ZN(n8408) );
  XNOR2_X1 U10517 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8407) );
  NAND2_X1 U10518 ( .A1(n9592), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8205) );
  XNOR2_X1 U10519 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8422) );
  XNOR2_X1 U10520 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8457) );
  NAND2_X1 U10521 ( .A1(n10070), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8208) );
  XNOR2_X1 U10522 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n8474) );
  NAND2_X1 U10523 ( .A1(n8476), .A2(n8474), .ZN(n8209) );
  AOI22_X1 U10524 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n10005), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n10053), .ZN(n8489) );
  AOI22_X1 U10525 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n10097), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n10144), .ZN(n8504) );
  NAND2_X1 U10526 ( .A1(n8506), .A2(n8504), .ZN(n8212) );
  AOI22_X1 U10527 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n10390), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n10457), .ZN(n8522) );
  NAND2_X1 U10528 ( .A1(n8538), .A2(n8539), .ZN(n8216) );
  NAND2_X1 U10529 ( .A1(n8553), .A2(n11022), .ZN(n8219) );
  NAND2_X1 U10530 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n8217), .ZN(n8218) );
  INV_X1 U10531 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12382) );
  AOI22_X1 U10532 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n11145), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n12382), .ZN(n8564) );
  INV_X1 U10533 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9689) );
  AOI22_X1 U10534 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_22__SCAN_IN), .B1(n11391), .B2(n9689), .ZN(n8579) );
  XNOR2_X1 U10535 ( .A(n8580), .B(n8579), .ZN(n10807) );
  AND3_X2 U10536 ( .A1(n8272), .A2(n8259), .A3(n8369), .ZN(n8222) );
  NOR2_X2 U10537 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n8221) );
  NOR2_X2 U10538 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8220) );
  NOR2_X1 U10539 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n8229) );
  NOR2_X1 U10540 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n8228) );
  AND2_X4 U10541 ( .A1(n10307), .A2(n9504), .ZN(n8353) );
  NAND2_X1 U10542 ( .A1(n10807), .A2(n8353), .ZN(n8237) );
  OR2_X1 U10543 ( .A1(n9361), .A2(n8235), .ZN(n8236) );
  NOR2_X1 U10544 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8376) );
  NAND2_X1 U10545 ( .A1(n8376), .A2(n10472), .ZN(n8264) );
  NAND2_X1 U10546 ( .A1(n8571), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8238) );
  NAND2_X1 U10547 ( .A1(n8583), .A2(n8238), .ZN(n12722) );
  INV_X1 U10548 ( .A(n8239), .ZN(n8241) );
  NAND2_X1 U10549 ( .A1(n8241), .A2(n8240), .ZN(n8243) );
  XNOR2_X2 U10550 ( .A(n8242), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8246) );
  AND2_X2 U10551 ( .A1(n8246), .A2(n8245), .ZN(n8344) );
  NAND2_X1 U10552 ( .A1(n12722), .A2(n8484), .ZN(n8249) );
  INV_X1 U10553 ( .A(n12087), .ZN(n8673) );
  AOI22_X1 U10554 ( .A1(n8673), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n12082), 
        .B2(P3_REG1_REG_22__SCAN_IN), .ZN(n8248) );
  NAND2_X1 U10555 ( .A1(n12083), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8247) );
  NAND2_X1 U10556 ( .A1(n8305), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8254) );
  OR2_X1 U10557 ( .A1(n8376), .A2(n10472), .ZN(n8250) );
  NAND2_X1 U10558 ( .A1(n8264), .A2(n8250), .ZN(n10721) );
  NAND2_X1 U10559 ( .A1(n8484), .A2(n10721), .ZN(n8253) );
  NAND2_X1 U10560 ( .A1(n12082), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8252) );
  INV_X1 U10561 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10720) );
  OR2_X1 U10562 ( .A1(n12087), .A2(n10720), .ZN(n8251) );
  XNOR2_X1 U10563 ( .A(n8256), .B(n7165), .ZN(n9520) );
  NAND2_X1 U10564 ( .A1(n8353), .A2(n9520), .ZN(n8263) );
  OR2_X1 U10565 ( .A1(n9361), .A2(SI_5_), .ZN(n8262) );
  NOR2_X1 U10566 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8258) );
  AND2_X1 U10567 ( .A1(n10322), .A2(n8258), .ZN(n8385) );
  OR2_X1 U10568 ( .A1(n8387), .A2(n8723), .ZN(n8260) );
  XNOR2_X1 U10569 ( .A(n8272), .B(n8260), .ZN(n10648) );
  OR2_X1 U10570 ( .A1(n10307), .A2(n14661), .ZN(n8261) );
  INV_X1 U10571 ( .A(n10722), .ZN(n14794) );
  NAND2_X1 U10572 ( .A1(n10926), .A2(n14794), .ZN(n10909) );
  INV_X1 U10573 ( .A(n10909), .ZN(n8322) );
  NAND2_X1 U10574 ( .A1(n8305), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8269) );
  NAND2_X1 U10575 ( .A1(n8264), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8265) );
  NAND2_X1 U10576 ( .A1(n8278), .A2(n8265), .ZN(n10941) );
  NAND2_X1 U10577 ( .A1(n8484), .A2(n10941), .ZN(n8268) );
  NAND2_X1 U10578 ( .A1(n12082), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8267) );
  INV_X1 U10579 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10929) );
  OR2_X1 U10580 ( .A1(n12087), .A2(n10929), .ZN(n8266) );
  INV_X1 U10581 ( .A(SI_6_), .ZN(n9509) );
  XNOR2_X1 U10582 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8270) );
  XNOR2_X1 U10583 ( .A(n8271), .B(n8270), .ZN(n9508) );
  NAND2_X1 U10584 ( .A1(n8353), .A2(n9508), .ZN(n8277) );
  NAND2_X1 U10585 ( .A1(n8387), .A2(n8272), .ZN(n8274) );
  NAND2_X1 U10586 ( .A1(n8274), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8273) );
  MUX2_X1 U10587 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8273), .S(
        P3_IR_REG_6__SCAN_IN), .Z(n8275) );
  NAND2_X1 U10588 ( .A1(n8275), .A2(n8300), .ZN(n10637) );
  OR2_X1 U10589 ( .A1(n10307), .A2(n10637), .ZN(n8276) );
  OAI211_X1 U10590 ( .C1(n9361), .C2(n9509), .A(n8277), .B(n8276), .ZN(n10933)
         );
  NAND2_X1 U10591 ( .A1(n10818), .A2(n10933), .ZN(n12197) );
  INV_X1 U10592 ( .A(n10818), .ZN(n12554) );
  INV_X1 U10593 ( .A(n10933), .ZN(n14799) );
  NAND2_X1 U10594 ( .A1(n12554), .A2(n14799), .ZN(n12196) );
  AND2_X1 U10595 ( .A1(n8278), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8279) );
  OR2_X1 U10596 ( .A1(n8279), .A2(n8291), .ZN(n10918) );
  NAND2_X1 U10597 ( .A1(n8344), .A2(n10918), .ZN(n8283) );
  NAND2_X1 U10598 ( .A1(n12083), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8282) );
  INV_X1 U10599 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10612) );
  OR2_X1 U10600 ( .A1(n8345), .A2(n10612), .ZN(n8281) );
  XNOR2_X1 U10601 ( .A(n8285), .B(n8284), .ZN(n9516) );
  NAND2_X1 U10602 ( .A1(n8353), .A2(n9516), .ZN(n8289) );
  NAND2_X1 U10603 ( .A1(n8300), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8287) );
  INV_X1 U10604 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8286) );
  XNOR2_X1 U10605 ( .A(n8287), .B(n8286), .ZN(n14697) );
  INV_X1 U10606 ( .A(n14697), .ZN(n10613) );
  OR2_X1 U10607 ( .A1(n10307), .A2(n10613), .ZN(n8288) );
  OAI211_X1 U10608 ( .C1(n9361), .C2(SI_7_), .A(n8289), .B(n8288), .ZN(n12201)
         );
  XNOR2_X1 U10609 ( .A(n12553), .B(n12201), .ZN(n10914) );
  INV_X1 U10610 ( .A(n10914), .ZN(n12199) );
  NAND2_X1 U10611 ( .A1(n8305), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8296) );
  NOR2_X1 U10612 ( .A1(n8291), .A2(n8290), .ZN(n8292) );
  OR2_X1 U10613 ( .A1(n8306), .A2(n8292), .ZN(n11061) );
  NAND2_X1 U10614 ( .A1(n8484), .A2(n11061), .ZN(n8295) );
  NAND2_X1 U10615 ( .A1(n12082), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8294) );
  INV_X1 U10616 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10618) );
  OR2_X1 U10617 ( .A1(n12087), .A2(n10618), .ZN(n8293) );
  INV_X1 U10618 ( .A(n8297), .ZN(n8298) );
  XNOR2_X1 U10619 ( .A(n8299), .B(n8298), .ZN(n9522) );
  NAND2_X1 U10620 ( .A1(n8353), .A2(n9522), .ZN(n8304) );
  OAI21_X1 U10621 ( .B1(n8300), .B2(P3_IR_REG_7__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8301) );
  XNOR2_X1 U10622 ( .A(n8301), .B(P3_IR_REG_8__SCAN_IN), .ZN(n14719) );
  OR2_X1 U10623 ( .A1(n10307), .A2(n10636), .ZN(n8303) );
  INV_X1 U10624 ( .A(SI_8_), .ZN(n9524) );
  OR2_X1 U10625 ( .A1(n9361), .A2(n9524), .ZN(n8302) );
  AND2_X1 U10626 ( .A1(n12207), .A2(n14815), .ZN(n11108) );
  INV_X1 U10627 ( .A(n11105), .ZN(n8320) );
  NAND2_X1 U10628 ( .A1(n8305), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8311) );
  OR2_X1 U10629 ( .A1(n8306), .A2(n10836), .ZN(n8307) );
  NAND2_X1 U10630 ( .A1(n8401), .A2(n8307), .ZN(n11119) );
  NAND2_X1 U10631 ( .A1(n8484), .A2(n11119), .ZN(n8310) );
  NAND2_X1 U10632 ( .A1(n12082), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8309) );
  INV_X1 U10633 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10624) );
  OR2_X1 U10634 ( .A1(n12087), .A2(n10624), .ZN(n8308) );
  XNOR2_X1 U10635 ( .A(n8313), .B(n8312), .ZN(n9525) );
  NAND2_X1 U10636 ( .A1(n8353), .A2(n9525), .ZN(n8319) );
  OR2_X1 U10637 ( .A1(n12096), .A2(SI_9_), .ZN(n8318) );
  NAND2_X1 U10638 ( .A1(n8314), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8316) );
  INV_X1 U10639 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8315) );
  XNOR2_X1 U10640 ( .A(n8316), .B(n8315), .ZN(n14739) );
  INV_X1 U10641 ( .A(n14739), .ZN(n10625) );
  OR2_X1 U10642 ( .A1(n10307), .A2(n10625), .ZN(n8317) );
  NAND2_X1 U10643 ( .A1(n11057), .A2(n10838), .ZN(n12213) );
  INV_X1 U10644 ( .A(n11057), .ZN(n12550) );
  INV_X1 U10645 ( .A(n10838), .ZN(n14820) );
  NAND2_X1 U10646 ( .A1(n12550), .A2(n14820), .ZN(n12214) );
  NAND2_X1 U10647 ( .A1(n12213), .A2(n12214), .ZN(n11113) );
  NAND2_X1 U10648 ( .A1(n8320), .A2(n11113), .ZN(n8321) );
  NOR2_X1 U10649 ( .A1(n8322), .A2(n8321), .ZN(n8398) );
  XNOR2_X1 U10650 ( .A(n8323), .B(n8338), .ZN(n9500) );
  INV_X1 U10651 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8324) );
  XNOR2_X1 U10652 ( .A(n8325), .B(n8324), .ZN(n10491) );
  OR2_X1 U10653 ( .A1(n10307), .A2(n10491), .ZN(n8326) );
  NAND2_X1 U10654 ( .A1(n8344), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8331) );
  INV_X1 U10655 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n14776) );
  OR2_X1 U10656 ( .A1(n8327), .A2(n14776), .ZN(n8333) );
  INV_X1 U10657 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n8328) );
  OR2_X1 U10658 ( .A1(n8676), .A2(n8328), .ZN(n8332) );
  INV_X1 U10659 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n8329) );
  NAND4_X1 U10660 ( .A1(n8331), .A2(n8333), .A3(n8332), .A4(n8330), .ZN(n12557) );
  NAND2_X1 U10661 ( .A1(n8305), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8337) );
  INV_X1 U10662 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n14605) );
  NAND2_X1 U10663 ( .A1(n8344), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8334) );
  INV_X1 U10664 ( .A(n8338), .ZN(n8340) );
  INV_X1 U10665 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8838) );
  NAND2_X1 U10666 ( .A1(n8838), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8339) );
  NAND2_X1 U10667 ( .A1(n8340), .A2(n8339), .ZN(n8341) );
  MUX2_X1 U10668 ( .A(SI_0_), .B(n8341), .S(n9504), .Z(n9498) );
  NAND2_X1 U10669 ( .A1(n9718), .A2(n12157), .ZN(n10202) );
  NAND2_X1 U10670 ( .A1(n9987), .A2(n10202), .ZN(n8343) );
  NAND2_X1 U10671 ( .A1(n8343), .A2(n9979), .ZN(n14759) );
  NAND2_X1 U10672 ( .A1(n6424), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8349) );
  NAND2_X1 U10673 ( .A1(n8344), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U10674 ( .A1(n8305), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8347) );
  INV_X1 U10675 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10333) );
  OR2_X1 U10676 ( .A1(n8345), .A2(n10333), .ZN(n8346) );
  INV_X1 U10677 ( .A(n8350), .ZN(n8351) );
  XNOR2_X1 U10678 ( .A(n8352), .B(n8351), .ZN(n9514) );
  NAND2_X1 U10679 ( .A1(n8353), .A2(n9514), .ZN(n8357) );
  OR2_X1 U10680 ( .A1(n12096), .A2(SI_2_), .ZN(n8356) );
  OR2_X1 U10681 ( .A1(n10307), .A2(n10334), .ZN(n8355) );
  NAND2_X1 U10682 ( .A1(n8358), .A2(n10056), .ZN(n12174) );
  INV_X1 U10683 ( .A(n10056), .ZN(n14754) );
  NAND2_X1 U10684 ( .A1(n14759), .A2(n12116), .ZN(n8360) );
  NAND2_X1 U10685 ( .A1(n8358), .A2(n14754), .ZN(n8359) );
  INV_X1 U10686 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n14786) );
  OR2_X1 U10687 ( .A1(n8327), .A2(n14786), .ZN(n8365) );
  INV_X1 U10688 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n8361) );
  NAND2_X1 U10689 ( .A1(n8484), .A2(n8361), .ZN(n8364) );
  NAND2_X1 U10690 ( .A1(n12082), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8363) );
  INV_X1 U10691 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10595) );
  OR2_X1 U10692 ( .A1(n12087), .A2(n10595), .ZN(n8362) );
  AND4_X2 U10693 ( .A1(n8365), .A2(n8364), .A3(n8363), .A4(n8362), .ZN(n14761)
         );
  INV_X1 U10694 ( .A(n8366), .ZN(n8367) );
  XNOR2_X1 U10695 ( .A(n8368), .B(n8367), .ZN(n9512) );
  NAND2_X1 U10696 ( .A1(n8353), .A2(n9512), .ZN(n8374) );
  OR2_X1 U10697 ( .A1(n12096), .A2(SI_3_), .ZN(n8373) );
  NAND2_X1 U10698 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n8370), .ZN(n8371) );
  XNOR2_X1 U10699 ( .A(n8369), .B(n8371), .ZN(n10644) );
  INV_X1 U10700 ( .A(n10644), .ZN(n14627) );
  OR2_X1 U10701 ( .A1(n10307), .A2(n14627), .ZN(n8372) );
  NAND2_X1 U10702 ( .A1(n14761), .A2(n10057), .ZN(n12176) );
  INV_X2 U10703 ( .A(n14761), .ZN(n12556) );
  INV_X1 U10704 ( .A(n10057), .ZN(n14782) );
  AND2_X2 U10705 ( .A1(n12176), .A2(n12179), .ZN(n12118) );
  NAND2_X1 U10706 ( .A1(n12556), .A2(n10057), .ZN(n8375) );
  INV_X1 U10707 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10730) );
  OR2_X1 U10708 ( .A1(n12087), .A2(n10730), .ZN(n8381) );
  NAND2_X1 U10709 ( .A1(n12083), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8380) );
  AND2_X1 U10710 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8377) );
  OR2_X1 U10711 ( .A1(n8377), .A2(n8376), .ZN(n10731) );
  NAND2_X1 U10712 ( .A1(n8484), .A2(n10731), .ZN(n8379) );
  NAND2_X1 U10713 ( .A1(n12082), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8378) );
  INV_X1 U10714 ( .A(n8382), .ZN(n8383) );
  XNOR2_X1 U10715 ( .A(n8384), .B(n8383), .ZN(n9518) );
  NAND2_X1 U10716 ( .A1(n8353), .A2(n9518), .ZN(n8390) );
  NOR2_X1 U10717 ( .A1(n8385), .A2(n8723), .ZN(n8386) );
  MUX2_X1 U10718 ( .A(n8723), .B(n8386), .S(P3_IR_REG_4__SCAN_IN), .Z(n8388)
         );
  OR2_X1 U10719 ( .A1(n10307), .A2(n14647), .ZN(n8389) );
  OAI211_X1 U10720 ( .C1(n9361), .C2(SI_4_), .A(n8390), .B(n8389), .ZN(n12182)
         );
  XNOR2_X1 U10721 ( .A(n12181), .B(n12182), .ZN(n12121) );
  INV_X1 U10722 ( .A(n12182), .ZN(n14791) );
  NAND2_X1 U10723 ( .A1(n12181), .A2(n14791), .ZN(n8391) );
  NAND2_X1 U10724 ( .A1(n10926), .A2(n10722), .ZN(n12190) );
  INV_X1 U10725 ( .A(n10926), .ZN(n12555) );
  NAND2_X1 U10726 ( .A1(n12555), .A2(n14794), .ZN(n12189) );
  INV_X1 U10727 ( .A(n12186), .ZN(n10716) );
  NAND2_X1 U10728 ( .A1(n10717), .A2(n10716), .ZN(n10715) );
  INV_X1 U10729 ( .A(n12201), .ZN(n14811) );
  NAND2_X1 U10730 ( .A1(n12553), .A2(n14811), .ZN(n8392) );
  NAND2_X1 U10731 ( .A1(n12554), .A2(n10933), .ZN(n10910) );
  OR2_X1 U10732 ( .A1(n12199), .A2(n10910), .ZN(n10912) );
  AND2_X1 U10733 ( .A1(n8392), .A2(n10912), .ZN(n11107) );
  INV_X1 U10734 ( .A(n11108), .ZN(n8393) );
  NAND2_X1 U10735 ( .A1(n8393), .A2(n11113), .ZN(n8394) );
  OR2_X1 U10736 ( .A1(n11107), .A2(n8394), .ZN(n8397) );
  INV_X1 U10737 ( .A(n11113), .ZN(n8395) );
  NAND2_X1 U10738 ( .A1(n12551), .A2(n12208), .ZN(n11109) );
  OR2_X1 U10739 ( .A1(n8395), .A2(n11109), .ZN(n8396) );
  AOI21_X1 U10740 ( .B1(n8398), .B2(n10715), .A(n7335), .ZN(n8400) );
  NAND2_X1 U10741 ( .A1(n12550), .A2(n10838), .ZN(n8399) );
  NAND2_X1 U10742 ( .A1(n8400), .A2(n8399), .ZN(n11031) );
  NAND2_X1 U10743 ( .A1(n12083), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8406) );
  NAND2_X1 U10744 ( .A1(n12082), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8405) );
  NAND2_X1 U10745 ( .A1(n8401), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U10746 ( .A1(n8415), .A2(n8402), .ZN(n10957) );
  NAND2_X1 U10747 ( .A1(n8484), .A2(n10957), .ZN(n8404) );
  INV_X1 U10748 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10629) );
  OR2_X1 U10749 ( .A1(n12087), .A2(n10629), .ZN(n8403) );
  XNOR2_X1 U10750 ( .A(n8408), .B(n8407), .ZN(n14030) );
  NAND2_X1 U10751 ( .A1(n8353), .A2(n14030), .ZN(n8413) );
  OR2_X1 U10752 ( .A1(n8409), .A2(n8723), .ZN(n8410) );
  XNOR2_X1 U10753 ( .A(n8410), .B(n8424), .ZN(n14033) );
  OR2_X1 U10754 ( .A1(n10307), .A2(n11198), .ZN(n8412) );
  OR2_X1 U10755 ( .A1(n9361), .A2(SI_10_), .ZN(n8411) );
  NAND2_X1 U10756 ( .A1(n11317), .A2(n10967), .ZN(n12218) );
  INV_X1 U10757 ( .A(n10967), .ZN(n14826) );
  NAND2_X1 U10758 ( .A1(n12549), .A2(n14826), .ZN(n12225) );
  NAND2_X1 U10759 ( .A1(n12218), .A2(n12225), .ZN(n11032) );
  AND2_X1 U10760 ( .A1(n12549), .A2(n10967), .ZN(n8414) );
  NAND2_X1 U10761 ( .A1(n12083), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8421) );
  AND2_X1 U10762 ( .A1(n8415), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8416) );
  OR2_X1 U10763 ( .A1(n8416), .A2(n8432), .ZN(n11321) );
  NAND2_X1 U10764 ( .A1(n8484), .A2(n11321), .ZN(n8420) );
  NAND2_X1 U10765 ( .A1(n12082), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8419) );
  INV_X1 U10766 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n8417) );
  OR2_X1 U10767 ( .A1(n12087), .A2(n8417), .ZN(n8418) );
  XNOR2_X1 U10768 ( .A(n8423), .B(n8422), .ZN(n9537) );
  NAND2_X1 U10769 ( .A1(n8353), .A2(n9537), .ZN(n8429) );
  OR2_X1 U10770 ( .A1(n9361), .A2(SI_11_), .ZN(n8428) );
  NAND2_X1 U10771 ( .A1(n8409), .A2(n8424), .ZN(n8438) );
  NAND2_X1 U10772 ( .A1(n8438), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8426) );
  XNOR2_X1 U10773 ( .A(n8426), .B(n8425), .ZN(n11302) );
  INV_X1 U10774 ( .A(n11302), .ZN(n11185) );
  OR2_X1 U10775 ( .A1(n10307), .A2(n11185), .ZN(n8427) );
  NAND2_X1 U10776 ( .A1(n12548), .A2(n14105), .ZN(n8430) );
  INV_X1 U10777 ( .A(n14105), .ZN(n11324) );
  NAND2_X1 U10778 ( .A1(n12083), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8437) );
  OR2_X1 U10779 ( .A1(n8432), .A2(n8431), .ZN(n8433) );
  NAND2_X1 U10780 ( .A1(n8466), .A2(n8433), .ZN(n11380) );
  NAND2_X1 U10781 ( .A1(n8484), .A2(n11380), .ZN(n8436) );
  NAND2_X1 U10782 ( .A1(n12082), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8435) );
  INV_X1 U10783 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11350) );
  OR2_X1 U10784 ( .A1(n12087), .A2(n11350), .ZN(n8434) );
  NAND2_X1 U10785 ( .A1(n8447), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8439) );
  XNOR2_X1 U10786 ( .A(n8439), .B(P3_IR_REG_12__SCAN_IN), .ZN(n11476) );
  OAI22_X1 U10787 ( .A1(n12096), .A2(n14938), .B1(n10307), .B2(n11469), .ZN(
        n8440) );
  INV_X1 U10788 ( .A(n8440), .ZN(n8445) );
  INV_X1 U10789 ( .A(n8441), .ZN(n8442) );
  XNOR2_X1 U10790 ( .A(n8443), .B(n8442), .ZN(n9550) );
  NAND2_X1 U10791 ( .A1(n9550), .A2(n8353), .ZN(n8444) );
  NAND2_X1 U10792 ( .A1(n8445), .A2(n8444), .ZN(n11385) );
  NAND2_X1 U10793 ( .A1(n11503), .A2(n11385), .ZN(n12233) );
  INV_X1 U10794 ( .A(n11385), .ZN(n14100) );
  NAND2_X1 U10795 ( .A1(n12547), .A2(n14100), .ZN(n12230) );
  NAND2_X1 U10796 ( .A1(n12233), .A2(n12230), .ZN(n11346) );
  XNOR2_X1 U10797 ( .A(n8446), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9575) );
  NAND2_X1 U10798 ( .A1(n9575), .A2(n8353), .ZN(n8451) );
  NOR2_X1 U10799 ( .A1(n8447), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n8460) );
  OR2_X1 U10800 ( .A1(n8460), .A2(n8723), .ZN(n8448) );
  INV_X1 U10801 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8459) );
  XNOR2_X1 U10802 ( .A(n8448), .B(n8459), .ZN(n11640) );
  INV_X1 U10803 ( .A(n11640), .ZN(n11626) );
  OAI22_X1 U10804 ( .A1(n12096), .A2(SI_13_), .B1(n11626), .B2(n10307), .ZN(
        n8449) );
  INV_X1 U10805 ( .A(n8449), .ZN(n8450) );
  NAND2_X1 U10806 ( .A1(n8451), .A2(n8450), .ZN(n14095) );
  INV_X1 U10807 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n8452) );
  OR2_X1 U10808 ( .A1(n12087), .A2(n8452), .ZN(n8456) );
  NAND2_X1 U10809 ( .A1(n12083), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8455) );
  XNOR2_X1 U10810 ( .A(n8466), .B(P3_REG3_REG_13__SCAN_IN), .ZN(n11506) );
  NAND2_X1 U10811 ( .A1(n8484), .A2(n11506), .ZN(n8454) );
  NAND2_X1 U10812 ( .A1(n12082), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8453) );
  NAND4_X1 U10813 ( .A1(n8456), .A2(n8455), .A3(n8454), .A4(n8453), .ZN(n12546) );
  OR2_X1 U10814 ( .A1(n14095), .A2(n12546), .ZN(n12236) );
  NAND2_X1 U10815 ( .A1(n14095), .A2(n12546), .ZN(n12235) );
  INV_X1 U10816 ( .A(n12546), .ZN(n11560) );
  NOR2_X1 U10817 ( .A1(n14095), .A2(n11560), .ZN(n11488) );
  XNOR2_X1 U10818 ( .A(n8458), .B(n8457), .ZN(n9587) );
  NAND2_X1 U10819 ( .A1(n9587), .A2(n8353), .ZN(n8465) );
  NAND2_X1 U10820 ( .A1(n8460), .A2(n8459), .ZN(n8477) );
  NAND2_X1 U10821 ( .A1(n8477), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8462) );
  INV_X1 U10822 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8461) );
  XNOR2_X1 U10823 ( .A(n8462), .B(n8461), .ZN(n12561) );
  INV_X1 U10824 ( .A(n12561), .ZN(n12565) );
  OAI22_X1 U10825 ( .A1(n12096), .A2(SI_14_), .B1(n12565), .B2(n10307), .ZN(
        n8463) );
  INV_X1 U10826 ( .A(n8463), .ZN(n8464) );
  INV_X1 U10827 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12564) );
  OR2_X1 U10828 ( .A1(n12087), .A2(n12564), .ZN(n8471) );
  NAND2_X1 U10829 ( .A1(n12083), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8470) );
  OAI21_X1 U10830 ( .B1(n8466), .B2(P3_REG3_REG_13__SCAN_IN), .A(
        P3_REG3_REG_14__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U10831 ( .A1(n8467), .A2(n8482), .ZN(n11566) );
  NAND2_X1 U10832 ( .A1(n8344), .A2(n11566), .ZN(n8469) );
  NAND2_X1 U10833 ( .A1(n12082), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8468) );
  NAND4_X1 U10834 ( .A1(n8471), .A2(n8470), .A3(n8469), .A4(n8468), .ZN(n12545) );
  OR2_X1 U10835 ( .A1(n11624), .A2(n12545), .ZN(n12241) );
  NAND2_X1 U10836 ( .A1(n11624), .A2(n12545), .ZN(n12240) );
  NAND2_X1 U10837 ( .A1(n12241), .A2(n12240), .ZN(n12234) );
  INV_X1 U10838 ( .A(n11624), .ZN(n8472) );
  NAND2_X1 U10839 ( .A1(n8472), .A2(n12545), .ZN(n8473) );
  NAND2_X1 U10840 ( .A1(n11490), .A2(n8473), .ZN(n11600) );
  INV_X1 U10841 ( .A(n8474), .ZN(n8475) );
  XNOR2_X1 U10842 ( .A(n8476), .B(n8475), .ZN(n9629) );
  NAND2_X1 U10843 ( .A1(n9629), .A2(n8353), .ZN(n8481) );
  OAI21_X1 U10844 ( .B1(n8477), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8478) );
  XNOR2_X1 U10845 ( .A(n8478), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12605) );
  OAI22_X1 U10846 ( .A1(n12096), .A2(n9631), .B1(n10307), .B2(n12593), .ZN(
        n8479) );
  INV_X1 U10847 ( .A(n8479), .ZN(n8480) );
  NAND2_X1 U10848 ( .A1(n8481), .A2(n8480), .ZN(n12246) );
  NAND2_X1 U10849 ( .A1(n12083), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8488) );
  AND2_X1 U10850 ( .A1(n8482), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8483) );
  OR2_X1 U10851 ( .A1(n8483), .A2(n8497), .ZN(n11679) );
  NAND2_X1 U10852 ( .A1(n8484), .A2(n11679), .ZN(n8487) );
  NAND2_X1 U10853 ( .A1(n12082), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8486) );
  INV_X1 U10854 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12560) );
  OR2_X1 U10855 ( .A1(n12087), .A2(n12560), .ZN(n8485) );
  XNOR2_X1 U10856 ( .A(n12246), .B(n12247), .ZN(n11599) );
  INV_X1 U10857 ( .A(n8489), .ZN(n8490) );
  XNOR2_X1 U10858 ( .A(n8491), .B(n8490), .ZN(n9785) );
  NAND2_X1 U10859 ( .A1(n9785), .A2(n8353), .ZN(n8496) );
  OR2_X1 U10860 ( .A1(n8492), .A2(n8723), .ZN(n8493) );
  XNOR2_X1 U10861 ( .A(n8493), .B(P3_IR_REG_16__SCAN_IN), .ZN(n14054) );
  OAI22_X1 U10862 ( .A1(n12096), .A2(n9787), .B1(n10307), .B2(n12609), .ZN(
        n8494) );
  INV_X1 U10863 ( .A(n8494), .ZN(n8495) );
  INV_X1 U10864 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12585) );
  OR2_X1 U10865 ( .A1(n12087), .A2(n12585), .ZN(n8502) );
  NAND2_X1 U10866 ( .A1(n12083), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8501) );
  NOR2_X1 U10867 ( .A1(n8497), .A2(n11816), .ZN(n8498) );
  OR2_X1 U10868 ( .A1(n8515), .A2(n8498), .ZN(n11819) );
  NAND2_X1 U10869 ( .A1(n8344), .A2(n11819), .ZN(n8500) );
  NAND2_X1 U10870 ( .A1(n12082), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8499) );
  NAND4_X1 U10871 ( .A1(n8502), .A2(n8501), .A3(n8500), .A4(n8499), .ZN(n12544) );
  INV_X1 U10872 ( .A(n8504), .ZN(n8505) );
  XNOR2_X1 U10873 ( .A(n8506), .B(n8505), .ZN(n14023) );
  NAND2_X1 U10874 ( .A1(n14023), .A2(n8353), .ZN(n8514) );
  NAND2_X1 U10875 ( .A1(n8507), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8508) );
  MUX2_X1 U10876 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8508), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n8510) );
  AND2_X1 U10877 ( .A1(n8510), .A2(n8540), .ZN(n14071) );
  OAI22_X1 U10878 ( .A1(n12096), .A2(n8511), .B1(n10307), .B2(n14025), .ZN(
        n8512) );
  INV_X1 U10879 ( .A(n8512), .ZN(n8513) );
  NAND2_X1 U10880 ( .A1(n12083), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8520) );
  OR2_X1 U10881 ( .A1(n8515), .A2(n12477), .ZN(n8516) );
  NAND2_X1 U10882 ( .A1(n8531), .A2(n8516), .ZN(n12481) );
  NAND2_X1 U10883 ( .A1(n8344), .A2(n12481), .ZN(n8519) );
  NAND2_X1 U10884 ( .A1(n12082), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8518) );
  INV_X1 U10885 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14082) );
  OR2_X1 U10886 ( .A1(n12087), .A2(n14082), .ZN(n8517) );
  OR2_X1 U10887 ( .A1(n12385), .A2(n12386), .ZN(n12149) );
  NAND2_X1 U10888 ( .A1(n12385), .A2(n12386), .ZN(n12148) );
  NAND2_X1 U10889 ( .A1(n12149), .A2(n12148), .ZN(n12126) );
  INV_X1 U10890 ( .A(n8522), .ZN(n8523) );
  XNOR2_X1 U10891 ( .A(n8524), .B(n8523), .ZN(n14039) );
  NAND2_X1 U10892 ( .A1(n14039), .A2(n8353), .ZN(n8530) );
  INV_X1 U10893 ( .A(SI_18_), .ZN(n8527) );
  NAND2_X1 U10894 ( .A1(n8540), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8526) );
  INV_X1 U10895 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8525) );
  XNOR2_X1 U10896 ( .A(n8526), .B(n8525), .ZN(n14041) );
  OAI22_X1 U10897 ( .A1(n12096), .A2(n8527), .B1(n10307), .B2(n14041), .ZN(
        n8528) );
  INV_X1 U10898 ( .A(n8528), .ZN(n8529) );
  NAND2_X1 U10899 ( .A1(n12083), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8536) );
  NAND2_X1 U10900 ( .A1(n12082), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8535) );
  NAND2_X1 U10901 ( .A1(n8531), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8532) );
  NAND2_X1 U10902 ( .A1(n8546), .A2(n8532), .ZN(n12769) );
  NAND2_X1 U10903 ( .A1(n8344), .A2(n12769), .ZN(n8534) );
  INV_X1 U10904 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12771) );
  OR2_X1 U10905 ( .A1(n12087), .A2(n12771), .ZN(n8533) );
  NAND2_X1 U10906 ( .A1(n12774), .A2(n12478), .ZN(n12151) );
  NAND2_X1 U10907 ( .A1(n12150), .A2(n12151), .ZN(n12777) );
  NAND2_X1 U10908 ( .A1(n12762), .A2(n12777), .ZN(n12761) );
  XNOR2_X1 U10909 ( .A(n8539), .B(n8538), .ZN(n10045) );
  NAND2_X1 U10910 ( .A1(n10045), .A2(n8353), .ZN(n8545) );
  INV_X1 U10911 ( .A(n8659), .ZN(n8541) );
  NAND2_X1 U10912 ( .A1(n8541), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8542) );
  XNOR2_X2 U10913 ( .A(n8542), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12623) );
  OAI22_X1 U10914 ( .A1(n12096), .A2(SI_19_), .B1(n12623), .B2(n10307), .ZN(
        n8543) );
  INV_X1 U10915 ( .A(n8543), .ZN(n8544) );
  NAND2_X1 U10916 ( .A1(n12083), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8552) );
  NAND2_X1 U10917 ( .A1(n12082), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8551) );
  AND2_X1 U10918 ( .A1(n8546), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8547) );
  OR2_X1 U10919 ( .A1(n8547), .A2(n8556), .ZN(n12754) );
  NAND2_X1 U10920 ( .A1(n8344), .A2(n12754), .ZN(n8550) );
  INV_X1 U10921 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n8548) );
  OR2_X1 U10922 ( .A1(n12087), .A2(n8548), .ZN(n8549) );
  AND2_X1 U10923 ( .A1(n12857), .A2(n12514), .ZN(n12107) );
  OR2_X1 U10924 ( .A1(n12857), .A2(n12514), .ZN(n12108) );
  XNOR2_X1 U10925 ( .A(n8553), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U10926 ( .A1(n10452), .A2(n8353), .ZN(n8555) );
  OR2_X1 U10927 ( .A1(n9361), .A2(n10453), .ZN(n8554) );
  NOR2_X1 U10928 ( .A1(n8556), .A2(n14920), .ZN(n8557) );
  OR2_X1 U10929 ( .A1(n8569), .A2(n8557), .ZN(n12744) );
  NAND2_X1 U10930 ( .A1(n12744), .A2(n8484), .ZN(n8562) );
  INV_X1 U10931 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n8558) );
  OR2_X1 U10932 ( .A1(n12087), .A2(n8558), .ZN(n8561) );
  NAND2_X1 U10933 ( .A1(n12083), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8560) );
  NAND2_X1 U10934 ( .A1(n12082), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8559) );
  NAND4_X1 U10935 ( .A1(n8562), .A2(n8561), .A3(n8560), .A4(n8559), .ZN(n12542) );
  NAND2_X1 U10936 ( .A1(n12853), .A2(n12542), .ZN(n12147) );
  INV_X1 U10937 ( .A(n12853), .ZN(n8563) );
  NAND2_X1 U10938 ( .A1(n8563), .A2(n12394), .ZN(n12146) );
  NAND2_X1 U10939 ( .A1(n12147), .A2(n12146), .ZN(n12738) );
  NAND2_X1 U10940 ( .A1(n12739), .A2(n12738), .ZN(n12737) );
  NAND2_X1 U10941 ( .A1(n12737), .A2(n7345), .ZN(n12727) );
  INV_X1 U10942 ( .A(n8564), .ZN(n8565) );
  XNOR2_X1 U10943 ( .A(n8566), .B(n8565), .ZN(n10533) );
  NAND2_X1 U10944 ( .A1(n10533), .A2(n8353), .ZN(n8568) );
  INV_X1 U10945 ( .A(SI_21_), .ZN(n10534) );
  OR2_X1 U10946 ( .A1(n9361), .A2(n10534), .ZN(n8567) );
  INV_X1 U10947 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12807) );
  OR2_X1 U10948 ( .A1(n8569), .A2(n12458), .ZN(n8570) );
  NAND2_X1 U10949 ( .A1(n8571), .A2(n8570), .ZN(n12732) );
  NAND2_X1 U10950 ( .A1(n12732), .A2(n8484), .ZN(n8576) );
  NAND2_X1 U10951 ( .A1(n12083), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8574) );
  INV_X1 U10952 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n8572) );
  OR2_X1 U10953 ( .A1(n12087), .A2(n8572), .ZN(n8573) );
  AND2_X1 U10954 ( .A1(n8574), .A2(n8573), .ZN(n8575) );
  OAI211_X1 U10955 ( .C1(n8676), .C2(n12807), .A(n8576), .B(n8575), .ZN(n12541) );
  AND2_X1 U10956 ( .A1(n12460), .A2(n12541), .ZN(n12110) );
  OR2_X1 U10957 ( .A1(n12460), .A2(n12541), .ZN(n12111) );
  INV_X1 U10958 ( .A(n8577), .ZN(n8578) );
  AOI22_X1 U10959 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_23__SCAN_IN), .B1(n11442), .B2(n14852), .ZN(n8589) );
  XNOR2_X1 U10960 ( .A(n8590), .B(n8589), .ZN(n11101) );
  NAND2_X1 U10961 ( .A1(n11101), .A2(n8353), .ZN(n8582) );
  OR2_X1 U10962 ( .A1(n9361), .A2(n11103), .ZN(n8581) );
  NAND2_X1 U10963 ( .A1(n8583), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8584) );
  NAND2_X1 U10964 ( .A1(n8594), .A2(n8584), .ZN(n12712) );
  NAND2_X1 U10965 ( .A1(n12712), .A2(n8484), .ZN(n8587) );
  AOI22_X1 U10966 ( .A1(n8673), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n12083), 
        .B2(P3_REG0_REG_23__SCAN_IN), .ZN(n8586) );
  NAND2_X1 U10967 ( .A1(n12082), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8585) );
  NAND2_X1 U10968 ( .A1(n12842), .A2(n12487), .ZN(n8588) );
  INV_X1 U10969 ( .A(n12842), .ZN(n12432) );
  NAND2_X1 U10970 ( .A1(n12432), .A2(n12539), .ZN(n12694) );
  NAND2_X1 U10971 ( .A1(n8588), .A2(n12694), .ZN(n12142) );
  INV_X1 U10972 ( .A(n12694), .ZN(n8602) );
  INV_X1 U10973 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11537) );
  NAND2_X1 U10974 ( .A1(n11442), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8591) );
  XNOR2_X1 U10975 ( .A(n14948), .B(n8604), .ZN(n8603) );
  XOR2_X1 U10976 ( .A(n11537), .B(n8603), .Z(n11465) );
  NAND2_X1 U10977 ( .A1(n11465), .A2(n8353), .ZN(n8593) );
  INV_X1 U10978 ( .A(SI_24_), .ZN(n11462) );
  OR2_X1 U10979 ( .A1(n12096), .A2(n11462), .ZN(n8592) );
  AND2_X1 U10980 ( .A1(n8594), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8595) );
  OR2_X1 U10981 ( .A1(n8595), .A2(n8611), .ZN(n12702) );
  NAND2_X1 U10982 ( .A1(n12702), .A2(n8344), .ZN(n8601) );
  INV_X1 U10983 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U10984 ( .A1(n12083), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U10985 ( .A1(n12082), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8596) );
  OAI211_X1 U10986 ( .C1(n8598), .C2(n12087), .A(n8597), .B(n8596), .ZN(n8599)
         );
  INV_X1 U10987 ( .A(n8599), .ZN(n8600) );
  NAND2_X1 U10988 ( .A1(n8601), .A2(n8600), .ZN(n12538) );
  INV_X1 U10989 ( .A(n12538), .ZN(n12407) );
  NAND2_X1 U10990 ( .A1(n12696), .A2(n7340), .ZN(n12683) );
  NAND2_X1 U10991 ( .A1(n8603), .A2(n11537), .ZN(n8606) );
  NAND2_X1 U10992 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n8604), .ZN(n8605) );
  AOI22_X1 U10993 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n11613), .B2(n11616), .ZN(n8607) );
  XNOR2_X1 U10994 ( .A(n8620), .B(n8607), .ZN(n11607) );
  NAND2_X1 U10995 ( .A1(n11607), .A2(n8353), .ZN(n8609) );
  OR2_X1 U10996 ( .A1(n9361), .A2(n11608), .ZN(n8608) );
  INV_X1 U10997 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8610) );
  NAND2_X1 U10998 ( .A1(n8611), .A2(n8610), .ZN(n8624) );
  OR2_X1 U10999 ( .A1(n8611), .A2(n8610), .ZN(n8612) );
  NAND2_X1 U11000 ( .A1(n8624), .A2(n8612), .ZN(n12689) );
  NAND2_X1 U11001 ( .A1(n12689), .A2(n8344), .ZN(n8617) );
  INV_X1 U11002 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n14849) );
  NAND2_X1 U11003 ( .A1(n8673), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8614) );
  NAND2_X1 U11004 ( .A1(n12082), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8613) );
  OAI211_X1 U11005 ( .C1(n8327), .C2(n14849), .A(n8614), .B(n8613), .ZN(n8615)
         );
  INV_X1 U11006 ( .A(n8615), .ZN(n8616) );
  NAND2_X1 U11007 ( .A1(n12469), .A2(n12670), .ZN(n12277) );
  NAND2_X1 U11008 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n11613), .ZN(n8619) );
  AOI22_X1 U11009 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n13442), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n6674), .ZN(n8621) );
  XNOR2_X1 U11010 ( .A(n8634), .B(n8621), .ZN(n11690) );
  NAND2_X1 U11011 ( .A1(n11690), .A2(n8353), .ZN(n8623) );
  NAND2_X1 U11012 ( .A1(n8624), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8625) );
  NAND2_X1 U11013 ( .A1(n8639), .A2(n8625), .ZN(n12675) );
  NAND2_X1 U11014 ( .A1(n12675), .A2(n8344), .ZN(n8631) );
  INV_X1 U11015 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U11016 ( .A1(n12083), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U11017 ( .A1(n12082), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8626) );
  OAI211_X1 U11018 ( .C1(n12087), .C2(n8628), .A(n8627), .B(n8626), .ZN(n8629)
         );
  INV_X1 U11019 ( .A(n8629), .ZN(n8630) );
  NOR2_X1 U11020 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n6674), .ZN(n8635) );
  AOI22_X1 U11021 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n14882), .B2(n11842), .ZN(n8636) );
  XNOR2_X1 U11022 ( .A(n8648), .B(n8636), .ZN(n12070) );
  NAND2_X1 U11023 ( .A1(n12070), .A2(n8353), .ZN(n8638) );
  INV_X1 U11024 ( .A(SI_27_), .ZN(n12071) );
  AND2_X1 U11025 ( .A1(n8639), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8640) );
  OR2_X1 U11026 ( .A1(n8640), .A2(n8653), .ZN(n12659) );
  NAND2_X1 U11027 ( .A1(n12659), .A2(n8344), .ZN(n8645) );
  INV_X1 U11028 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n12660) );
  NAND2_X1 U11029 ( .A1(n12082), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8642) );
  NAND2_X1 U11030 ( .A1(n12083), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8641) );
  OAI211_X1 U11031 ( .C1(n12087), .C2(n12660), .A(n8642), .B(n8641), .ZN(n8643) );
  INV_X1 U11032 ( .A(n8643), .ZN(n8644) );
  XNOR2_X1 U11033 ( .A(n12781), .B(n12536), .ZN(n12141) );
  INV_X1 U11034 ( .A(n12781), .ZN(n12279) );
  NAND2_X1 U11035 ( .A1(n12279), .A2(n12671), .ZN(n8647) );
  NAND2_X1 U11036 ( .A1(n12655), .A2(n8647), .ZN(n8670) );
  NAND2_X1 U11037 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n14882), .ZN(n8649) );
  AOI22_X1 U11038 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n13439), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n14011), .ZN(n8650) );
  XNOR2_X1 U11039 ( .A(n9358), .B(n8650), .ZN(n12878) );
  NAND2_X1 U11040 ( .A1(n12878), .A2(n8353), .ZN(n8652) );
  OR2_X1 U11041 ( .A1(n12096), .A2(n14863), .ZN(n8651) );
  INV_X1 U11042 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n12449) );
  NOR2_X1 U11043 ( .A1(n8653), .A2(n12449), .ZN(n8654) );
  INV_X1 U11044 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12647) );
  NAND2_X1 U11045 ( .A1(n12083), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8656) );
  NAND2_X1 U11046 ( .A1(n12082), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8655) );
  OAI211_X1 U11047 ( .C1(n12647), .C2(n12087), .A(n8656), .B(n8655), .ZN(n8657) );
  AOI21_X1 U11048 ( .B1(n12448), .B2(n8344), .A(n8657), .ZN(n12419) );
  NAND2_X1 U11049 ( .A1(n12652), .A2(n12419), .ZN(n12289) );
  NAND2_X1 U11050 ( .A1(n8713), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8661) );
  NAND2_X1 U11051 ( .A1(n12310), .A2(n12623), .ZN(n8758) );
  NAND2_X1 U11052 ( .A1(n8668), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8663) );
  XNOR2_X2 U11053 ( .A(n8663), .B(n8662), .ZN(n12163) );
  INV_X1 U11054 ( .A(n8664), .ZN(n8665) );
  NAND2_X1 U11055 ( .A1(n8665), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8667) );
  MUX2_X1 U11056 ( .A(n8667), .B(P3_IR_REG_31__SCAN_IN), .S(n8666), .Z(n8669)
         );
  NAND2_X1 U11057 ( .A1(n10207), .A2(n8757), .ZN(n12307) );
  AOI21_X1 U11058 ( .B1(n8670), .B2(n12445), .A(n14767), .ZN(n8684) );
  INV_X1 U11059 ( .A(n8670), .ZN(n8672) );
  INV_X1 U11060 ( .A(n12445), .ZN(n8671) );
  NAND2_X1 U11061 ( .A1(n8672), .A2(n8671), .ZN(n9357) );
  NAND2_X1 U11062 ( .A1(n12637), .A2(n8344), .ZN(n12090) );
  INV_X1 U11063 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8677) );
  NAND2_X1 U11064 ( .A1(n12083), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U11065 ( .A1(n8673), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8674) );
  OAI211_X1 U11066 ( .C1(n8677), .C2(n8676), .A(n8675), .B(n8674), .ZN(n8678)
         );
  INV_X1 U11067 ( .A(n8678), .ZN(n8679) );
  OR2_X1 U11068 ( .A1(n6630), .A2(n12073), .ZN(n10317) );
  NAND2_X1 U11069 ( .A1(n10307), .A2(n10317), .ZN(n8682) );
  OAI22_X1 U11070 ( .A1(n12451), .A2(n14760), .B1(n12671), .B2(n14762), .ZN(
        n8683) );
  AOI21_X1 U11071 ( .B1(n8684), .B2(n9357), .A(n8683), .ZN(n12654) );
  NOR2_X4 U11072 ( .A1(n9718), .A2(n10274), .ZN(n12164) );
  NAND2_X1 U11073 ( .A1(n12164), .A2(n12166), .ZN(n9985) );
  NAND2_X1 U11074 ( .A1(n9985), .A2(n12165), .ZN(n14753) );
  INV_X1 U11075 ( .A(n12116), .ZN(n14758) );
  NAND2_X1 U11076 ( .A1(n14753), .A2(n14758), .ZN(n14752) );
  NAND2_X1 U11077 ( .A1(n10444), .A2(n12118), .ZN(n8685) );
  NAND2_X1 U11078 ( .A1(n8685), .A2(n12176), .ZN(n10725) );
  INV_X1 U11079 ( .A(n12121), .ZN(n12178) );
  NAND2_X1 U11080 ( .A1(n10725), .A2(n12178), .ZN(n8687) );
  INV_X1 U11081 ( .A(n12181), .ZN(n12180) );
  NAND2_X1 U11082 ( .A1(n12180), .A2(n14791), .ZN(n8686) );
  NAND2_X1 U11083 ( .A1(n10714), .A2(n12186), .ZN(n8688) );
  INV_X1 U11084 ( .A(n12553), .ZN(n11058) );
  XNOR2_X1 U11085 ( .A(n12551), .B(n12208), .ZN(n12205) );
  NAND2_X1 U11086 ( .A1(n11012), .A2(n12205), .ZN(n8690) );
  NAND2_X1 U11087 ( .A1(n12207), .A2(n12208), .ZN(n8689) );
  NAND2_X1 U11088 ( .A1(n8691), .A2(n12218), .ZN(n11292) );
  NAND2_X1 U11089 ( .A1(n11315), .A2(n14105), .ZN(n12220) );
  NAND2_X1 U11090 ( .A1(n12548), .A2(n11324), .ZN(n12227) );
  NAND2_X1 U11091 ( .A1(n11292), .A2(n12226), .ZN(n8692) );
  INV_X1 U11092 ( .A(n11346), .ZN(n12124) );
  AND2_X1 U11093 ( .A1(n12124), .A2(n12235), .ZN(n11492) );
  INV_X1 U11094 ( .A(n12240), .ZN(n8696) );
  AND2_X1 U11095 ( .A1(n11492), .A2(n12240), .ZN(n8693) );
  NAND2_X1 U11096 ( .A1(n11345), .A2(n8693), .ZN(n8699) );
  INV_X1 U11097 ( .A(n12235), .ZN(n8695) );
  AND2_X1 U11098 ( .A1(n12236), .A2(n12233), .ZN(n8694) );
  NOR2_X1 U11099 ( .A1(n7341), .A2(n8697), .ZN(n8698) );
  NAND2_X1 U11100 ( .A1(n8699), .A2(n8698), .ZN(n11602) );
  NAND2_X1 U11101 ( .A1(n12246), .A2(n12247), .ZN(n12251) );
  XNOR2_X1 U11102 ( .A(n12254), .B(n12544), .ZN(n12127) );
  NAND2_X1 U11103 ( .A1(n12254), .A2(n12476), .ZN(n12252) );
  INV_X1 U11104 ( .A(n12126), .ZN(n12258) );
  NAND2_X1 U11105 ( .A1(n11801), .A2(n12258), .ZN(n8700) );
  NAND2_X1 U11106 ( .A1(n8700), .A2(n12148), .ZN(n12776) );
  INV_X1 U11107 ( .A(n12776), .ZN(n8701) );
  OR2_X1 U11108 ( .A1(n12857), .A2(n12766), .ZN(n12262) );
  NAND2_X1 U11109 ( .A1(n8702), .A2(n12262), .ZN(n12743) );
  NAND2_X1 U11110 ( .A1(n8703), .A2(n12147), .ZN(n12731) );
  INV_X1 U11111 ( .A(n12541), .ZN(n12396) );
  NOR2_X1 U11112 ( .A1(n12460), .A2(n12396), .ZN(n8704) );
  OAI21_X1 U11113 ( .B1(n12720), .B2(n12144), .A(n12143), .ZN(n12711) );
  NAND2_X1 U11114 ( .A1(n12842), .A2(n12539), .ZN(n12275) );
  NAND2_X1 U11115 ( .A1(n12491), .A2(n12407), .ZN(n12273) );
  INV_X1 U11116 ( .A(n12682), .ZN(n12687) );
  NAND2_X1 U11117 ( .A1(n12529), .A2(n12415), .ZN(n12283) );
  AND2_X1 U11118 ( .A1(n12781), .A2(n12671), .ZN(n12286) );
  OAI21_X1 U11119 ( .B1(n12161), .B2(n8757), .A(n12623), .ZN(n8706) );
  NAND2_X1 U11120 ( .A1(n8706), .A2(n12163), .ZN(n8709) );
  NAND2_X1 U11121 ( .A1(n12163), .A2(n10455), .ZN(n8707) );
  NAND2_X1 U11122 ( .A1(n12161), .A2(n8707), .ZN(n8708) );
  NAND2_X1 U11123 ( .A1(n8709), .A2(n8708), .ZN(n9991) );
  NAND2_X1 U11124 ( .A1(n12161), .A2(n12163), .ZN(n14827) );
  NAND2_X1 U11125 ( .A1(n10455), .A2(n12105), .ZN(n12309) );
  INV_X1 U11126 ( .A(n12309), .ZN(n12303) );
  AND2_X1 U11127 ( .A1(n14827), .A2(n12303), .ZN(n8710) );
  NAND2_X1 U11128 ( .A1(n9991), .A2(n8710), .ZN(n8712) );
  NOR2_X1 U11129 ( .A1(n10455), .A2(n12623), .ZN(n8711) );
  NAND2_X1 U11130 ( .A1(n12310), .A2(n8711), .ZN(n8747) );
  AND2_X1 U11131 ( .A1(n8712), .A2(n8747), .ZN(n14808) );
  INV_X1 U11132 ( .A(n12302), .ZN(n14756) );
  NAND2_X1 U11133 ( .A1(n12161), .A2(n14756), .ZN(n14821) );
  NOR2_X1 U11134 ( .A1(n8716), .A2(n8723), .ZN(n8717) );
  INV_X1 U11135 ( .A(n8718), .ZN(n8719) );
  INV_X1 U11136 ( .A(n11610), .ZN(n8726) );
  NAND2_X1 U11137 ( .A1(n8720), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8722) );
  INV_X1 U11138 ( .A(n11463), .ZN(n8725) );
  NAND3_X1 U11139 ( .A1(n8726), .A2(n8725), .A3(n8740), .ZN(n9964) );
  XNOR2_X1 U11140 ( .A(n11463), .B(P3_B_REG_SCAN_IN), .ZN(n8727) );
  NAND2_X1 U11141 ( .A1(n11610), .A2(n8727), .ZN(n8728) );
  NOR2_X1 U11142 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .ZN(
        n8732) );
  NOR4_X1 U11143 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n8731) );
  NOR4_X1 U11144 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8730) );
  NOR4_X1 U11145 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8729) );
  NAND4_X1 U11146 ( .A1(n8732), .A2(n8731), .A3(n8730), .A4(n8729), .ZN(n8738)
         );
  NOR4_X1 U11147 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8736) );
  NOR4_X1 U11148 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8735) );
  NOR4_X1 U11149 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8734) );
  NOR4_X1 U11150 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8733) );
  NAND4_X1 U11151 ( .A1(n8736), .A2(n8735), .A3(n8734), .A4(n8733), .ZN(n8737)
         );
  NOR2_X1 U11152 ( .A1(n8738), .A2(n8737), .ZN(n8739) );
  NOR2_X1 U11153 ( .A1(n9562), .A2(n8739), .ZN(n8759) );
  NOR2_X1 U11154 ( .A1(n12308), .A2(n8759), .ZN(n8746) );
  INV_X1 U11155 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9569) );
  NAND2_X1 U11156 ( .A1(n8742), .A2(n9569), .ZN(n8741) );
  NAND2_X1 U11157 ( .A1(n11693), .A2(n11610), .ZN(n9566) );
  INV_X1 U11158 ( .A(n10127), .ZN(n8744) );
  INV_X1 U11159 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9565) );
  NAND2_X1 U11160 ( .A1(n8742), .A2(n9565), .ZN(n8743) );
  NAND2_X1 U11161 ( .A1(n11693), .A2(n11463), .ZN(n9563) );
  NAND2_X1 U11162 ( .A1(n8744), .A2(n9975), .ZN(n8756) );
  INV_X1 U11163 ( .A(n9975), .ZN(n8745) );
  NAND2_X1 U11164 ( .A1(n8745), .A2(n10127), .ZN(n8760) );
  NAND2_X1 U11165 ( .A1(n12294), .A2(n8747), .ZN(n10126) );
  AND2_X1 U11166 ( .A1(n10129), .A2(n10126), .ZN(n8750) );
  OAI22_X1 U11167 ( .A1(n14827), .A2(n8757), .B1(n12623), .B2(n12161), .ZN(
        n8748) );
  AOI21_X1 U11168 ( .B1(n8748), .B2(n12309), .A(n12288), .ZN(n8749) );
  MUX2_X1 U11169 ( .A(n8750), .B(n8749), .S(n10127), .Z(n8751) );
  MUX2_X1 U11170 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n8764), .S(n14846), .Z(
        n8752) );
  INV_X1 U11171 ( .A(n8752), .ZN(n8755) );
  INV_X1 U11172 ( .A(n12826), .ZN(n8753) );
  NAND2_X1 U11173 ( .A1(n12652), .A2(n8753), .ZN(n8754) );
  NAND2_X1 U11174 ( .A1(n8755), .A2(n8754), .ZN(P3_U3487) );
  OR2_X1 U11175 ( .A1(n8756), .A2(n8759), .ZN(n10000) );
  NAND2_X1 U11176 ( .A1(n12163), .A2(n8757), .ZN(n12139) );
  OR2_X1 U11177 ( .A1(n12139), .A2(n8758), .ZN(n9992) );
  NAND2_X1 U11178 ( .A1(n12288), .A2(n12303), .ZN(n10133) );
  AND2_X1 U11179 ( .A1(n9992), .A2(n10133), .ZN(n8762) );
  INV_X1 U11180 ( .A(n9991), .ZN(n8761) );
  OAI22_X1 U11181 ( .A1(n10000), .A2(n8762), .B1(n9998), .B2(n8761), .ZN(n8763) );
  INV_X1 U11182 ( .A(n12865), .ZN(n8765) );
  NAND2_X1 U11183 ( .A1(n12652), .A2(n8765), .ZN(n8766) );
  NAND2_X1 U11184 ( .A1(n6535), .A2(n8766), .ZN(P3_U3455) );
  NOR2_X1 U11185 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n8768) );
  NOR2_X1 U11186 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), 
        .ZN(n8767) );
  OR2_X2 U11187 ( .A1(n8776), .A2(n6613), .ZN(n8773) );
  NAND2_X1 U11188 ( .A1(n8794), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8774) );
  INV_X1 U11189 ( .A(n8775), .ZN(n8777) );
  NOR2_X2 U11190 ( .A1(n8777), .A2(n8776), .ZN(n8782) );
  NAND2_X1 U11191 ( .A1(n8887), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n8909) );
  NOR2_X1 U11192 ( .A1(n8909), .A2(n8908), .ZN(n8928) );
  NAND2_X1 U11193 ( .A1(n8928), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8951) );
  OR2_X1 U11194 ( .A1(n8951), .A2(n8950), .ZN(n8962) );
  AND2_X1 U11195 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n8778) );
  INV_X1 U11196 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9035) );
  INV_X1 U11197 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9112) );
  NAND2_X1 U11198 ( .A1(n9128), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9156) );
  NAND2_X1 U11199 ( .A1(n9155), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9184) );
  NAND2_X1 U11200 ( .A1(n9171), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9199) );
  NAND2_X1 U11201 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n9183), .ZN(n9217) );
  INV_X1 U11202 ( .A(n9217), .ZN(n8779) );
  NAND2_X1 U11203 ( .A1(n8779), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9229) );
  INV_X1 U11204 ( .A(n9229), .ZN(n8780) );
  NAND2_X1 U11205 ( .A1(n8780), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9246) );
  INV_X1 U11206 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8781) );
  NOR2_X1 U11207 ( .A1(n9246), .A2(n8781), .ZN(n11883) );
  NAND2_X1 U11208 ( .A1(n6462), .A2(n11883), .ZN(n8787) );
  NAND2_X1 U11209 ( .A1(n6464), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8786) );
  NAND2_X1 U11210 ( .A1(n6466), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8785) );
  NAND2_X1 U11211 ( .A1(n9266), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8784) );
  AND4_X1 U11212 ( .A1(n8787), .A2(n8786), .A3(n8785), .A4(n8784), .ZN(n12372)
         );
  INV_X2 U11213 ( .A(n9270), .ZN(n9235) );
  NAND2_X1 U11214 ( .A1(n13433), .A2(n9262), .ZN(n8796) );
  NAND2_X1 U11215 ( .A1(n9271), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8795) );
  INV_X2 U11216 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8797) );
  XNOR2_X2 U11217 ( .A(n8814), .B(n8813), .ZN(n10556) );
  INV_X1 U11218 ( .A(n9076), .ZN(n8802) );
  NAND4_X1 U11219 ( .A1(n8813), .A2(n9101), .A3(n9085), .A4(n8797), .ZN(n8800)
         );
  INV_X1 U11220 ( .A(n8798), .ZN(n8799) );
  NAND2_X1 U11221 ( .A1(n8810), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8803) );
  MUX2_X1 U11222 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8803), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n8806) );
  NAND2_X1 U11223 ( .A1(n8806), .A2(n9334), .ZN(n9908) );
  XNOR2_X1 U11224 ( .A(n10556), .B(n9908), .ZN(n8818) );
  NAND2_X1 U11225 ( .A1(n6613), .A2(n6448), .ZN(n8809) );
  NAND2_X1 U11226 ( .A1(n8818), .A2(n12380), .ZN(n8817) );
  NAND2_X1 U11227 ( .A1(n8814), .A2(n8813), .ZN(n8815) );
  INV_X1 U11228 ( .A(n8818), .ZN(n9305) );
  INV_X1 U11229 ( .A(n11020), .ZN(n9302) );
  MUX2_X1 U11230 ( .A(n12372), .B(n13919), .S(n9238), .Z(n9257) );
  INV_X1 U11231 ( .A(n9257), .ZN(n9261) );
  NAND2_X1 U11232 ( .A1(n9539), .A2(n9235), .ZN(n8822) );
  INV_X1 U11233 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9542) );
  OR2_X1 U11234 ( .A1(n8916), .A2(n6613), .ZN(n8819) );
  XNOR2_X1 U11235 ( .A(n8915), .B(n8819), .ZN(n9609) );
  INV_X1 U11236 ( .A(n8820), .ZN(n8821) );
  OAI21_X1 U11237 ( .B1(n8887), .B2(P1_REG3_REG_5__SCAN_IN), .A(n8909), .ZN(
        n10547) );
  INV_X1 U11238 ( .A(n10547), .ZN(n10301) );
  NAND2_X1 U11239 ( .A1(n6462), .A2(n10301), .ZN(n8826) );
  NAND2_X1 U11240 ( .A1(n6425), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n8825) );
  NAND2_X1 U11241 ( .A1(n6465), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8824) );
  NAND2_X1 U11242 ( .A1(n8889), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8823) );
  MUX2_X1 U11243 ( .A(n10552), .B(n13594), .S(n9192), .Z(n8938) );
  INV_X1 U11244 ( .A(n9559), .ZN(n9053) );
  OR2_X1 U11245 ( .A1(n8828), .A2(n6613), .ZN(n8829) );
  NAND2_X1 U11246 ( .A1(n9053), .A2(n13623), .ZN(n8830) );
  NAND2_X1 U11247 ( .A1(n6425), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8833) );
  NAND2_X1 U11248 ( .A1(n8889), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8832) );
  NAND2_X1 U11249 ( .A1(n9274), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8831) );
  NAND2_X1 U11250 ( .A1(n9274), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8836) );
  NAND2_X1 U11251 ( .A1(n8888), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8835) );
  NAND2_X1 U11252 ( .A1(n8889), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8837) );
  NAND3_X2 U11253 ( .A1(n7337), .A2(n7338), .A3(n8837), .ZN(n13598) );
  INV_X1 U11254 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n13617) );
  NAND2_X1 U11255 ( .A1(n9504), .A2(SI_0_), .ZN(n8839) );
  NAND2_X1 U11256 ( .A1(n8839), .A2(n8838), .ZN(n8841) );
  NAND2_X1 U11257 ( .A1(n8841), .A2(n8840), .ZN(n14018) );
  MUX2_X1 U11258 ( .A(n13617), .B(n14018), .S(n9559), .Z(n8863) );
  INV_X1 U11259 ( .A(n8861), .ZN(n8860) );
  NAND2_X1 U11260 ( .A1(n9247), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8845) );
  NAND2_X1 U11261 ( .A1(n9274), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8843) );
  NAND2_X1 U11262 ( .A1(n6421), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8842) );
  BUF_X1 U11263 ( .A(n8846), .Z(n8847) );
  NOR2_X1 U11264 ( .A1(n9504), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8848) );
  NOR2_X1 U11265 ( .A1(n8847), .A2(n8848), .ZN(n8850) );
  NAND2_X1 U11266 ( .A1(n9506), .A2(n9504), .ZN(n8849) );
  NAND2_X1 U11267 ( .A1(n8850), .A2(n8849), .ZN(n8858) );
  INV_X1 U11268 ( .A(n9506), .ZN(n8851) );
  MUX2_X1 U11269 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8851), .S(n9505), .Z(n8852) );
  INV_X1 U11270 ( .A(n14009), .ZN(n9760) );
  NAND2_X1 U11271 ( .A1(n8852), .A2(n9760), .ZN(n8857) );
  NAND2_X1 U11272 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8853) );
  MUX2_X1 U11273 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8853), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n8855) );
  INV_X1 U11274 ( .A(n8828), .ZN(n8854) );
  INV_X1 U11275 ( .A(n13605), .ZN(n13602) );
  NAND3_X1 U11276 ( .A1(n8847), .A2(n13602), .A3(n14009), .ZN(n8856) );
  AND3_X2 U11277 ( .A1(n8858), .A2(n8857), .A3(n8856), .ZN(n14322) );
  INV_X1 U11278 ( .A(n14322), .ZN(n8859) );
  NAND2_X1 U11279 ( .A1(n8860), .A2(n9928), .ZN(n8862) );
  NAND2_X1 U11280 ( .A1(n9761), .A2(n14322), .ZN(n9284) );
  NAND2_X1 U11281 ( .A1(n8861), .A2(n9284), .ZN(n9929) );
  MUX2_X1 U11282 ( .A(n8862), .B(n9929), .S(n9238), .Z(n8867) );
  OAI21_X1 U11283 ( .B1(n13598), .B2(n10098), .A(n9926), .ZN(n9912) );
  INV_X1 U11284 ( .A(n9747), .ZN(n8864) );
  AND2_X1 U11285 ( .A1(n9912), .A2(n8864), .ZN(n8866) );
  MUX2_X1 U11286 ( .A(n9928), .B(n9284), .S(n9192), .Z(n8865) );
  OAI21_X1 U11287 ( .B1(n8867), .B2(n8866), .A(n8865), .ZN(n8869) );
  MUX2_X1 U11288 ( .A(n13597), .B(n13540), .S(n9192), .Z(n8868) );
  INV_X1 U11289 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8870) );
  NAND2_X1 U11290 ( .A1(n6463), .A2(n8870), .ZN(n8874) );
  NAND2_X1 U11291 ( .A1(n6425), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8873) );
  NAND2_X1 U11292 ( .A1(n8889), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8872) );
  NAND2_X1 U11293 ( .A1(n6465), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8871) );
  NAND4_X1 U11294 ( .A1(n8874), .A2(n8873), .A3(n8872), .A4(n8871), .ZN(n13596) );
  NAND2_X1 U11295 ( .A1(n9527), .A2(n9235), .ZN(n8881) );
  INV_X1 U11296 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9528) );
  NAND2_X1 U11297 ( .A1(n8875), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8876) );
  MUX2_X1 U11298 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8876), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n8878) );
  OAI22_X1 U11299 ( .A1(n6456), .A2(n9528), .B1(n9559), .B2(n9772), .ZN(n8879)
         );
  INV_X1 U11300 ( .A(n8879), .ZN(n8880) );
  NAND2_X1 U11301 ( .A1(n8881), .A2(n8880), .ZN(n14305) );
  NAND2_X1 U11302 ( .A1(n10175), .A2(n14305), .ZN(n10107) );
  NAND2_X1 U11303 ( .A1(n14328), .A2(n13596), .ZN(n8883) );
  NAND2_X1 U11304 ( .A1(n8882), .A2(n14298), .ZN(n8885) );
  MUX2_X1 U11305 ( .A(n8883), .B(n10107), .S(n9192), .Z(n8884) );
  NAND2_X1 U11306 ( .A1(n8885), .A2(n8884), .ZN(n8901) );
  NOR2_X1 U11307 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8886) );
  NOR2_X1 U11308 ( .A1(n8887), .A2(n8886), .ZN(n10462) );
  NAND2_X1 U11309 ( .A1(n6463), .A2(n10462), .ZN(n8892) );
  NAND2_X1 U11310 ( .A1(n6425), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8891) );
  NAND2_X1 U11311 ( .A1(n6466), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8890) );
  NAND2_X1 U11312 ( .A1(n9533), .A2(n9235), .ZN(n8898) );
  INV_X1 U11313 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9534) );
  NAND2_X1 U11314 ( .A1(n8877), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8894) );
  INV_X1 U11315 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8893) );
  XNOR2_X1 U11316 ( .A(n8894), .B(n8893), .ZN(n13640) );
  OAI22_X1 U11317 ( .A1(n8895), .A2(n9534), .B1(n9559), .B2(n13640), .ZN(n8896) );
  INV_X1 U11318 ( .A(n8896), .ZN(n8897) );
  NAND2_X2 U11319 ( .A1(n8898), .A2(n8897), .ZN(n14335) );
  MUX2_X1 U11320 ( .A(n13595), .B(n14335), .S(n9192), .Z(n8902) );
  NAND2_X1 U11321 ( .A1(n8901), .A2(n8902), .ZN(n8900) );
  MUX2_X1 U11322 ( .A(n14335), .B(n13595), .S(n9192), .Z(n8899) );
  NAND2_X1 U11323 ( .A1(n8900), .A2(n8899), .ZN(n8906) );
  INV_X1 U11324 ( .A(n8901), .ZN(n8904) );
  INV_X1 U11325 ( .A(n8902), .ZN(n8903) );
  NAND2_X1 U11326 ( .A1(n8904), .A2(n8903), .ZN(n8905) );
  MUX2_X1 U11327 ( .A(n13594), .B(n10552), .S(n9192), .Z(n8907) );
  AND2_X1 U11328 ( .A1(n8909), .A2(n8908), .ZN(n8910) );
  NOR2_X1 U11329 ( .A1(n8928), .A2(n8910), .ZN(n10884) );
  NAND2_X1 U11330 ( .A1(n6463), .A2(n10884), .ZN(n8914) );
  NAND2_X1 U11331 ( .A1(n6425), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8913) );
  NAND2_X1 U11332 ( .A1(n6466), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8912) );
  NAND2_X1 U11333 ( .A1(n8889), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8911) );
  NAND4_X1 U11334 ( .A1(n8914), .A2(n8913), .A3(n8912), .A4(n8911), .ZN(n13593) );
  NAND2_X1 U11335 ( .A1(n9552), .A2(n9262), .ZN(n8920) );
  AND2_X1 U11336 ( .A1(n8916), .A2(n8915), .ZN(n8922) );
  OR2_X1 U11337 ( .A1(n8922), .A2(n6613), .ZN(n8917) );
  XNOR2_X1 U11338 ( .A(n8917), .B(n8921), .ZN(n9717) );
  INV_X1 U11339 ( .A(n8918), .ZN(n8919) );
  MUX2_X1 U11340 ( .A(n13593), .B(n14346), .S(n9192), .Z(n8940) );
  NAND2_X1 U11341 ( .A1(n9555), .A2(n9262), .ZN(n8927) );
  NAND2_X1 U11342 ( .A1(n8922), .A2(n8921), .ZN(n8945) );
  NAND2_X1 U11343 ( .A1(n8945), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8924) );
  XNOR2_X1 U11344 ( .A(n8924), .B(n8923), .ZN(n9813) );
  INV_X1 U11345 ( .A(n8925), .ZN(n8926) );
  NAND2_X1 U11346 ( .A1(n8927), .A2(n8926), .ZN(n11045) );
  OR2_X1 U11347 ( .A1(n8928), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8929) );
  AND2_X1 U11348 ( .A1(n8951), .A2(n8929), .ZN(n11050) );
  NAND2_X1 U11349 ( .A1(n6463), .A2(n11050), .ZN(n8933) );
  NAND2_X1 U11350 ( .A1(n6425), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8932) );
  NAND2_X1 U11351 ( .A1(n9265), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8931) );
  NAND2_X1 U11352 ( .A1(n8889), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8930) );
  NAND4_X1 U11353 ( .A1(n8933), .A2(n8932), .A3(n8931), .A4(n8930), .ZN(n13592) );
  INV_X1 U11354 ( .A(n13592), .ZN(n8934) );
  OR2_X1 U11355 ( .A1(n11045), .A2(n8934), .ZN(n10763) );
  NAND2_X1 U11356 ( .A1(n11045), .A2(n8934), .ZN(n10764) );
  NAND2_X1 U11357 ( .A1(n10763), .A2(n10764), .ZN(n10754) );
  NAND3_X1 U11358 ( .A1(n10763), .A2(n9238), .A3(n14346), .ZN(n8936) );
  NAND3_X1 U11359 ( .A1(n10764), .A2(n9192), .A3(n13593), .ZN(n8935) );
  AND2_X1 U11360 ( .A1(n8936), .A2(n8935), .ZN(n8939) );
  OAI21_X1 U11361 ( .B1(n8940), .B2(n10754), .A(n8939), .ZN(n8937) );
  INV_X1 U11362 ( .A(n8939), .ZN(n8942) );
  INV_X1 U11363 ( .A(n8940), .ZN(n8941) );
  NAND2_X1 U11364 ( .A1(n8942), .A2(n8941), .ZN(n8944) );
  MUX2_X1 U11365 ( .A(n10764), .B(n10763), .S(n9192), .Z(n8943) );
  NAND2_X1 U11366 ( .A1(n9570), .A2(n9262), .ZN(n8949) );
  NAND2_X1 U11367 ( .A1(n9051), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8946) );
  XNOR2_X1 U11368 ( .A(n8946), .B(n6451), .ZN(n9617) );
  INV_X1 U11369 ( .A(n8947), .ZN(n8948) );
  NAND2_X1 U11370 ( .A1(n8949), .A2(n8948), .ZN(n11258) );
  NAND2_X1 U11371 ( .A1(n8951), .A2(n8950), .ZN(n8952) );
  AND2_X1 U11372 ( .A1(n8962), .A2(n8952), .ZN(n11253) );
  NAND2_X1 U11373 ( .A1(n6462), .A2(n11253), .ZN(n8956) );
  NAND2_X1 U11374 ( .A1(n6464), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8955) );
  NAND2_X1 U11375 ( .A1(n9265), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8954) );
  NAND2_X1 U11376 ( .A1(n8889), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8953) );
  NAND4_X1 U11377 ( .A1(n8956), .A2(n8955), .A3(n8954), .A4(n8953), .ZN(n13591) );
  NAND2_X1 U11378 ( .A1(n11258), .A2(n11246), .ZN(n9283) );
  OR2_X1 U11379 ( .A1(n11258), .A2(n11246), .ZN(n10788) );
  MUX2_X1 U11380 ( .A(n9283), .B(n10788), .S(n9238), .Z(n8957) );
  INV_X1 U11381 ( .A(n11258), .ZN(n14364) );
  MUX2_X1 U11382 ( .A(n11246), .B(n14364), .S(n9192), .Z(n8959) );
  OR2_X1 U11383 ( .A1(n11258), .A2(n13591), .ZN(n10786) );
  NAND2_X1 U11384 ( .A1(n8959), .A2(n10786), .ZN(n8960) );
  AND2_X1 U11385 ( .A1(n8962), .A2(n8961), .ZN(n8963) );
  NOR2_X1 U11386 ( .A1(n8996), .A2(n8963), .ZN(n11423) );
  NAND2_X1 U11387 ( .A1(n6463), .A2(n11423), .ZN(n8967) );
  NAND2_X1 U11388 ( .A1(n6464), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8966) );
  NAND2_X1 U11389 ( .A1(n9265), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8965) );
  NAND2_X1 U11390 ( .A1(n9266), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8964) );
  NAND4_X1 U11391 ( .A1(n8967), .A2(n8966), .A3(n8965), .A4(n8964), .ZN(n13590) );
  NAND2_X1 U11392 ( .A1(n9583), .A2(n9262), .ZN(n8972) );
  NAND2_X1 U11393 ( .A1(n8980), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8969) );
  INV_X1 U11394 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8968) );
  XNOR2_X1 U11395 ( .A(n8969), .B(n8968), .ZN(n9700) );
  INV_X1 U11396 ( .A(n8970), .ZN(n8971) );
  MUX2_X1 U11397 ( .A(n11577), .B(n11426), .S(n9192), .Z(n8974) );
  INV_X1 U11398 ( .A(n11426), .ZN(n10803) );
  MUX2_X1 U11399 ( .A(n13590), .B(n10803), .S(n9238), .Z(n8973) );
  INV_X1 U11400 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8975) );
  XNOR2_X1 U11401 ( .A(n8996), .B(n8975), .ZN(n14286) );
  NAND2_X1 U11402 ( .A1(n6462), .A2(n14286), .ZN(n8979) );
  NAND2_X1 U11403 ( .A1(n6464), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8978) );
  NAND2_X1 U11404 ( .A1(n9265), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n8977) );
  NAND2_X1 U11405 ( .A1(n9266), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8976) );
  NAND4_X1 U11406 ( .A1(n8979), .A2(n8978), .A3(n8977), .A4(n8976), .ZN(n14130) );
  NAND2_X1 U11407 ( .A1(n9589), .A2(n9235), .ZN(n8987) );
  NOR2_X1 U11408 ( .A1(n8983), .A2(n6613), .ZN(n8981) );
  MUX2_X1 U11409 ( .A(n6613), .B(n8981), .S(P1_IR_REG_10__SCAN_IN), .Z(n8985)
         );
  NAND2_X1 U11410 ( .A1(n8983), .A2(n8982), .ZN(n9015) );
  INV_X1 U11411 ( .A(n9015), .ZN(n8984) );
  NOR2_X1 U11412 ( .A1(n8985), .A2(n8984), .ZN(n10379) );
  AOI22_X1 U11413 ( .A1(n10379), .A2(n9053), .B1(n9271), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n8986) );
  NAND2_X1 U11414 ( .A1(n8987), .A2(n8986), .ZN(n14287) );
  MUX2_X1 U11415 ( .A(n14130), .B(n14287), .S(n9238), .Z(n8991) );
  NAND2_X1 U11416 ( .A1(n8990), .A2(n8991), .ZN(n8989) );
  MUX2_X1 U11417 ( .A(n14130), .B(n14287), .S(n9192), .Z(n8988) );
  NAND2_X1 U11418 ( .A1(n8989), .A2(n8988), .ZN(n8995) );
  INV_X1 U11419 ( .A(n8990), .ZN(n8993) );
  INV_X1 U11420 ( .A(n8991), .ZN(n8992) );
  NAND2_X1 U11421 ( .A1(n8993), .A2(n8992), .ZN(n8994) );
  NAND2_X1 U11422 ( .A1(n8995), .A2(n8994), .ZN(n9006) );
  AOI21_X1 U11423 ( .B1(n8996), .B2(P1_REG3_REG_10__SCAN_IN), .A(
        P1_REG3_REG_11__SCAN_IN), .ZN(n8997) );
  OR2_X1 U11424 ( .A1(n9009), .A2(n8997), .ZN(n14145) );
  INV_X1 U11425 ( .A(n14145), .ZN(n14169) );
  NAND2_X1 U11426 ( .A1(n6462), .A2(n14169), .ZN(n9001) );
  NAND2_X1 U11427 ( .A1(n6464), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9000) );
  NAND2_X1 U11428 ( .A1(n9265), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8999) );
  NAND2_X1 U11429 ( .A1(n8889), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8998) );
  NAND4_X1 U11430 ( .A1(n9001), .A2(n9000), .A3(n8999), .A4(n8998), .ZN(n14291) );
  NAND2_X1 U11431 ( .A1(n9624), .A2(n9262), .ZN(n9004) );
  NAND2_X1 U11432 ( .A1(n9015), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9002) );
  XNOR2_X1 U11433 ( .A(n9002), .B(P1_IR_REG_11__SCAN_IN), .ZN(n13674) );
  AOI22_X1 U11434 ( .A1(n13674), .A2(n9053), .B1(n9271), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n9003) );
  MUX2_X1 U11435 ( .A(n14291), .B(n14172), .S(n9192), .Z(n9007) );
  MUX2_X1 U11436 ( .A(n14291), .B(n14172), .S(n9238), .Z(n9005) );
  INV_X1 U11437 ( .A(n9007), .ZN(n9008) );
  OR2_X1 U11438 ( .A1(n9009), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9010) );
  AND2_X1 U11439 ( .A1(n9041), .A2(n9010), .ZN(n11795) );
  NAND2_X1 U11440 ( .A1(n6462), .A2(n11795), .ZN(n9014) );
  NAND2_X1 U11441 ( .A1(n6464), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9013) );
  NAND2_X1 U11442 ( .A1(n9265), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9012) );
  NAND2_X1 U11443 ( .A1(n9266), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9011) );
  NAND4_X1 U11444 ( .A1(n9014), .A2(n9013), .A3(n9012), .A4(n9011), .ZN(n14129) );
  NAND2_X1 U11445 ( .A1(n9782), .A2(n9262), .ZN(n9018) );
  NAND2_X1 U11446 ( .A1(n9016), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9028) );
  XNOR2_X1 U11447 ( .A(n9028), .B(P1_IR_REG_12__SCAN_IN), .ZN(n13694) );
  AOI22_X1 U11448 ( .A1(n13694), .A2(n9053), .B1(n9271), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n9017) );
  NAND2_X2 U11449 ( .A1(n9018), .A2(n9017), .ZN(n11787) );
  MUX2_X1 U11450 ( .A(n14129), .B(n11787), .S(n9238), .Z(n9022) );
  NAND2_X1 U11451 ( .A1(n9021), .A2(n9022), .ZN(n9020) );
  MUX2_X1 U11452 ( .A(n14129), .B(n11787), .S(n9192), .Z(n9019) );
  NAND2_X1 U11453 ( .A1(n9020), .A2(n9019), .ZN(n9026) );
  INV_X1 U11454 ( .A(n9022), .ZN(n9023) );
  NAND2_X1 U11455 ( .A1(n9024), .A2(n9023), .ZN(n9025) );
  NAND2_X1 U11456 ( .A1(n10050), .A2(n9262), .ZN(n9033) );
  INV_X1 U11457 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9027) );
  NAND2_X1 U11458 ( .A1(n9028), .A2(n9027), .ZN(n9029) );
  NAND2_X1 U11459 ( .A1(n9029), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9047) );
  INV_X1 U11460 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9046) );
  NAND2_X1 U11461 ( .A1(n9047), .A2(n9046), .ZN(n9030) );
  NAND2_X1 U11462 ( .A1(n9030), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9031) );
  AOI22_X1 U11463 ( .A1(n11392), .A2(n9053), .B1(n9271), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9032) );
  OAI21_X1 U11464 ( .B1(n9041), .B2(n9035), .A(n9034), .ZN(n9036) );
  NAND2_X1 U11465 ( .A1(n9036), .A2(n9056), .ZN(n14128) );
  INV_X1 U11466 ( .A(n14128), .ZN(n11331) );
  NAND2_X1 U11467 ( .A1(n6463), .A2(n11331), .ZN(n9040) );
  NAND2_X1 U11468 ( .A1(n6464), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9039) );
  NAND2_X1 U11469 ( .A1(n9266), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9038) );
  NAND2_X1 U11470 ( .A1(n9265), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9037) );
  NAND4_X1 U11471 ( .A1(n9040), .A2(n9039), .A3(n9038), .A4(n9037), .ZN(n13588) );
  INV_X1 U11472 ( .A(n13588), .ZN(n13571) );
  XNOR2_X1 U11473 ( .A(n14210), .B(n13571), .ZN(n9290) );
  XNOR2_X1 U11474 ( .A(n9041), .B(P1_REG3_REG_13__SCAN_IN), .ZN(n11838) );
  NAND2_X1 U11475 ( .A1(n6462), .A2(n11838), .ZN(n9045) );
  NAND2_X1 U11476 ( .A1(n6464), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9044) );
  NAND2_X1 U11477 ( .A1(n9266), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9043) );
  NAND2_X1 U11478 ( .A1(n9265), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9042) );
  NAND4_X1 U11479 ( .A1(n9045), .A2(n9044), .A3(n9043), .A4(n9042), .ZN(n13589) );
  NAND2_X1 U11480 ( .A1(n9827), .A2(n9235), .ZN(n9048) );
  XNOR2_X1 U11481 ( .A(n9047), .B(n9046), .ZN(n10415) );
  MUX2_X1 U11482 ( .A(n13589), .B(n11832), .S(n9192), .Z(n9064) );
  NAND2_X1 U11483 ( .A1(n10139), .A2(n9235), .ZN(n9055) );
  OAI21_X1 U11484 ( .B1(n9051), .B2(n9050), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9052) );
  XNOR2_X1 U11485 ( .A(n9052), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11402) );
  AOI22_X1 U11486 ( .A1(n9271), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9053), 
        .B2(n11402), .ZN(n9054) );
  AND2_X1 U11487 ( .A1(n9056), .A2(n14977), .ZN(n9057) );
  NOR2_X1 U11488 ( .A1(n9070), .A2(n9057), .ZN(n13575) );
  NAND2_X1 U11489 ( .A1(n6462), .A2(n13575), .ZN(n9061) );
  NAND2_X1 U11490 ( .A1(n6464), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9060) );
  NAND2_X1 U11491 ( .A1(n9265), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n9059) );
  NAND2_X1 U11492 ( .A1(n9266), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n9058) );
  NAND4_X1 U11493 ( .A1(n9061), .A2(n9060), .A3(n9059), .A4(n9058), .ZN(n13587) );
  INV_X1 U11494 ( .A(n13587), .ZN(n11908) );
  OR2_X1 U11495 ( .A1(n14210), .A2(n13571), .ZN(n11540) );
  NAND2_X1 U11496 ( .A1(n11656), .A2(n11540), .ZN(n9062) );
  NAND2_X1 U11497 ( .A1(n9062), .A2(n9192), .ZN(n9063) );
  MUX2_X1 U11498 ( .A(n11832), .B(n9065), .S(n9192), .Z(n9066) );
  NAND2_X1 U11499 ( .A1(n14210), .A2(n13571), .ZN(n11538) );
  NAND2_X1 U11500 ( .A1(n9281), .A2(n11538), .ZN(n9067) );
  OR2_X1 U11501 ( .A1(n11656), .A2(n9192), .ZN(n9068) );
  NAND2_X1 U11502 ( .A1(n9069), .A2(n9068), .ZN(n9082) );
  NOR2_X1 U11503 ( .A1(n9070), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9071) );
  OR2_X1 U11504 ( .A1(n9091), .A2(n9071), .ZN(n13504) );
  NAND2_X1 U11505 ( .A1(n9265), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9073) );
  NAND2_X1 U11506 ( .A1(n9266), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9072) );
  AND2_X1 U11507 ( .A1(n9073), .A2(n9072), .ZN(n9075) );
  NAND2_X1 U11508 ( .A1(n6464), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9074) );
  OAI211_X1 U11509 ( .C1(n13504), .C2(n9130), .A(n9075), .B(n9074), .ZN(n13586) );
  NAND2_X1 U11510 ( .A1(n10004), .A2(n9235), .ZN(n9080) );
  NAND2_X1 U11511 ( .A1(n9076), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9077) );
  XNOR2_X1 U11512 ( .A(n9077), .B(n8797), .ZN(n11591) );
  INV_X1 U11513 ( .A(n9078), .ZN(n9079) );
  MUX2_X1 U11514 ( .A(n13586), .B(n14195), .S(n9192), .Z(n9083) );
  MUX2_X1 U11515 ( .A(n13586), .B(n14195), .S(n9238), .Z(n9081) );
  NAND2_X1 U11516 ( .A1(n10096), .A2(n9235), .ZN(n9090) );
  NAND2_X1 U11517 ( .A1(n9084), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9086) );
  MUX2_X1 U11518 ( .A(n9086), .B(P1_IR_REG_31__SCAN_IN), .S(n9085), .Z(n9087)
         );
  AND2_X1 U11519 ( .A1(n9087), .A2(n6578), .ZN(n11589) );
  INV_X1 U11520 ( .A(n9088), .ZN(n9089) );
  NOR2_X1 U11521 ( .A1(n9091), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9092) );
  OR2_X1 U11522 ( .A1(n9097), .A2(n9092), .ZN(n13510) );
  AOI22_X1 U11523 ( .A1(n9266), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n9265), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U11524 ( .A1(n6464), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9093) );
  OAI211_X1 U11525 ( .C1(n13510), .C2(n9130), .A(n9094), .B(n9093), .ZN(n13585) );
  XNOR2_X1 U11526 ( .A(n14154), .B(n13585), .ZN(n14155) );
  INV_X1 U11527 ( .A(n13585), .ZN(n13891) );
  NAND2_X1 U11528 ( .A1(n14154), .A2(n13891), .ZN(n9095) );
  OR2_X1 U11529 ( .A1(n14154), .A2(n13891), .ZN(n11866) );
  MUX2_X1 U11530 ( .A(n9095), .B(n11866), .S(n9238), .Z(n9096) );
  OR2_X1 U11531 ( .A1(n9097), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9098) );
  NAND2_X1 U11532 ( .A1(n9113), .A2(n9098), .ZN(n13903) );
  AOI22_X1 U11533 ( .A1(n9266), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n9265), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n9100) );
  NAND2_X1 U11534 ( .A1(n6464), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9099) );
  OAI211_X1 U11535 ( .C1(n13903), .C2(n9130), .A(n9100), .B(n9099), .ZN(n13875) );
  XNOR2_X1 U11536 ( .A(n13875), .B(n9238), .ZN(n9107) );
  NAND2_X1 U11537 ( .A1(n10389), .A2(n9235), .ZN(n9105) );
  NAND2_X1 U11538 ( .A1(n6578), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9102) );
  XNOR2_X1 U11539 ( .A(n9102), .B(n9101), .ZN(n13711) );
  INV_X1 U11540 ( .A(n9103), .ZN(n9104) );
  XNOR2_X1 U11541 ( .A(n14180), .B(n9192), .ZN(n9106) );
  OAI21_X1 U11542 ( .B1(n9108), .B2(n9107), .A(n9106), .ZN(n9123) );
  NAND2_X1 U11543 ( .A1(n9108), .A2(n9107), .ZN(n9122) );
  NAND2_X1 U11544 ( .A1(n10555), .A2(n9262), .ZN(n9111) );
  INV_X1 U11545 ( .A(n9109), .ZN(n9110) );
  NAND2_X1 U11546 ( .A1(n9113), .A2(n9112), .ZN(n9114) );
  AND2_X1 U11547 ( .A1(n9127), .A2(n9114), .ZN(n13877) );
  NAND2_X1 U11548 ( .A1(n13877), .A2(n6462), .ZN(n9121) );
  INV_X1 U11549 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9118) );
  NAND2_X1 U11550 ( .A1(n9265), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9116) );
  NAND2_X1 U11551 ( .A1(n9266), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9115) );
  OAI211_X1 U11552 ( .C1(n9118), .C2(n9117), .A(n9116), .B(n9115), .ZN(n9119)
         );
  INV_X1 U11553 ( .A(n9119), .ZN(n9120) );
  OR2_X1 U11554 ( .A1(n13874), .A2(n13893), .ZN(n9124) );
  NAND2_X1 U11555 ( .A1(n13874), .A2(n13893), .ZN(n11871) );
  NAND3_X1 U11556 ( .A1(n9123), .A2(n9122), .A3(n13871), .ZN(n9126) );
  MUX2_X1 U11557 ( .A(n11871), .B(n9124), .S(n9192), .Z(n9125) );
  NAND2_X1 U11558 ( .A1(n9126), .A2(n9125), .ZN(n9141) );
  NAND2_X1 U11559 ( .A1(n9127), .A2(n11949), .ZN(n9129) );
  INV_X1 U11560 ( .A(n9128), .ZN(n9145) );
  NAND2_X1 U11561 ( .A1(n9129), .A2(n9145), .ZN(n13861) );
  OR2_X1 U11562 ( .A1(n13861), .A2(n9130), .ZN(n9136) );
  INV_X1 U11563 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9133) );
  NAND2_X1 U11564 ( .A1(n6466), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U11565 ( .A1(n9266), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9131) );
  OAI211_X1 U11566 ( .C1(n9133), .C2(n9117), .A(n9132), .B(n9131), .ZN(n9134)
         );
  INV_X1 U11567 ( .A(n9134), .ZN(n9135) );
  NAND2_X1 U11568 ( .A1(n10993), .A2(n9262), .ZN(n9138) );
  NAND2_X1 U11569 ( .A1(n9271), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9137) );
  MUX2_X1 U11570 ( .A(n13476), .B(n13971), .S(n9192), .Z(n9140) );
  INV_X1 U11571 ( .A(n13971), .ZN(n9280) );
  MUX2_X1 U11572 ( .A(n13876), .B(n9280), .S(n9238), .Z(n9139) );
  OAI21_X1 U11573 ( .B1(n9141), .B2(n9140), .A(n9139), .ZN(n9143) );
  NAND2_X1 U11574 ( .A1(n9141), .A2(n9140), .ZN(n9142) );
  INV_X1 U11575 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13484) );
  AOI21_X1 U11576 ( .B1(n13484), .B2(n9145), .A(n9144), .ZN(n13846) );
  NAND2_X1 U11577 ( .A1(n6463), .A2(n13846), .ZN(n9149) );
  NAND2_X1 U11578 ( .A1(n6464), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9148) );
  NAND2_X1 U11579 ( .A1(n6466), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9147) );
  NAND2_X1 U11580 ( .A1(n9266), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9146) );
  NAND4_X1 U11581 ( .A1(n9149), .A2(n9148), .A3(n9147), .A4(n9146), .ZN(n13828) );
  NAND2_X1 U11582 ( .A1(n11142), .A2(n9262), .ZN(n9151) );
  NAND2_X1 U11583 ( .A1(n9271), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9150) );
  MUX2_X1 U11584 ( .A(n13828), .B(n13965), .S(n9238), .Z(n9153) );
  MUX2_X1 U11585 ( .A(n13828), .B(n13965), .S(n9192), .Z(n9152) );
  INV_X1 U11586 ( .A(n9153), .ZN(n9154) );
  NAND2_X1 U11587 ( .A1(n6464), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n9160) );
  INV_X1 U11588 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13529) );
  AOI21_X1 U11589 ( .B1(n13529), .B2(n9156), .A(n9155), .ZN(n13833) );
  NAND2_X1 U11590 ( .A1(n6462), .A2(n13833), .ZN(n9159) );
  NAND2_X1 U11591 ( .A1(n9266), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9158) );
  NAND2_X1 U11592 ( .A1(n6466), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9157) );
  NAND4_X1 U11593 ( .A1(n9160), .A2(n9159), .A3(n9158), .A4(n9157), .ZN(n13583) );
  NAND2_X1 U11594 ( .A1(n9161), .A2(n9504), .ZN(n9162) );
  MUX2_X1 U11595 ( .A(n13583), .B(n13960), .S(n9192), .Z(n9166) );
  MUX2_X1 U11596 ( .A(n13583), .B(n13960), .S(n9238), .Z(n9163) );
  NAND2_X1 U11597 ( .A1(n9164), .A2(n9163), .ZN(n9170) );
  INV_X1 U11598 ( .A(n9165), .ZN(n9168) );
  INV_X1 U11599 ( .A(n9166), .ZN(n9167) );
  NAND2_X1 U11600 ( .A1(n9168), .A2(n9167), .ZN(n9169) );
  NAND2_X1 U11601 ( .A1(n9170), .A2(n9169), .ZN(n9180) );
  INV_X1 U11602 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13461) );
  AOI21_X1 U11603 ( .B1(n13461), .B2(n9172), .A(n9171), .ZN(n13817) );
  NAND2_X1 U11604 ( .A1(n6463), .A2(n13817), .ZN(n9176) );
  NAND2_X1 U11605 ( .A1(n6464), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9175) );
  NAND2_X1 U11606 ( .A1(n6466), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9174) );
  NAND2_X1 U11607 ( .A1(n9266), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9173) );
  NAND4_X1 U11608 ( .A1(n9176), .A2(n9175), .A3(n9174), .A4(n9173), .ZN(n13827) );
  NAND2_X1 U11609 ( .A1(n11444), .A2(n9262), .ZN(n9178) );
  NAND2_X1 U11610 ( .A1(n9271), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9177) );
  NAND2_X2 U11611 ( .A1(n9178), .A2(n9177), .ZN(n13952) );
  MUX2_X1 U11612 ( .A(n13827), .B(n13952), .S(n9238), .Z(n9181) );
  MUX2_X1 U11613 ( .A(n13827), .B(n13952), .S(n9192), .Z(n9179) );
  INV_X1 U11614 ( .A(n9181), .ZN(n9182) );
  INV_X1 U11615 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9185) );
  AOI21_X1 U11616 ( .B1(n9185), .B2(n9184), .A(n9183), .ZN(n13804) );
  NAND2_X1 U11617 ( .A1(n6462), .A2(n13804), .ZN(n9189) );
  NAND2_X1 U11618 ( .A1(n6464), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9188) );
  NAND2_X1 U11619 ( .A1(n6466), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9187) );
  NAND2_X1 U11620 ( .A1(n9266), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9186) );
  NAND4_X1 U11621 ( .A1(n9189), .A2(n9188), .A3(n9187), .A4(n9186), .ZN(n13779) );
  NAND2_X1 U11622 ( .A1(n11531), .A2(n9262), .ZN(n9191) );
  NAND2_X1 U11623 ( .A1(n9271), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9190) );
  MUX2_X1 U11624 ( .A(n13779), .B(n13805), .S(n9192), .Z(n9196) );
  MUX2_X1 U11625 ( .A(n13779), .B(n13805), .S(n9238), .Z(n9193) );
  NAND2_X1 U11626 ( .A1(n9194), .A2(n9193), .ZN(n9198) );
  NAND2_X1 U11627 ( .A1(n9198), .A2(n9197), .ZN(n9210) );
  INV_X1 U11628 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9200) );
  NAND2_X1 U11629 ( .A1(n9200), .A2(n9199), .ZN(n9201) );
  AND2_X1 U11630 ( .A1(n9201), .A2(n9217), .ZN(n13782) );
  NAND2_X1 U11631 ( .A1(n6463), .A2(n13782), .ZN(n9205) );
  NAND2_X1 U11632 ( .A1(n6464), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9204) );
  NAND2_X1 U11633 ( .A1(n6466), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9203) );
  NAND2_X1 U11634 ( .A1(n9266), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9202) );
  NAND4_X1 U11635 ( .A1(n9205), .A2(n9204), .A3(n9203), .A4(n9202), .ZN(n13799) );
  NAND2_X1 U11636 ( .A1(n11611), .A2(n9262), .ZN(n9207) );
  NAND2_X1 U11637 ( .A1(n9271), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9206) );
  MUX2_X1 U11638 ( .A(n13799), .B(n13942), .S(n9238), .Z(n9211) );
  NAND2_X1 U11639 ( .A1(n9210), .A2(n9211), .ZN(n9209) );
  MUX2_X1 U11640 ( .A(n13799), .B(n13942), .S(n9192), .Z(n9208) );
  NAND2_X1 U11641 ( .A1(n9209), .A2(n9208), .ZN(n9215) );
  NAND2_X1 U11642 ( .A1(n9213), .A2(n9212), .ZN(n9214) );
  NAND2_X1 U11643 ( .A1(n9215), .A2(n9214), .ZN(n9226) );
  INV_X1 U11644 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9216) );
  NAND2_X1 U11645 ( .A1(n9217), .A2(n9216), .ZN(n9218) );
  NAND2_X1 U11646 ( .A1(n6463), .A2(n13768), .ZN(n9222) );
  NAND2_X1 U11647 ( .A1(n6464), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U11648 ( .A1(n6466), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9220) );
  NAND2_X1 U11649 ( .A1(n9266), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9219) );
  NAND4_X1 U11650 ( .A1(n9222), .A2(n9221), .A3(n9220), .A4(n9219), .ZN(n13778) );
  NAND2_X1 U11651 ( .A1(n13441), .A2(n9262), .ZN(n9224) );
  NAND2_X1 U11652 ( .A1(n9271), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9223) );
  MUX2_X1 U11653 ( .A(n13778), .B(n13562), .S(n9192), .Z(n9227) );
  MUX2_X1 U11654 ( .A(n13778), .B(n13562), .S(n9238), .Z(n9225) );
  INV_X1 U11655 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9228) );
  NAND2_X1 U11656 ( .A1(n9229), .A2(n9228), .ZN(n9230) );
  NAND2_X1 U11657 ( .A1(n6462), .A2(n13449), .ZN(n9234) );
  NAND2_X1 U11658 ( .A1(n6464), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9233) );
  NAND2_X1 U11659 ( .A1(n9266), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9232) );
  NAND2_X1 U11660 ( .A1(n6466), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9231) );
  NAND4_X1 U11661 ( .A1(n9234), .A2(n9233), .A3(n9232), .A4(n9231), .ZN(n13765) );
  NAND2_X1 U11662 ( .A1(n11841), .A2(n9235), .ZN(n9237) );
  NAND2_X1 U11663 ( .A1(n9271), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9236) );
  MUX2_X1 U11664 ( .A(n13765), .B(n13454), .S(n9238), .Z(n9242) );
  MUX2_X1 U11665 ( .A(n13765), .B(n13454), .S(n9192), .Z(n9239) );
  NAND2_X1 U11666 ( .A1(n9240), .A2(n9239), .ZN(n9245) );
  INV_X1 U11667 ( .A(n9241), .ZN(n9244) );
  INV_X1 U11668 ( .A(n9242), .ZN(n9243) );
  NAND2_X1 U11669 ( .A1(n6464), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9251) );
  XNOR2_X1 U11670 ( .A(n9246), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n13748) );
  NAND2_X1 U11671 ( .A1(n6463), .A2(n13748), .ZN(n9250) );
  NAND2_X1 U11672 ( .A1(n9266), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9249) );
  NAND2_X1 U11673 ( .A1(n6465), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9248) );
  NAND4_X1 U11674 ( .A1(n9251), .A2(n9250), .A3(n9249), .A4(n9248), .ZN(n13582) );
  NAND2_X1 U11675 ( .A1(n9271), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9252) );
  MUX2_X1 U11676 ( .A(n13582), .B(n13927), .S(n9192), .Z(n9254) );
  MUX2_X1 U11677 ( .A(n13582), .B(n13927), .S(n9238), .Z(n9255) );
  INV_X1 U11678 ( .A(n12372), .ZN(n13581) );
  MUX2_X1 U11679 ( .A(n13581), .B(n11880), .S(n9192), .Z(n9256) );
  NAND2_X1 U11680 ( .A1(n9271), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n9263) );
  NAND2_X1 U11681 ( .A1(n6464), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n9269) );
  NAND2_X1 U11682 ( .A1(n6465), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9268) );
  NAND2_X1 U11683 ( .A1(n9266), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9267) );
  AND3_X1 U11684 ( .A1(n9269), .A2(n9268), .A3(n9267), .ZN(n9300) );
  XNOR2_X1 U11685 ( .A(n13732), .B(n9300), .ZN(n9324) );
  INV_X1 U11686 ( .A(n9324), .ZN(n9333) );
  NAND2_X1 U11687 ( .A1(n9271), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9272) );
  NAND2_X1 U11688 ( .A1(n6464), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9277) );
  NAND2_X1 U11689 ( .A1(n6466), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9276) );
  NAND2_X1 U11690 ( .A1(n9266), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9275) );
  AND3_X1 U11691 ( .A1(n9277), .A2(n9276), .A3(n9275), .ZN(n9306) );
  INV_X1 U11692 ( .A(n9306), .ZN(n13580) );
  XNOR2_X1 U11693 ( .A(n13738), .B(n13580), .ZN(n9297) );
  XOR2_X1 U11694 ( .A(n13582), .B(n13927), .Z(n13746) );
  XNOR2_X1 U11695 ( .A(n13454), .B(n13560), .ZN(n12049) );
  NAND2_X1 U11696 ( .A1(n13562), .A2(n13493), .ZN(n12044) );
  OR2_X1 U11697 ( .A1(n13562), .A2(n13493), .ZN(n9278) );
  NAND2_X1 U11698 ( .A1(n12044), .A2(n9278), .ZN(n13760) );
  NAND2_X1 U11699 ( .A1(n13942), .A2(n13799), .ZN(n11859) );
  OR2_X1 U11700 ( .A1(n13942), .A2(n13799), .ZN(n9279) );
  NAND2_X1 U11701 ( .A1(n11859), .A2(n9279), .ZN(n13785) );
  INV_X1 U11702 ( .A(n13828), .ZN(n13531) );
  XNOR2_X1 U11703 ( .A(n13965), .B(n13531), .ZN(n13842) );
  XNOR2_X1 U11704 ( .A(n9280), .B(n13876), .ZN(n13859) );
  NAND2_X1 U11705 ( .A1(n11656), .A2(n9281), .ZN(n11547) );
  INV_X1 U11706 ( .A(n14155), .ZN(n14147) );
  XNOR2_X1 U11707 ( .A(n14195), .B(n13586), .ZN(n11653) );
  INV_X1 U11708 ( .A(n14130), .ZN(n11572) );
  OR2_X1 U11709 ( .A1(n14287), .A2(n11572), .ZN(n11232) );
  NAND2_X1 U11710 ( .A1(n14287), .A2(n11572), .ZN(n9282) );
  NAND2_X1 U11711 ( .A1(n11232), .A2(n9282), .ZN(n14289) );
  XNOR2_X1 U11712 ( .A(n14172), .B(n11792), .ZN(n14171) );
  XNOR2_X1 U11713 ( .A(n10803), .B(n11577), .ZN(n11222) );
  AND2_X1 U11714 ( .A1(n10788), .A2(n9283), .ZN(n10758) );
  AND2_X2 U11715 ( .A1(n9928), .A2(n9284), .ZN(n10092) );
  NAND4_X1 U11716 ( .A1(n10092), .A2(n14298), .A3(n9912), .A4(n10103), .ZN(
        n9285) );
  NOR4_X1 U11717 ( .A1(n10148), .A2(n10223), .A3(n9285), .A4(n10754), .ZN(
        n9286) );
  XNOR2_X1 U11718 ( .A(n14346), .B(n13593), .ZN(n10353) );
  NAND3_X1 U11719 ( .A1(n10758), .A2(n9286), .A3(n10353), .ZN(n9287) );
  NOR4_X1 U11720 ( .A1(n14289), .A2(n14171), .A3(n11222), .A4(n9287), .ZN(
        n9288) );
  XNOR2_X1 U11721 ( .A(n11832), .B(n13589), .ZN(n11336) );
  XNOR2_X1 U11722 ( .A(n11787), .B(n14129), .ZN(n11261) );
  NAND4_X1 U11723 ( .A1(n11653), .A2(n9288), .A3(n11336), .A4(n11261), .ZN(
        n9289) );
  NOR4_X1 U11724 ( .A1(n11547), .A2(n9290), .A3(n14147), .A4(n9289), .ZN(n9291) );
  XNOR2_X1 U11725 ( .A(n14180), .B(n13875), .ZN(n13897) );
  NAND4_X1 U11726 ( .A1(n13859), .A2(n13871), .A3(n9291), .A4(n13897), .ZN(
        n9292) );
  NOR3_X1 U11727 ( .A1(n13837), .A2(n13842), .A3(n9292), .ZN(n9293) );
  XNOR2_X1 U11728 ( .A(n13805), .B(n13779), .ZN(n13793) );
  NAND4_X1 U11729 ( .A1(n13785), .A2(n9293), .A3(n13813), .A4(n13793), .ZN(
        n9294) );
  NOR4_X1 U11730 ( .A1(n13746), .A2(n12049), .A3(n13760), .A4(n9294), .ZN(
        n9295) );
  XNOR2_X1 U11731 ( .A(n11880), .B(n13581), .ZN(n11878) );
  NAND2_X1 U11732 ( .A1(n9333), .A2(n7356), .ZN(n9298) );
  NAND2_X1 U11733 ( .A1(n9302), .A2(n12380), .ZN(n9762) );
  INV_X1 U11734 ( .A(n9300), .ZN(n13734) );
  MUX2_X1 U11735 ( .A(n13734), .B(n9238), .S(n13732), .Z(n9301) );
  NAND2_X1 U11736 ( .A1(n9238), .A2(n13734), .ZN(n9308) );
  OR2_X1 U11737 ( .A1(n9747), .A2(n10556), .ZN(n9304) );
  OAI21_X1 U11738 ( .B1(n14017), .B2(n9302), .A(n9911), .ZN(n9303) );
  AND2_X1 U11739 ( .A1(n9304), .A2(n9303), .ZN(n9320) );
  NAND2_X1 U11740 ( .A1(n9305), .A2(n12380), .ZN(n9307) );
  AOI21_X1 U11741 ( .B1(n9308), .B2(n9307), .A(n9306), .ZN(n9309) );
  AOI21_X1 U11742 ( .B1(n13738), .B2(n9192), .A(n9309), .ZN(n9326) );
  INV_X1 U11743 ( .A(n9326), .ZN(n9330) );
  NAND2_X1 U11744 ( .A1(n9334), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9310) );
  AND2_X1 U11745 ( .A1(n9743), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9561) );
  INV_X1 U11746 ( .A(n9561), .ZN(n11445) );
  NOR2_X1 U11747 ( .A1(n9330), .A2(n11445), .ZN(n9319) );
  NAND2_X1 U11748 ( .A1(n13738), .A2(n9238), .ZN(n9316) );
  INV_X1 U11749 ( .A(n9311), .ZN(n9312) );
  NAND2_X1 U11750 ( .A1(n9312), .A2(n13734), .ZN(n9313) );
  NAND2_X1 U11751 ( .A1(n9314), .A2(n13580), .ZN(n9315) );
  NAND2_X1 U11752 ( .A1(n9316), .A2(n9315), .ZN(n9321) );
  INV_X1 U11753 ( .A(n9321), .ZN(n9332) );
  INV_X1 U11754 ( .A(n9320), .ZN(n9317) );
  NAND2_X1 U11755 ( .A1(n9317), .A2(n9762), .ZN(n9323) );
  NOR3_X1 U11756 ( .A1(n9332), .A2(n11445), .A3(n9323), .ZN(n9327) );
  NAND2_X1 U11757 ( .A1(n9320), .A2(n9561), .ZN(n9329) );
  AOI211_X1 U11758 ( .C1(n9326), .C2(n9321), .A(n9329), .B(n9324), .ZN(n9322)
         );
  NAND2_X1 U11759 ( .A1(n9355), .A2(n9322), .ZN(n9353) );
  NAND3_X1 U11760 ( .A1(n9328), .A2(n9327), .A3(n9326), .ZN(n9350) );
  INV_X1 U11761 ( .A(n9329), .ZN(n9331) );
  NAND4_X1 U11762 ( .A1(n9333), .A2(n9332), .A3(n9331), .A4(n9330), .ZN(n9349)
         );
  AND2_X1 U11763 ( .A1(n11020), .A2(n10556), .ZN(n9757) );
  NAND2_X1 U11764 ( .A1(n9341), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9336) );
  MUX2_X1 U11765 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9336), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n9337) );
  INV_X1 U11766 ( .A(n9338), .ZN(n9339) );
  NAND2_X1 U11767 ( .A1(n9339), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9340) );
  MUX2_X1 U11768 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9340), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9342) );
  NAND2_X1 U11769 ( .A1(n9342), .A2(n9341), .ZN(n11614) );
  NOR2_X1 U11770 ( .A1(n14015), .A2(n11614), .ZN(n9343) );
  NAND2_X1 U11771 ( .A1(n9344), .A2(n9754), .ZN(n9744) );
  INV_X1 U11772 ( .A(n8847), .ZN(n9599) );
  INV_X1 U11773 ( .A(n9911), .ZN(n9346) );
  AND2_X2 U11774 ( .A1(n9346), .A2(n9760), .ZN(n14131) );
  NAND3_X1 U11775 ( .A1(n10034), .A2(n9599), .A3(n14131), .ZN(n9347) );
  OAI211_X1 U11776 ( .C1(n14017), .C2(n11445), .A(n9347), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9348) );
  OAI211_X1 U11777 ( .C1(n9355), .C2(n9354), .A(n9353), .B(n9352), .ZN(
        P1_U3242) );
  NAND2_X1 U11778 ( .A1(n9357), .A2(n7366), .ZN(n9365) );
  NOR2_X1 U11779 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n14011), .ZN(n9359) );
  OAI22_X1 U11780 ( .A1(n9359), .A2(n9358), .B1(P2_DATAO_REG_28__SCAN_IN), 
        .B2(n13439), .ZN(n12064) );
  AOI22_X1 U11781 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n14007), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n13434), .ZN(n12065) );
  INV_X1 U11782 ( .A(n12065), .ZN(n9360) );
  XNOR2_X1 U11783 ( .A(n12064), .B(n9360), .ZN(n12873) );
  NAND2_X1 U11784 ( .A1(n12873), .A2(n8353), .ZN(n9363) );
  OR2_X1 U11785 ( .A1(n9361), .A2(n12875), .ZN(n9362) );
  NAND2_X1 U11786 ( .A1(n9363), .A2(n9362), .ZN(n9377) );
  NAND2_X1 U11787 ( .A1(n9377), .A2(n12451), .ZN(n12292) );
  NAND2_X1 U11788 ( .A1(n12297), .A2(n12292), .ZN(n12135) );
  INV_X1 U11789 ( .A(n12135), .ZN(n9364) );
  XNOR2_X1 U11790 ( .A(n9365), .B(n9364), .ZN(n9366) );
  NAND2_X1 U11791 ( .A1(n9366), .A2(n12768), .ZN(n9374) );
  INV_X1 U11792 ( .A(n12419), .ZN(n12535) );
  INV_X1 U11793 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n12644) );
  NAND2_X1 U11794 ( .A1(n12082), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9368) );
  NAND2_X1 U11795 ( .A1(n12083), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9367) );
  OAI211_X1 U11796 ( .C1(n12087), .C2(n12644), .A(n9368), .B(n9367), .ZN(n9369) );
  INV_X1 U11797 ( .A(n9369), .ZN(n9370) );
  NAND2_X1 U11798 ( .A1(n12090), .A2(n9370), .ZN(n12534) );
  INV_X1 U11799 ( .A(P3_B_REG_SCAN_IN), .ZN(n9371) );
  NOR2_X1 U11800 ( .A1(n6630), .A2(n9371), .ZN(n9372) );
  NOR2_X1 U11801 ( .A1(n14760), .A2(n9372), .ZN(n12638) );
  AOI22_X1 U11802 ( .A1(n12535), .A2(n12763), .B1(n12534), .B2(n12638), .ZN(
        n9373) );
  INV_X1 U11803 ( .A(n12291), .ZN(n9375) );
  NAND2_X1 U11804 ( .A1(n9495), .A2(n14846), .ZN(n9381) );
  INV_X1 U11805 ( .A(n9377), .ZN(n12075) );
  NOR2_X1 U11806 ( .A1(n12075), .A2(n12826), .ZN(n9378) );
  NOR2_X1 U11807 ( .A1(n9378), .A2(n9379), .ZN(n9380) );
  NAND2_X1 U11808 ( .A1(n9381), .A2(n9380), .ZN(P3_U3488) );
  INV_X1 U11809 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9462) );
  INV_X1 U11810 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n9382) );
  XOR2_X1 U11811 ( .A(n9382), .B(P1_ADDR_REG_14__SCAN_IN), .Z(n9463) );
  INV_X1 U11812 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9408) );
  INV_X1 U11813 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n9406) );
  XOR2_X1 U11814 ( .A(n9406), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n9459) );
  INV_X1 U11815 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n9404) );
  INV_X1 U11816 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9413) );
  XOR2_X1 U11817 ( .A(n9400), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n9451) );
  INV_X1 U11818 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14728) );
  INV_X1 U11819 ( .A(n9424), .ZN(n9423) );
  NOR2_X1 U11820 ( .A1(n9385), .A2(n9384), .ZN(n9386) );
  NOR2_X1 U11821 ( .A1(n9388), .A2(n14650), .ZN(n9390) );
  NOR2_X1 U11822 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n9418), .ZN(n9389) );
  INV_X1 U11823 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n14668) );
  NOR2_X1 U11824 ( .A1(n9391), .A2(n14668), .ZN(n9393) );
  INV_X1 U11825 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9439) );
  NOR2_X1 U11826 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n9439), .ZN(n9394) );
  NOR2_X1 U11827 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n9395), .ZN(n9397) );
  XNOR2_X1 U11828 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n9395), .ZN(n9443) );
  INV_X1 U11829 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9444) );
  INV_X1 U11830 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9601) );
  XNOR2_X1 U11831 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n9601), .ZN(n9416) );
  NAND2_X1 U11832 ( .A1(n9451), .A2(n9450), .ZN(n9399) );
  NOR2_X1 U11833 ( .A1(n9413), .A2(n9414), .ZN(n9402) );
  INV_X1 U11834 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n10662) );
  NAND2_X1 U11835 ( .A1(n9413), .A2(n9414), .ZN(n9401) );
  XNOR2_X1 U11836 ( .A(n9404), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n9411) );
  NAND2_X1 U11837 ( .A1(n9459), .A2(n9458), .ZN(n9405) );
  INV_X1 U11838 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14947) );
  NAND2_X1 U11839 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14947), .ZN(n9407) );
  XOR2_X1 U11840 ( .A(n9463), .B(n9464), .Z(n14257) );
  XNOR2_X1 U11841 ( .A(n14947), .B(P1_ADDR_REG_13__SCAN_IN), .ZN(n9409) );
  XOR2_X1 U11842 ( .A(n9410), .B(n9409), .Z(n14251) );
  INV_X1 U11843 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n9457) );
  XOR2_X1 U11844 ( .A(n9412), .B(n9411), .Z(n14245) );
  XOR2_X1 U11845 ( .A(n9413), .B(P3_ADDR_REG_10__SCAN_IN), .Z(n9415) );
  XNOR2_X1 U11846 ( .A(n9415), .B(n9414), .ZN(n14046) );
  XOR2_X1 U11847 ( .A(n9417), .B(n9416), .Z(n9449) );
  XNOR2_X1 U11848 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n9418), .ZN(n9419) );
  NAND2_X1 U11849 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n9419), .ZN(n9432) );
  XOR2_X1 U11850 ( .A(n9419), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n14996) );
  INV_X1 U11851 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9429) );
  XNOR2_X1 U11852 ( .A(n9421), .B(n9420), .ZN(n14027) );
  XNOR2_X1 U11853 ( .A(n9423), .B(n9422), .ZN(n9425) );
  NAND2_X1 U11854 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n9425), .ZN(n9427) );
  AOI21_X1 U11855 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14613), .A(n9424), .ZN(
        n14999) );
  INV_X1 U11856 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n14998) );
  NOR2_X1 U11857 ( .A1(n14999), .A2(n14998), .ZN(n15008) );
  XOR2_X1 U11858 ( .A(n9425), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n15007) );
  NAND2_X1 U11859 ( .A1(n15008), .A2(n15007), .ZN(n9426) );
  NAND2_X1 U11860 ( .A1(n9427), .A2(n9426), .ZN(n14028) );
  NAND2_X1 U11861 ( .A1(n14027), .A2(n14028), .ZN(n9428) );
  NOR2_X1 U11862 ( .A1(n14027), .A2(n14028), .ZN(n14026) );
  AOI21_X1 U11863 ( .B1(n9429), .B2(n9428), .A(n14026), .ZN(n15003) );
  XNOR2_X1 U11864 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n9430), .ZN(n15004) );
  NOR2_X1 U11865 ( .A1(n15003), .A2(n15004), .ZN(n9431) );
  INV_X1 U11866 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15005) );
  NAND2_X1 U11867 ( .A1(n15003), .A2(n15004), .ZN(n15002) );
  OAI21_X1 U11868 ( .B1(n9431), .B2(n15005), .A(n15002), .ZN(n14995) );
  INV_X1 U11869 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n13653) );
  NOR2_X1 U11870 ( .A1(n9435), .A2(n9434), .ZN(n9437) );
  NOR2_X1 U11871 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n14997), .ZN(n9436) );
  NAND2_X1 U11872 ( .A1(n9438), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9442) );
  XOR2_X1 U11873 ( .A(n9439), .B(P3_ADDR_REG_6__SCAN_IN), .Z(n9441) );
  XOR2_X1 U11874 ( .A(n9441), .B(n9440), .Z(n14034) );
  XOR2_X1 U11875 ( .A(n9444), .B(n9443), .Z(n15001) );
  NAND2_X1 U11876 ( .A1(n15000), .A2(n15001), .ZN(n9447) );
  NAND2_X1 U11877 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n9445), .ZN(n9446) );
  XNOR2_X1 U11878 ( .A(n9451), .B(n9450), .ZN(n9452) );
  NAND2_X1 U11879 ( .A1(n9454), .A2(n9452), .ZN(n9455) );
  INV_X1 U11880 ( .A(n9452), .ZN(n9453) );
  INV_X1 U11881 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14047) );
  NAND2_X1 U11882 ( .A1(n14244), .A2(n14245), .ZN(n9456) );
  XNOR2_X1 U11883 ( .A(n9459), .B(n9458), .ZN(n14248) );
  INV_X1 U11884 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14498) );
  NOR2_X1 U11885 ( .A1(n14251), .A2(n14252), .ZN(n9460) );
  INV_X1 U11886 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14253) );
  OAI21_X2 U11887 ( .B1(n9460), .B2(n14253), .A(n14250), .ZN(n14256) );
  NAND2_X1 U11888 ( .A1(n14257), .A2(n14256), .ZN(n9461) );
  NOR2_X1 U11889 ( .A1(n14257), .A2(n14256), .ZN(n14255) );
  AOI21_X1 U11890 ( .B1(n9462), .B2(n9461), .A(n14255), .ZN(n9468) );
  INV_X1 U11891 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14279) );
  XOR2_X1 U11892 ( .A(n14279), .B(P3_ADDR_REG_15__SCAN_IN), .Z(n9467) );
  INV_X1 U11893 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9466) );
  NAND2_X1 U11894 ( .A1(n9464), .A2(n9463), .ZN(n9465) );
  XOR2_X1 U11895 ( .A(n9467), .B(n9471), .Z(n9469) );
  NOR2_X1 U11896 ( .A1(n9468), .A2(n9469), .ZN(n14260) );
  NOR2_X1 U11897 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n14259), .ZN(n9470) );
  NOR2_X1 U11898 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14279), .ZN(n9472) );
  INV_X1 U11899 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n12574) );
  OAI22_X1 U11900 ( .A1(n9472), .A2(n9471), .B1(P1_ADDR_REG_15__SCAN_IN), .B2(
        n12574), .ZN(n9478) );
  INV_X1 U11901 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14929) );
  XNOR2_X1 U11902 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n14929), .ZN(n9473) );
  XOR2_X1 U11903 ( .A(n9478), .B(n9473), .Z(n9474) );
  NOR2_X1 U11904 ( .A1(n9475), .A2(n9474), .ZN(n14263) );
  AND2_X1 U11905 ( .A1(n14929), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n9479) );
  OAI22_X1 U11906 ( .A1(n9479), .A2(n9478), .B1(P3_ADDR_REG_16__SCAN_IN), .B2(
        n14929), .ZN(n9481) );
  XOR2_X1 U11907 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n9481), .Z(n9482) );
  XNOR2_X1 U11908 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n9482), .ZN(n14051) );
  INV_X1 U11909 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14052) );
  NAND2_X1 U11910 ( .A1(n14050), .A2(n14051), .ZN(n14049) );
  OAI21_X2 U11911 ( .B1(n9480), .B2(n14052), .A(n14049), .ZN(n9486) );
  INV_X1 U11912 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n9487) );
  NOR2_X1 U11913 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n9481), .ZN(n9484) );
  XNOR2_X1 U11914 ( .A(n9487), .B(n9488), .ZN(n9489) );
  XNOR2_X1 U11915 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(n9489), .ZN(n9485) );
  NOR2_X1 U11916 ( .A1(n9488), .A2(n9487), .ZN(n9491) );
  NOR2_X1 U11917 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9489), .ZN(n9490) );
  NOR2_X1 U11918 ( .A1(n9491), .A2(n9490), .ZN(n9493) );
  XNOR2_X1 U11919 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9492) );
  INV_X1 U11920 ( .A(n9964), .ZN(n9496) );
  OR2_X2 U11921 ( .A1(n9754), .A2(n9546), .ZN(n13615) );
  INV_X1 U11922 ( .A(n13615), .ZN(P1_U4016) );
  INV_X1 U11923 ( .A(n9634), .ZN(n9632) );
  OR3_X2 U11924 ( .A1(n9633), .A2(n9632), .A3(P2_U3088), .ZN(n13072) );
  INV_X1 U11925 ( .A(n13072), .ZN(P2_U3947) );
  NAND2_X1 U11926 ( .A1(n9498), .A2(P3_U3151), .ZN(n9499) );
  OAI21_X1 U11927 ( .B1(n10321), .B2(P3_U3151), .A(n9499), .ZN(P3_U3295) );
  AND2_X1 U11928 ( .A1(n9501), .A2(P2_U3088), .ZN(n13436) );
  INV_X2 U11929 ( .A(n13436), .ZN(n13444) );
  AND2_X1 U11930 ( .A1(n9504), .A2(P2_U3088), .ZN(n13431) );
  INV_X2 U11931 ( .A(n13431), .ZN(n12041) );
  OAI222_X1 U11932 ( .A1(n13444), .A2(n9506), .B1(n9647), .B2(P2_U3088), .C1(
        n7413), .C2(n12041), .ZN(P2_U3326) );
  INV_X1 U11933 ( .A(n14038), .ZN(n12880) );
  INV_X1 U11934 ( .A(n9500), .ZN(n9503) );
  AND2_X1 U11935 ( .A1(n9501), .A2(P3_U3151), .ZN(n14037) );
  INV_X2 U11936 ( .A(n14037), .ZN(n12874) );
  OAI222_X1 U11937 ( .A1(n12880), .A2(n9503), .B1(n12874), .B2(n9502), .C1(
        P3_U3151), .C2(n10491), .ZN(P3_U3294) );
  NOR2_X1 U11938 ( .A1(n9504), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14000) );
  INV_X2 U11939 ( .A(n14000), .ZN(n14012) );
  INV_X1 U11940 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9507) );
  AND2_X1 U11941 ( .A1(n9505), .A2(P1_U3086), .ZN(n11443) );
  OAI222_X1 U11942 ( .A1(P1_U3086), .A2(n13605), .B1(n14012), .B2(n9507), .C1(
        n14014), .C2(n9506), .ZN(P1_U3354) );
  INV_X1 U11943 ( .A(n9508), .ZN(n9510) );
  OAI222_X1 U11944 ( .A1(P3_U3151), .A2(n10637), .B1(n12880), .B2(n9510), .C1(
        n9509), .C2(n12874), .ZN(P3_U3289) );
  INV_X1 U11945 ( .A(SI_3_), .ZN(n9511) );
  OAI222_X1 U11946 ( .A1(n10644), .A2(P3_U3151), .B1(n12880), .B2(n9512), .C1(
        n9511), .C2(n12874), .ZN(P3_U3292) );
  INV_X1 U11947 ( .A(SI_2_), .ZN(n9513) );
  OAI222_X1 U11948 ( .A1(n10641), .A2(P3_U3151), .B1(n12880), .B2(n9514), .C1(
        n9513), .C2(n12874), .ZN(P3_U3293) );
  INV_X1 U11949 ( .A(SI_7_), .ZN(n9515) );
  OAI222_X1 U11950 ( .A1(n14697), .A2(P3_U3151), .B1(n12880), .B2(n9516), .C1(
        n9515), .C2(n12874), .ZN(P3_U3288) );
  INV_X1 U11951 ( .A(n14647), .ZN(n10639) );
  INV_X1 U11952 ( .A(SI_4_), .ZN(n9517) );
  OAI222_X1 U11953 ( .A1(n10639), .A2(P3_U3151), .B1(n12880), .B2(n9518), .C1(
        n9517), .C2(n12874), .ZN(P3_U3291) );
  INV_X1 U11954 ( .A(SI_5_), .ZN(n9519) );
  OAI222_X1 U11955 ( .A1(n10648), .A2(P3_U3151), .B1(n12880), .B2(n9520), .C1(
        n9519), .C2(n12874), .ZN(P3_U3290) );
  INV_X1 U11956 ( .A(n13623), .ZN(n9594) );
  OAI222_X1 U11957 ( .A1(n14012), .A2(n9521), .B1(n14014), .B2(n9529), .C1(
        P1_U3086), .C2(n9594), .ZN(P1_U3353) );
  INV_X1 U11958 ( .A(n9522), .ZN(n9523) );
  OAI222_X1 U11959 ( .A1(P3_U3151), .A2(n10636), .B1(n12874), .B2(n9524), .C1(
        n12880), .C2(n9523), .ZN(P3_U3287) );
  INV_X1 U11960 ( .A(SI_9_), .ZN(n9526) );
  OAI222_X1 U11961 ( .A1(P3_U3151), .A2(n14739), .B1(n12874), .B2(n9526), .C1(
        n12880), .C2(n9525), .ZN(P3_U3286) );
  INV_X1 U11962 ( .A(n9527), .ZN(n9531) );
  OAI222_X1 U11963 ( .A1(n14012), .A2(n9528), .B1(n14014), .B2(n9531), .C1(
        P1_U3086), .C2(n9772), .ZN(P1_U3352) );
  OAI222_X1 U11964 ( .A1(n12041), .A2(n9530), .B1(n13444), .B2(n9529), .C1(
        P2_U3088), .C2(n9653), .ZN(P2_U3325) );
  INV_X1 U11965 ( .A(n9656), .ZN(n14425) );
  OAI222_X1 U11966 ( .A1(n12041), .A2(n9532), .B1(n13444), .B2(n9531), .C1(
        P2_U3088), .C2(n14425), .ZN(P2_U3324) );
  INV_X1 U11967 ( .A(n9533), .ZN(n9535) );
  OAI222_X1 U11968 ( .A1(n14012), .A2(n9534), .B1(n14014), .B2(n9535), .C1(
        P1_U3086), .C2(n13640), .ZN(P1_U3351) );
  INV_X1 U11969 ( .A(n9659), .ZN(n9799) );
  OAI222_X1 U11970 ( .A1(n12041), .A2(n9536), .B1(n13444), .B2(n9535), .C1(
        P2_U3088), .C2(n9799), .ZN(P2_U3323) );
  OAI222_X1 U11971 ( .A1(P3_U3151), .A2(n11302), .B1(n12874), .B2(n9538), .C1(
        n12880), .C2(n9537), .ZN(P3_U3284) );
  INV_X1 U11972 ( .A(n9539), .ZN(n9541) );
  OAI222_X1 U11973 ( .A1(n12041), .A2(n9540), .B1(n13444), .B2(n9541), .C1(
        P2_U3088), .C2(n9672), .ZN(P2_U3322) );
  OAI222_X1 U11974 ( .A1(n14012), .A2(n9542), .B1(n14014), .B2(n9541), .C1(
        P1_U3086), .C2(n9609), .ZN(P1_U3350) );
  NAND2_X1 U11975 ( .A1(n11614), .A2(P1_B_REG_SCAN_IN), .ZN(n9543) );
  OR2_X1 U11976 ( .A1(n11534), .A2(n9543), .ZN(n9545) );
  INV_X1 U11977 ( .A(P1_B_REG_SCAN_IN), .ZN(n11881) );
  NAND2_X1 U11978 ( .A1(n11534), .A2(n11881), .ZN(n9544) );
  INV_X1 U11979 ( .A(n9763), .ZN(n9766) );
  OR2_X1 U11980 ( .A1(n9740), .A2(n9766), .ZN(n14320) );
  INV_X1 U11981 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9728) );
  AND2_X1 U11982 ( .A1(n14015), .A2(n11614), .ZN(n9727) );
  AOI22_X1 U11983 ( .A1(n14320), .A2(n9728), .B1(n9549), .B2(n9727), .ZN(
        P1_U3446) );
  INV_X1 U11984 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9739) );
  INV_X1 U11985 ( .A(n9741), .ZN(n9548) );
  AOI22_X1 U11986 ( .A1(n14320), .A2(n9739), .B1(n9549), .B2(n9548), .ZN(
        P1_U3445) );
  INV_X1 U11987 ( .A(n9550), .ZN(n9551) );
  OAI222_X1 U11988 ( .A1(P3_U3151), .A2(n11469), .B1(n12874), .B2(n14938), 
        .C1(n12880), .C2(n9551), .ZN(P3_U3283) );
  INV_X1 U11989 ( .A(n9552), .ZN(n9553) );
  OAI222_X1 U11990 ( .A1(n14012), .A2(n14864), .B1(n14014), .B2(n9553), .C1(
        P1_U3086), .C2(n9717), .ZN(P1_U3349) );
  INV_X1 U11991 ( .A(n9947), .ZN(n9687) );
  OAI222_X1 U11992 ( .A1(n12041), .A2(n9554), .B1(n13444), .B2(n9553), .C1(
        P2_U3088), .C2(n9687), .ZN(P2_U3321) );
  INV_X1 U11993 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9556) );
  INV_X1 U11994 ( .A(n9555), .ZN(n9557) );
  INV_X1 U11995 ( .A(n9951), .ZN(n14440) );
  OAI222_X1 U11996 ( .A1(n12041), .A2(n9556), .B1(n13444), .B2(n9557), .C1(
        P2_U3088), .C2(n14440), .ZN(P2_U3320) );
  OAI222_X1 U11997 ( .A1(n14012), .A2(n9558), .B1(n14014), .B2(n9557), .C1(
        P1_U3086), .C2(n9813), .ZN(P1_U3348) );
  OR2_X1 U11998 ( .A1(n9911), .A2(n9743), .ZN(n9560) );
  NAND2_X1 U11999 ( .A1(n9560), .A2(n9559), .ZN(n9576) );
  AND2_X1 U12000 ( .A1(n9576), .A2(n9577), .ZN(n13708) );
  NOR2_X1 U12001 ( .A1(n13708), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12002 ( .A(n9563), .ZN(n9564) );
  AOI22_X1 U12003 ( .A1(n14965), .A2(n9565), .B1(n9564), .B2(n9567), .ZN(
        P3_U3376) );
  INV_X1 U12004 ( .A(n9566), .ZN(n9568) );
  AOI22_X1 U12005 ( .A1(n14965), .A2(n9569), .B1(n9568), .B2(n9567), .ZN(
        P3_U3377) );
  INV_X1 U12006 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9571) );
  INV_X1 U12007 ( .A(n9570), .ZN(n9572) );
  INV_X1 U12008 ( .A(n9954), .ZN(n14451) );
  OAI222_X1 U12009 ( .A1(n12041), .A2(n9571), .B1(n13444), .B2(n9572), .C1(
        P2_U3088), .C2(n14451), .ZN(P2_U3319) );
  OAI222_X1 U12010 ( .A1(n14012), .A2(n9573), .B1(n14014), .B2(n9572), .C1(
        P1_U3086), .C2(n9617), .ZN(P1_U3347) );
  OAI222_X1 U12011 ( .A1(n11640), .A2(P3_U3151), .B1(n12880), .B2(n9575), .C1(
        n9574), .C2(n12874), .ZN(P3_U3282) );
  AND2_X1 U12012 ( .A1(n14965), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12013 ( .A1(n14965), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12014 ( .A1(n14965), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12015 ( .A1(n14965), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12016 ( .A1(n14965), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12017 ( .A1(n14965), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12018 ( .A1(n14965), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12019 ( .A1(n14965), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12020 ( .A1(n14965), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12021 ( .A1(n14965), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12022 ( .A1(n14965), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12023 ( .A1(n14965), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12024 ( .A1(n14965), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12025 ( .A1(n14965), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12026 ( .A1(n14965), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U12027 ( .A1(n14965), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12028 ( .A1(n14965), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12029 ( .A1(n14965), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12030 ( .A1(n14965), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12031 ( .A1(n14965), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12032 ( .A1(n14965), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12033 ( .A1(n14965), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12034 ( .A1(n14965), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12035 ( .A1(n14965), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12036 ( .A1(n14965), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12037 ( .A1(n14965), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12038 ( .A1(n14965), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12039 ( .A1(n14965), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12040 ( .A1(n14965), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  INV_X1 U12041 ( .A(n13708), .ZN(n14278) );
  INV_X1 U12042 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9582) );
  INV_X1 U12043 ( .A(n9576), .ZN(n9578) );
  AND2_X1 U12044 ( .A1(n9578), .A2(n9577), .ZN(n9614) );
  INV_X1 U12045 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9753) );
  OAI21_X1 U12046 ( .B1(n8847), .B2(P1_REG2_REG_0__SCAN_IN), .A(n9760), .ZN(
        n13616) );
  AOI21_X1 U12047 ( .B1(n8847), .B2(n9753), .A(n13616), .ZN(n9579) );
  XNOR2_X1 U12048 ( .A(n9579), .B(n13617), .ZN(n9580) );
  AOI22_X1 U12049 ( .A1(n9614), .A2(n9580), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9581) );
  OAI21_X1 U12050 ( .B1(n14278), .B2(n9582), .A(n9581), .ZN(P1_U3243) );
  INV_X1 U12051 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9584) );
  INV_X1 U12052 ( .A(n9583), .ZN(n9585) );
  INV_X1 U12053 ( .A(n10424), .ZN(n10433) );
  OAI222_X1 U12054 ( .A1(n12041), .A2(n9584), .B1(n13444), .B2(n9585), .C1(
        P2_U3088), .C2(n10433), .ZN(P2_U3318) );
  OAI222_X1 U12055 ( .A1(n14012), .A2(n9586), .B1(n14014), .B2(n9585), .C1(
        P1_U3086), .C2(n9700), .ZN(P1_U3346) );
  OAI222_X1 U12056 ( .A1(P3_U3151), .A2(n12561), .B1(n12874), .B2(n9588), .C1(
        n12880), .C2(n9587), .ZN(P3_U3281) );
  INV_X1 U12057 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9590) );
  INV_X1 U12058 ( .A(n9589), .ZN(n9591) );
  INV_X1 U12059 ( .A(n10434), .ZN(n14465) );
  OAI222_X1 U12060 ( .A1(n12041), .A2(n9590), .B1(n13444), .B2(n9591), .C1(
        P2_U3088), .C2(n14465), .ZN(P2_U3317) );
  INV_X1 U12061 ( .A(n10379), .ZN(n10372) );
  OAI222_X1 U12062 ( .A1(n14012), .A2(n9592), .B1(n14014), .B2(n9591), .C1(
        P1_U3086), .C2(n10372), .ZN(P1_U3345) );
  INV_X1 U12063 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9593) );
  MUX2_X1 U12064 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9593), .S(n9617), .Z(n9598)
         );
  INV_X1 U12065 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n14385) );
  INV_X1 U12066 ( .A(n9717), .ZN(n9610) );
  INV_X1 U12067 ( .A(n9609), .ZN(n13655) );
  INV_X1 U12068 ( .A(n13640), .ZN(n9607) );
  INV_X1 U12069 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n14379) );
  MUX2_X1 U12070 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n14379), .S(n13605), .Z(
        n13603) );
  OR3_X1 U12071 ( .A1(n13603), .A2(n9753), .A3(n13617), .ZN(n13628) );
  NAND2_X1 U12072 ( .A1(n13602), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n13627) );
  INV_X1 U12073 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9940) );
  MUX2_X1 U12074 ( .A(n9940), .B(P1_REG1_REG_2__SCAN_IN), .S(n13623), .Z(
        n13626) );
  NOR2_X1 U12075 ( .A1(n9594), .A2(n9940), .ZN(n9774) );
  INV_X1 U12076 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9595) );
  MUX2_X1 U12077 ( .A(n9595), .B(P1_REG1_REG_3__SCAN_IN), .S(n9772), .Z(n9773)
         );
  OAI21_X1 U12078 ( .B1(n13625), .B2(n9774), .A(n9773), .ZN(n13636) );
  INV_X1 U12079 ( .A(n9772), .ZN(n9596) );
  NAND2_X1 U12080 ( .A1(n9596), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n13635) );
  INV_X1 U12081 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n14877) );
  MUX2_X1 U12082 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n14877), .S(n13640), .Z(
        n13634) );
  AOI21_X1 U12083 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9607), .A(n13638), .ZN(
        n13657) );
  INV_X1 U12084 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10233) );
  MUX2_X1 U12085 ( .A(n10233), .B(P1_REG1_REG_5__SCAN_IN), .S(n9609), .Z(
        n13658) );
  NAND2_X1 U12086 ( .A1(n13657), .A2(n13658), .ZN(n13656) );
  OAI21_X1 U12087 ( .B1(n13655), .B2(P1_REG1_REG_5__SCAN_IN), .A(n13656), .ZN(
        n9708) );
  INV_X1 U12088 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14383) );
  MUX2_X1 U12089 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n14383), .S(n9717), .Z(n9707) );
  AOI21_X1 U12090 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n9610), .A(n9706), .ZN(
        n9806) );
  MUX2_X1 U12091 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n14385), .S(n9813), .Z(n9805) );
  OAI21_X1 U12092 ( .B1(n14385), .B2(n9813), .A(n9807), .ZN(n9597) );
  NOR2_X1 U12093 ( .A1(n9597), .A2(n9598), .ZN(n9697) );
  AOI21_X1 U12094 ( .B1(n9598), .B2(n9597), .A(n9697), .ZN(n9623) );
  NOR2_X2 U12095 ( .A1(n9600), .A2(n9599), .ZN(n13726) );
  INV_X1 U12096 ( .A(n9617), .ZN(n9694) );
  NAND2_X1 U12097 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11254) );
  OAI21_X1 U12098 ( .B1(n14278), .B2(n9601), .A(n11254), .ZN(n9602) );
  AOI21_X1 U12099 ( .B1(n9694), .B2(n13723), .A(n9602), .ZN(n9622) );
  NAND2_X1 U12100 ( .A1(n13602), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9604) );
  INV_X1 U12101 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n13606) );
  NAND2_X1 U12102 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13614) );
  AOI21_X1 U12103 ( .B1(n13605), .B2(n13606), .A(n13614), .ZN(n9603) );
  NAND2_X1 U12104 ( .A1(n9604), .A2(n9603), .ZN(n13609) );
  NAND2_X1 U12105 ( .A1(n13609), .A2(n9604), .ZN(n13621) );
  INV_X1 U12106 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9605) );
  XNOR2_X1 U12107 ( .A(n13623), .B(n9605), .ZN(n13620) );
  AOI22_X1 U12108 ( .A1(n13621), .A2(n13620), .B1(P1_REG2_REG_2__SCAN_IN), 
        .B2(n13623), .ZN(n9778) );
  INV_X1 U12109 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9606) );
  MUX2_X1 U12110 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9606), .S(n9772), .Z(n9777)
         );
  NOR2_X1 U12111 ( .A1(n9778), .A2(n9777), .ZN(n13643) );
  NOR2_X1 U12112 ( .A1(n9772), .A2(n9606), .ZN(n13642) );
  INV_X1 U12113 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10118) );
  MUX2_X1 U12114 ( .A(n10118), .B(P1_REG2_REG_4__SCAN_IN), .S(n13640), .Z(
        n13641) );
  OAI21_X1 U12115 ( .B1(n13643), .B2(n13642), .A(n13641), .ZN(n13663) );
  NAND2_X1 U12116 ( .A1(n9607), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n13662) );
  INV_X1 U12117 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9608) );
  MUX2_X1 U12118 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9608), .S(n9609), .Z(n13661) );
  AOI21_X1 U12119 ( .B1(n13663), .B2(n13662), .A(n13661), .ZN(n13660) );
  NOR2_X1 U12120 ( .A1(n9609), .A2(n9608), .ZN(n9710) );
  INV_X1 U12121 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10154) );
  MUX2_X1 U12122 ( .A(n10154), .B(P1_REG2_REG_6__SCAN_IN), .S(n9717), .Z(n9709) );
  OAI21_X1 U12123 ( .B1(n13660), .B2(n9710), .A(n9709), .ZN(n9802) );
  NAND2_X1 U12124 ( .A1(n9610), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9801) );
  INV_X1 U12125 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10363) );
  MUX2_X1 U12126 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10363), .S(n9813), .Z(n9800) );
  AOI21_X1 U12127 ( .B1(n9802), .B2(n9801), .A(n9800), .ZN(n9615) );
  NOR2_X1 U12128 ( .A1(n9813), .A2(n10363), .ZN(n9616) );
  INV_X1 U12129 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9611) );
  MUX2_X1 U12130 ( .A(n9611), .B(P1_REG2_REG_8__SCAN_IN), .S(n9617), .Z(n9612)
         );
  OAI21_X1 U12131 ( .B1(n9615), .B2(n9616), .A(n9612), .ZN(n9692) );
  NOR2_X1 U12132 ( .A1(n8847), .A2(n14009), .ZN(n9613) );
  NAND2_X1 U12133 ( .A1(n9614), .A2(n9613), .ZN(n14270) );
  INV_X1 U12134 ( .A(n9615), .ZN(n9804) );
  INV_X1 U12135 ( .A(n9616), .ZN(n9619) );
  MUX2_X1 U12136 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n9611), .S(n9617), .Z(n9618)
         );
  NAND3_X1 U12137 ( .A1(n9804), .A2(n9619), .A3(n9618), .ZN(n9620) );
  NAND3_X1 U12138 ( .A1(n9692), .A2(n13725), .A3(n9620), .ZN(n9621) );
  OAI211_X1 U12139 ( .C1(n9623), .C2(n14272), .A(n9622), .B(n9621), .ZN(
        P1_U3251) );
  INV_X2 U12140 ( .A(n11443), .ZN(n14014) );
  INV_X1 U12141 ( .A(n9624), .ZN(n9626) );
  INV_X1 U12142 ( .A(n13674), .ZN(n10380) );
  OAI222_X1 U12143 ( .A1(n14012), .A2(n9625), .B1(n14014), .B2(n9626), .C1(
        P1_U3086), .C2(n10380), .ZN(P1_U3344) );
  INV_X1 U12144 ( .A(n10441), .ZN(n10422) );
  OAI222_X1 U12145 ( .A1(n12041), .A2(n9627), .B1(n13444), .B2(n9626), .C1(
        P2_U3088), .C2(n10422), .ZN(P2_U3316) );
  INV_X1 U12146 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n14897) );
  NAND2_X1 U12147 ( .A1(n12181), .A2(P3_U3897), .ZN(n9628) );
  OAI21_X1 U12148 ( .B1(P3_U3897), .B2(n14897), .A(n9628), .ZN(P3_U3495) );
  INV_X1 U12149 ( .A(n9629), .ZN(n9630) );
  OAI222_X1 U12150 ( .A1(P3_U3151), .A2(n12593), .B1(n12874), .B2(n9631), .C1(
        n12880), .C2(n9630), .ZN(P3_U3280) );
  OR2_X1 U12151 ( .A1(n9633), .A2(n9632), .ZN(n9637) );
  NAND2_X1 U12152 ( .A1(n9634), .A2(n10017), .ZN(n9635) );
  NAND2_X1 U12153 ( .A1(n9635), .A2(n7434), .ZN(n9636) );
  NAND2_X1 U12154 ( .A1(n9664), .A2(n8181), .ZN(n14392) );
  OR2_X1 U12155 ( .A1(n9664), .A2(P2_U3088), .ZN(n14497) );
  OR2_X1 U12156 ( .A1(n8181), .A2(P2_U3088), .ZN(n13437) );
  NOR2_X1 U12157 ( .A1(n13437), .A2(n8183), .ZN(n9638) );
  INV_X1 U12158 ( .A(n9653), .ZN(n14411) );
  INV_X1 U12159 ( .A(n9647), .ZN(n14395) );
  INV_X1 U12160 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10996) );
  MUX2_X1 U12161 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10996), .S(n9653), .Z(
        n14416) );
  NOR2_X1 U12162 ( .A1(n14417), .A2(n14416), .ZN(n14415) );
  INV_X1 U12163 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9639) );
  MUX2_X1 U12164 ( .A(n9639), .B(P2_REG2_REG_3__SCAN_IN), .S(n9656), .Z(n14428) );
  INV_X1 U12165 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9640) );
  MUX2_X1 U12166 ( .A(n9640), .B(P2_REG2_REG_4__SCAN_IN), .S(n9659), .Z(n9792)
         );
  AOI21_X1 U12167 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n9659), .A(n9791), .ZN(
        n9643) );
  INV_X1 U12168 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9641) );
  MUX2_X1 U12169 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n9641), .S(n9672), .Z(n9642)
         );
  NAND2_X1 U12170 ( .A1(n9643), .A2(n9642), .ZN(n9644) );
  NAND3_X1 U12171 ( .A1(n14526), .A2(n9682), .A3(n9644), .ZN(n9668) );
  INV_X1 U12172 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9645) );
  MUX2_X1 U12173 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9645), .S(n9656), .Z(n14432) );
  XNOR2_X1 U12174 ( .A(n9653), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n14412) );
  INV_X1 U12175 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9646) );
  OR2_X1 U12176 ( .A1(n9647), .A2(n9646), .ZN(n9651) );
  NAND2_X1 U12177 ( .A1(n9647), .A2(n9646), .ZN(n9648) );
  NAND2_X1 U12178 ( .A1(n9651), .A2(n9648), .ZN(n14396) );
  INV_X1 U12179 ( .A(n14396), .ZN(n9650) );
  AND2_X1 U12180 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9649) );
  NAND2_X1 U12181 ( .A1(n9650), .A2(n9649), .ZN(n14400) );
  NAND2_X1 U12182 ( .A1(n14400), .A2(n9651), .ZN(n14413) );
  NAND2_X1 U12183 ( .A1(n14412), .A2(n14413), .ZN(n9655) );
  INV_X1 U12184 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9652) );
  OR2_X1 U12185 ( .A1(n9653), .A2(n9652), .ZN(n9654) );
  NAND2_X1 U12186 ( .A1(n9655), .A2(n9654), .ZN(n14433) );
  NAND2_X1 U12187 ( .A1(n14432), .A2(n14433), .ZN(n14431) );
  NAND2_X1 U12188 ( .A1(n9656), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9657) );
  NAND2_X1 U12189 ( .A1(n14431), .A2(n9657), .ZN(n9790) );
  INV_X1 U12190 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9658) );
  MUX2_X1 U12191 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9658), .S(n9659), .Z(n9789)
         );
  NAND2_X1 U12192 ( .A1(n9790), .A2(n9789), .ZN(n9788) );
  NAND2_X1 U12193 ( .A1(n9659), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9660) );
  NAND2_X1 U12194 ( .A1(n9788), .A2(n9660), .ZN(n9666) );
  INV_X1 U12195 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9661) );
  MUX2_X1 U12196 ( .A(n9661), .B(P2_REG1_REG_5__SCAN_IN), .S(n9672), .Z(n9665)
         );
  INV_X1 U12197 ( .A(n8183), .ZN(n9662) );
  NOR2_X1 U12198 ( .A1(n13437), .A2(n9662), .ZN(n9663) );
  NAND2_X1 U12199 ( .A1(n9664), .A2(n9663), .ZN(n14483) );
  NAND2_X1 U12200 ( .A1(n9666), .A2(n9665), .ZN(n9674) );
  OAI211_X1 U12201 ( .C1(n9666), .C2(n9665), .A(n14542), .B(n9674), .ZN(n9667)
         );
  NAND2_X1 U12202 ( .A1(n9668), .A2(n9667), .ZN(n9670) );
  NAND2_X1 U12203 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10264) );
  INV_X1 U12204 ( .A(n10264), .ZN(n9669) );
  AOI211_X1 U12205 ( .C1(n14540), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n9670), .B(
        n9669), .ZN(n9671) );
  OAI21_X1 U12206 ( .B1(n9672), .B2(n14547), .A(n9671), .ZN(P2_U3219) );
  NAND2_X1 U12207 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n10693) );
  NAND2_X1 U12208 ( .A1(n9679), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9673) );
  NAND2_X1 U12209 ( .A1(n9674), .A2(n9673), .ZN(n9677) );
  INV_X1 U12210 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9675) );
  MUX2_X1 U12211 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9675), .S(n9947), .Z(n9676)
         );
  NAND2_X1 U12212 ( .A1(n9677), .A2(n9676), .ZN(n9949) );
  OAI211_X1 U12213 ( .C1(n9677), .C2(n9676), .A(n14542), .B(n9949), .ZN(n9678)
         );
  NAND2_X1 U12214 ( .A1(n10693), .A2(n9678), .ZN(n9685) );
  NAND2_X1 U12215 ( .A1(n9679), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9681) );
  MUX2_X1 U12216 ( .A(n10676), .B(P2_REG2_REG_6__SCAN_IN), .S(n9947), .Z(n9680) );
  AND3_X1 U12217 ( .A1(n9682), .A2(n9681), .A3(n9680), .ZN(n9683) );
  NOR3_X1 U12218 ( .A1(n9941), .A2(n9683), .A3(n14536), .ZN(n9684) );
  AOI211_X1 U12219 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n14540), .A(n9685), .B(
        n9684), .ZN(n9686) );
  OAI21_X1 U12220 ( .B1(n9687), .B2(n14547), .A(n9686), .ZN(P2_U3220) );
  NAND2_X1 U12221 ( .A1(n13012), .A2(P2_U3947), .ZN(n9688) );
  OAI21_X1 U12222 ( .B1(P2_U3947), .B2(n9689), .A(n9688), .ZN(P2_U3553) );
  NAND2_X1 U12223 ( .A1(n9694), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9691) );
  INV_X1 U12224 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10799) );
  MUX2_X1 U12225 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10799), .S(n9700), .Z(n9690) );
  AOI21_X1 U12226 ( .B1(n9692), .B2(n9691), .A(n9690), .ZN(n9818) );
  NAND3_X1 U12227 ( .A1(n9692), .A2(n9691), .A3(n9690), .ZN(n9693) );
  NAND2_X1 U12228 ( .A1(n9693), .A2(n13725), .ZN(n9705) );
  NOR2_X1 U12229 ( .A1(n9694), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9695) );
  INV_X1 U12230 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n11029) );
  MUX2_X1 U12231 ( .A(n11029), .B(P1_REG1_REG_9__SCAN_IN), .S(n9700), .Z(n9696) );
  INV_X1 U12232 ( .A(n9814), .ZN(n9699) );
  NOR3_X1 U12233 ( .A1(n9697), .A2(n9696), .A3(n9695), .ZN(n9698) );
  OAI21_X1 U12234 ( .B1(n9699), .B2(n9698), .A(n13726), .ZN(n9704) );
  INV_X1 U12235 ( .A(n9700), .ZN(n9819) );
  INV_X1 U12236 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9701) );
  NAND2_X1 U12237 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11420) );
  OAI21_X1 U12238 ( .B1(n14278), .B2(n9701), .A(n11420), .ZN(n9702) );
  AOI21_X1 U12239 ( .B1(n9819), .B2(n13723), .A(n9702), .ZN(n9703) );
  OAI211_X1 U12240 ( .C1(n9818), .C2(n9705), .A(n9704), .B(n9703), .ZN(
        P1_U3252) );
  AOI211_X1 U12241 ( .C1(n9708), .C2(n9707), .A(n9706), .B(n14272), .ZN(n9714)
         );
  INV_X1 U12242 ( .A(n9802), .ZN(n9712) );
  NOR3_X1 U12243 ( .A1(n13660), .A2(n9710), .A3(n9709), .ZN(n9711) );
  NOR3_X1 U12244 ( .A1(n14270), .A2(n9712), .A3(n9711), .ZN(n9713) );
  NOR2_X1 U12245 ( .A1(n9714), .A2(n9713), .ZN(n9716) );
  NOR2_X1 U12246 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8908), .ZN(n10883) );
  AOI21_X1 U12247 ( .B1(n13708), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10883), .ZN(
        n9715) );
  OAI211_X1 U12248 ( .C1(n9717), .C2(n14274), .A(n9716), .B(n9715), .ZN(
        P1_U3249) );
  INV_X1 U12249 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n14954) );
  NAND2_X1 U12250 ( .A1(n9718), .A2(P3_U3897), .ZN(n9719) );
  OAI21_X1 U12251 ( .B1(P3_U3897), .B2(n14954), .A(n9719), .ZN(P3_U3491) );
  INV_X1 U12252 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10220) );
  INV_X1 U12253 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n14398) );
  INV_X1 U12254 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9720) );
  NAND2_X1 U12255 ( .A1(n14526), .A2(n9720), .ZN(n9721) );
  OAI211_X1 U12256 ( .C1(n14483), .C2(P2_REG1_REG_0__SCAN_IN), .A(n14547), .B(
        n9721), .ZN(n9722) );
  INV_X1 U12257 ( .A(n9722), .ZN(n9724) );
  AOI22_X1 U12258 ( .A1(n14542), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n14526), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n9723) );
  MUX2_X1 U12259 ( .A(n9724), .B(n9723), .S(n14397), .Z(n9726) );
  NAND2_X1 U12260 ( .A1(n14540), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n9725) );
  OAI211_X1 U12261 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10220), .A(n9726), .B(
        n9725), .ZN(P2_U3214) );
  AOI21_X1 U12262 ( .B1(n9740), .B2(n9728), .A(n9727), .ZN(n9903) );
  NOR2_X1 U12263 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .ZN(
        n14980) );
  NOR4_X1 U12264 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n9731) );
  NOR4_X1 U12265 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n9730) );
  NOR4_X1 U12266 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n9729) );
  AND4_X1 U12267 ( .A1(n14980), .A2(n9731), .A3(n9730), .A4(n9729), .ZN(n9737)
         );
  NOR4_X1 U12268 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9735) );
  NOR4_X1 U12269 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n9734) );
  NOR4_X1 U12270 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9733) );
  NOR4_X1 U12271 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9732) );
  AND4_X1 U12272 ( .A1(n9735), .A2(n9734), .A3(n9733), .A4(n9732), .ZN(n9736)
         );
  NAND2_X1 U12273 ( .A1(n9737), .A2(n9736), .ZN(n9738) );
  NAND2_X1 U12274 ( .A1(n9740), .A2(n9738), .ZN(n9904) );
  NAND2_X1 U12275 ( .A1(n9903), .A2(n9904), .ZN(n10033) );
  NAND2_X1 U12276 ( .A1(n9740), .A2(n9739), .ZN(n9742) );
  NAND2_X1 U12277 ( .A1(n9742), .A2(n9741), .ZN(n9916) );
  OR2_X1 U12278 ( .A1(n10033), .A2(n9916), .ZN(n9765) );
  NAND2_X1 U12279 ( .A1(n14310), .A2(n11272), .ZN(n9905) );
  NAND2_X1 U12280 ( .A1(n9765), .A2(n9905), .ZN(n9746) );
  NOR2_X1 U12281 ( .A1(n9744), .A2(n9743), .ZN(n9745) );
  NAND2_X1 U12282 ( .A1(n9746), .A2(n9745), .ZN(n10171) );
  OR2_X1 U12283 ( .A1(n10171), .A2(P1_U3086), .ZN(n13542) );
  INV_X1 U12284 ( .A(n13542), .ZN(n9843) );
  INV_X1 U12285 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9770) );
  INV_X1 U12286 ( .A(n9754), .ZN(n9748) );
  AND2_X1 U12287 ( .A1(n9748), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n9749) );
  NAND2_X1 U12288 ( .A1(n10179), .A2(n13598), .ZN(n9752) );
  INV_X2 U12289 ( .A(n11942), .ZN(n12363) );
  NAND2_X1 U12290 ( .A1(n12363), .A2(n10098), .ZN(n9751) );
  OAI21_X1 U12291 ( .B1(n9755), .B2(n9836), .A(n9835), .ZN(n13613) );
  INV_X1 U12292 ( .A(n9756), .ZN(n9914) );
  NAND3_X1 U12293 ( .A1(n14371), .A2(n9763), .A3(n9911), .ZN(n9758) );
  NAND2_X1 U12294 ( .A1(n13613), .A2(n14139), .ZN(n9769) );
  INV_X1 U12295 ( .A(n9765), .ZN(n9759) );
  INV_X2 U12296 ( .A(n13892), .ZN(n14292) );
  NAND2_X1 U12297 ( .A1(n14141), .A2(n14292), .ZN(n13570) );
  INV_X1 U12298 ( .A(n13570), .ZN(n13541) );
  NOR2_X1 U12299 ( .A1(n9762), .A2(n14017), .ZN(n10036) );
  NAND2_X1 U12300 ( .A1(n10036), .A2(n9763), .ZN(n9764) );
  OR2_X1 U12301 ( .A1(n9765), .A2(n9764), .ZN(n9767) );
  AOI22_X1 U12302 ( .A1(n13541), .A2(n9761), .B1(n10098), .B2(n14142), .ZN(
        n9768) );
  OAI211_X1 U12303 ( .C1(n9843), .C2(n9770), .A(n9769), .B(n9768), .ZN(
        P1_U3232) );
  NAND2_X1 U12304 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10172) );
  NAND2_X1 U12305 ( .A1(n13708), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n9771) );
  OAI211_X1 U12306 ( .C1(n14274), .C2(n9772), .A(n10172), .B(n9771), .ZN(n9781) );
  INV_X1 U12307 ( .A(n13636), .ZN(n9776) );
  NOR3_X1 U12308 ( .A1(n13625), .A2(n9774), .A3(n9773), .ZN(n9775) );
  NOR3_X1 U12309 ( .A1(n14272), .A2(n9776), .A3(n9775), .ZN(n9780) );
  AOI211_X1 U12310 ( .C1(n9778), .C2(n9777), .A(n13643), .B(n14270), .ZN(n9779) );
  OR3_X1 U12311 ( .A1(n9781), .A2(n9780), .A3(n9779), .ZN(P1_U3246) );
  INV_X1 U12312 ( .A(n9782), .ZN(n9784) );
  INV_X1 U12313 ( .A(n14494), .ZN(n11454) );
  OAI222_X1 U12314 ( .A1(n13444), .A2(n9784), .B1(n11454), .B2(P2_U3088), .C1(
        n9783), .C2(n12041), .ZN(P2_U3315) );
  INV_X1 U12315 ( .A(n13694), .ZN(n10381) );
  OAI222_X1 U12316 ( .A1(n14012), .A2(n6680), .B1(n14014), .B2(n9784), .C1(
        n10381), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U12317 ( .A(n9785), .ZN(n9786) );
  OAI222_X1 U12318 ( .A1(P3_U3151), .A2(n12609), .B1(n12874), .B2(n9787), .C1(
        n12880), .C2(n9786), .ZN(P3_U3279) );
  OAI211_X1 U12319 ( .C1(n9790), .C2(n9789), .A(n14542), .B(n9788), .ZN(n9796)
         );
  AOI211_X1 U12320 ( .C1(n9793), .C2(n9792), .A(n9791), .B(n14536), .ZN(n9794)
         );
  INV_X1 U12321 ( .A(n9794), .ZN(n9795) );
  NAND2_X1 U12322 ( .A1(n9796), .A2(n9795), .ZN(n9797) );
  AND2_X1 U12323 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10495) );
  AOI211_X1 U12324 ( .C1(n14540), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n9797), .B(
        n10495), .ZN(n9798) );
  OAI21_X1 U12325 ( .B1(n9799), .B2(n14547), .A(n9798), .ZN(P2_U3218) );
  NAND3_X1 U12326 ( .A1(n9802), .A2(n9801), .A3(n9800), .ZN(n9803) );
  NAND3_X1 U12327 ( .A1(n13725), .A2(n9804), .A3(n9803), .ZN(n9812) );
  NAND2_X1 U12328 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11048) );
  AOI21_X1 U12329 ( .B1(n9806), .B2(n9805), .A(n14272), .ZN(n9808) );
  NAND2_X1 U12330 ( .A1(n9808), .A2(n9807), .ZN(n9809) );
  NAND2_X1 U12331 ( .A1(n11048), .A2(n9809), .ZN(n9810) );
  AOI21_X1 U12332 ( .B1(n13708), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n9810), .ZN(
        n9811) );
  OAI211_X1 U12333 ( .C1(n14274), .C2(n9813), .A(n9812), .B(n9811), .ZN(
        P1_U3250) );
  OAI21_X1 U12334 ( .B1(n9819), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9814), .ZN(
        n9816) );
  INV_X1 U12335 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14389) );
  MUX2_X1 U12336 ( .A(n14389), .B(P1_REG1_REG_10__SCAN_IN), .S(n10379), .Z(
        n9815) );
  AOI211_X1 U12337 ( .C1(n9816), .C2(n9815), .A(n14272), .B(n10378), .ZN(n9817) );
  INV_X1 U12338 ( .A(n9817), .ZN(n9826) );
  NAND2_X1 U12339 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n11579)
         );
  AOI21_X1 U12340 ( .B1(n9819), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9818), .ZN(
        n9821) );
  INV_X1 U12341 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10371) );
  MUX2_X1 U12342 ( .A(n10371), .B(P1_REG2_REG_10__SCAN_IN), .S(n10379), .Z(
        n9820) );
  NOR2_X1 U12343 ( .A1(n9821), .A2(n9820), .ZN(n13677) );
  AOI211_X1 U12344 ( .C1(n9821), .C2(n9820), .A(n13677), .B(n14270), .ZN(n9822) );
  INV_X1 U12345 ( .A(n9822), .ZN(n9823) );
  NAND2_X1 U12346 ( .A1(n11579), .A2(n9823), .ZN(n9824) );
  AOI21_X1 U12347 ( .B1(n13708), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n9824), .ZN(
        n9825) );
  OAI211_X1 U12348 ( .C1(n14274), .C2(n10372), .A(n9826), .B(n9825), .ZN(
        P1_U3253) );
  INV_X1 U12349 ( .A(n9827), .ZN(n9885) );
  OAI222_X1 U12350 ( .A1(n13444), .A2(n9885), .B1(n14510), .B2(P2_U3088), .C1(
        n9828), .C2(n12041), .ZN(P2_U3314) );
  INV_X1 U12351 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n13599) );
  NAND2_X1 U12352 ( .A1(n10556), .A2(n14017), .ZN(n9829) );
  NAND2_X1 U12353 ( .A1(n9747), .A2(n9829), .ZN(n9834) );
  XNOR2_X1 U12354 ( .A(n9830), .B(n9834), .ZN(n9832) );
  OAI22_X1 U12355 ( .A1(n11940), .A2(n10080), .B1(n14322), .B2(n11941), .ZN(
        n9831) );
  AND2_X1 U12356 ( .A1(n9832), .A2(n9831), .ZN(n9833) );
  NOR2_X1 U12357 ( .A1(n9832), .A2(n9831), .ZN(n10176) );
  OAI21_X1 U12358 ( .B1(n10541), .B2(n9836), .A(n9835), .ZN(n9837) );
  OAI21_X1 U12359 ( .B1(n9838), .B2(n9837), .A(n10178), .ZN(n9839) );
  NAND2_X1 U12360 ( .A1(n9839), .A2(n14139), .ZN(n9842) );
  NAND2_X1 U12361 ( .A1(n14292), .A2(n13597), .ZN(n10084) );
  OAI22_X1 U12362 ( .A1(n13513), .A2(n10084), .B1(n13579), .B2(n14322), .ZN(
        n9840) );
  AOI21_X1 U12363 ( .B1(n13557), .B2(n13598), .A(n9840), .ZN(n9841) );
  OAI211_X1 U12364 ( .C1(n9843), .C2(n13599), .A(n9842), .B(n9841), .ZN(
        P1_U3222) );
  INV_X1 U12365 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n14891) );
  INV_X1 U12366 ( .A(n12247), .ZN(n11683) );
  NAND2_X1 U12367 ( .A1(n11683), .A2(P3_U3897), .ZN(n9844) );
  OAI21_X1 U12368 ( .B1(P3_U3897), .B2(n14891), .A(n9844), .ZN(P3_U3506) );
  INV_X1 U12369 ( .A(P2_B_REG_SCAN_IN), .ZN(n12016) );
  XNOR2_X1 U12370 ( .A(n11532), .B(n12016), .ZN(n9845) );
  NAND2_X1 U12371 ( .A1(n9845), .A2(n11612), .ZN(n9846) );
  INV_X1 U12372 ( .A(n13443), .ZN(n9862) );
  NOR4_X1 U12373 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n9850) );
  NOR4_X1 U12374 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n9849) );
  NOR4_X1 U12375 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9848) );
  NOR4_X1 U12376 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9847) );
  AND4_X1 U12377 ( .A1(n9850), .A2(n9849), .A3(n9848), .A4(n9847), .ZN(n9856)
         );
  NOR2_X1 U12378 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .ZN(
        n9854) );
  NOR4_X1 U12379 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n9853) );
  NOR4_X1 U12380 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n9852) );
  NOR4_X1 U12381 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n9851) );
  AND4_X1 U12382 ( .A1(n9854), .A2(n9853), .A3(n9852), .A4(n9851), .ZN(n9855)
         );
  NAND2_X1 U12383 ( .A1(n9856), .A2(n9855), .ZN(n9857) );
  INV_X1 U12384 ( .A(n10006), .ZN(n9861) );
  INV_X1 U12385 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14554) );
  NAND2_X1 U12386 ( .A1(n14548), .A2(n14554), .ZN(n9859) );
  NAND2_X1 U12387 ( .A1(n11612), .A2(n13443), .ZN(n9858) );
  NAND2_X1 U12388 ( .A1(n9859), .A2(n9858), .ZN(n14555) );
  OR2_X2 U12389 ( .A1(n9866), .A2(n9860), .ZN(n9876) );
  NAND3_X1 U12390 ( .A1(n9861), .A2(n14555), .A3(n10011), .ZN(n9921) );
  INV_X1 U12391 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14552) );
  NAND2_X1 U12392 ( .A1(n14548), .A2(n14552), .ZN(n9864) );
  OR2_X1 U12393 ( .A1(n11532), .A2(n9862), .ZN(n9863) );
  NAND2_X1 U12394 ( .A1(n10017), .A2(n10013), .ZN(n10008) );
  AND2_X1 U12395 ( .A1(n14556), .A2(n10008), .ZN(n9865) );
  NAND2_X1 U12396 ( .A1(n10007), .A2(n9865), .ZN(n10190) );
  INV_X1 U12397 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9881) );
  INV_X1 U12398 ( .A(n10025), .ZN(n10212) );
  NAND2_X1 U12399 ( .A1(n9869), .A2(n10212), .ZN(n10024) );
  XNOR2_X1 U12400 ( .A(n9891), .B(n10024), .ZN(n11009) );
  XNOR2_X1 U12401 ( .A(n10215), .B(n9891), .ZN(n9875) );
  NAND2_X1 U12402 ( .A1(n9866), .A2(n9870), .ZN(n9871) );
  NAND2_X1 U12403 ( .A1(n10017), .A2(n8181), .ZN(n12997) );
  NAND2_X1 U12404 ( .A1(n13037), .A2(n8146), .ZN(n9874) );
  NAND2_X1 U12405 ( .A1(n13038), .A2(n9869), .ZN(n9873) );
  AND2_X1 U12406 ( .A1(n9874), .A2(n9873), .ZN(n10014) );
  OAI21_X1 U12407 ( .B1(n9875), .B2(n13268), .A(n10014), .ZN(n11007) );
  INV_X1 U12408 ( .A(n11007), .ZN(n9879) );
  NOR2_X4 U12409 ( .A1(n9876), .A2(n10010), .ZN(n13379) );
  NAND2_X1 U12410 ( .A1(n11003), .A2(n10025), .ZN(n9889) );
  OAI211_X1 U12411 ( .C1(n11003), .C2(n10025), .A(n13379), .B(n9889), .ZN(
        n11004) );
  INV_X1 U12412 ( .A(n11004), .ZN(n9877) );
  AOI21_X1 U12413 ( .B1(n14567), .B2(n10026), .A(n9877), .ZN(n9878) );
  OAI211_X1 U12414 ( .C1(n14571), .C2(n11009), .A(n9879), .B(n9878), .ZN(n9922) );
  NAND2_X1 U12415 ( .A1(n10992), .A2(n9922), .ZN(n9880) );
  OAI21_X1 U12416 ( .B1(n10992), .B2(n9881), .A(n9880), .ZN(P2_U3433) );
  INV_X1 U12417 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9884) );
  AOI21_X1 U12418 ( .B1(n13268), .B2(n9868), .A(n10199), .ZN(n9882) );
  AND2_X1 U12419 ( .A1(n8148), .A2(n13037), .ZN(n10217) );
  NOR2_X1 U12420 ( .A1(n9882), .A2(n10217), .ZN(n10194) );
  NAND2_X1 U12421 ( .A1(n10212), .A2(n10023), .ZN(n10214) );
  OAI211_X1 U12422 ( .C1(n10199), .C2(n13341), .A(n10194), .B(n10214), .ZN(
        n9924) );
  NAND2_X1 U12423 ( .A1(n10992), .A2(n9924), .ZN(n9883) );
  OAI21_X1 U12424 ( .B1(n10992), .B2(n9884), .A(n9883), .ZN(P2_U3430) );
  OAI222_X1 U12425 ( .A1(n14012), .A2(n9886), .B1(n14014), .B2(n9885), .C1(
        n10415), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U12426 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9902) );
  INV_X1 U12427 ( .A(n10024), .ZN(n9888) );
  OR2_X1 U12428 ( .A1(n8148), .A2(n10026), .ZN(n9887) );
  XNOR2_X1 U12429 ( .A(n10280), .B(n10278), .ZN(n11002) );
  NAND2_X1 U12430 ( .A1(n9889), .A2(n8145), .ZN(n9890) );
  NAND3_X1 U12431 ( .A1(n10773), .A2(n13379), .A3(n9890), .ZN(n10997) );
  INV_X1 U12432 ( .A(n10997), .ZN(n9899) );
  INV_X1 U12433 ( .A(n10215), .ZN(n9892) );
  NAND2_X1 U12434 ( .A1(n9892), .A2(n9891), .ZN(n9893) );
  NAND2_X1 U12435 ( .A1(n9893), .A2(n7339), .ZN(n9894) );
  NAND2_X1 U12436 ( .A1(n9894), .A2(n10278), .ZN(n10287) );
  OAI21_X1 U12437 ( .B1(n10278), .B2(n9894), .A(n10287), .ZN(n9895) );
  NAND2_X1 U12438 ( .A1(n9895), .A2(n13284), .ZN(n9898) );
  NAND2_X1 U12439 ( .A1(n13037), .A2(n8149), .ZN(n9897) );
  NAND2_X1 U12440 ( .A1(n13038), .A2(n8148), .ZN(n9896) );
  AND2_X1 U12441 ( .A1(n9897), .A2(n9896), .ZN(n11955) );
  NAND2_X1 U12442 ( .A1(n9898), .A2(n11955), .ZN(n11000) );
  AOI211_X1 U12443 ( .C1(n14567), .C2(n8145), .A(n9899), .B(n11000), .ZN(n9900) );
  OAI21_X1 U12444 ( .B1(n14571), .B2(n11002), .A(n9900), .ZN(n13406) );
  NAND2_X1 U12445 ( .A1(n13406), .A2(n10992), .ZN(n9901) );
  OAI21_X1 U12446 ( .B1(n10992), .B2(n9902), .A(n9901), .ZN(P2_U3436) );
  INV_X1 U12447 ( .A(n9903), .ZN(n9906) );
  AND3_X1 U12448 ( .A1(n9906), .A2(n9905), .A3(n9904), .ZN(n9907) );
  AND2_X1 U12449 ( .A1(n9907), .A2(n10034), .ZN(n9917) );
  OR2_X1 U12450 ( .A1(n12380), .A2(n11020), .ZN(n9910) );
  OR2_X1 U12451 ( .A1(n9908), .A2(n10556), .ZN(n9909) );
  AOI21_X1 U12452 ( .B1(n14357), .B2(n14349), .A(n9912), .ZN(n9913) );
  AOI21_X1 U12453 ( .B1(n14292), .B2(n9761), .A(n9913), .ZN(n10102) );
  OAI21_X1 U12454 ( .B1(n8863), .B2(n9914), .A(n10102), .ZN(n9918) );
  NAND2_X1 U12455 ( .A1(n9918), .A2(n14391), .ZN(n9915) );
  OAI21_X1 U12456 ( .B1(n14391), .B2(n9753), .A(n9915), .ZN(P1_U3528) );
  INV_X1 U12457 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n14922) );
  NAND2_X1 U12458 ( .A1(n9918), .A2(n14378), .ZN(n9919) );
  OAI21_X1 U12459 ( .B1(n14378), .B2(n14922), .A(n9919), .ZN(P1_U3459) );
  INV_X1 U12460 ( .A(n10008), .ZN(n9920) );
  NAND2_X1 U12461 ( .A1(n10988), .A2(n9922), .ZN(n9923) );
  OAI21_X1 U12462 ( .B1(n10988), .B2(n9646), .A(n9923), .ZN(P2_U3500) );
  NAND2_X1 U12463 ( .A1(n10988), .A2(n9924), .ZN(n9925) );
  OAI21_X1 U12464 ( .B1(n10988), .B2(n14398), .A(n9925), .ZN(P2_U3499) );
  INV_X1 U12465 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9937) );
  INV_X1 U12466 ( .A(n13540), .ZN(n10111) );
  INV_X1 U12467 ( .A(n9926), .ZN(n10091) );
  NAND2_X1 U12468 ( .A1(n10080), .A2(n14322), .ZN(n9927) );
  XNOR2_X1 U12469 ( .A(n10110), .B(n10109), .ZN(n9933) );
  NAND2_X1 U12470 ( .A1(n9929), .A2(n9928), .ZN(n10104) );
  XNOR2_X1 U12471 ( .A(n10104), .B(n10109), .ZN(n9931) );
  AOI22_X1 U12472 ( .A1(n14292), .A2(n13596), .B1(n14131), .B2(n9761), .ZN(
        n9930) );
  OAI21_X1 U12473 ( .B1(n9931), .B2(n14357), .A(n9930), .ZN(n9932) );
  AOI21_X1 U12474 ( .B1(n14375), .B2(n9933), .A(n9932), .ZN(n10043) );
  NAND2_X1 U12475 ( .A1(n8863), .A2(n14322), .ZN(n10079) );
  INV_X1 U12476 ( .A(n10079), .ZN(n9935) );
  INV_X1 U12477 ( .A(n14312), .ZN(n9934) );
  OAI211_X1 U12478 ( .C1(n10111), .C2(n9935), .A(n9934), .B(n14310), .ZN(
        n10038) );
  OAI211_X1 U12479 ( .C1(n10111), .C2(n14371), .A(n10043), .B(n10038), .ZN(
        n9938) );
  NAND2_X1 U12480 ( .A1(n9938), .A2(n14378), .ZN(n9936) );
  OAI21_X1 U12481 ( .B1(n14378), .B2(n9937), .A(n9936), .ZN(P1_U3465) );
  NAND2_X1 U12482 ( .A1(n9938), .A2(n14391), .ZN(n9939) );
  OAI21_X1 U12483 ( .B1(n14391), .B2(n9940), .A(n9939), .ZN(P1_U3530) );
  INV_X1 U12484 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9942) );
  MUX2_X1 U12485 ( .A(n9942), .B(P2_REG2_REG_7__SCAN_IN), .S(n9951), .Z(n14443) );
  AOI21_X1 U12486 ( .B1(n9951), .B2(P2_REG2_REG_7__SCAN_IN), .A(n14442), .ZN(
        n14459) );
  INV_X1 U12487 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9943) );
  MUX2_X1 U12488 ( .A(n9943), .B(P2_REG2_REG_8__SCAN_IN), .S(n9954), .Z(n14458) );
  NOR2_X1 U12489 ( .A1(n14459), .A2(n14458), .ZN(n14457) );
  AOI21_X1 U12490 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n9954), .A(n14457), .ZN(
        n9946) );
  INV_X1 U12491 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9944) );
  MUX2_X1 U12492 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n9944), .S(n10424), .Z(n9945) );
  NAND2_X1 U12493 ( .A1(n9946), .A2(n9945), .ZN(n10423) );
  OAI21_X1 U12494 ( .B1(n9946), .B2(n9945), .A(n10423), .ZN(n9962) );
  NAND2_X1 U12495 ( .A1(n9947), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U12496 ( .A1(n9949), .A2(n9948), .ZN(n14447) );
  INV_X1 U12497 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9950) );
  MUX2_X1 U12498 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9950), .S(n9951), .Z(n14446) );
  NAND2_X1 U12499 ( .A1(n14447), .A2(n14446), .ZN(n14445) );
  NAND2_X1 U12500 ( .A1(n9951), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U12501 ( .A1(n14445), .A2(n9952), .ZN(n14456) );
  INV_X1 U12502 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9953) );
  MUX2_X1 U12503 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9953), .S(n9954), .Z(n14455) );
  AND2_X1 U12504 ( .A1(n14456), .A2(n14455), .ZN(n14453) );
  AOI21_X1 U12505 ( .B1(n9954), .B2(P2_REG1_REG_8__SCAN_IN), .A(n14453), .ZN(
        n9956) );
  INV_X1 U12506 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10858) );
  MUX2_X1 U12507 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10858), .S(n10424), .Z(
        n9955) );
  NOR2_X1 U12508 ( .A1(n9956), .A2(n9955), .ZN(n9957) );
  AND2_X1 U12509 ( .A1(n9956), .A2(n9955), .ZN(n10432) );
  OAI21_X1 U12510 ( .B1(n9957), .B2(n10432), .A(n14542), .ZN(n9960) );
  AND2_X1 U12511 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n9958) );
  AOI21_X1 U12512 ( .B1(n14540), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n9958), .ZN(
        n9959) );
  OAI211_X1 U12513 ( .C1(n14547), .C2(n10433), .A(n9960), .B(n9959), .ZN(n9961) );
  AOI21_X1 U12514 ( .B1(n9962), .B2(n14526), .A(n9961), .ZN(n9963) );
  INV_X1 U12515 ( .A(n9963), .ZN(P2_U3223) );
  INV_X1 U12516 ( .A(n9992), .ZN(n9966) );
  NAND2_X1 U12517 ( .A1(n10129), .A2(n9964), .ZN(n9965) );
  AOI21_X1 U12518 ( .B1(n9998), .B2(n9966), .A(n9965), .ZN(n9968) );
  NAND2_X1 U12519 ( .A1(n10000), .A2(n9991), .ZN(n9967) );
  NAND2_X1 U12520 ( .A1(n9968), .A2(n9967), .ZN(n9969) );
  NAND2_X1 U12521 ( .A1(n9969), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9973) );
  NOR2_X1 U12522 ( .A1(n12308), .A2(n10133), .ZN(n9971) );
  OR2_X1 U12523 ( .A1(n10305), .A2(P3_U3151), .ZN(n12313) );
  INV_X1 U12524 ( .A(n12313), .ZN(n9970) );
  AOI21_X1 U12525 ( .B1(n9998), .B2(n9971), .A(n9970), .ZN(n9972) );
  NOR2_X1 U12526 ( .A1(n12523), .A2(P3_U3151), .ZN(n10078) );
  INV_X1 U12527 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10208) );
  INV_X1 U12528 ( .A(n12139), .ZN(n9974) );
  NAND2_X1 U12529 ( .A1(n9975), .A2(n9974), .ZN(n9978) );
  NAND2_X1 U12530 ( .A1(n12163), .A2(n12623), .ZN(n9976) );
  NAND2_X1 U12531 ( .A1(n9976), .A2(n10455), .ZN(n9977) );
  NAND2_X1 U12532 ( .A1(n9979), .A2(n6419), .ZN(n9981) );
  NAND3_X1 U12533 ( .A1(n12557), .A2(n6420), .A3(n9982), .ZN(n9983) );
  NAND2_X1 U12534 ( .A1(n10202), .A2(n6420), .ZN(n9984) );
  NAND2_X1 U12535 ( .A1(n9985), .A2(n9984), .ZN(n9986) );
  INV_X1 U12536 ( .A(n12164), .ZN(n9988) );
  NAND3_X1 U12537 ( .A1(n9988), .A2(n9987), .A3(n12444), .ZN(n9989) );
  OAI211_X1 U12538 ( .C1(n9990), .C2(n10202), .A(n10055), .B(n9989), .ZN(n9996) );
  NAND2_X1 U12539 ( .A1(n9991), .A2(n14827), .ZN(n9993) );
  OAI22_X1 U12540 ( .A1(n10000), .A2(n9993), .B1(n9998), .B2(n9992), .ZN(n9995) );
  NAND2_X1 U12541 ( .A1(n9996), .A2(n12509), .ZN(n10003) );
  OR2_X1 U12542 ( .A1(n12308), .A2(n12309), .ZN(n9997) );
  NOR2_X1 U12543 ( .A1(n9998), .A2(n9997), .ZN(n10474) );
  NAND2_X1 U12544 ( .A1(n10474), .A2(n12763), .ZN(n12475) );
  INV_X1 U12545 ( .A(n12475), .ZN(n12522) );
  OR2_X1 U12546 ( .A1(n12308), .A2(n14827), .ZN(n9999) );
  AOI21_X2 U12547 ( .B1(n10000), .B2(n12302), .A(n9999), .ZN(n12528) );
  NAND2_X1 U12548 ( .A1(n10474), .A2(n12765), .ZN(n12526) );
  OAI22_X1 U12549 ( .A1(n10200), .A2(n12518), .B1(n8358), .B2(n12526), .ZN(
        n10001) );
  AOI21_X1 U12550 ( .B1(n12522), .B2(n9718), .A(n10001), .ZN(n10002) );
  OAI211_X1 U12551 ( .C1(n10078), .C2(n10208), .A(n10003), .B(n10002), .ZN(
        P3_U3162) );
  INV_X1 U12552 ( .A(n10004), .ZN(n10052) );
  OAI222_X1 U12553 ( .A1(n13444), .A2(n10052), .B1(n13083), .B2(P2_U3088), 
        .C1(n10005), .C2(n12041), .ZN(P2_U3311) );
  OAI21_X1 U12554 ( .B1(n10191), .B2(n10007), .A(n10011), .ZN(n10009) );
  NAND2_X1 U12555 ( .A1(n10009), .A2(n10008), .ZN(n10260) );
  NOR2_X1 U12556 ( .A1(n10260), .A2(n14553), .ZN(n11954) );
  INV_X1 U12557 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n14393) );
  NAND2_X1 U12558 ( .A1(n10023), .A2(n10010), .ZN(n10573) );
  NOR2_X2 U12559 ( .A1(n10016), .A2(n10013), .ZN(n12999) );
  INV_X1 U12560 ( .A(n10014), .ZN(n10015) );
  AOI22_X1 U12561 ( .A1(n6418), .A2(n10026), .B1(n12999), .B2(n10015), .ZN(
        n10031) );
  INV_X1 U12562 ( .A(n10016), .ZN(n10020) );
  INV_X1 U12563 ( .A(n10017), .ZN(n10018) );
  NAND2_X2 U12564 ( .A1(n13379), .A2(n13093), .ZN(n10256) );
  NAND2_X1 U12565 ( .A1(n10256), .A2(n8148), .ZN(n10237) );
  NAND2_X1 U12566 ( .A1(n10027), .A2(n10028), .ZN(n10240) );
  OAI21_X1 U12567 ( .B1(n10028), .B2(n10027), .A(n10240), .ZN(n10029) );
  NAND2_X1 U12568 ( .A1(n13035), .A2(n10029), .ZN(n10030) );
  OAI211_X1 U12569 ( .C1(n11954), .C2(n14393), .A(n10031), .B(n10030), .ZN(
        P2_U3194) );
  NOR2_X1 U12570 ( .A1(n10033), .A2(n10032), .ZN(n10035) );
  NAND2_X1 U12571 ( .A1(n10035), .A2(n10034), .ZN(n11885) );
  INV_X1 U12572 ( .A(n10036), .ZN(n10037) );
  AOI22_X1 U12573 ( .A1(n14284), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n14285), .ZN(n10040) );
  OR2_X1 U12574 ( .A1(n14160), .A2(n10038), .ZN(n10039) );
  OAI211_X1 U12575 ( .C1(n13883), .C2(n10111), .A(n10040), .B(n10039), .ZN(
        n10041) );
  INV_X1 U12576 ( .A(n10041), .ZN(n10042) );
  OAI21_X1 U12577 ( .B1(n10043), .B2(n14318), .A(n10042), .ZN(P1_U3291) );
  OAI222_X1 U12578 ( .A1(n12880), .A2(n10045), .B1(n12874), .B2(n10044), .C1(
        P3_U3151), .C2(n12105), .ZN(P3_U3276) );
  AND2_X1 U12579 ( .A1(n9718), .A2(n10274), .ZN(n12114) );
  NOR2_X1 U12580 ( .A1(n12164), .A2(n12114), .ZN(n10135) );
  INV_X1 U12581 ( .A(n10078), .ZN(n10046) );
  NAND2_X1 U12582 ( .A1(n10046), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10049) );
  INV_X1 U12583 ( .A(n12526), .ZN(n10047) );
  AOI22_X1 U12584 ( .A1(n12557), .A2(n10047), .B1(n12528), .B2(n12157), .ZN(
        n10048) );
  OAI211_X1 U12585 ( .C1(n10135), .C2(n12531), .A(n10049), .B(n10048), .ZN(
        P3_U3172) );
  INV_X1 U12586 ( .A(n10050), .ZN(n10069) );
  INV_X1 U12587 ( .A(n11731), .ZN(n11742) );
  OAI222_X1 U12588 ( .A1(n13444), .A2(n10069), .B1(n11742), .B2(P2_U3088), 
        .C1(n10051), .C2(n12041), .ZN(P2_U3313) );
  OAI222_X1 U12589 ( .A1(n14012), .A2(n10053), .B1(n14014), .B2(n10052), .C1(
        n11591), .C2(P1_U3086), .ZN(P1_U3339) );
  NAND2_X1 U12590 ( .A1(n10055), .A2(n10054), .ZN(n10071) );
  XNOR2_X1 U12591 ( .A(n10056), .B(n6420), .ZN(n10058) );
  XNOR2_X1 U12592 ( .A(n10058), .B(n8358), .ZN(n10072) );
  NAND2_X1 U12593 ( .A1(n10071), .A2(n10072), .ZN(n10061) );
  XNOR2_X1 U12594 ( .A(n10057), .B(n6419), .ZN(n10394) );
  XNOR2_X1 U12595 ( .A(n10394), .B(n14761), .ZN(n10062) );
  INV_X1 U12596 ( .A(n10058), .ZN(n10059) );
  NAND2_X1 U12597 ( .A1(n10059), .A2(n8358), .ZN(n10063) );
  AND2_X1 U12598 ( .A1(n10062), .A2(n10063), .ZN(n10060) );
  NAND2_X1 U12599 ( .A1(n10396), .A2(n12509), .ZN(n10068) );
  AOI21_X1 U12600 ( .B1(n10061), .B2(n10063), .A(n10062), .ZN(n10067) );
  OAI22_X1 U12601 ( .A1(n12518), .A2(n14782), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n8361), .ZN(n10065) );
  OAI22_X1 U12602 ( .A1(n12180), .A2(n12526), .B1(n8358), .B2(n12475), .ZN(
        n10064) );
  AOI211_X1 U12603 ( .C1(n8361), .C2(n12523), .A(n10065), .B(n10064), .ZN(
        n10066) );
  OAI21_X1 U12604 ( .B1(n10068), .B2(n10067), .A(n10066), .ZN(P3_U3158) );
  INV_X1 U12605 ( .A(n11392), .ZN(n11401) );
  OAI222_X1 U12606 ( .A1(n14012), .A2(n10070), .B1(n14014), .B2(n10069), .C1(
        n11401), .C2(P1_U3086), .ZN(P1_U3341) );
  INV_X1 U12607 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10077) );
  OAI21_X1 U12608 ( .B1(n10072), .B2(n10071), .A(n10061), .ZN(n10073) );
  NAND2_X1 U12609 ( .A1(n10073), .A2(n12509), .ZN(n10076) );
  OAI22_X1 U12610 ( .A1(n12518), .A2(n14754), .B1(n14761), .B2(n12526), .ZN(
        n10074) );
  AOI21_X1 U12611 ( .B1(n12522), .B2(n12557), .A(n10074), .ZN(n10075) );
  OAI211_X1 U12612 ( .C1(n10078), .C2(n10077), .A(n10076), .B(n10075), .ZN(
        P3_U3177) );
  OAI21_X1 U12613 ( .B1(n14322), .B2(n8863), .A(n10079), .ZN(n10087) );
  XNOR2_X1 U12614 ( .A(n10087), .B(n10080), .ZN(n10083) );
  INV_X1 U12615 ( .A(n10092), .ZN(n10081) );
  NOR2_X1 U12616 ( .A1(n10081), .A2(n14131), .ZN(n10082) );
  MUX2_X1 U12617 ( .A(n10083), .B(n10082), .S(n13598), .Z(n10086) );
  AOI21_X1 U12618 ( .B1(n14131), .B2(n13598), .A(n14353), .ZN(n10085) );
  OAI21_X1 U12619 ( .B1(n10086), .B2(n10085), .A(n10084), .ZN(n14323) );
  INV_X1 U12620 ( .A(n14323), .ZN(n10095) );
  INV_X1 U12621 ( .A(n10087), .ZN(n10088) );
  NAND2_X1 U12622 ( .A1(n10088), .A2(n14310), .ZN(n14321) );
  OAI22_X1 U12623 ( .A1(n14160), .A2(n14321), .B1(n13599), .B2(n14302), .ZN(
        n10090) );
  NOR2_X1 U12624 ( .A1(n13883), .A2(n14322), .ZN(n10089) );
  AOI211_X1 U12625 ( .C1(n13880), .C2(P1_REG2_REG_1__SCAN_IN), .A(n10090), .B(
        n10089), .ZN(n10094) );
  XNOR2_X1 U12626 ( .A(n10092), .B(n10091), .ZN(n14325) );
  NAND2_X1 U12627 ( .A1(n14315), .A2(n14325), .ZN(n10093) );
  OAI211_X1 U12628 ( .C1(n14318), .C2(n10095), .A(n10094), .B(n10093), .ZN(
        P1_U3292) );
  INV_X1 U12629 ( .A(n10096), .ZN(n10143) );
  INV_X1 U12630 ( .A(n14520), .ZN(n13085) );
  OAI222_X1 U12631 ( .A1(n13444), .A2(n10143), .B1(n13085), .B2(P2_U3088), 
        .C1(n10097), .C2(n12041), .ZN(P2_U3310) );
  OR2_X1 U12632 ( .A1(n14160), .A2(n14182), .ZN(n13907) );
  INV_X1 U12633 ( .A(n13907), .ZN(n10099) );
  OAI21_X1 U12634 ( .B1(n14306), .B2(n10099), .A(n10098), .ZN(n10101) );
  AOI22_X1 U12635 ( .A1(n14284), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n14285), .ZN(n10100) );
  OAI211_X1 U12636 ( .C1(n14318), .C2(n10102), .A(n10101), .B(n10100), .ZN(
        P1_U3293) );
  INV_X1 U12637 ( .A(n10148), .ZN(n10159) );
  NAND2_X1 U12638 ( .A1(n10104), .A2(n10103), .ZN(n10106) );
  NAND2_X1 U12639 ( .A1(n6611), .A2(n13540), .ZN(n10105) );
  NAND2_X1 U12640 ( .A1(n10106), .A2(n10105), .ZN(n14297) );
  NAND2_X1 U12641 ( .A1(n14297), .A2(n14298), .ZN(n10108) );
  XNOR2_X1 U12642 ( .A(n10159), .B(n10160), .ZN(n14341) );
  INV_X1 U12643 ( .A(n14341), .ZN(n10125) );
  INV_X1 U12644 ( .A(n13885), .ZN(n13868) );
  NAND2_X1 U12645 ( .A1(n6611), .A2(n10111), .ZN(n10112) );
  NAND2_X1 U12646 ( .A1(n10113), .A2(n10112), .ZN(n14307) );
  NAND2_X1 U12647 ( .A1(n10175), .A2(n14328), .ZN(n10114) );
  XNOR2_X1 U12648 ( .A(n10149), .B(n10148), .ZN(n14334) );
  INV_X1 U12649 ( .A(n14335), .ZN(n10121) );
  OAI211_X1 U12650 ( .C1(n14309), .C2(n10121), .A(n14310), .B(n10228), .ZN(
        n14337) );
  NOR2_X1 U12651 ( .A1(n14337), .A2(n14160), .ZN(n10123) );
  NAND2_X1 U12652 ( .A1(n14292), .A2(n13594), .ZN(n10117) );
  NAND2_X1 U12653 ( .A1(n14131), .A2(n13596), .ZN(n10116) );
  AND2_X1 U12654 ( .A1(n10117), .A2(n10116), .ZN(n14338) );
  MUX2_X1 U12655 ( .A(n14338), .B(n10118), .S(n14318), .Z(n10120) );
  NAND2_X1 U12656 ( .A1(n14285), .A2(n10462), .ZN(n10119) );
  OAI211_X1 U12657 ( .C1(n10121), .C2(n13883), .A(n10120), .B(n10119), .ZN(
        n10122) );
  AOI211_X1 U12658 ( .C1(n14334), .C2(n14315), .A(n10123), .B(n10122), .ZN(
        n10124) );
  OAI21_X1 U12659 ( .B1(n10125), .B2(n13868), .A(n10124), .ZN(P1_U3289) );
  XNOR2_X1 U12660 ( .A(n10127), .B(n10126), .ZN(n10128) );
  NAND3_X1 U12661 ( .A1(n10130), .A2(n10129), .A3(n10128), .ZN(n10136) );
  OR2_X1 U12662 ( .A1(n14756), .A2(n14827), .ZN(n10131) );
  OR2_X1 U12663 ( .A1(n12302), .A2(n14827), .ZN(n10132) );
  NAND2_X1 U12664 ( .A1(n10133), .A2(n14827), .ZN(n10134) );
  INV_X1 U12665 ( .A(n12557), .ZN(n14763) );
  OAI22_X1 U12666 ( .A1(n10135), .A2(n10134), .B1(n14763), .B2(n14760), .ZN(
        n10276) );
  AOI21_X1 U12667 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n12755), .A(n10276), .ZN(
        n10137) );
  MUX2_X1 U12668 ( .A(n14605), .B(n10137), .S(n14770), .Z(n10138) );
  OAI21_X1 U12669 ( .B1(n10274), .B2(n12757), .A(n10138), .ZN(P3_U3233) );
  INV_X1 U12670 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10140) );
  INV_X1 U12671 ( .A(n10139), .ZN(n10141) );
  INV_X1 U12672 ( .A(n11402), .ZN(n14273) );
  OAI222_X1 U12673 ( .A1(n14012), .A2(n10140), .B1(n14014), .B2(n10141), .C1(
        P1_U3086), .C2(n14273), .ZN(P1_U3340) );
  INV_X1 U12674 ( .A(n14511), .ZN(n11744) );
  OAI222_X1 U12675 ( .A1(n12041), .A2(n10142), .B1(n13444), .B2(n10141), .C1(
        P2_U3088), .C2(n11744), .ZN(P2_U3312) );
  OAI222_X1 U12676 ( .A1(n14012), .A2(n10144), .B1(n14014), .B2(n10143), .C1(
        n13702), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U12677 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10145) );
  OAI22_X1 U12678 ( .A1(n12865), .A2(n10274), .B1(n14833), .B2(n10145), .ZN(
        n10146) );
  AOI21_X1 U12679 ( .B1(n10276), .B2(n14833), .A(n10146), .ZN(n10147) );
  INV_X1 U12680 ( .A(n10147), .ZN(P3_U3390) );
  OR2_X1 U12681 ( .A1(n13595), .A2(n14335), .ZN(n10150) );
  OR2_X1 U12682 ( .A1(n10552), .A2(n13594), .ZN(n10151) );
  XNOR2_X1 U12683 ( .A(n10355), .B(n10353), .ZN(n14350) );
  OAI211_X1 U12684 ( .C1(n10229), .C2(n10887), .A(n10358), .B(n14310), .ZN(
        n14347) );
  INV_X1 U12685 ( .A(n14347), .ZN(n10158) );
  NAND2_X1 U12686 ( .A1(n14292), .A2(n13592), .ZN(n10153) );
  NAND2_X1 U12687 ( .A1(n14131), .A2(n13594), .ZN(n10152) );
  AND2_X1 U12688 ( .A1(n10153), .A2(n10152), .ZN(n14343) );
  MUX2_X1 U12689 ( .A(n14343), .B(n10154), .S(n14318), .Z(n10156) );
  NAND2_X1 U12690 ( .A1(n14285), .A2(n10884), .ZN(n10155) );
  OAI211_X1 U12691 ( .C1(n10887), .C2(n13883), .A(n10156), .B(n10155), .ZN(
        n10157) );
  AOI21_X1 U12692 ( .B1(n14314), .B2(n10158), .A(n10157), .ZN(n10168) );
  NAND2_X1 U12693 ( .A1(n14335), .A2(n10161), .ZN(n10162) );
  INV_X1 U12694 ( .A(n10223), .ZN(n10163) );
  NAND2_X1 U12695 ( .A1(n10552), .A2(n10164), .ZN(n10165) );
  XNOR2_X1 U12696 ( .A(n10352), .B(n10353), .ZN(n14352) );
  NAND2_X1 U12697 ( .A1(n14352), .A2(n13885), .ZN(n10167) );
  OAI211_X1 U12698 ( .C1(n14350), .C2(n13887), .A(n10168), .B(n10167), .ZN(
        P1_U3287) );
  NAND2_X1 U12699 ( .A1(n14292), .A2(n13595), .ZN(n10170) );
  NAND2_X1 U12700 ( .A1(n14131), .A2(n13597), .ZN(n10169) );
  AND2_X1 U12701 ( .A1(n10170), .A2(n10169), .ZN(n14299) );
  NAND2_X1 U12702 ( .A1(n13576), .A2(n8870), .ZN(n10173) );
  OAI211_X1 U12703 ( .C1(n14299), .C2(n13513), .A(n10173), .B(n10172), .ZN(
        n10188) );
  OAI22_X1 U12704 ( .A1(n10175), .A2(n11941), .B1(n14328), .B2(n11942), .ZN(
        n10174) );
  XNOR2_X1 U12705 ( .A(n10174), .B(n9834), .ZN(n10459) );
  OAI22_X1 U12706 ( .A1(n11940), .A2(n10175), .B1(n14328), .B2(n11941), .ZN(
        n10458) );
  XNOR2_X1 U12707 ( .A(n10459), .B(n10458), .ZN(n10186) );
  INV_X1 U12708 ( .A(n10176), .ZN(n10177) );
  AOI22_X1 U12709 ( .A1(n10179), .A2(n13597), .B1(n12363), .B2(n13540), .ZN(
        n10181) );
  XNOR2_X1 U12710 ( .A(n10181), .B(n9834), .ZN(n10183) );
  AOI211_X1 U12711 ( .C1(n10186), .C2(n10185), .A(n13564), .B(n7026), .ZN(
        n10187) );
  AOI211_X1 U12712 ( .C1(n14305), .C2(n14142), .A(n10188), .B(n10187), .ZN(
        n10189) );
  INV_X1 U12713 ( .A(n10189), .ZN(P1_U3218) );
  OR2_X1 U12714 ( .A1(n10191), .A2(n10190), .ZN(n10192) );
  NAND2_X1 U12715 ( .A1(n10195), .A2(n11143), .ZN(n10560) );
  INV_X1 U12716 ( .A(n10560), .ZN(n10193) );
  NAND2_X1 U12717 ( .A1(n13257), .A2(n10193), .ZN(n13185) );
  OAI21_X1 U12718 ( .B1(n10195), .B2(n10214), .A(n10194), .ZN(n10196) );
  INV_X1 U12719 ( .A(n13245), .ZN(n13291) );
  AOI22_X1 U12720 ( .A1(n13257), .A2(n10196), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n13291), .ZN(n10198) );
  NAND2_X1 U12721 ( .A1(n13304), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10197) );
  OAI211_X1 U12722 ( .C1(n13185), .C2(n10199), .A(n10198), .B(n10197), .ZN(
        P2_U3265) );
  NOR2_X1 U12723 ( .A1(n10200), .A2(n14827), .ZN(n14774) );
  XNOR2_X1 U12724 ( .A(n9987), .B(n12164), .ZN(n10206) );
  AOI22_X1 U12725 ( .A1(n10201), .A2(n12765), .B1(n12763), .B2(n9718), .ZN(
        n10205) );
  XNOR2_X1 U12726 ( .A(n9987), .B(n10202), .ZN(n10203) );
  NAND2_X1 U12727 ( .A1(n10203), .A2(n12768), .ZN(n10204) );
  OAI211_X1 U12728 ( .C1(n10206), .C2(n14808), .A(n10205), .B(n10204), .ZN(
        n14773) );
  AOI21_X1 U12729 ( .B1(n14774), .B2(n12302), .A(n14773), .ZN(n10211) );
  INV_X1 U12730 ( .A(n10206), .ZN(n14775) );
  NAND2_X1 U12731 ( .A1(n10207), .A2(n14756), .ZN(n10712) );
  INV_X1 U12732 ( .A(n10712), .ZN(n14769) );
  NAND2_X1 U12733 ( .A1(n14770), .A2(n14769), .ZN(n11124) );
  INV_X1 U12734 ( .A(n11124), .ZN(n12678) );
  OAI22_X1 U12735 ( .A1(n14770), .A2(n8329), .B1(n10208), .B2(n14755), .ZN(
        n10209) );
  AOI21_X1 U12736 ( .B1(n14775), .B2(n12678), .A(n10209), .ZN(n10210) );
  OAI21_X1 U12737 ( .B1(n10211), .B2(n14772), .A(n10210), .ZN(P3_U3232) );
  INV_X1 U12738 ( .A(n10256), .ZN(n11970) );
  OR2_X1 U12739 ( .A1(n13023), .A2(n11970), .ZN(n11989) );
  NAND2_X1 U12740 ( .A1(n13013), .A2(n9869), .ZN(n10213) );
  INV_X1 U12741 ( .A(n6418), .ZN(n13045) );
  MUX2_X1 U12742 ( .A(n10213), .B(n13045), .S(n10212), .Z(n10219) );
  AOI21_X1 U12743 ( .B1(n10215), .B2(n10214), .A(n13023), .ZN(n10216) );
  AOI21_X1 U12744 ( .B1(n10217), .B2(n12999), .A(n10216), .ZN(n10218) );
  OAI211_X1 U12745 ( .C1(n11954), .C2(n10220), .A(n10219), .B(n10218), .ZN(
        P2_U3204) );
  XNOR2_X1 U12746 ( .A(n10221), .B(n10223), .ZN(n10227) );
  XNOR2_X1 U12747 ( .A(n10222), .B(n10223), .ZN(n10225) );
  AOI22_X1 U12748 ( .A1(n14292), .A2(n13593), .B1(n14131), .B2(n13595), .ZN(
        n10224) );
  OAI21_X1 U12749 ( .B1(n10225), .B2(n14357), .A(n10224), .ZN(n10226) );
  AOI21_X1 U12750 ( .B1(n14375), .B2(n10227), .A(n10226), .ZN(n10300) );
  INV_X1 U12751 ( .A(n10228), .ZN(n10231) );
  INV_X1 U12752 ( .A(n10229), .ZN(n10230) );
  OAI211_X1 U12753 ( .C1(n6883), .C2(n10231), .A(n10230), .B(n14310), .ZN(
        n10304) );
  OAI211_X1 U12754 ( .C1(n6883), .C2(n14371), .A(n10300), .B(n10304), .ZN(
        n10234) );
  NAND2_X1 U12755 ( .A1(n10234), .A2(n14391), .ZN(n10232) );
  OAI21_X1 U12756 ( .B1(n14391), .B2(n10233), .A(n10232), .ZN(P1_U3533) );
  INV_X1 U12757 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10236) );
  NAND2_X1 U12758 ( .A1(n10234), .A2(n14378), .ZN(n10235) );
  OAI21_X1 U12759 ( .B1(n14378), .B2(n10236), .A(n10235), .ZN(P1_U3474) );
  INV_X1 U12760 ( .A(n11956), .ZN(n10238) );
  NAND2_X1 U12761 ( .A1(n10238), .A2(n10237), .ZN(n10239) );
  NAND2_X1 U12762 ( .A1(n10240), .A2(n10239), .ZN(n10241) );
  XNOR2_X1 U12763 ( .A(n12921), .B(n8145), .ZN(n10242) );
  NAND2_X1 U12764 ( .A1(n6458), .A2(n8146), .ZN(n10243) );
  XNOR2_X1 U12765 ( .A(n10242), .B(n10243), .ZN(n11957) );
  INV_X1 U12766 ( .A(n10242), .ZN(n10244) );
  NAND2_X1 U12767 ( .A1(n10244), .A2(n10243), .ZN(n10245) );
  XNOR2_X1 U12768 ( .A(n12921), .B(n10772), .ZN(n10246) );
  AND2_X1 U12769 ( .A1(n10256), .A2(n8149), .ZN(n10247) );
  NAND2_X1 U12770 ( .A1(n10246), .A2(n10247), .ZN(n10251) );
  INV_X1 U12771 ( .A(n10246), .ZN(n10499) );
  INV_X1 U12772 ( .A(n10247), .ZN(n10248) );
  NAND2_X1 U12773 ( .A1(n10499), .A2(n10248), .ZN(n10249) );
  NAND2_X1 U12774 ( .A1(n10251), .A2(n10249), .ZN(n10345) );
  XNOR2_X1 U12775 ( .A(n14566), .B(n12921), .ZN(n10265) );
  BUF_X1 U12776 ( .A(n10256), .Z(n12916) );
  XNOR2_X1 U12777 ( .A(n10265), .B(n10253), .ZN(n10498) );
  AND2_X1 U12778 ( .A1(n10498), .A2(n10251), .ZN(n10252) );
  INV_X1 U12779 ( .A(n10265), .ZN(n10254) );
  NAND2_X1 U12780 ( .A1(n10254), .A2(n10253), .ZN(n10255) );
  NAND2_X1 U12781 ( .A1(n10266), .A2(n10255), .ZN(n10257) );
  XNOR2_X1 U12782 ( .A(n10507), .B(n12948), .ZN(n10699) );
  NAND2_X1 U12783 ( .A1(n12916), .A2(n13070), .ZN(n10700) );
  XNOR2_X1 U12784 ( .A(n10699), .B(n10700), .ZN(n10267) );
  NAND2_X1 U12785 ( .A1(n10257), .A2(n10267), .ZN(n10703) );
  INV_X1 U12786 ( .A(n10258), .ZN(n10259) );
  OR2_X1 U12787 ( .A1(n10260), .A2(n10259), .ZN(n10261) );
  INV_X1 U12788 ( .A(n13015), .ZN(n13042) );
  INV_X1 U12789 ( .A(n10684), .ZN(n10272) );
  INV_X1 U12790 ( .A(n13069), .ZN(n10517) );
  OAI22_X1 U12791 ( .A1(n10262), .A2(n12995), .B1(n10517), .B2(n12997), .ZN(
        n10293) );
  NAND2_X1 U12792 ( .A1(n12999), .A2(n10293), .ZN(n10263) );
  OAI211_X1 U12793 ( .C1(n13045), .C2(n6923), .A(n10264), .B(n10263), .ZN(
        n10271) );
  AOI22_X1 U12794 ( .A1(n13013), .A2(n13071), .B1(n13035), .B2(n10265), .ZN(
        n10269) );
  INV_X1 U12795 ( .A(n10266), .ZN(n10268) );
  NOR3_X1 U12796 ( .A1(n10269), .A2(n10268), .A3(n10267), .ZN(n10270) );
  AOI211_X1 U12797 ( .C1(n13042), .C2(n10272), .A(n10271), .B(n10270), .ZN(
        n10273) );
  OAI21_X1 U12798 ( .B1(n10703), .B2(n13023), .A(n10273), .ZN(P2_U3199) );
  INV_X1 U12799 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10309) );
  OAI22_X1 U12800 ( .A1(n12826), .A2(n10274), .B1(n14846), .B2(n10309), .ZN(
        n10275) );
  AOI21_X1 U12801 ( .B1(n10276), .B2(n14846), .A(n10275), .ZN(n10277) );
  INV_X1 U12802 ( .A(n10277), .ZN(P3_U3459) );
  INV_X1 U12803 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10297) );
  INV_X1 U12804 ( .A(n10278), .ZN(n10279) );
  OR2_X1 U12805 ( .A1(n8146), .A2(n8145), .ZN(n10281) );
  NAND2_X1 U12806 ( .A1(n10282), .A2(n14561), .ZN(n10283) );
  NAND2_X1 U12807 ( .A1(n10284), .A2(n10283), .ZN(n10563) );
  INV_X1 U12808 ( .A(n10562), .ZN(n10566) );
  OR2_X1 U12809 ( .A1(n13071), .A2(n14566), .ZN(n10285) );
  XNOR2_X1 U12810 ( .A(n10506), .B(n10504), .ZN(n10689) );
  INV_X1 U12811 ( .A(n10288), .ZN(n10779) );
  NAND2_X1 U12812 ( .A1(n10778), .A2(n10779), .ZN(n10564) );
  NAND2_X1 U12813 ( .A1(n10564), .A2(n10565), .ZN(n10289) );
  NAND2_X1 U12814 ( .A1(n10289), .A2(n10562), .ZN(n10568) );
  NAND2_X1 U12815 ( .A1(n10568), .A2(n10290), .ZN(n10291) );
  NAND2_X1 U12816 ( .A1(n10291), .A2(n10504), .ZN(n10516) );
  OAI21_X1 U12817 ( .B1(n10504), .B2(n10291), .A(n10516), .ZN(n10294) );
  NOR2_X1 U12818 ( .A1(n10689), .A2(n9868), .ZN(n10292) );
  AOI211_X1 U12819 ( .C1(n13284), .C2(n10294), .A(n10293), .B(n10292), .ZN(
        n10683) );
  INV_X1 U12820 ( .A(n10525), .ZN(n10678) );
  AOI211_X1 U12821 ( .C1(n10507), .C2(n10571), .A(n13289), .B(n10678), .ZN(
        n10686) );
  AOI21_X1 U12822 ( .B1(n14567), .B2(n10507), .A(n10686), .ZN(n10295) );
  OAI211_X1 U12823 ( .C1(n10689), .C2(n13341), .A(n10683), .B(n10295), .ZN(
        n10298) );
  NAND2_X1 U12824 ( .A1(n10298), .A2(n10992), .ZN(n10296) );
  OAI21_X1 U12825 ( .B1(n10992), .B2(n10297), .A(n10296), .ZN(P2_U3445) );
  NAND2_X1 U12826 ( .A1(n10298), .A2(n10988), .ZN(n10299) );
  OAI21_X1 U12827 ( .B1(n10988), .B2(n9661), .A(n10299), .ZN(P2_U3504) );
  MUX2_X1 U12828 ( .A(n9608), .B(n10300), .S(n14303), .Z(n10303) );
  AOI22_X1 U12829 ( .A1(n14306), .A2(n10552), .B1(n10301), .B2(n14285), .ZN(
        n10302) );
  OAI211_X1 U12830 ( .C1(n14160), .C2(n10304), .A(n10303), .B(n10302), .ZN(
        P1_U3288) );
  NAND2_X1 U12831 ( .A1(n12308), .A2(n12313), .ZN(n10315) );
  NAND2_X1 U12832 ( .A1(n12288), .A2(n10305), .ZN(n10306) );
  AND2_X1 U12833 ( .A1(n10307), .A2(n10306), .ZN(n10314) );
  AND2_X1 U12834 ( .A1(n10315), .A2(n10314), .ZN(n10319) );
  MUX2_X1 U12835 ( .A(n12552), .B(n10308), .S(n6630), .Z(n14740) );
  INV_X1 U12836 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n14835) );
  AND2_X1 U12837 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10321), .ZN(n10310) );
  OR2_X1 U12838 ( .A1(n10491), .A2(n10310), .ZN(n10311) );
  AND2_X1 U12839 ( .A1(n10311), .A2(n7342), .ZN(n10483) );
  NAND2_X1 U12840 ( .A1(P3_REG1_REG_1__SCAN_IN), .A2(n10483), .ZN(n10482) );
  NAND2_X1 U12841 ( .A1(n7342), .A2(n10482), .ZN(n10312) );
  OAI21_X1 U12842 ( .B1(n10313), .B2(n10312), .A(n10642), .ZN(n10329) );
  INV_X1 U12843 ( .A(n10314), .ZN(n10316) );
  OAI22_X1 U12844 ( .A1(n14727), .A2(n14923), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10077), .ZN(n10328) );
  INV_X1 U12845 ( .A(n10317), .ZN(n10318) );
  NAND2_X1 U12846 ( .A1(n10322), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10320) );
  OAI221_X1 U12847 ( .B1(n10491), .B2(P3_REG2_REG_0__SCAN_IN), .C1(n10491), 
        .C2(n10321), .A(n10320), .ZN(n10481) );
  NAND2_X1 U12848 ( .A1(P3_REG2_REG_2__SCAN_IN), .A2(n10641), .ZN(n10323) );
  OAI21_X1 U12849 ( .B1(P3_REG2_REG_2__SCAN_IN), .B2(n10641), .A(n10323), .ZN(
        n10324) );
  AOI21_X1 U12850 ( .B1(n10325), .B2(n10324), .A(n10579), .ZN(n10326) );
  NOR2_X1 U12851 ( .A1(n14750), .A2(n10326), .ZN(n10327) );
  AOI211_X1 U12852 ( .C1(n14746), .C2(n10329), .A(n10328), .B(n10327), .ZN(
        n10342) );
  MUX2_X1 U12853 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n8681), .Z(n10330) );
  NOR2_X1 U12854 ( .A1(n10330), .A2(n10491), .ZN(n10332) );
  AOI21_X1 U12855 ( .B1(n10330), .B2(n10491), .A(n10332), .ZN(n10479) );
  MUX2_X1 U12856 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n8681), .Z(n10331) );
  NOR2_X1 U12857 ( .A1(n10331), .A2(n10321), .ZN(n14610) );
  NAND2_X1 U12858 ( .A1(n10479), .A2(n14610), .ZN(n10478) );
  INV_X1 U12859 ( .A(n10332), .ZN(n10339) );
  MUX2_X1 U12860 ( .A(n10333), .B(n14835), .S(n8681), .Z(n10335) );
  NAND2_X1 U12861 ( .A1(n10335), .A2(n10334), .ZN(n10593) );
  INV_X1 U12862 ( .A(n10335), .ZN(n10336) );
  NAND2_X1 U12863 ( .A1(n10336), .A2(n10641), .ZN(n10337) );
  NAND2_X1 U12864 ( .A1(n10593), .A2(n10337), .ZN(n10338) );
  AOI21_X1 U12865 ( .B1(n10478), .B2(n10339), .A(n10338), .ZN(n14623) );
  AND3_X1 U12866 ( .A1(n10478), .A2(n10339), .A3(n10338), .ZN(n10340) );
  NAND2_X1 U12867 ( .A1(P3_U3897), .A2(n6630), .ZN(n14709) );
  OAI21_X1 U12868 ( .B1(n14623), .B2(n10340), .A(n14735), .ZN(n10341) );
  OAI211_X1 U12869 ( .C1(n14740), .C2(n10641), .A(n10342), .B(n10341), .ZN(
        P3_U3184) );
  INV_X1 U12870 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10343) );
  NOR2_X1 U12871 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10343), .ZN(n14423) );
  AOI22_X1 U12872 ( .A1(n13038), .A2(n8146), .B1(n13037), .B2(n13071), .ZN(
        n10780) );
  NOR2_X1 U12873 ( .A1(n13040), .A2(n10780), .ZN(n10344) );
  AOI211_X1 U12874 ( .C1(n10772), .C2(n6418), .A(n14423), .B(n10344), .ZN(
        n10349) );
  AOI21_X1 U12875 ( .B1(n10346), .B2(n10345), .A(n13023), .ZN(n10347) );
  NAND2_X1 U12876 ( .A1(n10347), .A2(n10492), .ZN(n10348) );
  OAI211_X1 U12877 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n13015), .A(n10349), .B(
        n10348), .ZN(P2_U3190) );
  NAND2_X1 U12878 ( .A1(n12552), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n10350) );
  OAI21_X1 U12879 ( .B1(n12451), .B2(n12552), .A(n10350), .ZN(P3_U3520) );
  INV_X1 U12880 ( .A(n13593), .ZN(n10549) );
  AND2_X1 U12881 ( .A1(n14346), .A2(n10549), .ZN(n10351) );
  XOR2_X1 U12882 ( .A(n10754), .B(n10766), .Z(n14358) );
  INV_X1 U12883 ( .A(n10353), .ZN(n10354) );
  NAND2_X1 U12884 ( .A1(n10355), .A2(n10354), .ZN(n10357) );
  OR2_X1 U12885 ( .A1(n14346), .A2(n13593), .ZN(n10356) );
  XNOR2_X1 U12886 ( .A(n10755), .B(n10754), .ZN(n14361) );
  AOI21_X1 U12887 ( .B1(n10358), .B2(n11045), .A(n14182), .ZN(n10359) );
  NAND2_X1 U12888 ( .A1(n10359), .A2(n10759), .ZN(n14356) );
  NAND2_X1 U12889 ( .A1(n14292), .A2(n13591), .ZN(n10361) );
  NAND2_X1 U12890 ( .A1(n14131), .A2(n13593), .ZN(n10360) );
  AND2_X1 U12891 ( .A1(n10361), .A2(n10360), .ZN(n14355) );
  INV_X1 U12892 ( .A(n11050), .ZN(n10362) );
  OAI22_X1 U12893 ( .A1(n13880), .A2(n14355), .B1(n10362), .B2(n14302), .ZN(
        n10365) );
  NOR2_X1 U12894 ( .A1(n14303), .A2(n10363), .ZN(n10364) );
  AOI211_X1 U12895 ( .C1(n14306), .C2(n11045), .A(n10365), .B(n10364), .ZN(
        n10366) );
  OAI21_X1 U12896 ( .B1(n14160), .B2(n14356), .A(n10366), .ZN(n10367) );
  AOI21_X1 U12897 ( .B1(n14361), .B2(n14315), .A(n10367), .ZN(n10368) );
  OAI21_X1 U12898 ( .B1(n14358), .B2(n13868), .A(n10368), .ZN(P1_U3286) );
  INV_X1 U12899 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10369) );
  MUX2_X1 U12900 ( .A(n10369), .B(P1_REG2_REG_13__SCAN_IN), .S(n10415), .Z(
        n10377) );
  OR2_X1 U12901 ( .A1(n13694), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10375) );
  INV_X1 U12902 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10370) );
  AOI22_X1 U12903 ( .A1(n13694), .A2(n10370), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n10381), .ZN(n13691) );
  INV_X1 U12904 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10373) );
  NOR2_X1 U12905 ( .A1(n10372), .A2(n10371), .ZN(n13676) );
  MUX2_X1 U12906 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10373), .S(n13674), .Z(
        n13675) );
  OAI21_X1 U12907 ( .B1(n13677), .B2(n13676), .A(n13675), .ZN(n13679) );
  OAI21_X1 U12908 ( .B1(n10373), .B2(n10380), .A(n13679), .ZN(n13692) );
  NOR2_X1 U12909 ( .A1(n13691), .A2(n13692), .ZN(n13690) );
  INV_X1 U12910 ( .A(n13690), .ZN(n10374) );
  AND2_X1 U12911 ( .A1(n10375), .A2(n10374), .ZN(n10376) );
  NAND2_X1 U12912 ( .A1(n10377), .A2(n10376), .ZN(n10414) );
  OAI211_X1 U12913 ( .C1(n10377), .C2(n10376), .A(n10414), .B(n13725), .ZN(
        n10388) );
  NAND2_X1 U12914 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n11835)
         );
  INV_X1 U12915 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11372) );
  AOI21_X1 U12916 ( .B1(n10379), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10378), 
        .ZN(n13669) );
  INV_X1 U12917 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n14228) );
  MUX2_X1 U12918 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n14228), .S(n13674), .Z(
        n13670) );
  NAND2_X1 U12919 ( .A1(n13669), .A2(n13670), .ZN(n13685) );
  NAND2_X1 U12920 ( .A1(n10380), .A2(n14228), .ZN(n13683) );
  MUX2_X1 U12921 ( .A(n11372), .B(P1_REG1_REG_12__SCAN_IN), .S(n13694), .Z(
        n13684) );
  AOI21_X1 U12922 ( .B1(n13685), .B2(n13683), .A(n13684), .ZN(n13687) );
  INV_X1 U12923 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10382) );
  MUX2_X1 U12924 ( .A(n10382), .B(P1_REG1_REG_13__SCAN_IN), .S(n10415), .Z(
        n10383) );
  NAND2_X1 U12925 ( .A1(n10384), .A2(n10383), .ZN(n10407) );
  OAI211_X1 U12926 ( .C1(n10384), .C2(n10383), .A(n13726), .B(n10407), .ZN(
        n10385) );
  NAND2_X1 U12927 ( .A1(n11835), .A2(n10385), .ZN(n10386) );
  AOI21_X1 U12928 ( .B1(n13708), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10386), 
        .ZN(n10387) );
  OAI211_X1 U12929 ( .C1(n14274), .C2(n10415), .A(n10388), .B(n10387), .ZN(
        P1_U3256) );
  INV_X1 U12930 ( .A(n10389), .ZN(n10456) );
  INV_X1 U12931 ( .A(n13087), .ZN(n14546) );
  OAI222_X1 U12932 ( .A1(n13444), .A2(n10456), .B1(n14546), .B2(P2_U3088), 
        .C1(n10390), .C2(n12041), .ZN(P2_U3309) );
  NAND2_X1 U12933 ( .A1(n12556), .A2(n12763), .ZN(n10392) );
  NAND2_X1 U12934 ( .A1(n12555), .A2(n12765), .ZN(n10391) );
  AND2_X1 U12935 ( .A1(n10392), .A2(n10391), .ZN(n10728) );
  AOI22_X1 U12936 ( .A1(n12528), .A2(n14791), .B1(P3_REG3_REG_4__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10393) );
  OAI21_X1 U12937 ( .B1(n10728), .B2(n12503), .A(n10393), .ZN(n10405) );
  NAND2_X1 U12938 ( .A1(n12556), .A2(n10394), .ZN(n10395) );
  XNOR2_X1 U12939 ( .A(n12182), .B(n6420), .ZN(n10397) );
  NAND2_X1 U12940 ( .A1(n12180), .A2(n10397), .ZN(n10467) );
  INV_X1 U12941 ( .A(n10397), .ZN(n10398) );
  NAND2_X1 U12942 ( .A1(n10398), .A2(n12181), .ZN(n10399) );
  NAND2_X1 U12943 ( .A1(n10467), .A2(n10399), .ZN(n10401) );
  NAND2_X1 U12944 ( .A1(n10402), .A2(n10401), .ZN(n10403) );
  AOI21_X1 U12945 ( .B1(n10468), .B2(n10403), .A(n12531), .ZN(n10404) );
  AOI211_X1 U12946 ( .C1(n10731), .C2(n12523), .A(n10405), .B(n10404), .ZN(
        n10406) );
  INV_X1 U12947 ( .A(n10406), .ZN(P3_U3170) );
  INV_X1 U12948 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14216) );
  AOI22_X1 U12949 ( .A1(n11392), .A2(n14216), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n11401), .ZN(n10409) );
  OAI21_X1 U12950 ( .B1(n10415), .B2(n10382), .A(n10407), .ZN(n10408) );
  NOR2_X1 U12951 ( .A1(n10409), .A2(n10408), .ZN(n11400) );
  AOI21_X1 U12952 ( .B1(n10409), .B2(n10408), .A(n11400), .ZN(n10420) );
  NAND2_X1 U12953 ( .A1(n13708), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n10410) );
  NAND2_X1 U12954 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14126)
         );
  NAND2_X1 U12955 ( .A1(n10410), .A2(n14126), .ZN(n10411) );
  AOI21_X1 U12956 ( .B1(n11392), .B2(n13723), .A(n10411), .ZN(n10419) );
  INV_X1 U12957 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10412) );
  MUX2_X1 U12958 ( .A(n10412), .B(P1_REG2_REG_14__SCAN_IN), .S(n11392), .Z(
        n10413) );
  INV_X1 U12959 ( .A(n10413), .ZN(n10417) );
  OAI21_X1 U12960 ( .B1(n10415), .B2(n10369), .A(n10414), .ZN(n10416) );
  NAND2_X1 U12961 ( .A1(n10417), .A2(n10416), .ZN(n11393) );
  OAI211_X1 U12962 ( .C1(n10417), .C2(n10416), .A(n13725), .B(n11393), .ZN(
        n10418) );
  OAI211_X1 U12963 ( .C1(n10420), .C2(n14272), .A(n10419), .B(n10418), .ZN(
        P1_U3257) );
  INV_X1 U12964 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10421) );
  OR2_X1 U12965 ( .A1(n10422), .A2(n10421), .ZN(n10426) );
  NAND2_X1 U12966 ( .A1(n10422), .A2(n10421), .ZN(n14487) );
  OAI21_X1 U12967 ( .B1(n10424), .B2(P2_REG2_REG_9__SCAN_IN), .A(n10423), .ZN(
        n14472) );
  INV_X1 U12968 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10425) );
  MUX2_X1 U12969 ( .A(n10425), .B(P2_REG2_REG_10__SCAN_IN), .S(n10434), .Z(
        n14473) );
  AOI21_X1 U12970 ( .B1(n10426), .B2(n14487), .A(n10427), .ZN(n10429) );
  INV_X1 U12971 ( .A(n14489), .ZN(n10428) );
  OAI21_X1 U12972 ( .B1(n10429), .B2(n10428), .A(n14526), .ZN(n10443) );
  INV_X1 U12973 ( .A(n14547), .ZN(n14521) );
  OAI22_X1 U12974 ( .A1(n14497), .A2(n9457), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7649), .ZN(n10440) );
  INV_X1 U12975 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10431) );
  NAND2_X1 U12976 ( .A1(n10434), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10437) );
  OAI21_X1 U12977 ( .B1(n10441), .B2(n10431), .A(n10437), .ZN(n10430) );
  AOI21_X1 U12978 ( .B1(n10441), .B2(n10431), .A(n10430), .ZN(n10438) );
  AOI21_X1 U12979 ( .B1(n10858), .B2(n10433), .A(n10432), .ZN(n14470) );
  INV_X1 U12980 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10435) );
  MUX2_X1 U12981 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n10435), .S(n10434), .Z(
        n14469) );
  NAND2_X1 U12982 ( .A1(n14470), .A2(n14469), .ZN(n14468) );
  NAND2_X1 U12983 ( .A1(n10441), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n11447) );
  OAI21_X1 U12984 ( .B1(n10441), .B2(P2_REG1_REG_11__SCAN_IN), .A(n11447), 
        .ZN(n10436) );
  AOI21_X1 U12985 ( .B1(n14468), .B2(n10437), .A(n10436), .ZN(n14482) );
  AOI211_X1 U12986 ( .C1(n10438), .C2(n14468), .A(n14483), .B(n14482), .ZN(
        n10439) );
  AOI211_X1 U12987 ( .C1(n14521), .C2(n10441), .A(n10440), .B(n10439), .ZN(
        n10442) );
  NAND2_X1 U12988 ( .A1(n10443), .A2(n10442), .ZN(P2_U3225) );
  XOR2_X1 U12989 ( .A(n10444), .B(n12118), .Z(n14783) );
  AOI22_X1 U12990 ( .A1(n10201), .A2(n12763), .B1(n12765), .B2(n12181), .ZN(
        n10448) );
  INV_X1 U12991 ( .A(n12118), .ZN(n10446) );
  OAI211_X1 U12992 ( .C1(n6603), .C2(n10446), .A(n12768), .B(n10445), .ZN(
        n10447) );
  OAI211_X1 U12993 ( .C1(n14783), .C2(n14808), .A(n10448), .B(n10447), .ZN(
        n14785) );
  NAND2_X1 U12994 ( .A1(n14785), .A2(n14770), .ZN(n10451) );
  OAI22_X1 U12995 ( .A1(n12757), .A2(n14782), .B1(n14755), .B2(
        P3_REG3_REG_3__SCAN_IN), .ZN(n10449) );
  AOI21_X1 U12996 ( .B1(n14772), .B2(P3_REG2_REG_3__SCAN_IN), .A(n10449), .ZN(
        n10450) );
  OAI211_X1 U12997 ( .C1(n14783), .C2(n11124), .A(n10451), .B(n10450), .ZN(
        P3_U3230) );
  INV_X1 U12998 ( .A(n10452), .ZN(n10454) );
  OAI222_X1 U12999 ( .A1(P3_U3151), .A2(n10455), .B1(n12880), .B2(n10454), 
        .C1(n10453), .C2(n12874), .ZN(P3_U3275) );
  OAI222_X1 U13000 ( .A1(n14012), .A2(n10457), .B1(n14014), .B2(n10456), .C1(
        n13711), .C2(P1_U3086), .ZN(P1_U3337) );
  AOI22_X1 U13001 ( .A1(n12364), .A2(n13595), .B1(n14335), .B2(n12365), .ZN(
        n10536) );
  INV_X1 U13002 ( .A(n10536), .ZN(n10460) );
  AOI22_X1 U13003 ( .A1(n14335), .A2(n12363), .B1(n12365), .B2(n13595), .ZN(
        n10461) );
  XOR2_X1 U13004 ( .A(n12366), .B(n10461), .Z(n10537) );
  XNOR2_X1 U13005 ( .A(n10538), .B(n10537), .ZN(n10466) );
  NAND2_X1 U13006 ( .A1(n13576), .A2(n10462), .ZN(n10463) );
  NAND2_X1 U13007 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n13639) );
  OAI211_X1 U13008 ( .C1(n14338), .C2(n13513), .A(n10463), .B(n13639), .ZN(
        n10464) );
  AOI21_X1 U13009 ( .B1(n14335), .B2(n14142), .A(n10464), .ZN(n10465) );
  OAI21_X1 U13010 ( .B1(n10466), .B2(n13564), .A(n10465), .ZN(P1_U3230) );
  INV_X1 U13011 ( .A(n10721), .ZN(n10477) );
  XNOR2_X1 U13012 ( .A(n10722), .B(n6420), .ZN(n10809) );
  XNOR2_X1 U13013 ( .A(n10809), .B(n10926), .ZN(n10470) );
  NAND2_X1 U13014 ( .A1(n10468), .A2(n10467), .ZN(n10469) );
  OAI21_X1 U13015 ( .B1(n10470), .B2(n10469), .A(n10823), .ZN(n10471) );
  NAND2_X1 U13016 ( .A1(n10471), .A2(n12509), .ZN(n10476) );
  OAI22_X1 U13017 ( .A1(n12180), .A2(n14762), .B1(n10818), .B2(n14760), .ZN(
        n10718) );
  OAI22_X1 U13018 ( .A1(n12518), .A2(n14794), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10472), .ZN(n10473) );
  AOI21_X1 U13019 ( .B1(n10718), .B2(n10474), .A(n10473), .ZN(n10475) );
  OAI211_X1 U13020 ( .C1(n10477), .C2(n12450), .A(n10476), .B(n10475), .ZN(
        P3_U3167) );
  OAI21_X1 U13021 ( .B1(n14610), .B2(n10479), .A(n10478), .ZN(n10489) );
  AOI21_X1 U13022 ( .B1(n10481), .B2(n8329), .A(n10480), .ZN(n10487) );
  OAI21_X1 U13023 ( .B1(n10483), .B2(P3_REG1_REG_1__SCAN_IN), .A(n10482), .ZN(
        n10484) );
  NAND2_X1 U13024 ( .A1(n14746), .A2(n10484), .ZN(n10486) );
  AOI22_X1 U13025 ( .A1(n14743), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10485) );
  OAI211_X1 U13026 ( .C1(n10487), .C2(n14750), .A(n10486), .B(n10485), .ZN(
        n10488) );
  AOI21_X1 U13027 ( .B1(n14735), .B2(n10489), .A(n10488), .ZN(n10490) );
  OAI21_X1 U13028 ( .B1(n10491), .B2(n14740), .A(n10490), .ZN(P3_U3183) );
  OAI21_X1 U13029 ( .B1(n10498), .B2(n10492), .A(n10266), .ZN(n10502) );
  NAND2_X1 U13030 ( .A1(n13037), .A2(n13070), .ZN(n10494) );
  NAND2_X1 U13031 ( .A1(n13038), .A2(n8149), .ZN(n10493) );
  NAND2_X1 U13032 ( .A1(n10494), .A2(n10493), .ZN(n10569) );
  AOI21_X1 U13033 ( .B1(n12999), .B2(n10569), .A(n10495), .ZN(n10497) );
  NAND2_X1 U13034 ( .A1(n6418), .A2(n14566), .ZN(n10496) );
  OAI211_X1 U13035 ( .C1(n13015), .C2(n10575), .A(n10497), .B(n10496), .ZN(
        n10501) );
  NOR4_X1 U13036 ( .A1(n11989), .A2(n10282), .A3(n10499), .A4(n10498), .ZN(
        n10500) );
  AOI211_X1 U13037 ( .C1(n13035), .C2(n10502), .A(n10501), .B(n10500), .ZN(
        n10503) );
  INV_X1 U13038 ( .A(n10503), .ZN(P2_U3202) );
  OR2_X1 U13039 ( .A1(n10507), .A2(n13070), .ZN(n10508) );
  INV_X1 U13040 ( .A(n10670), .ZN(n10509) );
  NAND2_X1 U13041 ( .A1(n10668), .A2(n10509), .ZN(n10511) );
  OR2_X1 U13042 ( .A1(n10694), .A2(n13069), .ZN(n10510) );
  OR2_X1 U13043 ( .A1(n10953), .A2(n13068), .ZN(n10512) );
  NAND2_X1 U13044 ( .A1(n10513), .A2(n10522), .ZN(n10514) );
  NAND2_X1 U13045 ( .A1(n10975), .A2(n10514), .ZN(n10894) );
  NAND2_X1 U13046 ( .A1(n10516), .A2(n10515), .ZN(n10671) );
  NAND2_X1 U13047 ( .A1(n10671), .A2(n10670), .ZN(n10669) );
  NAND2_X1 U13048 ( .A1(n10694), .A2(n10517), .ZN(n10518) );
  OR2_X1 U13049 ( .A1(n10953), .A2(n10742), .ZN(n10519) );
  NAND2_X1 U13050 ( .A1(n10943), .A2(n10519), .ZN(n10521) );
  NAND2_X1 U13051 ( .A1(n10953), .A2(n10742), .ZN(n10520) );
  AOI21_X1 U13052 ( .B1(n10523), .B2(n6977), .A(n13268), .ZN(n10524) );
  INV_X1 U13053 ( .A(n13066), .ZN(n10979) );
  OAI22_X1 U13054 ( .A1(n10742), .A2(n12995), .B1(n10979), .B2(n12997), .ZN(
        n10747) );
  AOI21_X1 U13055 ( .B1(n10524), .B2(n10847), .A(n10747), .ZN(n10897) );
  INV_X1 U13056 ( .A(n10890), .ZN(n10526) );
  INV_X1 U13057 ( .A(n10953), .ZN(n14583) );
  AND2_X2 U13058 ( .A1(n14583), .A2(n10950), .ZN(n10948) );
  NAND2_X1 U13059 ( .A1(n10526), .A2(n10948), .ZN(n10855) );
  OR2_X1 U13060 ( .A1(n10526), .A2(n10948), .ZN(n10527) );
  AND3_X1 U13061 ( .A1(n10855), .A2(n13379), .A3(n10527), .ZN(n10891) );
  AOI21_X1 U13062 ( .B1(n14567), .B2(n10890), .A(n10891), .ZN(n10528) );
  OAI211_X1 U13063 ( .C1(n14571), .C2(n10894), .A(n10897), .B(n10528), .ZN(
        n10530) );
  NAND2_X1 U13064 ( .A1(n10530), .A2(n10988), .ZN(n10529) );
  OAI21_X1 U13065 ( .B1(n10988), .B2(n9953), .A(n10529), .ZN(P2_U3507) );
  INV_X1 U13066 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10532) );
  NAND2_X1 U13067 ( .A1(n10530), .A2(n10992), .ZN(n10531) );
  OAI21_X1 U13068 ( .B1(n10992), .B2(n10532), .A(n10531), .ZN(P2_U3454) );
  INV_X1 U13069 ( .A(n10533), .ZN(n10535) );
  OAI222_X1 U13070 ( .A1(n12880), .A2(n10535), .B1(n12874), .B2(n10534), .C1(
        P3_U3151), .C2(n12163), .ZN(P3_U3274) );
  AOI22_X1 U13071 ( .A1(n10538), .A2(n10537), .B1(n7029), .B2(n10460), .ZN(
        n10876) );
  NAND2_X1 U13072 ( .A1(n10552), .A2(n12363), .ZN(n10540) );
  NAND2_X1 U13073 ( .A1(n12365), .A2(n13594), .ZN(n10539) );
  NAND2_X1 U13074 ( .A1(n10540), .A2(n10539), .ZN(n10542) );
  XNOR2_X1 U13075 ( .A(n10542), .B(n10541), .ZN(n10544) );
  AOI22_X1 U13076 ( .A1(n10552), .A2(n12365), .B1(n12364), .B2(n13594), .ZN(
        n10543) );
  AND2_X1 U13077 ( .A1(n10544), .A2(n10543), .ZN(n10875) );
  INV_X1 U13078 ( .A(n10875), .ZN(n10545) );
  OR2_X1 U13079 ( .A1(n10544), .A2(n10543), .ZN(n10874) );
  NAND2_X1 U13080 ( .A1(n10545), .A2(n10874), .ZN(n10546) );
  XNOR2_X1 U13081 ( .A(n10876), .B(n10546), .ZN(n10554) );
  NOR2_X1 U13082 ( .A1(n14146), .A2(n10547), .ZN(n10551) );
  NAND2_X1 U13083 ( .A1(n13557), .A2(n13595), .ZN(n10548) );
  NAND2_X1 U13084 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n13652) );
  OAI211_X1 U13085 ( .C1(n10549), .C2(n13570), .A(n10548), .B(n13652), .ZN(
        n10550) );
  AOI211_X1 U13086 ( .C1(n10552), .C2(n14142), .A(n10551), .B(n10550), .ZN(
        n10553) );
  OAI21_X1 U13087 ( .B1(n10554), .B2(n13564), .A(n10553), .ZN(P1_U3227) );
  INV_X1 U13088 ( .A(n10555), .ZN(n10558) );
  OAI222_X1 U13089 ( .A1(n14012), .A2(n10557), .B1(n14014), .B2(n10558), .C1(
        P1_U3086), .C2(n10556), .ZN(P1_U3336) );
  OAI222_X1 U13090 ( .A1(n12041), .A2(n10559), .B1(n13444), .B2(n10558), .C1(
        P2_U3088), .C2(n13093), .ZN(P2_U3308) );
  NAND2_X1 U13091 ( .A1(n9868), .A2(n10560), .ZN(n10561) );
  XNOR2_X1 U13092 ( .A(n10563), .B(n10562), .ZN(n14570) );
  NAND3_X1 U13093 ( .A1(n10564), .A2(n10566), .A3(n10565), .ZN(n10567) );
  AOI21_X1 U13094 ( .B1(n10568), .B2(n10567), .A(n13268), .ZN(n10570) );
  NOR2_X1 U13095 ( .A1(n10570), .A2(n10569), .ZN(n14568) );
  MUX2_X1 U13096 ( .A(n9640), .B(n14568), .S(n13257), .Z(n10578) );
  INV_X1 U13097 ( .A(n10776), .ZN(n10572) );
  AOI211_X1 U13098 ( .C1(n14566), .C2(n10572), .A(n13289), .B(n6924), .ZN(
        n14565) );
  INV_X1 U13099 ( .A(n10573), .ZN(n10574) );
  OAI22_X1 U13100 ( .A1(n13294), .A2(n8141), .B1(n13245), .B2(n10575), .ZN(
        n10576) );
  AOI21_X1 U13101 ( .B1(n13302), .B2(n14565), .A(n10576), .ZN(n10577) );
  OAI211_X1 U13102 ( .C1(n13299), .C2(n14570), .A(n10578), .B(n10577), .ZN(
        P2_U3261) );
  NOR2_X1 U13103 ( .A1(n14627), .A2(n10580), .ZN(n10581) );
  XNOR2_X1 U13104 ( .A(n10580), .B(n14627), .ZN(n14615) );
  NOR2_X1 U13105 ( .A1(n10595), .A2(n14615), .ZN(n14614) );
  NOR2_X1 U13106 ( .A1(n10581), .A2(n14614), .ZN(n14633) );
  OR2_X1 U13107 ( .A1(n14647), .A2(n10730), .ZN(n10583) );
  NAND2_X1 U13108 ( .A1(n14647), .A2(n10730), .ZN(n10582) );
  NAND2_X1 U13109 ( .A1(n10583), .A2(n10582), .ZN(n14632) );
  AND2_X2 U13110 ( .A1(n14630), .A2(n10583), .ZN(n10584) );
  XNOR2_X1 U13111 ( .A(n10584), .B(n14661), .ZN(n14652) );
  NOR2_X1 U13112 ( .A1(n14661), .A2(n10584), .ZN(n10585) );
  NAND2_X1 U13113 ( .A1(n10637), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10586) );
  OAI21_X1 U13114 ( .B1(n10637), .B2(P3_REG2_REG_6__SCAN_IN), .A(n10586), .ZN(
        n14669) );
  NOR2_X1 U13115 ( .A1(n10613), .A2(n10587), .ZN(n10588) );
  NOR2_X1 U13116 ( .A1(n10612), .A2(n14689), .ZN(n14688) );
  NAND2_X1 U13117 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n10636), .ZN(n10589) );
  OAI21_X1 U13118 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n10636), .A(n10589), .ZN(
        n14713) );
  NOR2_X1 U13119 ( .A1(n14714), .A2(n14713), .ZN(n14712) );
  NOR2_X1 U13120 ( .A1(n10625), .A2(n10590), .ZN(n10591) );
  AOI22_X1 U13121 ( .A1(n11198), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n10629), 
        .B2(n14033), .ZN(n10592) );
  AOI21_X1 U13122 ( .B1(n6595), .B2(n10592), .A(n11184), .ZN(n10667) );
  INV_X1 U13123 ( .A(n10593), .ZN(n14622) );
  INV_X1 U13124 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10594) );
  MUX2_X1 U13125 ( .A(n10595), .B(n10594), .S(n8681), .Z(n10596) );
  NAND2_X1 U13126 ( .A1(n10596), .A2(n14627), .ZN(n14641) );
  INV_X1 U13127 ( .A(n10596), .ZN(n10597) );
  NAND2_X1 U13128 ( .A1(n10597), .A2(n10644), .ZN(n10598) );
  AND2_X1 U13129 ( .A1(n14641), .A2(n10598), .ZN(n14621) );
  OAI21_X1 U13130 ( .B1(n14623), .B2(n14622), .A(n14621), .ZN(n14642) );
  INV_X1 U13131 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10640) );
  MUX2_X1 U13132 ( .A(n10730), .B(n10640), .S(n8681), .Z(n10599) );
  NAND2_X1 U13133 ( .A1(n10599), .A2(n14647), .ZN(n10602) );
  INV_X1 U13134 ( .A(n10599), .ZN(n10600) );
  NAND2_X1 U13135 ( .A1(n10600), .A2(n10639), .ZN(n10601) );
  NAND2_X1 U13136 ( .A1(n10602), .A2(n10601), .ZN(n14640) );
  AOI21_X1 U13137 ( .B1(n14642), .B2(n14641), .A(n14640), .ZN(n14655) );
  INV_X1 U13138 ( .A(n10602), .ZN(n14654) );
  INV_X1 U13139 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10603) );
  MUX2_X1 U13140 ( .A(n10720), .B(n10603), .S(n12073), .Z(n10604) );
  NAND2_X1 U13141 ( .A1(n10604), .A2(n14661), .ZN(n14678) );
  INV_X1 U13142 ( .A(n10604), .ZN(n10605) );
  NAND2_X1 U13143 ( .A1(n10605), .A2(n10648), .ZN(n10606) );
  AND2_X1 U13144 ( .A1(n14678), .A2(n10606), .ZN(n14653) );
  OAI21_X1 U13145 ( .B1(n14655), .B2(n14654), .A(n14653), .ZN(n14679) );
  INV_X1 U13146 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10638) );
  MUX2_X1 U13147 ( .A(n10929), .B(n10638), .S(n12073), .Z(n10607) );
  INV_X1 U13148 ( .A(n10637), .ZN(n14684) );
  NAND2_X1 U13149 ( .A1(n10607), .A2(n14684), .ZN(n10610) );
  INV_X1 U13150 ( .A(n10607), .ZN(n10608) );
  NAND2_X1 U13151 ( .A1(n10608), .A2(n10637), .ZN(n10609) );
  NAND2_X1 U13152 ( .A1(n10610), .A2(n10609), .ZN(n14677) );
  AOI21_X1 U13153 ( .B1(n14679), .B2(n14678), .A(n14677), .ZN(n14693) );
  INV_X1 U13154 ( .A(n10610), .ZN(n14692) );
  INV_X1 U13155 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n10611) );
  MUX2_X1 U13156 ( .A(n10612), .B(n10611), .S(n12073), .Z(n10614) );
  NAND2_X1 U13157 ( .A1(n10614), .A2(n10613), .ZN(n14707) );
  INV_X1 U13158 ( .A(n10614), .ZN(n10615) );
  NAND2_X1 U13159 ( .A1(n10615), .A2(n14697), .ZN(n10616) );
  AND2_X1 U13160 ( .A1(n14707), .A2(n10616), .ZN(n14691) );
  OAI21_X1 U13161 ( .B1(n14693), .B2(n14692), .A(n14691), .ZN(n14708) );
  INV_X1 U13162 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n10617) );
  MUX2_X1 U13163 ( .A(n10618), .B(n10617), .S(n12073), .Z(n10619) );
  NAND2_X1 U13164 ( .A1(n10619), .A2(n14719), .ZN(n10622) );
  INV_X1 U13165 ( .A(n10619), .ZN(n10620) );
  NAND2_X1 U13166 ( .A1(n10620), .A2(n10636), .ZN(n10621) );
  NAND2_X1 U13167 ( .A1(n10622), .A2(n10621), .ZN(n14706) );
  AOI21_X1 U13168 ( .B1(n14708), .B2(n14707), .A(n14706), .ZN(n14734) );
  INV_X1 U13169 ( .A(n10622), .ZN(n14733) );
  INV_X1 U13170 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n10623) );
  MUX2_X1 U13171 ( .A(n10624), .B(n10623), .S(n12073), .Z(n10626) );
  NAND2_X1 U13172 ( .A1(n10626), .A2(n10625), .ZN(n10634) );
  INV_X1 U13173 ( .A(n10626), .ZN(n10627) );
  NAND2_X1 U13174 ( .A1(n10627), .A2(n14739), .ZN(n10628) );
  AND2_X1 U13175 ( .A1(n10634), .A2(n10628), .ZN(n14732) );
  INV_X1 U13176 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n10657) );
  MUX2_X1 U13177 ( .A(n10629), .B(n10657), .S(n12073), .Z(n10630) );
  NAND2_X1 U13178 ( .A1(n10630), .A2(n11198), .ZN(n11190) );
  INV_X1 U13179 ( .A(n10630), .ZN(n10631) );
  NAND2_X1 U13180 ( .A1(n10631), .A2(n14033), .ZN(n10632) );
  NAND2_X1 U13181 ( .A1(n11190), .A2(n10632), .ZN(n10633) );
  AND3_X1 U13182 ( .A1(n14731), .A2(n10634), .A3(n10633), .ZN(n10635) );
  OAI21_X1 U13183 ( .B1(n11191), .B2(n10635), .A(n14735), .ZN(n10666) );
  NAND2_X1 U13184 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n10636), .ZN(n10654) );
  AOI22_X1 U13185 ( .A1(n14719), .A2(n10617), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n10636), .ZN(n14717) );
  NAND2_X1 U13186 ( .A1(n10637), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10651) );
  MUX2_X1 U13187 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n10638), .S(n10637), .Z(
        n14672) );
  NAND2_X1 U13188 ( .A1(n10639), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10647) );
  MUX2_X1 U13189 ( .A(n10640), .B(P3_REG1_REG_4__SCAN_IN), .S(n14647), .Z(
        n14635) );
  NAND2_X1 U13190 ( .A1(P3_REG1_REG_2__SCAN_IN), .A2(n10641), .ZN(n10643) );
  NAND2_X1 U13191 ( .A1(n10643), .A2(n10642), .ZN(n10645) );
  NAND2_X1 U13192 ( .A1(n10644), .A2(n10645), .ZN(n10646) );
  XOR2_X1 U13193 ( .A(n10645), .B(n10644), .Z(n14617) );
  NAND2_X1 U13194 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(n14617), .ZN(n14616) );
  NAND2_X1 U13195 ( .A1(n10648), .A2(n10649), .ZN(n10650) );
  NAND2_X1 U13196 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n14659), .ZN(n14658) );
  NAND2_X1 U13197 ( .A1(n14697), .A2(n10652), .ZN(n10653) );
  NAND2_X1 U13198 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n14701), .ZN(n14700) );
  NAND2_X1 U13199 ( .A1(n14739), .A2(n10655), .ZN(n10656) );
  NAND2_X1 U13200 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n14745), .ZN(n14744) );
  NOR2_X1 U13201 ( .A1(n11198), .A2(n10657), .ZN(n10658) );
  AOI21_X1 U13202 ( .B1(n11198), .B2(n10657), .A(n10658), .ZN(n10659) );
  OAI21_X1 U13203 ( .B1(n10660), .B2(n10659), .A(n11197), .ZN(n10664) );
  NAND2_X1 U13204 ( .A1(n14718), .A2(n11198), .ZN(n10661) );
  NAND2_X1 U13205 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n10964)
         );
  OAI211_X1 U13206 ( .C1(n10662), .C2(n14727), .A(n10661), .B(n10964), .ZN(
        n10663) );
  AOI21_X1 U13207 ( .B1(n10664), .B2(n14746), .A(n10663), .ZN(n10665) );
  OAI211_X1 U13208 ( .C1(n10667), .C2(n14750), .A(n10666), .B(n10665), .ZN(
        P3_U3192) );
  XNOR2_X1 U13209 ( .A(n10668), .B(n10670), .ZN(n14574) );
  INV_X1 U13210 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10676) );
  OAI21_X1 U13211 ( .B1(n10671), .B2(n10670), .A(n10669), .ZN(n10673) );
  OAI22_X1 U13212 ( .A1(n10672), .A2(n12995), .B1(n10742), .B2(n12997), .ZN(
        n10691) );
  AOI21_X1 U13213 ( .B1(n10673), .B2(n13284), .A(n10691), .ZN(n10674) );
  OAI21_X1 U13214 ( .B1(n9868), .B2(n14574), .A(n10674), .ZN(n14577) );
  INV_X1 U13215 ( .A(n14577), .ZN(n10675) );
  MUX2_X1 U13216 ( .A(n10676), .B(n10675), .S(n13257), .Z(n10682) );
  INV_X1 U13217 ( .A(n10694), .ZN(n14576) );
  INV_X1 U13218 ( .A(n10950), .ZN(n10677) );
  OAI211_X1 U13219 ( .C1(n14576), .C2(n10678), .A(n10677), .B(n13379), .ZN(
        n14575) );
  INV_X1 U13220 ( .A(n14575), .ZN(n10680) );
  OAI22_X1 U13221 ( .A1(n13294), .A2(n14576), .B1(n13245), .B2(n10690), .ZN(
        n10679) );
  AOI21_X1 U13222 ( .B1(n13302), .B2(n10680), .A(n10679), .ZN(n10681) );
  OAI211_X1 U13223 ( .C1(n14574), .C2(n13185), .A(n10682), .B(n10681), .ZN(
        P2_U3259) );
  MUX2_X1 U13224 ( .A(n9641), .B(n10683), .S(n13257), .Z(n10688) );
  OAI22_X1 U13225 ( .A1(n13294), .A2(n6923), .B1(n10684), .B2(n13245), .ZN(
        n10685) );
  AOI21_X1 U13226 ( .B1(n13302), .B2(n10686), .A(n10685), .ZN(n10687) );
  OAI211_X1 U13227 ( .C1(n10689), .C2(n13185), .A(n10688), .B(n10687), .ZN(
        P2_U3260) );
  INV_X1 U13228 ( .A(n10690), .ZN(n10710) );
  NAND2_X1 U13229 ( .A1(n12999), .A2(n10691), .ZN(n10692) );
  OAI211_X1 U13230 ( .C1(n13045), .C2(n14576), .A(n10693), .B(n10692), .ZN(
        n10709) );
  XNOR2_X1 U13231 ( .A(n10694), .B(n12948), .ZN(n10865) );
  AND2_X1 U13232 ( .A1(n12916), .A2(n13069), .ZN(n10695) );
  NAND2_X1 U13233 ( .A1(n10865), .A2(n10695), .ZN(n10734) );
  INV_X1 U13234 ( .A(n10865), .ZN(n10697) );
  INV_X1 U13235 ( .A(n10695), .ZN(n10696) );
  NAND2_X1 U13236 ( .A1(n10697), .A2(n10696), .ZN(n10698) );
  NAND2_X1 U13237 ( .A1(n10734), .A2(n10698), .ZN(n10707) );
  INV_X1 U13238 ( .A(n10699), .ZN(n10701) );
  NAND2_X1 U13239 ( .A1(n10701), .A2(n10700), .ZN(n10702) );
  NAND2_X1 U13240 ( .A1(n10703), .A2(n10702), .ZN(n10706) );
  INV_X1 U13241 ( .A(n10706), .ZN(n10705) );
  INV_X1 U13242 ( .A(n10707), .ZN(n10704) );
  NAND2_X1 U13243 ( .A1(n10705), .A2(n10704), .ZN(n10735) );
  INV_X1 U13244 ( .A(n10735), .ZN(n10867) );
  AOI211_X1 U13245 ( .C1(n10707), .C2(n10706), .A(n13023), .B(n10867), .ZN(
        n10708) );
  AOI211_X1 U13246 ( .C1(n13042), .C2(n10710), .A(n10709), .B(n10708), .ZN(
        n10711) );
  INV_X1 U13247 ( .A(n10711), .ZN(P2_U3211) );
  NAND2_X1 U13248 ( .A1(n14808), .A2(n10712), .ZN(n10713) );
  XOR2_X1 U13249 ( .A(n10714), .B(n12186), .Z(n14795) );
  OAI21_X1 U13250 ( .B1(n10717), .B2(n10716), .A(n10715), .ZN(n10719) );
  AOI21_X1 U13251 ( .B1(n10719), .B2(n12768), .A(n10718), .ZN(n14793) );
  MUX2_X1 U13252 ( .A(n10720), .B(n14793), .S(n14770), .Z(n10724) );
  AOI22_X1 U13253 ( .A1(n12773), .A2(n10722), .B1(n12755), .B2(n10721), .ZN(
        n10723) );
  OAI211_X1 U13254 ( .C1(n12663), .C2(n14795), .A(n10724), .B(n10723), .ZN(
        P3_U3228) );
  XNOR2_X1 U13255 ( .A(n10725), .B(n12121), .ZN(n14787) );
  OAI211_X1 U13256 ( .C1(n10727), .C2(n12121), .A(n10726), .B(n12768), .ZN(
        n10729) );
  AND2_X1 U13257 ( .A1(n10729), .A2(n10728), .ZN(n14788) );
  MUX2_X1 U13258 ( .A(n14788), .B(n10730), .S(n14772), .Z(n10733) );
  AOI22_X1 U13259 ( .A1(n12773), .A2(n14791), .B1(n12755), .B2(n10731), .ZN(
        n10732) );
  OAI211_X1 U13260 ( .C1(n12663), .C2(n14787), .A(n10733), .B(n10732), .ZN(
        P3_U3229) );
  XNOR2_X1 U13261 ( .A(n10953), .B(n12948), .ZN(n10736) );
  AND2_X1 U13262 ( .A1(n12916), .A2(n13068), .ZN(n10737) );
  NAND2_X1 U13263 ( .A1(n10736), .A2(n10737), .ZN(n10744) );
  INV_X1 U13264 ( .A(n10736), .ZN(n10741) );
  INV_X1 U13265 ( .A(n10737), .ZN(n10738) );
  NAND2_X1 U13266 ( .A1(n10741), .A2(n10738), .ZN(n10739) );
  AND2_X1 U13267 ( .A1(n10744), .A2(n10739), .ZN(n10866) );
  INV_X1 U13268 ( .A(n10746), .ZN(n10868) );
  NOR3_X1 U13269 ( .A1(n11989), .A2(n10742), .A3(n10741), .ZN(n10743) );
  AOI21_X1 U13270 ( .B1(n10868), .B2(n13035), .A(n10743), .ZN(n10753) );
  XNOR2_X1 U13271 ( .A(n10890), .B(n12948), .ZN(n10902) );
  NAND2_X1 U13272 ( .A1(n12916), .A2(n13067), .ZN(n10898) );
  AOI22_X1 U13273 ( .A1(n12999), .A2(n10747), .B1(P2_REG3_REG_8__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10749) );
  NAND2_X1 U13274 ( .A1(n6418), .A2(n10890), .ZN(n10748) );
  OAI211_X1 U13275 ( .C1(n13015), .C2(n10888), .A(n10749), .B(n10748), .ZN(
        n10750) );
  AOI21_X1 U13276 ( .B1(n6593), .B2(n13035), .A(n10750), .ZN(n10751) );
  OAI21_X1 U13277 ( .B1(n10753), .B2(n10752), .A(n10751), .ZN(P2_U3193) );
  NAND2_X1 U13278 ( .A1(n10755), .A2(n10754), .ZN(n10757) );
  OR2_X1 U13279 ( .A1(n11045), .A2(n13592), .ZN(n10756) );
  XNOR2_X1 U13280 ( .A(n10785), .B(n10789), .ZN(n14367) );
  INV_X1 U13281 ( .A(n10759), .ZN(n10761) );
  INV_X1 U13282 ( .A(n10800), .ZN(n10760) );
  OAI211_X1 U13283 ( .C1(n14364), .C2(n10761), .A(n10760), .B(n14310), .ZN(
        n14363) );
  AOI22_X1 U13284 ( .A1(n11258), .A2(n14306), .B1(n11253), .B2(n14285), .ZN(
        n10762) );
  OAI21_X1 U13285 ( .B1(n14363), .B2(n14160), .A(n10762), .ZN(n10769) );
  INV_X1 U13286 ( .A(n10763), .ZN(n10765) );
  XNOR2_X1 U13287 ( .A(n10790), .B(n10789), .ZN(n10767) );
  AOI22_X1 U13288 ( .A1(n14292), .A2(n13590), .B1(n14131), .B2(n13592), .ZN(
        n11256) );
  OAI21_X1 U13289 ( .B1(n10767), .B2(n14357), .A(n11256), .ZN(n14365) );
  MUX2_X1 U13290 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n14365), .S(n14303), .Z(
        n10768) );
  AOI211_X1 U13291 ( .C1(n14315), .C2(n14367), .A(n10769), .B(n10768), .ZN(
        n10770) );
  INV_X1 U13292 ( .A(n10770), .ZN(P1_U3285) );
  XNOR2_X1 U13293 ( .A(n10779), .B(n10771), .ZN(n14557) );
  NAND2_X1 U13294 ( .A1(n10773), .A2(n10772), .ZN(n10774) );
  NAND2_X1 U13295 ( .A1(n10774), .A2(n13379), .ZN(n10775) );
  NOR2_X1 U13296 ( .A1(n10776), .A2(n10775), .ZN(n14558) );
  OAI22_X1 U13297 ( .A1(n13294), .A2(n14561), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13245), .ZN(n10777) );
  AOI21_X1 U13298 ( .B1(n13302), .B2(n14558), .A(n10777), .ZN(n10784) );
  OAI21_X1 U13299 ( .B1(n10779), .B2(n10778), .A(n10564), .ZN(n10782) );
  INV_X1 U13300 ( .A(n10780), .ZN(n10781) );
  AOI21_X1 U13301 ( .B1(n10782), .B2(n13284), .A(n10781), .ZN(n14560) );
  MUX2_X1 U13302 ( .A(n9639), .B(n14560), .S(n13257), .Z(n10783) );
  OAI211_X1 U13303 ( .C1(n14557), .C2(n13299), .A(n10784), .B(n10783), .ZN(
        P2_U3262) );
  NAND2_X1 U13304 ( .A1(n10785), .A2(n10789), .ZN(n10787) );
  NAND2_X1 U13305 ( .A1(n10787), .A2(n10786), .ZN(n11223) );
  XNOR2_X1 U13306 ( .A(n11223), .B(n11222), .ZN(n10797) );
  INV_X1 U13307 ( .A(n14131), .ZN(n13890) );
  OAI22_X1 U13308 ( .A1(n13890), .A2(n11246), .B1(n11572), .B2(n13892), .ZN(
        n10796) );
  NAND2_X1 U13309 ( .A1(n10792), .A2(n10791), .ZN(n11230) );
  NAND2_X1 U13310 ( .A1(n10793), .A2(n11222), .ZN(n10794) );
  AOI21_X1 U13311 ( .B1(n11230), .B2(n10794), .A(n14357), .ZN(n10795) );
  AOI211_X1 U13312 ( .C1(n10797), .C2(n14375), .A(n10796), .B(n10795), .ZN(
        n11024) );
  INV_X1 U13313 ( .A(n11423), .ZN(n10798) );
  OAI22_X1 U13314 ( .A1(n14303), .A2(n10799), .B1(n10798), .B2(n14302), .ZN(
        n10802) );
  NAND2_X1 U13315 ( .A1(n10800), .A2(n11426), .ZN(n14290) );
  OAI211_X1 U13316 ( .C1(n10800), .C2(n11426), .A(n14310), .B(n14290), .ZN(
        n11023) );
  NOR2_X1 U13317 ( .A1(n11023), .A2(n14160), .ZN(n10801) );
  AOI211_X1 U13318 ( .C1(n14306), .C2(n10803), .A(n10802), .B(n10801), .ZN(
        n10804) );
  OAI21_X1 U13319 ( .B1(n11024), .B2(n14284), .A(n10804), .ZN(P1_U3284) );
  NOR2_X1 U13320 ( .A1(n12874), .A2(SI_22_), .ZN(n10805) );
  AOI21_X1 U13321 ( .B1(n12161), .B2(P3_STATE_REG_SCAN_IN), .A(n10805), .ZN(
        n10806) );
  OAI21_X1 U13322 ( .B1(n10807), .B2(n12880), .A(n10806), .ZN(n10808) );
  INV_X1 U13323 ( .A(n10808), .ZN(P3_U3273) );
  INV_X1 U13324 ( .A(n10809), .ZN(n10810) );
  NAND2_X1 U13325 ( .A1(n10810), .A2(n10926), .ZN(n10820) );
  NAND2_X1 U13326 ( .A1(n10823), .A2(n10820), .ZN(n10937) );
  XNOR2_X1 U13327 ( .A(n10933), .B(n12444), .ZN(n10817) );
  XNOR2_X1 U13328 ( .A(n10817), .B(n10818), .ZN(n10938) );
  NOR2_X1 U13329 ( .A1(n10937), .A2(n10938), .ZN(n10936) );
  NOR2_X1 U13330 ( .A1(n10818), .A2(n10817), .ZN(n10825) );
  NOR2_X1 U13331 ( .A1(n10936), .A2(n10825), .ZN(n11054) );
  XNOR2_X1 U13332 ( .A(n10914), .B(n12444), .ZN(n10824) );
  XNOR2_X1 U13333 ( .A(n11054), .B(n10824), .ZN(n10816) );
  NAND2_X1 U13334 ( .A1(n12554), .A2(n12763), .ZN(n10812) );
  NAND2_X1 U13335 ( .A1(n12551), .A2(n12765), .ZN(n10811) );
  AND2_X1 U13336 ( .A1(n10812), .A2(n10811), .ZN(n10916) );
  AOI22_X1 U13337 ( .A1(n12528), .A2(n14811), .B1(P3_REG3_REG_7__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10813) );
  OAI21_X1 U13338 ( .B1(n10916), .B2(n12503), .A(n10813), .ZN(n10814) );
  AOI21_X1 U13339 ( .B1(n10918), .B2(n12523), .A(n10814), .ZN(n10815) );
  OAI21_X1 U13340 ( .B1(n10816), .B2(n12531), .A(n10815), .ZN(P3_U3153) );
  XNOR2_X1 U13341 ( .A(n10838), .B(n12444), .ZN(n10958) );
  XNOR2_X1 U13342 ( .A(n10958), .B(n11057), .ZN(n10835) );
  XNOR2_X1 U13343 ( .A(n14815), .B(n12444), .ZN(n10828) );
  XNOR2_X1 U13344 ( .A(n10828), .B(n12207), .ZN(n10826) );
  NAND2_X1 U13345 ( .A1(n10818), .A2(n10817), .ZN(n10819) );
  NAND3_X1 U13346 ( .A1(n10826), .A2(n10820), .A3(n10819), .ZN(n10821) );
  NOR2_X1 U13347 ( .A1(n10824), .A2(n10821), .ZN(n10822) );
  INV_X1 U13348 ( .A(n10826), .ZN(n11055) );
  OAI21_X1 U13349 ( .B1(n11058), .B2(n11055), .A(n10824), .ZN(n10830) );
  INV_X1 U13350 ( .A(n10824), .ZN(n11053) );
  NAND2_X1 U13351 ( .A1(n10826), .A2(n10825), .ZN(n10827) );
  NAND2_X1 U13352 ( .A1(n11053), .A2(n10827), .ZN(n10829) );
  AOI22_X1 U13353 ( .A1(n10830), .A2(n10829), .B1(n10828), .B2(n12551), .ZN(
        n10831) );
  INV_X1 U13354 ( .A(n10835), .ZN(n10832) );
  INV_X1 U13355 ( .A(n10961), .ZN(n10833) );
  AOI21_X1 U13356 ( .B1(n10835), .B2(n10834), .A(n10833), .ZN(n10841) );
  NOR2_X1 U13357 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10836), .ZN(n14742) );
  OAI22_X1 U13358 ( .A1(n12207), .A2(n12475), .B1(n11317), .B2(n12526), .ZN(
        n10837) );
  AOI211_X1 U13359 ( .C1(n12528), .C2(n10838), .A(n14742), .B(n10837), .ZN(
        n10840) );
  NAND2_X1 U13360 ( .A1(n12523), .A2(n11119), .ZN(n10839) );
  OAI211_X1 U13361 ( .C1(n10841), .C2(n12531), .A(n10840), .B(n10839), .ZN(
        P3_U3171) );
  NAND2_X1 U13362 ( .A1(n10890), .A2(n13067), .ZN(n10970) );
  NAND2_X1 U13363 ( .A1(n10975), .A2(n10970), .ZN(n10842) );
  INV_X1 U13364 ( .A(n10849), .ZN(n10972) );
  NAND2_X1 U13365 ( .A1(n10842), .A2(n10972), .ZN(n10844) );
  OR2_X1 U13366 ( .A1(n10842), .A2(n10972), .ZN(n10843) );
  NAND2_X1 U13367 ( .A1(n10844), .A2(n10843), .ZN(n11095) );
  INV_X1 U13368 ( .A(n13067), .ZN(n10845) );
  OR2_X1 U13369 ( .A1(n10890), .A2(n10845), .ZN(n10846) );
  INV_X1 U13370 ( .A(n10850), .ZN(n10848) );
  AOI21_X1 U13371 ( .B1(n10848), .B2(n10972), .A(n13268), .ZN(n10853) );
  NAND2_X1 U13372 ( .A1(n13037), .A2(n13065), .ZN(n10852) );
  NAND2_X1 U13373 ( .A1(n13038), .A2(n13067), .ZN(n10851) );
  NAND2_X1 U13374 ( .A1(n10852), .A2(n10851), .ZN(n10900) );
  AOI21_X1 U13375 ( .B1(n10853), .B2(n10981), .A(n10900), .ZN(n11100) );
  INV_X1 U13376 ( .A(n10985), .ZN(n10854) );
  AOI211_X1 U13377 ( .C1(n11090), .C2(n10855), .A(n13289), .B(n10854), .ZN(
        n11098) );
  AOI21_X1 U13378 ( .B1(n14567), .B2(n11090), .A(n11098), .ZN(n10856) );
  OAI211_X1 U13379 ( .C1(n14571), .C2(n11095), .A(n11100), .B(n10856), .ZN(
        n10859) );
  NAND2_X1 U13380 ( .A1(n10859), .A2(n10988), .ZN(n10857) );
  OAI21_X1 U13381 ( .B1(n10988), .B2(n10858), .A(n10857), .ZN(P2_U3508) );
  INV_X1 U13382 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10861) );
  NAND2_X1 U13383 ( .A1(n10859), .A2(n10992), .ZN(n10860) );
  OAI21_X1 U13384 ( .B1(n10992), .B2(n10861), .A(n10860), .ZN(P2_U3457) );
  NAND2_X1 U13385 ( .A1(n13037), .A2(n13067), .ZN(n10863) );
  NAND2_X1 U13386 ( .A1(n13038), .A2(n13069), .ZN(n10862) );
  NAND2_X1 U13387 ( .A1(n10863), .A2(n10862), .ZN(n10944) );
  AND2_X1 U13388 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n14437) );
  AOI21_X1 U13389 ( .B1(n12999), .B2(n10944), .A(n14437), .ZN(n10864) );
  OAI21_X1 U13390 ( .B1(n13015), .B2(n10951), .A(n10864), .ZN(n10872) );
  NAND3_X1 U13391 ( .A1(n13013), .A2(n13069), .A3(n10865), .ZN(n10870) );
  OAI21_X1 U13392 ( .B1(n10867), .B2(n10866), .A(n13035), .ZN(n10869) );
  AOI21_X1 U13393 ( .B1(n10870), .B2(n10869), .A(n10868), .ZN(n10871) );
  AOI211_X1 U13394 ( .C1(n10953), .C2(n6418), .A(n10872), .B(n10871), .ZN(
        n10873) );
  INV_X1 U13395 ( .A(n10873), .ZN(P2_U3185) );
  NAND2_X1 U13396 ( .A1(n14346), .A2(n12363), .ZN(n10878) );
  NAND2_X1 U13397 ( .A1(n12365), .A2(n13593), .ZN(n10877) );
  NAND2_X1 U13398 ( .A1(n10878), .A2(n10877), .ZN(n10879) );
  XNOR2_X1 U13399 ( .A(n10879), .B(n12366), .ZN(n11038) );
  AOI22_X1 U13400 ( .A1(n14346), .A2(n12365), .B1(n12364), .B2(n13593), .ZN(
        n11039) );
  XNOR2_X1 U13401 ( .A(n11038), .B(n11039), .ZN(n10880) );
  OAI211_X1 U13402 ( .C1(n10881), .C2(n10880), .A(n11041), .B(n14139), .ZN(
        n10886) );
  NOR2_X1 U13403 ( .A1(n13513), .A2(n14343), .ZN(n10882) );
  AOI211_X1 U13404 ( .C1(n13576), .C2(n10884), .A(n10883), .B(n10882), .ZN(
        n10885) );
  OAI211_X1 U13405 ( .C1(n10887), .C2(n13579), .A(n10886), .B(n10885), .ZN(
        P1_U3239) );
  OAI22_X1 U13406 ( .A1(n13257), .A2(n9943), .B1(n10888), .B2(n13245), .ZN(
        n10889) );
  AOI21_X1 U13407 ( .B1(n13241), .B2(n10890), .A(n10889), .ZN(n10893) );
  NAND2_X1 U13408 ( .A1(n10891), .A2(n13302), .ZN(n10892) );
  OAI211_X1 U13409 ( .C1(n10894), .C2(n13299), .A(n10893), .B(n10892), .ZN(
        n10895) );
  INV_X1 U13410 ( .A(n10895), .ZN(n10896) );
  OAI21_X1 U13411 ( .B1(n10897), .B2(n13304), .A(n10896), .ZN(P2_U3257) );
  INV_X1 U13412 ( .A(n10902), .ZN(n10899) );
  XNOR2_X1 U13413 ( .A(n11090), .B(n12948), .ZN(n11151) );
  NAND2_X1 U13414 ( .A1(n12916), .A2(n13066), .ZN(n11152) );
  XNOR2_X1 U13415 ( .A(n11151), .B(n11152), .ZN(n10903) );
  AOI22_X1 U13416 ( .A1(n12999), .A2(n10900), .B1(P2_REG3_REG_9__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10901) );
  OAI21_X1 U13417 ( .B1(n13015), .B2(n11091), .A(n10901), .ZN(n10906) );
  AOI22_X1 U13418 ( .A1(n13013), .A2(n13067), .B1(n13035), .B2(n10902), .ZN(
        n10904) );
  NOR3_X1 U13419 ( .A1(n6593), .A2(n10904), .A3(n10903), .ZN(n10905) );
  AOI211_X1 U13420 ( .C1(n11090), .C2(n6418), .A(n10906), .B(n10905), .ZN(
        n10907) );
  OAI21_X1 U13421 ( .B1(n11155), .B2(n13023), .A(n10907), .ZN(P2_U3203) );
  XNOR2_X1 U13422 ( .A(n10908), .B(n10914), .ZN(n14807) );
  NAND2_X1 U13423 ( .A1(n10715), .A2(n10909), .ZN(n11106) );
  OR2_X1 U13424 ( .A1(n11106), .A2(n12113), .ZN(n10927) );
  NAND2_X1 U13425 ( .A1(n10927), .A2(n10910), .ZN(n10915) );
  OR2_X1 U13426 ( .A1(n11106), .A2(n10911), .ZN(n11010) );
  AND2_X1 U13427 ( .A1(n11010), .A2(n10912), .ZN(n10913) );
  OAI211_X1 U13428 ( .C1(n10915), .C2(n10914), .A(n10913), .B(n12768), .ZN(
        n10917) );
  NAND2_X1 U13429 ( .A1(n10917), .A2(n10916), .ZN(n14810) );
  NAND2_X1 U13430 ( .A1(n14810), .A2(n14770), .ZN(n10922) );
  INV_X1 U13431 ( .A(n10918), .ZN(n10919) );
  OAI22_X1 U13432 ( .A1(n12757), .A2(n12201), .B1(n10919), .B2(n14755), .ZN(
        n10920) );
  AOI21_X1 U13433 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n14772), .A(n10920), .ZN(
        n10921) );
  OAI211_X1 U13434 ( .C1(n12663), .C2(n14807), .A(n10922), .B(n10921), .ZN(
        P3_U3226) );
  OR2_X1 U13435 ( .A1(n10923), .A2(n12113), .ZN(n10924) );
  AOI21_X1 U13436 ( .B1(n11106), .B2(n12113), .A(n14767), .ZN(n10928) );
  OAI22_X1 U13437 ( .A1(n11058), .A2(n14760), .B1(n10926), .B2(n14762), .ZN(
        n10932) );
  AOI21_X1 U13438 ( .B1(n10928), .B2(n10927), .A(n10932), .ZN(n14801) );
  MUX2_X1 U13439 ( .A(n14801), .B(n10929), .S(n14772), .Z(n10931) );
  AOI22_X1 U13440 ( .A1(n12773), .A2(n10933), .B1(n12755), .B2(n10941), .ZN(
        n10930) );
  OAI211_X1 U13441 ( .C1(n12663), .C2(n14800), .A(n10931), .B(n10930), .ZN(
        P3_U3227) );
  INV_X1 U13442 ( .A(n10932), .ZN(n10935) );
  AOI22_X1 U13443 ( .A1(n12528), .A2(n10933), .B1(P3_REG3_REG_6__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10934) );
  OAI21_X1 U13444 ( .B1(n10935), .B2(n12503), .A(n10934), .ZN(n10940) );
  AOI211_X1 U13445 ( .C1(n10938), .C2(n10937), .A(n12531), .B(n10936), .ZN(
        n10939) );
  AOI211_X1 U13446 ( .C1(n10941), .C2(n12523), .A(n10940), .B(n10939), .ZN(
        n10942) );
  INV_X1 U13447 ( .A(n10942), .ZN(P3_U3179) );
  XOR2_X1 U13448 ( .A(n10943), .B(n10946), .Z(n10945) );
  AOI21_X1 U13449 ( .B1(n10945), .B2(n13284), .A(n10944), .ZN(n14584) );
  XNOR2_X1 U13450 ( .A(n10947), .B(n10946), .ZN(n14587) );
  INV_X1 U13451 ( .A(n13299), .ZN(n13232) );
  INV_X1 U13452 ( .A(n10948), .ZN(n10949) );
  OAI211_X1 U13453 ( .C1(n14583), .C2(n10950), .A(n10949), .B(n13379), .ZN(
        n14582) );
  OAI22_X1 U13454 ( .A1(n13257), .A2(n9942), .B1(n10951), .B2(n13245), .ZN(
        n10952) );
  AOI21_X1 U13455 ( .B1(n13241), .B2(n10953), .A(n10952), .ZN(n10954) );
  OAI21_X1 U13456 ( .B1(n13170), .B2(n14582), .A(n10954), .ZN(n10955) );
  AOI21_X1 U13457 ( .B1(n14587), .B2(n13232), .A(n10955), .ZN(n10956) );
  OAI21_X1 U13458 ( .B1(n14584), .B2(n13304), .A(n10956), .ZN(P2_U3258) );
  INV_X1 U13459 ( .A(n10957), .ZN(n11034) );
  NAND2_X1 U13460 ( .A1(n10958), .A2(n11057), .ZN(n10959) );
  AND2_X1 U13461 ( .A1(n10961), .A2(n10959), .ZN(n10963) );
  XNOR2_X1 U13462 ( .A(n10967), .B(n6420), .ZN(n11312) );
  XNOR2_X1 U13463 ( .A(n11312), .B(n11317), .ZN(n10962) );
  AND2_X1 U13464 ( .A1(n10962), .A2(n10959), .ZN(n10960) );
  OAI211_X1 U13465 ( .C1(n10963), .C2(n10962), .A(n12509), .B(n11314), .ZN(
        n10969) );
  NAND2_X1 U13466 ( .A1(n12550), .A2(n12522), .ZN(n10965) );
  OAI211_X1 U13467 ( .C1(n11315), .C2(n12526), .A(n10965), .B(n10964), .ZN(
        n10966) );
  AOI21_X1 U13468 ( .B1(n10967), .B2(n12528), .A(n10966), .ZN(n10968) );
  OAI211_X1 U13469 ( .C1(n11034), .C2(n12450), .A(n10969), .B(n10968), .ZN(
        P3_U3157) );
  NAND2_X1 U13470 ( .A1(n11090), .A2(n13066), .ZN(n10971) );
  AND2_X1 U13471 ( .A1(n10970), .A2(n10971), .ZN(n10974) );
  INV_X1 U13472 ( .A(n10971), .ZN(n10973) );
  INV_X1 U13473 ( .A(n10982), .ZN(n10976) );
  NAND2_X1 U13474 ( .A1(n10977), .A2(n10976), .ZN(n11065) );
  OR2_X1 U13475 ( .A1(n10977), .A2(n10976), .ZN(n10978) );
  NAND2_X1 U13476 ( .A1(n11065), .A2(n10978), .ZN(n11084) );
  OR2_X1 U13477 ( .A1(n11090), .A2(n10979), .ZN(n10980) );
  OAI211_X1 U13478 ( .C1(n10983), .C2(n10982), .A(n11067), .B(n13284), .ZN(
        n10984) );
  AOI22_X1 U13479 ( .A1(n13038), .A2(n13066), .B1(n13037), .B2(n13064), .ZN(
        n11161) );
  AND2_X1 U13480 ( .A1(n10984), .A2(n11161), .ZN(n11089) );
  NOR2_X2 U13481 ( .A1(n11146), .A2(n10985), .ZN(n11076) );
  AOI211_X1 U13482 ( .C1(n11146), .C2(n10985), .A(n13289), .B(n11076), .ZN(
        n11087) );
  AOI21_X1 U13483 ( .B1(n14567), .B2(n11146), .A(n11087), .ZN(n10986) );
  OAI211_X1 U13484 ( .C1(n14571), .C2(n11084), .A(n11089), .B(n10986), .ZN(
        n10989) );
  NAND2_X1 U13485 ( .A1(n10989), .A2(n10988), .ZN(n10987) );
  OAI21_X1 U13486 ( .B1(n10988), .B2(n10435), .A(n10987), .ZN(P2_U3509) );
  INV_X1 U13487 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10991) );
  NAND2_X1 U13488 ( .A1(n10989), .A2(n10992), .ZN(n10990) );
  OAI21_X1 U13489 ( .B1(n10992), .B2(n10991), .A(n10990), .ZN(P2_U3460) );
  INV_X1 U13490 ( .A(n10993), .ZN(n11021) );
  OAI222_X1 U13491 ( .A1(n13444), .A2(n11021), .B1(n10995), .B2(P2_U3088), 
        .C1(n10994), .C2(n12041), .ZN(P2_U3307) );
  INV_X1 U13492 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n14408) );
  OAI22_X1 U13493 ( .A1(n13257), .A2(n10996), .B1(n14408), .B2(n13245), .ZN(
        n10999) );
  AOI211_X1 U13494 ( .C1(n13257), .C2(n11000), .A(n10999), .B(n10998), .ZN(
        n11001) );
  OAI21_X1 U13495 ( .B1(n13299), .B2(n11002), .A(n11001), .ZN(P2_U3263) );
  OAI22_X1 U13496 ( .A1(n13257), .A2(n6771), .B1(n14393), .B2(n13245), .ZN(
        n11006) );
  OAI22_X1 U13497 ( .A1(n13170), .A2(n11004), .B1(n11003), .B2(n13294), .ZN(
        n11005) );
  AOI211_X1 U13498 ( .C1(n13257), .C2(n11007), .A(n11006), .B(n11005), .ZN(
        n11008) );
  OAI21_X1 U13499 ( .B1(n13299), .B2(n11009), .A(n11008), .ZN(P2_U3264) );
  NAND2_X1 U13500 ( .A1(n11010), .A2(n11107), .ZN(n11011) );
  INV_X1 U13501 ( .A(n12205), .ZN(n12122) );
  XNOR2_X1 U13502 ( .A(n11011), .B(n12122), .ZN(n11015) );
  XNOR2_X1 U13503 ( .A(n11012), .B(n12205), .ZN(n14814) );
  INV_X1 U13504 ( .A(n14808), .ZN(n14805) );
  OAI22_X1 U13505 ( .A1(n11058), .A2(n14762), .B1(n11057), .B2(n14760), .ZN(
        n11013) );
  AOI21_X1 U13506 ( .B1(n14814), .B2(n14805), .A(n11013), .ZN(n11014) );
  OAI21_X1 U13507 ( .B1(n11015), .B2(n14767), .A(n11014), .ZN(n14818) );
  INV_X1 U13508 ( .A(n14818), .ZN(n11019) );
  AOI22_X1 U13509 ( .A1(n12773), .A2(n12208), .B1(n12755), .B2(n11061), .ZN(
        n11016) );
  OAI21_X1 U13510 ( .B1(n10618), .B2(n14770), .A(n11016), .ZN(n11017) );
  AOI21_X1 U13511 ( .B1(n14814), .B2(n12678), .A(n11017), .ZN(n11018) );
  OAI21_X1 U13512 ( .B1(n11019), .B2(n14772), .A(n11018), .ZN(P3_U3225) );
  OAI222_X1 U13513 ( .A1(n14012), .A2(n11022), .B1(n14014), .B2(n11021), .C1(
        n11020), .C2(P1_U3086), .ZN(P1_U3335) );
  INV_X1 U13514 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11026) );
  OAI211_X1 U13515 ( .C1(n11426), .C2(n14371), .A(n11024), .B(n11023), .ZN(
        n11027) );
  NAND2_X1 U13516 ( .A1(n11027), .A2(n14378), .ZN(n11025) );
  OAI21_X1 U13517 ( .B1(n14378), .B2(n11026), .A(n11025), .ZN(P1_U3486) );
  NAND2_X1 U13518 ( .A1(n11027), .A2(n14391), .ZN(n11028) );
  OAI21_X1 U13519 ( .B1(n14391), .B2(n11029), .A(n11028), .ZN(P1_U3537) );
  INV_X1 U13520 ( .A(n11032), .ZN(n12216) );
  XNOR2_X1 U13521 ( .A(n11030), .B(n12216), .ZN(n14829) );
  XNOR2_X1 U13522 ( .A(n11031), .B(n11032), .ZN(n11033) );
  OAI222_X1 U13523 ( .A1(n14760), .A2(n11315), .B1(n14762), .B2(n11057), .C1(
        n11033), .C2(n14767), .ZN(n14831) );
  NAND2_X1 U13524 ( .A1(n14831), .A2(n14770), .ZN(n11037) );
  OAI22_X1 U13525 ( .A1(n12757), .A2(n14826), .B1(n11034), .B2(n14755), .ZN(
        n11035) );
  AOI21_X1 U13526 ( .B1(n14772), .B2(P3_REG2_REG_10__SCAN_IN), .A(n11035), 
        .ZN(n11036) );
  OAI211_X1 U13527 ( .C1(n14829), .C2(n12663), .A(n11037), .B(n11036), .ZN(
        P3_U3223) );
  INV_X1 U13528 ( .A(n11038), .ZN(n11040) );
  NAND2_X1 U13529 ( .A1(n11045), .A2(n12363), .ZN(n11043) );
  NAND2_X1 U13530 ( .A1(n12365), .A2(n13592), .ZN(n11042) );
  NAND2_X1 U13531 ( .A1(n11043), .A2(n11042), .ZN(n11044) );
  XNOR2_X1 U13532 ( .A(n11044), .B(n12366), .ZN(n11247) );
  AOI22_X1 U13533 ( .A1(n11045), .A2(n12365), .B1(n12364), .B2(n13592), .ZN(
        n11248) );
  XNOR2_X1 U13534 ( .A(n11247), .B(n11248), .ZN(n11046) );
  OAI211_X1 U13535 ( .C1(n11047), .C2(n11046), .A(n11250), .B(n14139), .ZN(
        n11052) );
  OAI21_X1 U13536 ( .B1(n13513), .B2(n14355), .A(n11048), .ZN(n11049) );
  AOI21_X1 U13537 ( .B1(n11050), .B2(n13576), .A(n11049), .ZN(n11051) );
  OAI211_X1 U13538 ( .C1(n6881), .C2(n13579), .A(n11052), .B(n11051), .ZN(
        P1_U3213) );
  MUX2_X1 U13539 ( .A(n11058), .B(n11054), .S(n11053), .Z(n11056) );
  XNOR2_X1 U13540 ( .A(n11056), .B(n11055), .ZN(n11063) );
  NAND2_X1 U13541 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n14725) );
  OAI21_X1 U13542 ( .B1(n12518), .B2(n14815), .A(n14725), .ZN(n11060) );
  OAI22_X1 U13543 ( .A1(n11058), .A2(n12475), .B1(n11057), .B2(n12526), .ZN(
        n11059) );
  AOI211_X1 U13544 ( .C1(n11061), .C2(n12523), .A(n11060), .B(n11059), .ZN(
        n11062) );
  OAI21_X1 U13545 ( .B1(n11063), .B2(n12531), .A(n11062), .ZN(P3_U3161) );
  NAND2_X1 U13546 ( .A1(n11146), .A2(n13065), .ZN(n11064) );
  NAND2_X1 U13547 ( .A1(n11065), .A2(n11064), .ZN(n11125) );
  XNOR2_X1 U13548 ( .A(n11125), .B(n11068), .ZN(n14590) );
  INV_X1 U13549 ( .A(n14590), .ZN(n11081) );
  INV_X1 U13550 ( .A(n13065), .ZN(n11167) );
  OR2_X1 U13551 ( .A1(n11146), .A2(n11167), .ZN(n11066) );
  INV_X1 U13552 ( .A(n11068), .ZN(n11069) );
  NAND2_X1 U13553 ( .A1(n11070), .A2(n11069), .ZN(n11071) );
  NAND2_X1 U13554 ( .A1(n11131), .A2(n11071), .ZN(n11072) );
  NAND2_X1 U13555 ( .A1(n11072), .A2(n13284), .ZN(n11075) );
  NAND2_X1 U13556 ( .A1(n13037), .A2(n13063), .ZN(n11074) );
  NAND2_X1 U13557 ( .A1(n13038), .A2(n13065), .ZN(n11073) );
  AND2_X1 U13558 ( .A1(n11074), .A2(n11073), .ZN(n11175) );
  NAND2_X1 U13559 ( .A1(n11075), .A2(n11175), .ZN(n14596) );
  INV_X1 U13560 ( .A(n11174), .ZN(n14593) );
  NAND2_X1 U13561 ( .A1(n14593), .A2(n11076), .ZN(n11137) );
  OAI211_X1 U13562 ( .C1(n14593), .C2(n11076), .A(n13379), .B(n11137), .ZN(
        n14591) );
  OAI22_X1 U13563 ( .A1(n13257), .A2(n10421), .B1(n11179), .B2(n13245), .ZN(
        n11077) );
  AOI21_X1 U13564 ( .B1(n11174), .B2(n13241), .A(n11077), .ZN(n11078) );
  OAI21_X1 U13565 ( .B1(n14591), .B2(n13170), .A(n11078), .ZN(n11079) );
  AOI21_X1 U13566 ( .B1(n14596), .B2(n13257), .A(n11079), .ZN(n11080) );
  OAI21_X1 U13567 ( .B1(n11081), .B2(n13299), .A(n11080), .ZN(P2_U3254) );
  INV_X1 U13568 ( .A(n11146), .ZN(n11166) );
  INV_X1 U13569 ( .A(n11082), .ZN(n11163) );
  AOI22_X1 U13570 ( .A1(n13304), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11163), 
        .B2(n13291), .ZN(n11083) );
  OAI21_X1 U13571 ( .B1(n11166), .B2(n13294), .A(n11083), .ZN(n11086) );
  NOR2_X1 U13572 ( .A1(n11084), .A2(n13299), .ZN(n11085) );
  AOI211_X1 U13573 ( .C1(n11087), .C2(n13302), .A(n11086), .B(n11085), .ZN(
        n11088) );
  OAI21_X1 U13574 ( .B1(n13304), .B2(n11089), .A(n11088), .ZN(P2_U3255) );
  INV_X1 U13575 ( .A(n11090), .ZN(n11094) );
  INV_X1 U13576 ( .A(n11091), .ZN(n11092) );
  AOI22_X1 U13577 ( .A1(n13304), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n11092), 
        .B2(n13291), .ZN(n11093) );
  OAI21_X1 U13578 ( .B1(n11094), .B2(n13294), .A(n11093), .ZN(n11097) );
  NOR2_X1 U13579 ( .A1(n11095), .A2(n13299), .ZN(n11096) );
  AOI211_X1 U13580 ( .C1(n11098), .C2(n13302), .A(n11097), .B(n11096), .ZN(
        n11099) );
  OAI21_X1 U13581 ( .B1(n13304), .B2(n11100), .A(n11099), .ZN(P2_U3256) );
  NAND2_X1 U13582 ( .A1(n11101), .A2(n14038), .ZN(n11102) );
  OAI211_X1 U13583 ( .C1(n11103), .C2(n12874), .A(n11102), .B(n12313), .ZN(
        P3_U3272) );
  XNOR2_X1 U13584 ( .A(n11104), .B(n8395), .ZN(n11116) );
  INV_X1 U13585 ( .A(n11116), .ZN(n14822) );
  OR2_X1 U13586 ( .A1(n11106), .A2(n11105), .ZN(n11112) );
  OR2_X1 U13587 ( .A1(n11108), .A2(n11107), .ZN(n11110) );
  AND2_X1 U13588 ( .A1(n11110), .A2(n11109), .ZN(n11111) );
  NAND2_X1 U13589 ( .A1(n11112), .A2(n11111), .ZN(n11114) );
  XNOR2_X1 U13590 ( .A(n11114), .B(n11113), .ZN(n11118) );
  OAI22_X1 U13591 ( .A1(n12207), .A2(n14762), .B1(n11317), .B2(n14760), .ZN(
        n11115) );
  AOI21_X1 U13592 ( .B1(n11116), .B2(n14805), .A(n11115), .ZN(n11117) );
  OAI21_X1 U13593 ( .B1(n11118), .B2(n14767), .A(n11117), .ZN(n14824) );
  NAND2_X1 U13594 ( .A1(n14824), .A2(n14770), .ZN(n11123) );
  INV_X1 U13595 ( .A(n11119), .ZN(n11120) );
  OAI22_X1 U13596 ( .A1(n12757), .A2(n14820), .B1(n11120), .B2(n14755), .ZN(
        n11121) );
  AOI21_X1 U13597 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n14772), .A(n11121), .ZN(
        n11122) );
  OAI211_X1 U13598 ( .C1(n14822), .C2(n11124), .A(n11123), .B(n11122), .ZN(
        P3_U3224) );
  OAI21_X1 U13599 ( .B1(n11125), .B2(n13064), .A(n11174), .ZN(n11127) );
  NAND2_X1 U13600 ( .A1(n11125), .A2(n13064), .ZN(n11126) );
  NAND2_X1 U13601 ( .A1(n11127), .A2(n11126), .ZN(n11210) );
  XNOR2_X1 U13602 ( .A(n11210), .B(n11128), .ZN(n13405) );
  INV_X1 U13603 ( .A(n11128), .ZN(n11132) );
  INV_X1 U13604 ( .A(n13064), .ZN(n11129) );
  NAND2_X1 U13605 ( .A1(n11174), .A2(n11129), .ZN(n11133) );
  AND2_X1 U13606 ( .A1(n11132), .A2(n11133), .ZN(n11130) );
  NAND2_X1 U13607 ( .A1(n11212), .A2(n13284), .ZN(n11135) );
  AOI21_X1 U13608 ( .B1(n11131), .B2(n11133), .A(n11132), .ZN(n11134) );
  AOI22_X1 U13609 ( .A1(n13038), .A2(n13064), .B1(n13037), .B2(n13062), .ZN(
        n11278) );
  OAI21_X1 U13610 ( .B1(n11135), .B2(n11134), .A(n11278), .ZN(n13401) );
  NAND2_X1 U13611 ( .A1(n13401), .A2(n13257), .ZN(n11141) );
  AOI211_X1 U13612 ( .C1(n13403), .C2(n11137), .A(n13289), .B(n11136), .ZN(
        n13402) );
  NOR2_X1 U13613 ( .A1(n7020), .A2(n13294), .ZN(n11139) );
  OAI22_X1 U13614 ( .A1(n13257), .A2(n11453), .B1(n11281), .B2(n13245), .ZN(
        n11138) );
  AOI211_X1 U13615 ( .C1(n13402), .C2(n13302), .A(n11139), .B(n11138), .ZN(
        n11140) );
  OAI211_X1 U13616 ( .C1(n13405), .C2(n13299), .A(n11141), .B(n11140), .ZN(
        P2_U3253) );
  INV_X1 U13617 ( .A(n11142), .ZN(n12381) );
  INV_X1 U13618 ( .A(n11143), .ZN(n11144) );
  OAI222_X1 U13619 ( .A1(n12041), .A2(n11145), .B1(n13444), .B2(n12381), .C1(
        P2_U3088), .C2(n11144), .ZN(P2_U3306) );
  XNOR2_X1 U13620 ( .A(n12948), .B(n11146), .ZN(n11147) );
  AND2_X1 U13621 ( .A1(n12916), .A2(n13065), .ZN(n11148) );
  NAND2_X1 U13622 ( .A1(n11147), .A2(n11148), .ZN(n11171) );
  INV_X1 U13623 ( .A(n11147), .ZN(n11168) );
  INV_X1 U13624 ( .A(n11148), .ZN(n11149) );
  NAND2_X1 U13625 ( .A1(n11168), .A2(n11149), .ZN(n11150) );
  NAND2_X1 U13626 ( .A1(n11171), .A2(n11150), .ZN(n11159) );
  INV_X1 U13627 ( .A(n11151), .ZN(n11153) );
  NAND2_X1 U13628 ( .A1(n11153), .A2(n11152), .ZN(n11154) );
  NAND2_X1 U13629 ( .A1(n11155), .A2(n11154), .ZN(n11158) );
  INV_X1 U13630 ( .A(n11159), .ZN(n11156) );
  INV_X1 U13631 ( .A(n11173), .ZN(n11170) );
  AOI211_X1 U13632 ( .C1(n11159), .C2(n11158), .A(n13023), .B(n11170), .ZN(
        n11160) );
  INV_X1 U13633 ( .A(n11160), .ZN(n11165) );
  OAI22_X1 U13634 ( .A1(n13040), .A2(n11161), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14937), .ZN(n11162) );
  AOI21_X1 U13635 ( .B1(n11163), .B2(n13042), .A(n11162), .ZN(n11164) );
  OAI211_X1 U13636 ( .C1(n11166), .C2(n13045), .A(n11165), .B(n11164), .ZN(
        P2_U3189) );
  NOR3_X1 U13637 ( .A1(n11168), .A2(n11167), .A3(n11989), .ZN(n11169) );
  AOI21_X1 U13638 ( .B1(n11170), .B2(n13035), .A(n11169), .ZN(n11183) );
  XNOR2_X1 U13639 ( .A(n11174), .B(n12948), .ZN(n11282) );
  NAND2_X1 U13640 ( .A1(n12916), .A2(n13064), .ZN(n11276) );
  XNOR2_X1 U13641 ( .A(n11282), .B(n11276), .ZN(n11182) );
  NAND2_X1 U13642 ( .A1(n11174), .A2(n6418), .ZN(n11178) );
  INV_X1 U13643 ( .A(n11175), .ZN(n11176) );
  AOI22_X1 U13644 ( .A1(n12999), .A2(n11176), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11177) );
  OAI211_X1 U13645 ( .C1(n13015), .C2(n11179), .A(n11178), .B(n11177), .ZN(
        n11180) );
  AOI21_X1 U13646 ( .B1(n6576), .B2(n13035), .A(n11180), .ZN(n11181) );
  OAI21_X1 U13647 ( .B1(n11183), .B2(n11182), .A(n11181), .ZN(P2_U3208) );
  NOR2_X1 U13648 ( .A1(n11185), .A2(n11186), .ZN(n11187) );
  NAND2_X1 U13649 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n11469), .ZN(n11188) );
  OAI21_X1 U13650 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n11469), .A(n11188), 
        .ZN(n11189) );
  AOI21_X1 U13651 ( .B1(n6579), .B2(n11189), .A(n11467), .ZN(n11209) );
  MUX2_X1 U13652 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12073), .Z(n11192) );
  XNOR2_X1 U13653 ( .A(n11192), .B(n11302), .ZN(n11304) );
  NOR2_X1 U13654 ( .A1(n11192), .A2(n11302), .ZN(n11194) );
  MUX2_X1 U13655 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12073), .Z(n11475) );
  XNOR2_X1 U13656 ( .A(n11475), .B(n11469), .ZN(n11193) );
  NOR3_X1 U13657 ( .A1(n11303), .A2(n11194), .A3(n11193), .ZN(n11480) );
  INV_X1 U13658 ( .A(n11480), .ZN(n11196) );
  OAI21_X1 U13659 ( .B1(n11303), .B2(n11194), .A(n11193), .ZN(n11195) );
  NAND3_X1 U13660 ( .A1(n11196), .A2(n14735), .A3(n11195), .ZN(n11208) );
  INV_X1 U13661 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14104) );
  AOI22_X1 U13662 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n11469), .B1(n11476), 
        .B2(n14104), .ZN(n11202) );
  NAND2_X1 U13663 ( .A1(n11302), .A2(n11199), .ZN(n11200) );
  NAND2_X1 U13664 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n11299), .ZN(n11298) );
  OAI21_X1 U13665 ( .B1(n11202), .B2(n11201), .A(n11470), .ZN(n11206) );
  NAND2_X1 U13666 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P3_U3151), .ZN(n11382)
         );
  INV_X1 U13667 ( .A(n11382), .ZN(n11203) );
  AOI21_X1 U13668 ( .B1(n14743), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11203), 
        .ZN(n11204) );
  OAI21_X1 U13669 ( .B1(n14740), .B2(n11469), .A(n11204), .ZN(n11205) );
  AOI21_X1 U13670 ( .B1(n11206), .B2(n14746), .A(n11205), .ZN(n11207) );
  OAI211_X1 U13671 ( .C1(n11209), .C2(n14750), .A(n11208), .B(n11207), .ZN(
        P3_U3194) );
  XNOR2_X1 U13672 ( .A(n11435), .B(n11213), .ZN(n13400) );
  NAND2_X1 U13673 ( .A1(n11212), .A2(n11211), .ZN(n11214) );
  OAI211_X1 U13674 ( .C1(n11214), .C2(n11213), .A(n11428), .B(n13284), .ZN(
        n11215) );
  AOI22_X1 U13675 ( .A1(n13038), .A2(n13063), .B1(n13037), .B2(n13061), .ZN(
        n11526) );
  NAND2_X1 U13676 ( .A1(n11215), .A2(n11526), .ZN(n13396) );
  NAND2_X1 U13677 ( .A1(n13396), .A2(n13257), .ZN(n11221) );
  INV_X1 U13678 ( .A(n11432), .ZN(n11216) );
  AOI211_X1 U13679 ( .C1(n13398), .C2(n11217), .A(n13289), .B(n11216), .ZN(
        n13397) );
  NOR2_X1 U13680 ( .A1(n6931), .A2(n13294), .ZN(n11219) );
  INV_X1 U13681 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11455) );
  OAI22_X1 U13682 ( .A1(n13257), .A2(n11455), .B1(n11524), .B2(n13245), .ZN(
        n11218) );
  AOI211_X1 U13683 ( .C1(n13397), .C2(n13302), .A(n11219), .B(n11218), .ZN(
        n11220) );
  OAI211_X1 U13684 ( .C1(n13400), .C2(n13299), .A(n11221), .B(n11220), .ZN(
        P2_U3252) );
  NAND2_X1 U13685 ( .A1(n11223), .A2(n11222), .ZN(n11225) );
  NAND2_X1 U13686 ( .A1(n11426), .A2(n11577), .ZN(n11224) );
  NAND2_X1 U13687 ( .A1(n11225), .A2(n11224), .ZN(n14288) );
  NAND2_X1 U13688 ( .A1(n14288), .A2(n14289), .ZN(n11227) );
  OR2_X1 U13689 ( .A1(n14287), .A2(n14130), .ZN(n11226) );
  OR2_X1 U13690 ( .A1(n14172), .A2(n14291), .ZN(n11228) );
  XNOR2_X1 U13691 ( .A(n11263), .B(n11261), .ZN(n11238) );
  AOI22_X1 U13692 ( .A1(n14292), .A2(n13589), .B1(n14131), .B2(n14291), .ZN(
        n11237) );
  OR2_X1 U13693 ( .A1(n11426), .A2(n13590), .ZN(n11229) );
  INV_X1 U13694 ( .A(n14289), .ZN(n11231) );
  INV_X1 U13695 ( .A(n14171), .ZN(n11233) );
  NAND2_X1 U13696 ( .A1(n14164), .A2(n11233), .ZN(n14167) );
  OR2_X1 U13697 ( .A1(n14172), .A2(n11792), .ZN(n11234) );
  NAND2_X1 U13698 ( .A1(n14167), .A2(n11234), .ZN(n11235) );
  OAI211_X1 U13699 ( .C1(n11235), .C2(n11261), .A(n11266), .B(n14353), .ZN(
        n11236) );
  OAI211_X1 U13700 ( .C1(n11238), .C2(n14349), .A(n11237), .B(n11236), .ZN(
        n11365) );
  NAND2_X1 U13701 ( .A1(n11787), .A2(n14174), .ZN(n11239) );
  NAND2_X1 U13702 ( .A1(n11239), .A2(n14310), .ZN(n11240) );
  OR2_X1 U13703 ( .A1(n11327), .A2(n11240), .ZN(n11366) );
  AOI22_X1 U13704 ( .A1(n14284), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n11795), 
        .B2(n14285), .ZN(n11242) );
  NAND2_X1 U13705 ( .A1(n11787), .A2(n14306), .ZN(n11241) );
  OAI211_X1 U13706 ( .C1(n11366), .C2(n14160), .A(n11242), .B(n11241), .ZN(
        n11243) );
  AOI21_X1 U13707 ( .B1(n11365), .B2(n14303), .A(n11243), .ZN(n11244) );
  INV_X1 U13708 ( .A(n11244), .ZN(P1_U3281) );
  OAI22_X1 U13709 ( .A1(n14364), .A2(n11942), .B1(n11246), .B2(n11941), .ZN(
        n11245) );
  XNOR2_X1 U13710 ( .A(n11245), .B(n12366), .ZN(n11412) );
  OAI22_X1 U13711 ( .A1(n14364), .A2(n11941), .B1(n11246), .B2(n11940), .ZN(
        n11413) );
  XNOR2_X1 U13712 ( .A(n11412), .B(n11413), .ZN(n11252) );
  INV_X1 U13713 ( .A(n11247), .ZN(n11249) );
  AOI21_X1 U13714 ( .B1(n11252), .B2(n11251), .A(n11416), .ZN(n11260) );
  NAND2_X1 U13715 ( .A1(n13576), .A2(n11253), .ZN(n11255) );
  OAI211_X1 U13716 ( .C1(n11256), .C2(n13513), .A(n11255), .B(n11254), .ZN(
        n11257) );
  AOI21_X1 U13717 ( .B1(n11258), .B2(n14142), .A(n11257), .ZN(n11259) );
  OAI21_X1 U13718 ( .B1(n11260), .B2(n13564), .A(n11259), .ZN(P1_U3221) );
  INV_X1 U13719 ( .A(n11261), .ZN(n11262) );
  XNOR2_X1 U13720 ( .A(n11338), .B(n11336), .ZN(n14217) );
  INV_X1 U13721 ( .A(n14129), .ZN(n11264) );
  OR2_X1 U13722 ( .A1(n11787), .A2(n11264), .ZN(n11265) );
  NAND2_X1 U13723 ( .A1(n11266), .A2(n11265), .ZN(n11267) );
  NAND2_X1 U13724 ( .A1(n11267), .A2(n11336), .ZN(n11326) );
  OAI211_X1 U13725 ( .C1(n11267), .C2(n11336), .A(n11326), .B(n14353), .ZN(
        n11269) );
  AOI22_X1 U13726 ( .A1(n14292), .A2(n13588), .B1(n14131), .B2(n14129), .ZN(
        n11268) );
  NAND2_X1 U13727 ( .A1(n11269), .A2(n11268), .ZN(n14222) );
  XNOR2_X1 U13728 ( .A(n11327), .B(n11832), .ZN(n11270) );
  NAND2_X1 U13729 ( .A1(n11270), .A2(n14310), .ZN(n14218) );
  INV_X1 U13730 ( .A(n11838), .ZN(n11271) );
  OAI22_X1 U13731 ( .A1(n14218), .A2(n11272), .B1(n14302), .B2(n11271), .ZN(
        n11273) );
  OAI21_X1 U13732 ( .B1(n14222), .B2(n11273), .A(n14303), .ZN(n11275) );
  AOI22_X1 U13733 ( .A1(n11832), .A2(n14306), .B1(n13880), .B2(
        P1_REG2_REG_13__SCAN_IN), .ZN(n11274) );
  OAI211_X1 U13734 ( .C1(n13887), .C2(n14217), .A(n11275), .B(n11274), .ZN(
        P1_U3280) );
  INV_X1 U13735 ( .A(n11282), .ZN(n11277) );
  XNOR2_X1 U13736 ( .A(n13403), .B(n12948), .ZN(n11516) );
  NAND2_X1 U13737 ( .A1(n12916), .A2(n13063), .ZN(n11517) );
  XNOR2_X1 U13738 ( .A(n11516), .B(n11517), .ZN(n11283) );
  INV_X1 U13739 ( .A(n11278), .ZN(n11279) );
  AOI22_X1 U13740 ( .A1(n12999), .A2(n11279), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11280) );
  OAI21_X1 U13741 ( .B1(n13015), .B2(n11281), .A(n11280), .ZN(n11286) );
  AOI22_X1 U13742 ( .A1(n11282), .A2(n13035), .B1(n13013), .B2(n13064), .ZN(
        n11284) );
  NOR3_X1 U13743 ( .A1(n6576), .A2(n11284), .A3(n11283), .ZN(n11285) );
  AOI211_X1 U13744 ( .C1(n13403), .C2(n6418), .A(n11286), .B(n11285), .ZN(
        n11287) );
  OAI21_X1 U13745 ( .B1(n11520), .B2(n13023), .A(n11287), .ZN(P2_U3196) );
  INV_X1 U13746 ( .A(n12226), .ZN(n11288) );
  XNOR2_X1 U13747 ( .A(n11289), .B(n11288), .ZN(n11291) );
  OAI22_X1 U13748 ( .A1(n11317), .A2(n14762), .B1(n11503), .B2(n14760), .ZN(
        n11290) );
  AOI21_X1 U13749 ( .B1(n11291), .B2(n12768), .A(n11290), .ZN(n14109) );
  XNOR2_X1 U13750 ( .A(n11292), .B(n12226), .ZN(n14107) );
  AOI22_X1 U13751 ( .A1(n14772), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n12755), 
        .B2(n11321), .ZN(n11293) );
  OAI21_X1 U13752 ( .B1(n11324), .B2(n12757), .A(n11293), .ZN(n11294) );
  AOI21_X1 U13753 ( .B1(n14107), .B2(n12778), .A(n11294), .ZN(n11295) );
  OAI21_X1 U13754 ( .B1(n14109), .B2(n14772), .A(n11295), .ZN(P3_U3222) );
  AOI21_X1 U13755 ( .B1(n8417), .B2(n11297), .A(n11296), .ZN(n11311) );
  OAI21_X1 U13756 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n11299), .A(n11298), 
        .ZN(n11309) );
  INV_X1 U13757 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11318) );
  NOR2_X1 U13758 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11318), .ZN(n11300) );
  AOI21_X1 U13759 ( .B1(n14743), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11300), 
        .ZN(n11301) );
  OAI21_X1 U13760 ( .B1(n14740), .B2(n11302), .A(n11301), .ZN(n11308) );
  AOI21_X1 U13761 ( .B1(n11305), .B2(n11304), .A(n11303), .ZN(n11306) );
  NOR2_X1 U13762 ( .A1(n11306), .A2(n14709), .ZN(n11307) );
  AOI211_X1 U13763 ( .C1(n14746), .C2(n11309), .A(n11308), .B(n11307), .ZN(
        n11310) );
  OAI21_X1 U13764 ( .B1(n11311), .B2(n14750), .A(n11310), .ZN(P3_U3193) );
  NAND2_X1 U13765 ( .A1(n12549), .A2(n11312), .ZN(n11313) );
  XNOR2_X1 U13766 ( .A(n14105), .B(n6420), .ZN(n11375) );
  XOR2_X1 U13767 ( .A(n11376), .B(n11375), .Z(n11377) );
  XNOR2_X1 U13768 ( .A(n11377), .B(n11315), .ZN(n11316) );
  NAND2_X1 U13769 ( .A1(n11316), .A2(n12509), .ZN(n11323) );
  NOR2_X1 U13770 ( .A1(n11317), .A2(n12475), .ZN(n11320) );
  OAI22_X1 U13771 ( .A1(n11503), .A2(n12526), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11318), .ZN(n11319) );
  AOI211_X1 U13772 ( .C1(n11321), .C2(n12523), .A(n11320), .B(n11319), .ZN(
        n11322) );
  OAI211_X1 U13773 ( .C1(n12518), .C2(n11324), .A(n11323), .B(n11322), .ZN(
        P3_U3176) );
  INV_X1 U13774 ( .A(n13589), .ZN(n11791) );
  OR2_X1 U13775 ( .A1(n11832), .A2(n11791), .ZN(n11325) );
  NAND2_X1 U13776 ( .A1(n11326), .A2(n11325), .ZN(n11539) );
  XNOR2_X1 U13777 ( .A(n11539), .B(n11341), .ZN(n14214) );
  INV_X1 U13778 ( .A(n11832), .ZN(n14219) );
  AOI211_X1 U13779 ( .C1(n14210), .C2(n11328), .A(n14182), .B(n6892), .ZN(
        n14208) );
  INV_X1 U13780 ( .A(n14210), .ZN(n11334) );
  NAND2_X1 U13781 ( .A1(n14292), .A2(n13587), .ZN(n11330) );
  NAND2_X1 U13782 ( .A1(n14131), .A2(n13589), .ZN(n11329) );
  NAND2_X1 U13783 ( .A1(n11330), .A2(n11329), .ZN(n14209) );
  AOI22_X1 U13784 ( .A1(n14303), .A2(n14209), .B1(n11331), .B2(n14285), .ZN(
        n11333) );
  NAND2_X1 U13785 ( .A1(n14284), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11332) );
  OAI211_X1 U13786 ( .C1(n11334), .C2(n13883), .A(n11333), .B(n11332), .ZN(
        n11335) );
  AOI21_X1 U13787 ( .B1(n14208), .B2(n14314), .A(n11335), .ZN(n11344) );
  INV_X1 U13788 ( .A(n11336), .ZN(n11337) );
  NAND2_X1 U13789 ( .A1(n11338), .A2(n11337), .ZN(n11340) );
  OR2_X1 U13790 ( .A1(n11832), .A2(n13589), .ZN(n11339) );
  NAND2_X1 U13791 ( .A1(n11342), .A2(n11341), .ZN(n14211) );
  NAND3_X1 U13792 ( .A1(n11546), .A2(n14211), .A3(n14315), .ZN(n11343) );
  OAI211_X1 U13793 ( .C1(n14214), .C2(n13868), .A(n11344), .B(n11343), .ZN(
        P1_U3279) );
  XNOR2_X1 U13794 ( .A(n11345), .B(n11346), .ZN(n14101) );
  XNOR2_X1 U13795 ( .A(n6600), .B(n11346), .ZN(n11348) );
  AND2_X1 U13796 ( .A1(n12546), .A2(n12765), .ZN(n11347) );
  AOI21_X1 U13797 ( .B1(n12548), .B2(n12763), .A(n11347), .ZN(n11383) );
  OAI21_X1 U13798 ( .B1(n11348), .B2(n14767), .A(n11383), .ZN(n14103) );
  NAND2_X1 U13799 ( .A1(n14103), .A2(n14770), .ZN(n11353) );
  INV_X1 U13800 ( .A(n11380), .ZN(n11349) );
  OAI22_X1 U13801 ( .A1(n14770), .A2(n11350), .B1(n11349), .B2(n14755), .ZN(
        n11351) );
  AOI21_X1 U13802 ( .B1(n12773), .B2(n11385), .A(n11351), .ZN(n11352) );
  OAI211_X1 U13803 ( .C1(n12663), .C2(n14101), .A(n11353), .B(n11352), .ZN(
        P3_U3221) );
  XNOR2_X1 U13804 ( .A(n11385), .B(n12444), .ZN(n11356) );
  NOR2_X1 U13805 ( .A1(n11356), .A2(n11503), .ZN(n11373) );
  INV_X1 U13806 ( .A(n11373), .ZN(n11355) );
  NAND2_X1 U13807 ( .A1(n12548), .A2(n11375), .ZN(n11354) );
  INV_X1 U13808 ( .A(n11356), .ZN(n11357) );
  NOR2_X1 U13809 ( .A1(n11357), .A2(n12547), .ZN(n11374) );
  XNOR2_X1 U13810 ( .A(n14095), .B(n12444), .ZN(n11557) );
  XNOR2_X1 U13811 ( .A(n11557), .B(n11560), .ZN(n11359) );
  XNOR2_X1 U13812 ( .A(n11558), .B(n11359), .ZN(n11364) );
  INV_X1 U13813 ( .A(n14095), .ZN(n11509) );
  AOI22_X1 U13814 ( .A1(n12547), .A2(n12522), .B1(P3_REG3_REG_13__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11361) );
  NAND2_X1 U13815 ( .A1(n12523), .A2(n11506), .ZN(n11360) );
  OAI211_X1 U13816 ( .C1(n11672), .C2(n12526), .A(n11361), .B(n11360), .ZN(
        n11362) );
  AOI21_X1 U13817 ( .B1(n11509), .B2(n12528), .A(n11362), .ZN(n11363) );
  OAI21_X1 U13818 ( .B1(n11364), .B2(n12531), .A(n11363), .ZN(P3_U3174) );
  INV_X1 U13819 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11369) );
  INV_X1 U13820 ( .A(n11787), .ZN(n11798) );
  INV_X1 U13821 ( .A(n11365), .ZN(n11367) );
  OAI211_X1 U13822 ( .C1(n11798), .C2(n14371), .A(n11367), .B(n11366), .ZN(
        n11370) );
  NAND2_X1 U13823 ( .A1(n11370), .A2(n14378), .ZN(n11368) );
  OAI21_X1 U13824 ( .B1(n14378), .B2(n11369), .A(n11368), .ZN(P1_U3495) );
  NAND2_X1 U13825 ( .A1(n11370), .A2(n14391), .ZN(n11371) );
  OAI21_X1 U13826 ( .B1(n14391), .B2(n11372), .A(n11371), .ZN(P1_U3540) );
  NOR2_X1 U13827 ( .A1(n11374), .A2(n11373), .ZN(n11379) );
  AOI22_X1 U13828 ( .A1(n11377), .A2(n12548), .B1(n11376), .B2(n11375), .ZN(
        n11378) );
  XOR2_X1 U13829 ( .A(n11379), .B(n11378), .Z(n11387) );
  NAND2_X1 U13830 ( .A1(n12523), .A2(n11380), .ZN(n11381) );
  OAI211_X1 U13831 ( .C1(n11383), .C2(n12503), .A(n11382), .B(n11381), .ZN(
        n11384) );
  AOI21_X1 U13832 ( .B1(n12528), .B2(n11385), .A(n11384), .ZN(n11386) );
  OAI21_X1 U13833 ( .B1(n11387), .B2(n12531), .A(n11386), .ZN(P3_U3164) );
  INV_X1 U13834 ( .A(n11388), .ZN(n11390) );
  INV_X1 U13835 ( .A(n9866), .ZN(n11389) );
  OAI222_X1 U13836 ( .A1(n12041), .A2(n11391), .B1(n13444), .B2(n11390), .C1(
        P2_U3088), .C2(n11389), .ZN(P2_U3305) );
  NAND2_X1 U13837 ( .A1(n11392), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11394) );
  NAND2_X1 U13838 ( .A1(n11394), .A2(n11393), .ZN(n11395) );
  NOR2_X1 U13839 ( .A1(n11402), .A2(n11395), .ZN(n11396) );
  XOR2_X1 U13840 ( .A(n11395), .B(n14273), .Z(n14268) );
  NOR2_X1 U13841 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14268), .ZN(n14267) );
  NOR2_X1 U13842 ( .A1(n11396), .A2(n14267), .ZN(n11399) );
  INV_X1 U13843 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11663) );
  NOR2_X1 U13844 ( .A1(n11591), .A2(n11663), .ZN(n11397) );
  AOI21_X1 U13845 ( .B1(n11663), .B2(n11591), .A(n11397), .ZN(n11398) );
  NAND2_X1 U13846 ( .A1(n11398), .A2(n11399), .ZN(n11585) );
  OAI211_X1 U13847 ( .C1(n11399), .C2(n11398), .A(n13725), .B(n11585), .ZN(
        n11411) );
  NAND2_X1 U13848 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13501)
         );
  NOR2_X1 U13849 ( .A1(n11402), .A2(n11403), .ZN(n11404) );
  XOR2_X1 U13850 ( .A(n14273), .B(n11403), .Z(n14266) );
  NOR2_X1 U13851 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14266), .ZN(n14265) );
  INV_X1 U13852 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14201) );
  NOR2_X1 U13853 ( .A1(n11591), .A2(n14201), .ZN(n11405) );
  AOI21_X1 U13854 ( .B1(n14201), .B2(n11591), .A(n11405), .ZN(n11406) );
  NAND2_X1 U13855 ( .A1(n11406), .A2(n11407), .ZN(n11590) );
  OAI211_X1 U13856 ( .C1(n11407), .C2(n11406), .A(n13726), .B(n11590), .ZN(
        n11408) );
  NAND2_X1 U13857 ( .A1(n13501), .A2(n11408), .ZN(n11409) );
  AOI21_X1 U13858 ( .B1(n13708), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11409), 
        .ZN(n11410) );
  OAI211_X1 U13859 ( .C1(n14274), .C2(n11591), .A(n11411), .B(n11410), .ZN(
        P1_U3259) );
  INV_X1 U13860 ( .A(n11412), .ZN(n11415) );
  INV_X1 U13861 ( .A(n11413), .ZN(n11414) );
  OAI22_X1 U13862 ( .A1(n11426), .A2(n11941), .B1(n11577), .B2(n11940), .ZN(
        n11569) );
  OAI22_X1 U13863 ( .A1(n11426), .A2(n11942), .B1(n11577), .B2(n11941), .ZN(
        n11417) );
  XNOR2_X1 U13864 ( .A(n11417), .B(n12366), .ZN(n11570) );
  XOR2_X1 U13865 ( .A(n11569), .B(n11570), .Z(n11418) );
  OAI211_X1 U13866 ( .C1(n11419), .C2(n11418), .A(n11571), .B(n14139), .ZN(
        n11425) );
  NAND2_X1 U13867 ( .A1(n13557), .A2(n13591), .ZN(n11421) );
  OAI211_X1 U13868 ( .C1(n11572), .C2(n13570), .A(n11421), .B(n11420), .ZN(
        n11422) );
  AOI21_X1 U13869 ( .B1(n11423), .B2(n13576), .A(n11422), .ZN(n11424) );
  OAI211_X1 U13870 ( .C1(n11426), .C2(n13579), .A(n11425), .B(n11424), .ZN(
        P1_U3231) );
  INV_X1 U13871 ( .A(n13062), .ZN(n11990) );
  XOR2_X1 U13872 ( .A(n11723), .B(n11436), .Z(n11431) );
  NAND2_X1 U13873 ( .A1(n13037), .A2(n13060), .ZN(n11430) );
  NAND2_X1 U13874 ( .A1(n13038), .A2(n13062), .ZN(n11429) );
  NAND2_X1 U13875 ( .A1(n11430), .A2(n11429), .ZN(n11985) );
  AOI21_X1 U13876 ( .B1(n11431), .B2(n13284), .A(n11985), .ZN(n13394) );
  INV_X1 U13877 ( .A(n11714), .ZN(n11712) );
  AOI211_X1 U13878 ( .C1(n13392), .C2(n11432), .A(n13289), .B(n11714), .ZN(
        n13391) );
  INV_X1 U13879 ( .A(n13392), .ZN(n11721) );
  AOI22_X1 U13880 ( .A1(n13304), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11984), 
        .B2(n13291), .ZN(n11433) );
  OAI21_X1 U13881 ( .B1(n11721), .B2(n13294), .A(n11433), .ZN(n11438) );
  NOR2_X1 U13882 ( .A1(n13398), .A2(n13062), .ZN(n11434) );
  XOR2_X1 U13883 ( .A(n11709), .B(n11436), .Z(n13395) );
  NOR2_X1 U13884 ( .A1(n13395), .A2(n13299), .ZN(n11437) );
  AOI211_X1 U13885 ( .C1(n13391), .C2(n13302), .A(n11438), .B(n11437), .ZN(
        n11439) );
  OAI21_X1 U13886 ( .B1(n13304), .B2(n13394), .A(n11439), .ZN(P2_U3251) );
  NAND2_X1 U13887 ( .A1(n11444), .A2(n13436), .ZN(n11441) );
  OAI211_X1 U13888 ( .C1(n11442), .C2(n12041), .A(n11441), .B(n11440), .ZN(
        P2_U3304) );
  NAND2_X1 U13889 ( .A1(n11444), .A2(n11443), .ZN(n11446) );
  OAI211_X1 U13890 ( .C1(n14852), .C2(n14012), .A(n11446), .B(n11445), .ZN(
        P1_U3332) );
  NAND2_X1 U13891 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n11987)
         );
  XNOR2_X1 U13892 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n11742), .ZN(n11451) );
  INV_X1 U13893 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11449) );
  INV_X1 U13894 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11448) );
  INV_X1 U13895 ( .A(n11447), .ZN(n14481) );
  XNOR2_X1 U13896 ( .A(n14494), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n14480) );
  NOR3_X1 U13897 ( .A1(n14482), .A2(n14481), .A3(n14480), .ZN(n14479) );
  AOI21_X1 U13898 ( .B1(n11454), .B2(n11448), .A(n14479), .ZN(n14507) );
  XNOR2_X1 U13899 ( .A(n14510), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n14506) );
  NAND2_X1 U13900 ( .A1(n14507), .A2(n14506), .ZN(n14505) );
  OAI21_X1 U13901 ( .B1(n14510), .B2(n11449), .A(n14505), .ZN(n11450) );
  NAND2_X1 U13902 ( .A1(n11451), .A2(n11450), .ZN(n11740) );
  OAI211_X1 U13903 ( .C1(n11451), .C2(n11450), .A(n14542), .B(n11740), .ZN(
        n11452) );
  NAND2_X1 U13904 ( .A1(n11987), .A2(n11452), .ZN(n11460) );
  MUX2_X1 U13905 ( .A(n11453), .B(P2_REG2_REG_12__SCAN_IN), .S(n14494), .Z(
        n14488) );
  AOI21_X1 U13906 ( .B1(n11454), .B2(n11453), .A(n14486), .ZN(n14501) );
  NOR2_X1 U13907 ( .A1(n14510), .A2(n11455), .ZN(n11456) );
  AOI21_X1 U13908 ( .B1(n11455), .B2(n14510), .A(n11456), .ZN(n14500) );
  NAND2_X1 U13909 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n11457), .ZN(n11732) );
  OAI211_X1 U13910 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n11457), .A(n14526), 
        .B(n11732), .ZN(n11458) );
  INV_X1 U13911 ( .A(n11458), .ZN(n11459) );
  AOI211_X1 U13912 ( .C1(P2_ADDR_REG_14__SCAN_IN), .C2(n14540), .A(n11460), 
        .B(n11459), .ZN(n11461) );
  OAI21_X1 U13913 ( .B1(n11742), .B2(n14547), .A(n11461), .ZN(P2_U3228) );
  OAI22_X1 U13914 ( .A1(n11463), .A2(P3_U3151), .B1(n11462), .B2(n12874), .ZN(
        n11464) );
  AOI21_X1 U13915 ( .B1(n11465), .B2(n14038), .A(n11464), .ZN(n11466) );
  INV_X1 U13916 ( .A(n11466), .ZN(P3_U3271) );
  AOI21_X1 U13917 ( .B1(n8452), .B2(n11468), .A(n11627), .ZN(n11487) );
  NAND2_X1 U13918 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n11469), .ZN(n11471) );
  NAND2_X1 U13919 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n11472), .ZN(n11631) );
  OAI21_X1 U13920 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n11472), .A(n11631), 
        .ZN(n11485) );
  INV_X1 U13921 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n14911) );
  NOR2_X1 U13922 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14911), .ZN(n11473) );
  AOI21_X1 U13923 ( .B1(n14743), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n11473), 
        .ZN(n11474) );
  OAI21_X1 U13924 ( .B1(n14740), .B2(n11640), .A(n11474), .ZN(n11484) );
  INV_X1 U13925 ( .A(n11475), .ZN(n11477) );
  NOR2_X1 U13926 ( .A1(n11477), .A2(n11476), .ZN(n11479) );
  MUX2_X1 U13927 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12073), .Z(n11641) );
  XNOR2_X1 U13928 ( .A(n11641), .B(n11640), .ZN(n11478) );
  INV_X1 U13929 ( .A(n11643), .ZN(n11482) );
  OAI21_X1 U13930 ( .B1(n11480), .B2(n11479), .A(n11478), .ZN(n11481) );
  AOI21_X1 U13931 ( .B1(n11482), .B2(n11481), .A(n14709), .ZN(n11483) );
  AOI211_X1 U13932 ( .C1(n11485), .C2(n14746), .A(n11484), .B(n11483), .ZN(
        n11486) );
  OAI21_X1 U13933 ( .B1(n11487), .B2(n14750), .A(n11486), .ZN(P3_U3195) );
  OR3_X1 U13934 ( .A1(n6588), .A2(n11488), .A3(n12234), .ZN(n11489) );
  NAND3_X1 U13935 ( .A1(n11490), .A2(n12768), .A3(n11489), .ZN(n11491) );
  AOI22_X1 U13936 ( .A1(n11683), .A2(n12765), .B1(n12763), .B2(n12546), .ZN(
        n11564) );
  NAND2_X1 U13937 ( .A1(n11491), .A2(n11564), .ZN(n11617) );
  INV_X1 U13938 ( .A(n11617), .ZN(n11499) );
  NAND2_X1 U13939 ( .A1(n11345), .A2(n11492), .ZN(n11494) );
  AND2_X1 U13940 ( .A1(n11494), .A2(n11493), .ZN(n11495) );
  XNOR2_X1 U13941 ( .A(n11495), .B(n12234), .ZN(n11618) );
  AOI22_X1 U13942 ( .A1(n14772), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n12755), 
        .B2(n11566), .ZN(n11496) );
  OAI21_X1 U13943 ( .B1(n11624), .B2(n12757), .A(n11496), .ZN(n11497) );
  AOI21_X1 U13944 ( .B1(n11618), .B2(n12778), .A(n11497), .ZN(n11498) );
  OAI21_X1 U13945 ( .B1(n11499), .B2(n14772), .A(n11498), .ZN(P3_U3219) );
  NAND2_X1 U13946 ( .A1(n11345), .A2(n12124), .ZN(n11500) );
  NAND2_X1 U13947 ( .A1(n11500), .A2(n12233), .ZN(n11501) );
  XOR2_X1 U13948 ( .A(n12232), .B(n11501), .Z(n14096) );
  AOI211_X1 U13949 ( .C1(n12232), .C2(n11502), .A(n14767), .B(n6588), .ZN(
        n11505) );
  OAI22_X1 U13950 ( .A1(n11672), .A2(n14760), .B1(n11503), .B2(n14762), .ZN(
        n11504) );
  OR2_X1 U13951 ( .A1(n11505), .A2(n11504), .ZN(n14098) );
  NAND2_X1 U13952 ( .A1(n14098), .A2(n14770), .ZN(n11511) );
  INV_X1 U13953 ( .A(n11506), .ZN(n11507) );
  OAI22_X1 U13954 ( .A1(n14770), .A2(n8452), .B1(n11507), .B2(n14755), .ZN(
        n11508) );
  AOI21_X1 U13955 ( .B1(n11509), .B2(n12773), .A(n11508), .ZN(n11510) );
  OAI211_X1 U13956 ( .C1(n14096), .C2(n12663), .A(n11511), .B(n11510), .ZN(
        P3_U3220) );
  XNOR2_X1 U13957 ( .A(n13398), .B(n12948), .ZN(n11512) );
  AND2_X1 U13958 ( .A1(n12916), .A2(n13062), .ZN(n11513) );
  NAND2_X1 U13959 ( .A1(n11512), .A2(n11513), .ZN(n11694) );
  INV_X1 U13960 ( .A(n11512), .ZN(n11991) );
  INV_X1 U13961 ( .A(n11513), .ZN(n11514) );
  NAND2_X1 U13962 ( .A1(n11991), .A2(n11514), .ZN(n11515) );
  NAND2_X1 U13963 ( .A1(n11694), .A2(n11515), .ZN(n11522) );
  INV_X1 U13964 ( .A(n11516), .ZN(n11518) );
  NAND2_X1 U13965 ( .A1(n11518), .A2(n11517), .ZN(n11519) );
  INV_X1 U13966 ( .A(n11695), .ZN(n11993) );
  AOI211_X1 U13967 ( .C1(n11522), .C2(n11521), .A(n13023), .B(n11993), .ZN(
        n11523) );
  INV_X1 U13968 ( .A(n11523), .ZN(n11530) );
  INV_X1 U13969 ( .A(n11524), .ZN(n11528) );
  OAI22_X1 U13970 ( .A1(n13040), .A2(n11526), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11525), .ZN(n11527) );
  AOI21_X1 U13971 ( .B1(n11528), .B2(n13042), .A(n11527), .ZN(n11529) );
  OAI211_X1 U13972 ( .C1(n6931), .C2(n13045), .A(n11530), .B(n11529), .ZN(
        P2_U3206) );
  INV_X1 U13973 ( .A(n11531), .ZN(n11536) );
  INV_X1 U13974 ( .A(n11532), .ZN(n11533) );
  OAI222_X1 U13975 ( .A1(n12041), .A2(n14948), .B1(n13444), .B2(n11536), .C1(
        P2_U3088), .C2(n11533), .ZN(P2_U3303) );
  INV_X1 U13976 ( .A(n11534), .ZN(n11535) );
  OAI222_X1 U13977 ( .A1(n14012), .A2(n11537), .B1(n14014), .B2(n11536), .C1(
        n11535), .C2(P1_U3086), .ZN(P1_U3331) );
  NAND2_X1 U13978 ( .A1(n11539), .A2(n11538), .ZN(n11541) );
  XNOR2_X1 U13979 ( .A(n11655), .B(n11547), .ZN(n11542) );
  NAND2_X1 U13980 ( .A1(n11542), .A2(n14353), .ZN(n11544) );
  AOI22_X1 U13981 ( .A1(n14292), .A2(n13586), .B1(n14131), .B2(n13588), .ZN(
        n11543) );
  NAND2_X1 U13982 ( .A1(n11544), .A2(n11543), .ZN(n14206) );
  INV_X1 U13983 ( .A(n14206), .ZN(n11556) );
  NAND2_X1 U13984 ( .A1(n14210), .A2(n13588), .ZN(n11545) );
  INV_X1 U13985 ( .A(n11547), .ZN(n11654) );
  NAND2_X1 U13986 ( .A1(n11548), .A2(n11654), .ZN(n11549) );
  NAND2_X1 U13987 ( .A1(n11652), .A2(n11549), .ZN(n14202) );
  NAND2_X1 U13988 ( .A1(n11907), .A2(n11550), .ZN(n11551) );
  NAND3_X1 U13989 ( .A1(n11660), .A2(n14310), .A3(n11551), .ZN(n14203) );
  AOI22_X1 U13990 ( .A1(n14284), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n13575), 
        .B2(n14285), .ZN(n11553) );
  NAND2_X1 U13991 ( .A1(n11907), .A2(n14306), .ZN(n11552) );
  OAI211_X1 U13992 ( .C1(n14203), .C2(n14160), .A(n11553), .B(n11552), .ZN(
        n11554) );
  AOI21_X1 U13993 ( .B1(n14202), .B2(n14315), .A(n11554), .ZN(n11555) );
  OAI21_X1 U13994 ( .B1(n11556), .B2(n14284), .A(n11555), .ZN(P1_U3278) );
  INV_X1 U13995 ( .A(n11558), .ZN(n11561) );
  AOI21_X2 U13996 ( .B1(n11561), .B2(n11560), .A(n11559), .ZN(n11563) );
  XNOR2_X1 U13997 ( .A(n11624), .B(n12444), .ZN(n11669) );
  XNOR2_X1 U13998 ( .A(n11669), .B(n11672), .ZN(n11562) );
  NAND2_X1 U13999 ( .A1(n11563), .A2(n11562), .ZN(n11670) );
  OAI211_X1 U14000 ( .C1(n11563), .C2(n11562), .A(n11670), .B(n12509), .ZN(
        n11568) );
  INV_X1 U14001 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n11634) );
  OAI22_X1 U14002 ( .A1(n11564), .A2(n12503), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11634), .ZN(n11565) );
  AOI21_X1 U14003 ( .B1(n11566), .B2(n12523), .A(n11565), .ZN(n11567) );
  OAI211_X1 U14004 ( .C1(n12518), .C2(n11624), .A(n11568), .B(n11567), .ZN(
        P3_U3155) );
  INV_X1 U14005 ( .A(n14287), .ZN(n14372) );
  NOR2_X1 U14006 ( .A1(n11940), .A2(n11572), .ZN(n11573) );
  AOI21_X1 U14007 ( .B1(n14287), .B2(n12365), .A(n11573), .ZN(n11781) );
  AOI22_X1 U14008 ( .A1(n14287), .A2(n12363), .B1(n12365), .B2(n14130), .ZN(
        n11574) );
  XNOR2_X1 U14009 ( .A(n11574), .B(n12366), .ZN(n11782) );
  XOR2_X1 U14010 ( .A(n11781), .B(n11782), .Z(n11575) );
  OAI211_X1 U14011 ( .C1(n11576), .C2(n11575), .A(n14135), .B(n14139), .ZN(
        n11582) );
  NOR2_X1 U14012 ( .A1(n13890), .A2(n11577), .ZN(n14281) );
  NAND2_X1 U14013 ( .A1(n14141), .A2(n14281), .ZN(n11578) );
  OAI211_X1 U14014 ( .C1(n13570), .C2(n11792), .A(n11579), .B(n11578), .ZN(
        n11580) );
  AOI21_X1 U14015 ( .B1(n14286), .B2(n13576), .A(n11580), .ZN(n11581) );
  OAI211_X1 U14016 ( .C1(n14372), .C2(n13579), .A(n11582), .B(n11581), .ZN(
        P1_U3217) );
  INV_X1 U14017 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11584) );
  NAND2_X1 U14018 ( .A1(n11589), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n13700) );
  INV_X1 U14019 ( .A(n13700), .ZN(n11583) );
  AOI21_X1 U14020 ( .B1(n11584), .B2(n13702), .A(n11583), .ZN(n11587) );
  OAI21_X1 U14021 ( .B1(n11591), .B2(n11663), .A(n11585), .ZN(n11586) );
  NAND2_X1 U14022 ( .A1(n11587), .A2(n11586), .ZN(n13699) );
  OAI211_X1 U14023 ( .C1(n11587), .C2(n11586), .A(n13725), .B(n13699), .ZN(
        n11597) );
  NAND2_X1 U14024 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13512)
         );
  NOR2_X1 U14025 ( .A1(n11589), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n11588) );
  AOI21_X1 U14026 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n11589), .A(n11588), 
        .ZN(n11593) );
  OAI21_X1 U14027 ( .B1(n14201), .B2(n11591), .A(n11590), .ZN(n11592) );
  OAI211_X1 U14028 ( .C1(n11593), .C2(n11592), .A(n13701), .B(n13726), .ZN(
        n11594) );
  NAND2_X1 U14029 ( .A1(n13512), .A2(n11594), .ZN(n11595) );
  AOI21_X1 U14030 ( .B1(n13708), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n11595), 
        .ZN(n11596) );
  OAI211_X1 U14031 ( .C1(n14274), .C2(n13702), .A(n11597), .B(n11596), .ZN(
        P1_U3260) );
  OAI211_X1 U14032 ( .C1(n11600), .C2(n11599), .A(n11598), .B(n12768), .ZN(
        n11601) );
  AOI22_X1 U14033 ( .A1(n12765), .A2(n12544), .B1(n12545), .B2(n12763), .ZN(
        n11676) );
  NAND2_X1 U14034 ( .A1(n11601), .A2(n11676), .ZN(n11752) );
  INV_X1 U14035 ( .A(n11752), .ZN(n11606) );
  XNOR2_X1 U14036 ( .A(n11602), .B(n12244), .ZN(n11753) );
  AOI22_X1 U14037 ( .A1(n14772), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n12755), 
        .B2(n11679), .ZN(n11603) );
  OAI21_X1 U14038 ( .B1(n11759), .B2(n12757), .A(n11603), .ZN(n11604) );
  AOI21_X1 U14039 ( .B1(n11753), .B2(n12778), .A(n11604), .ZN(n11605) );
  OAI21_X1 U14040 ( .B1(n11606), .B2(n14772), .A(n11605), .ZN(P3_U3218) );
  INV_X1 U14041 ( .A(n11607), .ZN(n11609) );
  OAI222_X1 U14042 ( .A1(n11610), .A2(P3_U3151), .B1(n12880), .B2(n11609), 
        .C1(n11608), .C2(n12874), .ZN(P3_U3270) );
  INV_X1 U14043 ( .A(n11611), .ZN(n11615) );
  OAI222_X1 U14044 ( .A1(n12041), .A2(n11613), .B1(n13444), .B2(n11615), .C1(
        P2_U3088), .C2(n11612), .ZN(P2_U3302) );
  OAI222_X1 U14045 ( .A1(n14012), .A2(n11616), .B1(n14014), .B2(n11615), .C1(
        n11614), .C2(P1_U3086), .ZN(P1_U3330) );
  INV_X1 U14046 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n11619) );
  AOI21_X1 U14047 ( .B1(n14106), .B2(n11618), .A(n11617), .ZN(n11621) );
  MUX2_X1 U14048 ( .A(n11619), .B(n11621), .S(n14833), .Z(n11620) );
  OAI21_X1 U14049 ( .B1(n12865), .B2(n11624), .A(n11620), .ZN(P3_U3432) );
  INV_X1 U14050 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n11622) );
  MUX2_X1 U14051 ( .A(n11622), .B(n11621), .S(n14846), .Z(n11623) );
  OAI21_X1 U14052 ( .B1(n12826), .B2(n11624), .A(n11623), .ZN(P3_U3473) );
  NOR2_X1 U14053 ( .A1(n11626), .A2(n11625), .ZN(n11628) );
  XNOR2_X1 U14054 ( .A(n12561), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n11639) );
  AOI21_X1 U14055 ( .B1(n6585), .B2(n11639), .A(n12558), .ZN(n11650) );
  NOR2_X1 U14056 ( .A1(n12561), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n11629) );
  AOI21_X1 U14057 ( .B1(P3_REG1_REG_14__SCAN_IN), .B2(n12561), .A(n11629), 
        .ZN(n11637) );
  NAND2_X1 U14058 ( .A1(n11640), .A2(n11630), .ZN(n11632) );
  OAI21_X1 U14059 ( .B1(n11637), .B2(n11633), .A(n12562), .ZN(n11648) );
  NOR2_X1 U14060 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11634), .ZN(n11635) );
  AOI21_X1 U14061 ( .B1(n14743), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n11635), 
        .ZN(n11636) );
  OAI21_X1 U14062 ( .B1(n14740), .B2(n12561), .A(n11636), .ZN(n11647) );
  INV_X1 U14063 ( .A(n11637), .ZN(n11638) );
  MUX2_X1 U14064 ( .A(n11639), .B(n11638), .S(n12073), .Z(n11645) );
  NOR2_X1 U14065 ( .A1(n11641), .A2(n11640), .ZN(n11642) );
  OR2_X1 U14066 ( .A1(n11643), .A2(n11642), .ZN(n11644) );
  AOI211_X1 U14067 ( .C1(n11645), .C2(n11644), .A(n14709), .B(n12570), .ZN(
        n11646) );
  AOI211_X1 U14068 ( .C1(n11648), .C2(n14746), .A(n11647), .B(n11646), .ZN(
        n11649) );
  OAI21_X1 U14069 ( .B1(n11650), .B2(n14750), .A(n11649), .ZN(P3_U3196) );
  OR2_X1 U14070 ( .A1(n11907), .A2(n13587), .ZN(n11651) );
  XNOR2_X1 U14071 ( .A(n11843), .B(n11864), .ZN(n14194) );
  INV_X1 U14072 ( .A(n14194), .ZN(n11668) );
  XNOR2_X1 U14073 ( .A(n11865), .B(n11864), .ZN(n11657) );
  NAND2_X1 U14074 ( .A1(n11657), .A2(n14353), .ZN(n11659) );
  AOI22_X1 U14075 ( .A1(n13585), .A2(n14292), .B1(n14131), .B2(n13587), .ZN(
        n11658) );
  NAND2_X1 U14076 ( .A1(n11659), .A2(n11658), .ZN(n14200) );
  NAND2_X1 U14077 ( .A1(n11660), .A2(n14195), .ZN(n11661) );
  NAND2_X1 U14078 ( .A1(n11661), .A2(n14310), .ZN(n11662) );
  OR2_X1 U14079 ( .A1(n14159), .A2(n11662), .ZN(n14196) );
  OAI22_X1 U14080 ( .A1(n14303), .A2(n11663), .B1(n13504), .B2(n14302), .ZN(
        n11664) );
  AOI21_X1 U14081 ( .B1(n14195), .B2(n14306), .A(n11664), .ZN(n11665) );
  OAI21_X1 U14082 ( .B1(n14196), .B2(n14160), .A(n11665), .ZN(n11666) );
  AOI21_X1 U14083 ( .B1(n14200), .B2(n14303), .A(n11666), .ZN(n11667) );
  OAI21_X1 U14084 ( .B1(n13887), .B2(n11668), .A(n11667), .ZN(P1_U3277) );
  XNOR2_X1 U14085 ( .A(n12246), .B(n12444), .ZN(n11812) );
  XNOR2_X1 U14086 ( .A(n11812), .B(n12247), .ZN(n11674) );
  INV_X1 U14087 ( .A(n11669), .ZN(n11671) );
  OAI21_X1 U14088 ( .B1(n11672), .B2(n11671), .A(n11670), .ZN(n11673) );
  AOI21_X1 U14089 ( .B1(n11674), .B2(n11673), .A(n11814), .ZN(n11681) );
  INV_X1 U14090 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n11675) );
  OAI22_X1 U14091 ( .A1(n11676), .A2(n12503), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11675), .ZN(n11678) );
  NOR2_X1 U14092 ( .A1(n11759), .A2(n12518), .ZN(n11677) );
  AOI211_X1 U14093 ( .C1(n11679), .C2(n12523), .A(n11678), .B(n11677), .ZN(
        n11680) );
  OAI21_X1 U14094 ( .B1(n11681), .B2(n12531), .A(n11680), .ZN(P3_U3181) );
  XOR2_X1 U14095 ( .A(n11682), .B(n12127), .Z(n11684) );
  AOI22_X1 U14096 ( .A1(n12763), .A2(n11683), .B1(n12764), .B2(n12765), .ZN(
        n11817) );
  OAI21_X1 U14097 ( .B1(n11684), .B2(n14767), .A(n11817), .ZN(n11806) );
  INV_X1 U14098 ( .A(n11806), .ZN(n11689) );
  XNOR2_X1 U14099 ( .A(n11685), .B(n12127), .ZN(n11807) );
  AOI22_X1 U14100 ( .A1(n14772), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n12755), 
        .B2(n11819), .ZN(n11686) );
  OAI21_X1 U14101 ( .B1(n11822), .B2(n12757), .A(n11686), .ZN(n11687) );
  AOI21_X1 U14102 ( .B1(n11807), .B2(n12778), .A(n11687), .ZN(n11688) );
  OAI21_X1 U14103 ( .B1(n11689), .B2(n14772), .A(n11688), .ZN(P3_U3217) );
  INV_X1 U14104 ( .A(n11690), .ZN(n11692) );
  OAI222_X1 U14105 ( .A1(n11693), .A2(P3_U3151), .B1(n12880), .B2(n11692), 
        .C1(n11691), .C2(n12874), .ZN(P3_U3269) );
  XNOR2_X1 U14106 ( .A(n13392), .B(n12948), .ZN(n11696) );
  NAND2_X1 U14107 ( .A1(n12916), .A2(n13061), .ZN(n11697) );
  XNOR2_X1 U14108 ( .A(n11696), .B(n11697), .ZN(n11994) );
  INV_X1 U14109 ( .A(n11696), .ZN(n11698) );
  NAND2_X1 U14110 ( .A1(n11698), .A2(n11697), .ZN(n11699) );
  AOI22_X1 U14111 ( .A1(n11701), .A2(n13035), .B1(n13013), .B2(n13060), .ZN(
        n11707) );
  AND2_X1 U14112 ( .A1(n12916), .A2(n13060), .ZN(n11700) );
  INV_X1 U14113 ( .A(n11967), .ZN(n11706) );
  NOR2_X1 U14114 ( .A1(n13015), .A2(n11716), .ZN(n11704) );
  INV_X1 U14115 ( .A(n13061), .ZN(n11720) );
  OAI22_X1 U14116 ( .A1(n12001), .A2(n12997), .B1(n11720), .B2(n12995), .ZN(
        n11725) );
  INV_X1 U14117 ( .A(n11725), .ZN(n11702) );
  OAI22_X1 U14118 ( .A1(n13040), .A2(n11702), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7742), .ZN(n11703) );
  AOI211_X1 U14119 ( .C1(n13387), .C2(n6418), .A(n11704), .B(n11703), .ZN(
        n11705) );
  OAI21_X1 U14120 ( .B1(n11707), .B2(n11706), .A(n11705), .ZN(P2_U3213) );
  NAND2_X1 U14121 ( .A1(n11711), .A2(n11710), .ZN(n11769) );
  XNOR2_X1 U14122 ( .A(n11769), .B(n11719), .ZN(n13390) );
  AOI21_X1 U14123 ( .B1(n13387), .B2(n11712), .A(n13289), .ZN(n11715) );
  AND2_X1 U14124 ( .A1(n11715), .A2(n11760), .ZN(n13386) );
  INV_X1 U14125 ( .A(n11716), .ZN(n11717) );
  AOI22_X1 U14126 ( .A1(n13304), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n11717), 
        .B2(n13291), .ZN(n11718) );
  OAI21_X1 U14127 ( .B1(n11713), .B2(n13294), .A(n11718), .ZN(n11728) );
  INV_X1 U14128 ( .A(n11719), .ZN(n11768) );
  NAND2_X1 U14129 ( .A1(n13392), .A2(n11720), .ZN(n11722) );
  OAI21_X1 U14130 ( .B1(n11768), .B2(n11724), .A(n11762), .ZN(n11726) );
  AOI21_X1 U14131 ( .B1(n11726), .B2(n13284), .A(n11725), .ZN(n13389) );
  NOR2_X1 U14132 ( .A1(n13389), .A2(n13304), .ZN(n11727) );
  AOI211_X1 U14133 ( .C1(n13386), .C2(n13302), .A(n11728), .B(n11727), .ZN(
        n11729) );
  OAI21_X1 U14134 ( .B1(n13299), .B2(n13390), .A(n11729), .ZN(P2_U3250) );
  NAND2_X1 U14135 ( .A1(n11731), .A2(n11730), .ZN(n11733) );
  NAND2_X1 U14136 ( .A1(n14511), .A2(n11734), .ZN(n11735) );
  NOR2_X1 U14137 ( .A1(n11737), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11736) );
  AOI21_X1 U14138 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n11737), .A(n11736), 
        .ZN(n11738) );
  NAND2_X1 U14139 ( .A1(n11738), .A2(n11739), .ZN(n13075) );
  OAI211_X1 U14140 ( .C1(n11739), .C2(n11738), .A(n14526), .B(n13075), .ZN(
        n11751) );
  NAND2_X1 U14141 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n12978)
         );
  OAI21_X1 U14142 ( .B1(n11742), .B2(n11741), .A(n11740), .ZN(n11743) );
  NAND2_X1 U14143 ( .A1(n14511), .A2(n11743), .ZN(n11745) );
  XNOR2_X1 U14144 ( .A(n11744), .B(n11743), .ZN(n14515) );
  NAND2_X1 U14145 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n14515), .ZN(n14514) );
  NAND2_X1 U14146 ( .A1(n11745), .A2(n14514), .ZN(n11747) );
  XNOR2_X1 U14147 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13083), .ZN(n11746) );
  NAND2_X1 U14148 ( .A1(n11746), .A2(n11747), .ZN(n13081) );
  OAI211_X1 U14149 ( .C1(n11747), .C2(n11746), .A(n14542), .B(n13081), .ZN(
        n11748) );
  NAND2_X1 U14150 ( .A1(n12978), .A2(n11748), .ZN(n11749) );
  AOI21_X1 U14151 ( .B1(n14540), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n11749), 
        .ZN(n11750) );
  OAI211_X1 U14152 ( .C1(n14547), .C2(n13083), .A(n11751), .B(n11750), .ZN(
        P2_U3230) );
  INV_X1 U14153 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n11754) );
  AOI21_X1 U14154 ( .B1(n14106), .B2(n11753), .A(n11752), .ZN(n11756) );
  MUX2_X1 U14155 ( .A(n11754), .B(n11756), .S(n14833), .Z(n11755) );
  OAI21_X1 U14156 ( .B1(n11759), .B2(n12865), .A(n11755), .ZN(P3_U3435) );
  INV_X1 U14157 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n11757) );
  MUX2_X1 U14158 ( .A(n11757), .B(n11756), .S(n14846), .Z(n11758) );
  OAI21_X1 U14159 ( .B1(n11759), .B2(n12826), .A(n11758), .ZN(P3_U3474) );
  AOI21_X1 U14160 ( .B1(n13378), .B2(n11760), .A(n13286), .ZN(n13380) );
  NOR2_X1 U14161 ( .A1(n13245), .A2(n12979), .ZN(n11767) );
  NAND2_X1 U14162 ( .A1(n11762), .A2(n11761), .ZN(n12003) );
  INV_X1 U14163 ( .A(n11763), .ZN(n11771) );
  XNOR2_X1 U14164 ( .A(n12003), .B(n11771), .ZN(n11765) );
  OAI22_X1 U14165 ( .A1(n12004), .A2(n12997), .B1(n11764), .B2(n12995), .ZN(
        n12976) );
  AOI21_X1 U14166 ( .B1(n11765), .B2(n13284), .A(n12976), .ZN(n13385) );
  INV_X1 U14167 ( .A(n13385), .ZN(n11766) );
  AOI211_X1 U14168 ( .C1(n11970), .C2(n13380), .A(n11767), .B(n11766), .ZN(
        n11775) );
  AOI22_X1 U14169 ( .A1(n13378), .A2(n13241), .B1(n13304), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n11774) );
  OR2_X1 U14170 ( .A1(n13387), .A2(n13060), .ZN(n11770) );
  NAND2_X1 U14171 ( .A1(n11772), .A2(n11771), .ZN(n13381) );
  NAND3_X1 U14172 ( .A1(n13382), .A2(n13381), .A3(n13232), .ZN(n11773) );
  OAI211_X1 U14173 ( .C1(n11775), .C2(n13304), .A(n11774), .B(n11773), .ZN(
        P2_U3249) );
  NOR2_X1 U14174 ( .A1(n11940), .A2(n11792), .ZN(n11776) );
  AOI21_X1 U14175 ( .B1(n14172), .B2(n12365), .A(n11776), .ZN(n11780) );
  INV_X1 U14176 ( .A(n11780), .ZN(n11785) );
  NAND2_X1 U14177 ( .A1(n14172), .A2(n12363), .ZN(n11778) );
  NAND2_X1 U14178 ( .A1(n12365), .A2(n14291), .ZN(n11777) );
  NAND2_X1 U14179 ( .A1(n11778), .A2(n11777), .ZN(n11779) );
  XNOR2_X1 U14180 ( .A(n11779), .B(n12366), .ZN(n11784) );
  XNOR2_X1 U14181 ( .A(n11784), .B(n11780), .ZN(n14137) );
  OR2_X1 U14182 ( .A1(n11782), .A2(n11781), .ZN(n14134) );
  AOI22_X1 U14183 ( .A1(n11787), .A2(n12363), .B1(n12365), .B2(n14129), .ZN(
        n11786) );
  XNOR2_X1 U14184 ( .A(n11786), .B(n12366), .ZN(n11823) );
  AOI22_X1 U14185 ( .A1(n11787), .A2(n12365), .B1(n12364), .B2(n14129), .ZN(
        n11824) );
  XNOR2_X1 U14186 ( .A(n11823), .B(n11824), .ZN(n11789) );
  AOI21_X1 U14187 ( .B1(n11788), .B2(n11789), .A(n13564), .ZN(n11790) );
  NAND2_X1 U14188 ( .A1(n11790), .A2(n11828), .ZN(n11797) );
  INV_X1 U14189 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n13688) );
  OAI22_X1 U14190 ( .A1(n13570), .A2(n11791), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13688), .ZN(n11794) );
  INV_X1 U14191 ( .A(n13557), .ZN(n13572) );
  NOR2_X1 U14192 ( .A1(n13572), .A2(n11792), .ZN(n11793) );
  AOI211_X1 U14193 ( .C1(n13576), .C2(n11795), .A(n11794), .B(n11793), .ZN(
        n11796) );
  OAI211_X1 U14194 ( .C1(n11798), .C2(n13579), .A(n11797), .B(n11796), .ZN(
        P1_U3224) );
  XNOR2_X1 U14195 ( .A(n11799), .B(n12126), .ZN(n11800) );
  OAI222_X1 U14196 ( .A1(n14760), .A2(n12478), .B1(n14762), .B2(n12476), .C1(
        n11800), .C2(n14767), .ZN(n12822) );
  INV_X1 U14197 ( .A(n12822), .ZN(n11805) );
  XNOR2_X1 U14198 ( .A(n11801), .B(n12258), .ZN(n12823) );
  AOI22_X1 U14199 ( .A1(n14772), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n12755), 
        .B2(n12481), .ZN(n11802) );
  OAI21_X1 U14200 ( .B1(n12866), .B2(n12757), .A(n11802), .ZN(n11803) );
  AOI21_X1 U14201 ( .B1(n12823), .B2(n12778), .A(n11803), .ZN(n11804) );
  OAI21_X1 U14202 ( .B1(n11805), .B2(n14772), .A(n11804), .ZN(P3_U3216) );
  INV_X1 U14203 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n11808) );
  AOI21_X1 U14204 ( .B1(n14106), .B2(n11807), .A(n11806), .ZN(n11810) );
  MUX2_X1 U14205 ( .A(n11808), .B(n11810), .S(n14833), .Z(n11809) );
  OAI21_X1 U14206 ( .B1(n11822), .B2(n12865), .A(n11809), .ZN(P3_U3438) );
  INV_X1 U14207 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12591) );
  MUX2_X1 U14208 ( .A(n12591), .B(n11810), .S(n14846), .Z(n11811) );
  OAI21_X1 U14209 ( .B1(n11822), .B2(n12826), .A(n11811), .ZN(P3_U3475) );
  XNOR2_X1 U14210 ( .A(n12254), .B(n12444), .ZN(n12383) );
  XNOR2_X1 U14211 ( .A(n12383), .B(n12544), .ZN(n11815) );
  OAI211_X1 U14212 ( .C1(n6586), .C2(n11815), .A(n12384), .B(n12509), .ZN(
        n11821) );
  OAI22_X1 U14213 ( .A1(n11817), .A2(n12503), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11816), .ZN(n11818) );
  AOI21_X1 U14214 ( .B1(n11819), .B2(n12523), .A(n11818), .ZN(n11820) );
  OAI211_X1 U14215 ( .C1(n11822), .C2(n12518), .A(n11821), .B(n11820), .ZN(
        P3_U3166) );
  INV_X1 U14216 ( .A(n11823), .ZN(n11826) );
  INV_X1 U14217 ( .A(n11824), .ZN(n11825) );
  NAND2_X1 U14218 ( .A1(n11826), .A2(n11825), .ZN(n11827) );
  NAND2_X1 U14219 ( .A1(n11832), .A2(n12363), .ZN(n11830) );
  NAND2_X1 U14220 ( .A1(n12365), .A2(n13589), .ZN(n11829) );
  NAND2_X1 U14221 ( .A1(n11830), .A2(n11829), .ZN(n11831) );
  XNOR2_X1 U14222 ( .A(n11831), .B(n12366), .ZN(n11898) );
  AOI22_X1 U14223 ( .A1(n11832), .A2(n12365), .B1(n12364), .B2(n13589), .ZN(
        n11896) );
  XNOR2_X1 U14224 ( .A(n11898), .B(n11896), .ZN(n11833) );
  OAI211_X1 U14225 ( .C1(n11834), .C2(n11833), .A(n14121), .B(n14139), .ZN(
        n11840) );
  NAND2_X1 U14226 ( .A1(n13557), .A2(n14129), .ZN(n11836) );
  OAI211_X1 U14227 ( .C1(n13571), .C2(n13570), .A(n11836), .B(n11835), .ZN(
        n11837) );
  AOI21_X1 U14228 ( .B1(n11838), .B2(n13576), .A(n11837), .ZN(n11839) );
  OAI211_X1 U14229 ( .C1(n14219), .C2(n13579), .A(n11840), .B(n11839), .ZN(
        P1_U3234) );
  INV_X1 U14230 ( .A(n11841), .ZN(n13440) );
  OAI222_X1 U14231 ( .A1(n14012), .A2(n11842), .B1(n14014), .B2(n13440), .C1(
        n8847), .C2(P1_U3086), .ZN(P1_U3328) );
  NAND2_X1 U14232 ( .A1(n11843), .A2(n11864), .ZN(n11845) );
  OR2_X1 U14233 ( .A1(n14195), .A2(n13586), .ZN(n11844) );
  NAND2_X1 U14234 ( .A1(n11845), .A2(n11844), .ZN(n14156) );
  NAND2_X1 U14235 ( .A1(n14154), .A2(n13585), .ZN(n11846) );
  OR2_X1 U14236 ( .A1(n14180), .A2(n13875), .ZN(n11848) );
  INV_X1 U14237 ( .A(n13871), .ZN(n11870) );
  INV_X1 U14238 ( .A(n13893), .ZN(n13584) );
  OR2_X1 U14239 ( .A1(n13874), .A2(n13584), .ZN(n11849) );
  OR2_X1 U14240 ( .A1(n13971), .A2(n13476), .ZN(n11853) );
  INV_X1 U14241 ( .A(n13842), .ZN(n13850) );
  NAND2_X1 U14242 ( .A1(n13836), .A2(n13837), .ZN(n11855) );
  OR2_X1 U14243 ( .A1(n13960), .A2(n13583), .ZN(n11854) );
  NAND2_X1 U14244 ( .A1(n13952), .A2(n13827), .ZN(n11856) );
  INV_X1 U14245 ( .A(n13454), .ZN(n13930) );
  INV_X1 U14246 ( .A(n13582), .ZN(n13452) );
  INV_X1 U14247 ( .A(n11878), .ZN(n11861) );
  INV_X1 U14248 ( .A(n13586), .ZN(n13569) );
  NAND2_X1 U14249 ( .A1(n14195), .A2(n13569), .ZN(n11863) );
  NAND2_X1 U14250 ( .A1(n13888), .A2(n13897), .ZN(n11869) );
  INV_X1 U14251 ( .A(n13875), .ZN(n11867) );
  OR2_X1 U14252 ( .A1(n14180), .A2(n11867), .ZN(n11868) );
  NAND2_X1 U14253 ( .A1(n13971), .A2(n13876), .ZN(n11872) );
  NAND2_X1 U14254 ( .A1(n13854), .A2(n11872), .ZN(n13841) );
  NAND2_X1 U14255 ( .A1(n13841), .A2(n13850), .ZN(n11874) );
  OR2_X1 U14256 ( .A1(n13965), .A2(n13531), .ZN(n11873) );
  INV_X1 U14257 ( .A(n13583), .ZN(n11875) );
  NAND2_X1 U14258 ( .A1(n13960), .A2(n11875), .ZN(n11876) );
  INV_X1 U14259 ( .A(n13827), .ZN(n13530) );
  NAND2_X1 U14260 ( .A1(n13952), .A2(n13530), .ZN(n11877) );
  INV_X1 U14261 ( .A(n13793), .ZN(n13795) );
  INV_X1 U14262 ( .A(n13805), .ZN(n13947) );
  NAND2_X1 U14263 ( .A1(n13947), .A2(n13779), .ZN(n13775) );
  NAND3_X1 U14264 ( .A1(n13798), .A2(n13785), .A3(n13775), .ZN(n13776) );
  INV_X1 U14265 ( .A(n13942), .ZN(n13784) );
  NAND2_X1 U14266 ( .A1(n13776), .A2(n7352), .ZN(n13763) );
  INV_X1 U14267 ( .A(n13760), .ZN(n13762) );
  NAND2_X1 U14268 ( .A1(n14159), .A2(n14190), .ZN(n14158) );
  NOR2_X2 U14269 ( .A1(n6487), .A2(n13942), .ZN(n13781) );
  NAND2_X1 U14270 ( .A1(n13936), .A2(n13781), .ZN(n13764) );
  NOR2_X2 U14271 ( .A1(n11880), .A2(n13754), .ZN(n13739) );
  AOI211_X1 U14272 ( .C1(n11880), .C2(n13754), .A(n14182), .B(n13739), .ZN(
        n13921) );
  NAND2_X1 U14273 ( .A1(n13921), .A2(n14314), .ZN(n11889) );
  NOR2_X1 U14274 ( .A1(n8847), .A2(n11881), .ZN(n11882) );
  NOR2_X1 U14275 ( .A1(n13892), .A2(n11882), .ZN(n13735) );
  NAND2_X1 U14276 ( .A1(n13735), .A2(n13580), .ZN(n13918) );
  INV_X1 U14277 ( .A(n11883), .ZN(n11884) );
  OAI22_X1 U14278 ( .A1(n11885), .A2(n13918), .B1(n11884), .B2(n14302), .ZN(
        n11887) );
  NAND2_X1 U14279 ( .A1(n14131), .A2(n13582), .ZN(n13917) );
  NOR2_X1 U14280 ( .A1(n13880), .A2(n13917), .ZN(n11886) );
  AOI211_X1 U14281 ( .C1(n13880), .C2(P1_REG2_REG_29__SCAN_IN), .A(n11887), 
        .B(n11886), .ZN(n11888) );
  OAI211_X1 U14282 ( .C1(n13919), .C2(n13883), .A(n11889), .B(n11888), .ZN(
        n11890) );
  AOI21_X1 U14283 ( .B1(n13885), .B2(n13916), .A(n11890), .ZN(n11891) );
  OAI21_X1 U14284 ( .B1(n13923), .B2(n13887), .A(n11891), .ZN(P1_U3356) );
  NAND2_X1 U14285 ( .A1(n14210), .A2(n12363), .ZN(n11893) );
  NAND2_X1 U14286 ( .A1(n12365), .A2(n13588), .ZN(n11892) );
  NAND2_X1 U14287 ( .A1(n11893), .A2(n11892), .ZN(n11894) );
  XNOR2_X1 U14288 ( .A(n11894), .B(n12366), .ZN(n11902) );
  NOR2_X1 U14289 ( .A1(n11940), .A2(n13571), .ZN(n11895) );
  AOI21_X1 U14290 ( .B1(n14210), .B2(n12365), .A(n11895), .ZN(n11900) );
  XNOR2_X1 U14291 ( .A(n11902), .B(n11900), .ZN(n14123) );
  INV_X1 U14292 ( .A(n11896), .ZN(n11897) );
  NAND2_X1 U14293 ( .A1(n11898), .A2(n11897), .ZN(n14120) );
  INV_X1 U14294 ( .A(n11900), .ZN(n11901) );
  NAND2_X1 U14295 ( .A1(n11907), .A2(n12363), .ZN(n11905) );
  NAND2_X1 U14296 ( .A1(n12365), .A2(n13587), .ZN(n11904) );
  NAND2_X1 U14297 ( .A1(n11905), .A2(n11904), .ZN(n11906) );
  XNOR2_X1 U14298 ( .A(n11906), .B(n12366), .ZN(n11909) );
  OAI22_X1 U14299 ( .A1(n6891), .A2(n11941), .B1(n11908), .B2(n11940), .ZN(
        n13567) );
  INV_X1 U14300 ( .A(n11909), .ZN(n11910) );
  AOI22_X1 U14301 ( .A1(n14195), .A2(n12363), .B1(n12365), .B2(n13586), .ZN(
        n11912) );
  XNOR2_X1 U14302 ( .A(n11912), .B(n12366), .ZN(n11913) );
  AOI22_X1 U14303 ( .A1(n14195), .A2(n12365), .B1(n12364), .B2(n13586), .ZN(
        n11914) );
  XNOR2_X1 U14304 ( .A(n11913), .B(n11914), .ZN(n13500) );
  NAND2_X1 U14305 ( .A1(n14154), .A2(n12363), .ZN(n11917) );
  NAND2_X1 U14306 ( .A1(n13585), .A2(n12365), .ZN(n11916) );
  NAND2_X1 U14307 ( .A1(n11917), .A2(n11916), .ZN(n11918) );
  XNOR2_X1 U14308 ( .A(n11918), .B(n12366), .ZN(n11932) );
  AOI22_X1 U14309 ( .A1(n14154), .A2(n12365), .B1(n12364), .B2(n13585), .ZN(
        n11933) );
  XNOR2_X1 U14310 ( .A(n11932), .B(n11933), .ZN(n13508) );
  NAND2_X1 U14311 ( .A1(n14180), .A2(n12363), .ZN(n11920) );
  NAND2_X1 U14312 ( .A1(n13875), .A2(n12365), .ZN(n11919) );
  NAND2_X1 U14313 ( .A1(n11920), .A2(n11919), .ZN(n11921) );
  XNOR2_X1 U14314 ( .A(n11921), .B(n12366), .ZN(n11924) );
  INV_X1 U14315 ( .A(n11924), .ZN(n11922) );
  AOI22_X1 U14316 ( .A1(n14180), .A2(n12365), .B1(n12364), .B2(n13875), .ZN(
        n11923) );
  NAND2_X1 U14317 ( .A1(n11922), .A2(n11923), .ZN(n11935) );
  INV_X1 U14318 ( .A(n11935), .ZN(n11925) );
  XNOR2_X1 U14319 ( .A(n11924), .B(n11923), .ZN(n13549) );
  OR2_X1 U14320 ( .A1(n11925), .A2(n13549), .ZN(n11931) );
  AND2_X1 U14321 ( .A1(n13508), .A2(n11931), .ZN(n13467) );
  OAI22_X1 U14322 ( .A1(n13977), .A2(n11942), .B1(n13893), .B2(n11941), .ZN(
        n11926) );
  XNOR2_X1 U14323 ( .A(n11926), .B(n12366), .ZN(n11930) );
  OAI22_X1 U14324 ( .A1(n13977), .A2(n11941), .B1(n13893), .B2(n11940), .ZN(
        n11929) );
  NAND2_X1 U14325 ( .A1(n11930), .A2(n11929), .ZN(n11928) );
  AND2_X1 U14326 ( .A1(n13467), .A2(n11928), .ZN(n11927) );
  INV_X1 U14327 ( .A(n11928), .ZN(n11939) );
  XNOR2_X1 U14328 ( .A(n11930), .B(n11929), .ZN(n13469) );
  INV_X1 U14329 ( .A(n13469), .ZN(n11938) );
  INV_X1 U14330 ( .A(n11931), .ZN(n11937) );
  INV_X1 U14331 ( .A(n11932), .ZN(n11934) );
  NAND2_X1 U14332 ( .A1(n11934), .A2(n11933), .ZN(n13546) );
  AND2_X1 U14333 ( .A1(n13546), .A2(n11935), .ZN(n11936) );
  OR2_X1 U14334 ( .A1(n11937), .A2(n11936), .ZN(n13468) );
  AND2_X1 U14335 ( .A1(n11938), .A2(n13468), .ZN(n13471) );
  OR2_X1 U14336 ( .A1(n11939), .A2(n13471), .ZN(n11944) );
  AND2_X1 U14337 ( .A1(n11946), .A2(n11944), .ZN(n11948) );
  OAI22_X1 U14338 ( .A1(n13971), .A2(n11941), .B1(n13476), .B2(n11940), .ZN(
        n12314) );
  OAI22_X1 U14339 ( .A1(n13971), .A2(n11942), .B1(n13476), .B2(n11941), .ZN(
        n11943) );
  XNOR2_X1 U14340 ( .A(n11943), .B(n12366), .ZN(n12315) );
  XOR2_X1 U14341 ( .A(n12314), .B(n12315), .Z(n11947) );
  AND2_X1 U14342 ( .A1(n11947), .A2(n11944), .ZN(n11945) );
  OAI211_X1 U14343 ( .C1(n11948), .C2(n11947), .A(n12317), .B(n14139), .ZN(
        n11953) );
  INV_X1 U14344 ( .A(n13861), .ZN(n11951) );
  AOI22_X1 U14345 ( .A1(n13584), .A2(n14131), .B1(n14292), .B2(n13828), .ZN(
        n13969) );
  OAI22_X1 U14346 ( .A1(n13969), .A2(n13513), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11949), .ZN(n11950) );
  AOI21_X1 U14347 ( .B1(n11951), .B2(n13576), .A(n11950), .ZN(n11952) );
  OAI211_X1 U14348 ( .C1(n13971), .C2(n13579), .A(n11953), .B(n11952), .ZN(
        P1_U3233) );
  INV_X1 U14349 ( .A(n11954), .ZN(n11962) );
  AOI22_X1 U14350 ( .A1(n13013), .A2(n8148), .B1(n13035), .B2(n11956), .ZN(
        n11959) );
  INV_X1 U14351 ( .A(n10240), .ZN(n11958) );
  NOR3_X1 U14352 ( .A1(n11959), .A2(n11958), .A3(n11957), .ZN(n11960) );
  AOI211_X1 U14353 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n11962), .A(n11961), .B(
        n11960), .ZN(n11963) );
  OAI21_X1 U14354 ( .B1(n11964), .B2(n13023), .A(n11963), .ZN(P2_U3209) );
  XNOR2_X1 U14355 ( .A(n13378), .B(n12917), .ZN(n11979) );
  NAND2_X1 U14356 ( .A1(n6458), .A2(n13059), .ZN(n11968) );
  XNOR2_X1 U14357 ( .A(n11979), .B(n11968), .ZN(n12975) );
  NAND2_X1 U14358 ( .A1(n11979), .A2(n11968), .ZN(n11969) );
  NAND2_X1 U14359 ( .A1(n11977), .A2(n11969), .ZN(n11971) );
  XNOR2_X1 U14360 ( .A(n13295), .B(n12948), .ZN(n12883) );
  NOR2_X1 U14361 ( .A1(n12004), .A2(n11970), .ZN(n12881) );
  XNOR2_X1 U14362 ( .A(n12883), .B(n12881), .ZN(n11978) );
  INV_X1 U14363 ( .A(n13292), .ZN(n11975) );
  NAND2_X1 U14364 ( .A1(n13057), .A2(n13037), .ZN(n11973) );
  NAND2_X1 U14365 ( .A1(n13059), .A2(n13038), .ZN(n11972) );
  NAND2_X1 U14366 ( .A1(n11973), .A2(n11972), .ZN(n13283) );
  AOI22_X1 U14367 ( .A1(n12999), .A2(n13283), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11974) );
  OAI21_X1 U14368 ( .B1(n13015), .B2(n11975), .A(n11974), .ZN(n11976) );
  AOI21_X1 U14369 ( .B1(n13374), .B2(n6418), .A(n11976), .ZN(n11983) );
  INV_X1 U14370 ( .A(n11978), .ZN(n11981) );
  OAI22_X1 U14371 ( .A1(n11979), .A2(n13023), .B1(n12001), .B2(n11989), .ZN(
        n11980) );
  NAND3_X1 U14372 ( .A1(n11977), .A2(n11981), .A3(n11980), .ZN(n11982) );
  OAI211_X1 U14373 ( .C1(n12885), .C2(n13023), .A(n11983), .B(n11982), .ZN(
        P2_U3200) );
  INV_X1 U14374 ( .A(n11984), .ZN(n11988) );
  NAND2_X1 U14375 ( .A1(n12999), .A2(n11985), .ZN(n11986) );
  OAI211_X1 U14376 ( .C1(n13015), .C2(n11988), .A(n11987), .B(n11986), .ZN(
        n11997) );
  NOR3_X1 U14377 ( .A1(n11991), .A2(n11990), .A3(n11989), .ZN(n11992) );
  AOI21_X1 U14378 ( .B1(n11993), .B2(n13035), .A(n11992), .ZN(n11995) );
  NOR2_X1 U14379 ( .A1(n11995), .A2(n11994), .ZN(n11996) );
  AOI211_X1 U14380 ( .C1(n13392), .C2(n6418), .A(n11997), .B(n11996), .ZN(
        n11998) );
  OAI21_X1 U14381 ( .B1(n11999), .B2(n13023), .A(n11998), .ZN(P2_U3187) );
  INV_X1 U14382 ( .A(n13349), .ZN(n12008) );
  INV_X1 U14383 ( .A(n13369), .ZN(n13274) );
  NAND2_X1 U14384 ( .A1(n12000), .A2(n13059), .ZN(n12002) );
  AOI22_X1 U14385 ( .A1(n12003), .A2(n12002), .B1(n12001), .B2(n13378), .ZN(
        n13282) );
  INV_X1 U14386 ( .A(n13365), .ZN(n13262) );
  INV_X1 U14387 ( .A(n13246), .ZN(n13235) );
  INV_X1 U14388 ( .A(n13354), .ZN(n13230) );
  INV_X1 U14389 ( .A(n13344), .ZN(n12009) );
  INV_X1 U14390 ( .A(n13338), .ZN(n13184) );
  INV_X1 U14391 ( .A(n13161), .ZN(n13156) );
  INV_X1 U14392 ( .A(n12010), .ZN(n12011) );
  XNOR2_X1 U14393 ( .A(n12015), .B(n12038), .ZN(n12019) );
  OAI21_X1 U14394 ( .B1(n8183), .B2(n12016), .A(n13037), .ZN(n13100) );
  INV_X1 U14395 ( .A(n13046), .ZN(n12017) );
  OAI22_X1 U14396 ( .A1(n13100), .A2(n12017), .B1(n12922), .B2(n12995), .ZN(
        n12018) );
  OR2_X2 U14397 ( .A1(n13349), .A2(n13226), .ZN(n13207) );
  NOR2_X2 U14398 ( .A1(n13113), .A2(n13310), .ZN(n13107) );
  AOI211_X1 U14399 ( .C1(n13310), .C2(n13113), .A(n13289), .B(n13107), .ZN(
        n13309) );
  INV_X1 U14400 ( .A(n12020), .ZN(n12021) );
  AOI22_X1 U14401 ( .A1(n13304), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n12021), 
        .B2(n13291), .ZN(n12022) );
  OAI21_X1 U14402 ( .B1(n12023), .B2(n13294), .A(n12022), .ZN(n12040) );
  NAND2_X1 U14403 ( .A1(n13378), .A2(n13059), .ZN(n12024) );
  INV_X1 U14404 ( .A(n12025), .ZN(n12026) );
  NAND2_X1 U14405 ( .A1(n13296), .A2(n12026), .ZN(n13277) );
  INV_X1 U14406 ( .A(n13277), .ZN(n12028) );
  OR2_X1 U14407 ( .A1(n13365), .A2(n13056), .ZN(n12029) );
  OR2_X1 U14408 ( .A1(n13369), .A2(n13057), .ZN(n13251) );
  AND2_X1 U14409 ( .A1(n12029), .A2(n13251), .ZN(n12030) );
  NAND2_X1 U14410 ( .A1(n13365), .A2(n13056), .ZN(n12031) );
  AND2_X1 U14411 ( .A1(n13359), .A2(n13055), .ZN(n12032) );
  NAND2_X1 U14412 ( .A1(n13214), .A2(n13213), .ZN(n13212) );
  NAND2_X1 U14413 ( .A1(n13349), .A2(n13012), .ZN(n12033) );
  NAND2_X1 U14414 ( .A1(n13212), .A2(n12033), .ZN(n13199) );
  OR2_X1 U14415 ( .A1(n13344), .A2(n13053), .ZN(n12034) );
  NAND2_X1 U14416 ( .A1(n13344), .A2(n13053), .ZN(n12035) );
  NAND2_X1 U14417 ( .A1(n13150), .A2(n13050), .ZN(n12036) );
  OAI222_X1 U14418 ( .A1(n13444), .A2(n14004), .B1(n12042), .B2(P2_U3088), 
        .C1(n12066), .C2(n12041), .ZN(P2_U3297) );
  NOR2_X1 U14419 ( .A1(n12045), .A2(n14349), .ZN(n12051) );
  NAND3_X1 U14420 ( .A1(n12043), .A2(n12044), .A3(n14353), .ZN(n12048) );
  INV_X1 U14421 ( .A(n12045), .ZN(n12046) );
  NAND2_X1 U14422 ( .A1(n12048), .A2(n12047), .ZN(n12050) );
  OAI22_X1 U14423 ( .A1(n13890), .A2(n13493), .B1(n13452), .B2(n13892), .ZN(
        n12053) );
  INV_X1 U14424 ( .A(n12053), .ZN(n12054) );
  NOR2_X2 U14425 ( .A1(n12057), .A2(n12056), .ZN(n13933) );
  AOI21_X1 U14426 ( .B1(n13454), .B2(n13764), .A(n14182), .ZN(n12059) );
  NAND2_X1 U14427 ( .A1(n12059), .A2(n13753), .ZN(n13931) );
  AOI22_X1 U14428 ( .A1(n14284), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13449), 
        .B2(n14285), .ZN(n12061) );
  NAND2_X1 U14429 ( .A1(n13454), .A2(n14306), .ZN(n12060) );
  OAI211_X1 U14430 ( .C1(n13931), .C2(n14160), .A(n12061), .B(n12060), .ZN(
        n12062) );
  INV_X1 U14431 ( .A(n12062), .ZN(n12063) );
  OAI21_X1 U14432 ( .B1(n13933), .B2(n13880), .A(n12063), .ZN(P1_U3266) );
  AOI22_X1 U14433 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n14007), .B1(n12065), 
        .B2(n12064), .ZN(n12092) );
  INV_X1 U14434 ( .A(n12092), .ZN(n12067) );
  INV_X1 U14435 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14879) );
  AOI22_X1 U14436 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(
        P1_DATAO_REG_30__SCAN_IN), .B1(n12066), .B2(n14879), .ZN(n12091) );
  XNOR2_X1 U14437 ( .A(n12067), .B(n12091), .ZN(n12079) );
  INV_X1 U14438 ( .A(n12079), .ZN(n12068) );
  OAI222_X1 U14439 ( .A1(n12069), .A2(P3_U3151), .B1(n12874), .B2(n14880), 
        .C1(n12880), .C2(n12068), .ZN(P3_U3265) );
  INV_X1 U14440 ( .A(n12070), .ZN(n12072) );
  OAI222_X1 U14441 ( .A1(P3_U3151), .A2(n12073), .B1(n12880), .B2(n12072), 
        .C1(n12071), .C2(n12874), .ZN(P3_U3268) );
  AOI22_X1 U14442 ( .A1(n12637), .A2(n12755), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n14772), .ZN(n12074) );
  OAI21_X1 U14443 ( .B1(n12075), .B2(n12757), .A(n12074), .ZN(n12076) );
  AOI21_X1 U14444 ( .B1(n7365), .B2(n12778), .A(n12076), .ZN(n12077) );
  OAI21_X1 U14445 ( .B1(n12078), .B2(n14772), .A(n12077), .ZN(P3_U3204) );
  NAND2_X1 U14446 ( .A1(n8353), .A2(n12079), .ZN(n12081) );
  OR2_X1 U14447 ( .A1(n12096), .A2(n14880), .ZN(n12080) );
  INV_X1 U14448 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12086) );
  NAND2_X1 U14449 ( .A1(n6424), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12085) );
  NAND2_X1 U14450 ( .A1(n12083), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12084) );
  OAI211_X1 U14451 ( .C1(n12087), .C2(n12086), .A(n12085), .B(n12084), .ZN(
        n12088) );
  INV_X1 U14452 ( .A(n12088), .ZN(n12089) );
  INV_X1 U14453 ( .A(n12640), .ZN(n12533) );
  OAI21_X1 U14454 ( .B1(n14091), .B2(n12533), .A(n12292), .ZN(n12099) );
  INV_X1 U14455 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n12093) );
  AOI22_X1 U14456 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(
        P1_DATAO_REG_31__SCAN_IN), .B1(n12094), .B2(n12093), .ZN(n12095) );
  INV_X1 U14457 ( .A(SI_31_), .ZN(n12872) );
  OR2_X1 U14458 ( .A1(n12096), .A2(n12872), .ZN(n12097) );
  OAI22_X1 U14459 ( .A1(n14089), .A2(n12640), .B1(n14091), .B2(n12534), .ZN(
        n12136) );
  AOI211_X1 U14460 ( .C1(n12100), .C2(n12297), .A(n12099), .B(n12136), .ZN(
        n12104) );
  INV_X1 U14461 ( .A(n14089), .ZN(n12643) );
  NOR2_X1 U14462 ( .A1(n12643), .A2(n12533), .ZN(n12299) );
  NAND2_X1 U14463 ( .A1(n12141), .A2(n12669), .ZN(n12285) );
  INV_X1 U14464 ( .A(n12144), .ZN(n12106) );
  INV_X1 U14465 ( .A(n12107), .ZN(n12109) );
  NAND2_X1 U14466 ( .A1(n12109), .A2(n12108), .ZN(n12752) );
  INV_X1 U14467 ( .A(n12752), .ZN(n12131) );
  INV_X1 U14468 ( .A(n12110), .ZN(n12112) );
  NAND2_X1 U14469 ( .A1(n12112), .A2(n12111), .ZN(n12730) );
  INV_X1 U14470 ( .A(n12730), .ZN(n12130) );
  INV_X1 U14471 ( .A(n12777), .ZN(n12257) );
  INV_X1 U14472 ( .A(n12113), .ZN(n12115) );
  NOR4_X1 U14473 ( .A1(n12164), .A2(n12116), .A3(n12115), .A4(n12162), .ZN(
        n12117) );
  NAND2_X1 U14474 ( .A1(n12216), .A2(n12117), .ZN(n12120) );
  NAND4_X1 U14475 ( .A1(n12199), .A2(n12118), .A3(n12186), .A4(n8395), .ZN(
        n12119) );
  NOR4_X1 U14476 ( .A1(n12122), .A2(n12121), .A3(n12120), .A4(n12119), .ZN(
        n12123) );
  NAND4_X1 U14477 ( .A1(n12226), .A2(n12124), .A3(n12232), .A4(n12123), .ZN(
        n12125) );
  NOR3_X1 U14478 ( .A1(n12126), .A2(n12234), .A3(n12125), .ZN(n12128) );
  NAND4_X1 U14479 ( .A1(n12257), .A2(n12128), .A3(n12127), .A4(n12244), .ZN(
        n12129) );
  NOR4_X1 U14480 ( .A1(n12131), .A2(n12130), .A3(n12738), .A4(n12129), .ZN(
        n12132) );
  AND4_X1 U14481 ( .A1(n12721), .A2(n12142), .A3(n12132), .A4(n12695), .ZN(
        n12133) );
  NAND4_X1 U14482 ( .A1(n12445), .A2(n12687), .A3(n12296), .A4(n12133), .ZN(
        n12134) );
  INV_X1 U14483 ( .A(n12136), .ZN(n12300) );
  NAND2_X1 U14484 ( .A1(n12137), .A2(n12300), .ZN(n12138) );
  INV_X1 U14485 ( .A(n12285), .ZN(n12278) );
  INV_X1 U14486 ( .A(n12142), .ZN(n12710) );
  INV_X1 U14487 ( .A(n12143), .ZN(n12145) );
  MUX2_X1 U14488 ( .A(n12145), .B(n12144), .S(n12294), .Z(n12272) );
  INV_X1 U14489 ( .A(n12721), .ZN(n12271) );
  NAND2_X1 U14490 ( .A1(n12541), .A2(n12294), .ZN(n12269) );
  MUX2_X1 U14491 ( .A(n12147), .B(n12146), .S(n12294), .Z(n12266) );
  INV_X1 U14492 ( .A(n12738), .ZN(n12742) );
  OAI211_X1 U14493 ( .C1(n12777), .C2(n12148), .A(n12262), .B(n12151), .ZN(
        n12155) );
  NAND2_X1 U14494 ( .A1(n12150), .A2(n12149), .ZN(n12152) );
  NAND2_X1 U14495 ( .A1(n12152), .A2(n12151), .ZN(n12153) );
  NAND2_X1 U14496 ( .A1(n7355), .A2(n12153), .ZN(n12154) );
  MUX2_X1 U14497 ( .A(n12155), .B(n12154), .S(n12288), .Z(n12156) );
  INV_X1 U14498 ( .A(n12156), .ZN(n12261) );
  INV_X1 U14499 ( .A(n12165), .ZN(n12160) );
  NOR2_X1 U14500 ( .A1(n12157), .A2(n12310), .ZN(n12158) );
  AOI21_X1 U14501 ( .B1(n9718), .B2(n12158), .A(n12163), .ZN(n12159) );
  OAI22_X1 U14502 ( .A1(n12162), .A2(n12161), .B1(n12160), .B2(n12159), .ZN(
        n12170) );
  NAND2_X1 U14503 ( .A1(n12164), .A2(n12163), .ZN(n12169) );
  MUX2_X1 U14504 ( .A(n12166), .B(n12165), .S(n12288), .Z(n12167) );
  NAND2_X1 U14505 ( .A1(n12167), .A2(n14758), .ZN(n12168) );
  AOI21_X1 U14506 ( .B1(n12170), .B2(n12169), .A(n12168), .ZN(n12173) );
  AOI21_X1 U14507 ( .B1(n12179), .B2(n12171), .A(n12294), .ZN(n12172) );
  AOI21_X1 U14508 ( .B1(n12176), .B2(n12174), .A(n12288), .ZN(n12175) );
  OAI21_X1 U14509 ( .B1(n12288), .B2(n12179), .A(n12178), .ZN(n12187) );
  NAND2_X1 U14510 ( .A1(n12180), .A2(n12294), .ZN(n12184) );
  NAND2_X1 U14511 ( .A1(n12181), .A2(n12288), .ZN(n12183) );
  MUX2_X1 U14512 ( .A(n12184), .B(n12183), .S(n12182), .Z(n12185) );
  OAI211_X1 U14513 ( .C1(n12188), .C2(n12187), .A(n12186), .B(n12185), .ZN(
        n12195) );
  NAND2_X1 U14514 ( .A1(n12196), .A2(n12189), .ZN(n12192) );
  NAND2_X1 U14515 ( .A1(n12197), .A2(n12190), .ZN(n12191) );
  MUX2_X1 U14516 ( .A(n12192), .B(n12191), .S(n12288), .Z(n12193) );
  INV_X1 U14517 ( .A(n12193), .ZN(n12194) );
  NAND2_X1 U14518 ( .A1(n12195), .A2(n12194), .ZN(n12200) );
  MUX2_X1 U14519 ( .A(n12197), .B(n12196), .S(n12288), .Z(n12198) );
  NAND3_X1 U14520 ( .A1(n12200), .A2(n12199), .A3(n12198), .ZN(n12206) );
  OR2_X1 U14521 ( .A1(n12201), .A2(n12294), .ZN(n12203) );
  NAND2_X1 U14522 ( .A1(n12201), .A2(n12294), .ZN(n12202) );
  MUX2_X1 U14523 ( .A(n12203), .B(n12202), .S(n12553), .Z(n12204) );
  NAND3_X1 U14524 ( .A1(n12206), .A2(n12205), .A3(n12204), .ZN(n12212) );
  NAND2_X1 U14525 ( .A1(n12551), .A2(n12288), .ZN(n12210) );
  NAND2_X1 U14526 ( .A1(n12207), .A2(n12294), .ZN(n12209) );
  MUX2_X1 U14527 ( .A(n12210), .B(n12209), .S(n12208), .Z(n12211) );
  NAND3_X1 U14528 ( .A1(n12212), .A2(n8395), .A3(n12211), .ZN(n12217) );
  MUX2_X1 U14529 ( .A(n12214), .B(n12213), .S(n12288), .Z(n12215) );
  NAND4_X1 U14530 ( .A1(n12217), .A2(n12216), .A3(n12226), .A4(n12215), .ZN(
        n12224) );
  INV_X1 U14531 ( .A(n12218), .ZN(n12219) );
  NAND2_X1 U14532 ( .A1(n12226), .A2(n12219), .ZN(n12221) );
  NAND3_X1 U14533 ( .A1(n12221), .A2(n12233), .A3(n12220), .ZN(n12222) );
  NAND2_X1 U14534 ( .A1(n12222), .A2(n12294), .ZN(n12223) );
  NAND2_X1 U14535 ( .A1(n12224), .A2(n12223), .ZN(n12231) );
  NAND2_X1 U14536 ( .A1(n12226), .A2(n6806), .ZN(n12228) );
  NAND3_X1 U14537 ( .A1(n12228), .A2(n12227), .A3(n12230), .ZN(n12229) );
  AOI22_X1 U14538 ( .A1(n12231), .A2(n12230), .B1(n12288), .B2(n12229), .ZN(
        n12239) );
  OAI21_X1 U14539 ( .B1(n12233), .B2(n12294), .A(n12232), .ZN(n12238) );
  MUX2_X1 U14540 ( .A(n12236), .B(n12235), .S(n12288), .Z(n12237) );
  OAI211_X1 U14541 ( .C1(n12239), .C2(n12238), .A(n6825), .B(n12237), .ZN(
        n12243) );
  MUX2_X1 U14542 ( .A(n12241), .B(n12240), .S(n12294), .Z(n12242) );
  NAND2_X1 U14543 ( .A1(n12243), .A2(n12242), .ZN(n12245) );
  NAND2_X1 U14544 ( .A1(n12245), .A2(n12244), .ZN(n12250) );
  OAI22_X1 U14545 ( .A1(n12254), .A2(n12476), .B1(n12247), .B2(n12246), .ZN(
        n12248) );
  NAND2_X1 U14546 ( .A1(n12248), .A2(n12294), .ZN(n12249) );
  AOI21_X1 U14547 ( .B1(n12252), .B2(n12251), .A(n12294), .ZN(n12255) );
  NAND2_X1 U14548 ( .A1(n12544), .A2(n12288), .ZN(n12253) );
  OAI22_X1 U14549 ( .A1(n12256), .A2(n12255), .B1(n12254), .B2(n12253), .ZN(
        n12259) );
  NAND3_X1 U14550 ( .A1(n12259), .A2(n12258), .A3(n12257), .ZN(n12260) );
  NAND2_X1 U14551 ( .A1(n12261), .A2(n12260), .ZN(n12264) );
  MUX2_X1 U14552 ( .A(n7355), .B(n12262), .S(n12288), .Z(n12263) );
  NAND3_X1 U14553 ( .A1(n12742), .A2(n12264), .A3(n12263), .ZN(n12265) );
  NAND3_X1 U14554 ( .A1(n12266), .A2(n12265), .A3(n12730), .ZN(n12268) );
  NAND3_X1 U14555 ( .A1(n12460), .A2(n12396), .A3(n12288), .ZN(n12267) );
  OAI211_X1 U14556 ( .C1(n12460), .C2(n12269), .A(n12268), .B(n12267), .ZN(
        n12270) );
  XNOR2_X1 U14557 ( .A(n12273), .B(n12288), .ZN(n12274) );
  NAND2_X1 U14558 ( .A1(n12279), .A2(n12536), .ZN(n12280) );
  NAND2_X1 U14559 ( .A1(n7177), .A2(n12282), .ZN(n12284) );
  INV_X1 U14560 ( .A(n12286), .ZN(n12287) );
  NAND3_X1 U14561 ( .A1(n12289), .A2(n12288), .A3(n12287), .ZN(n12290) );
  OAI211_X1 U14562 ( .C1(n12295), .C2(n12294), .A(n12293), .B(n12292), .ZN(
        n12298) );
  NAND3_X1 U14563 ( .A1(n12298), .A2(n12297), .A3(n12296), .ZN(n12301) );
  AOI21_X1 U14564 ( .B1(n12301), .B2(n12300), .A(n12299), .ZN(n12304) );
  NOR2_X1 U14565 ( .A1(n12304), .A2(n12302), .ZN(n12306) );
  NOR4_X1 U14566 ( .A1(n14762), .A2(n12309), .A3(n12308), .A4(n6630), .ZN(
        n12312) );
  OAI21_X1 U14567 ( .B1(n12313), .B2(n12310), .A(P3_B_REG_SCAN_IN), .ZN(n12311) );
  NAND2_X1 U14568 ( .A1(n12315), .A2(n12314), .ZN(n12316) );
  AOI22_X1 U14569 ( .A1(n13965), .A2(n12363), .B1(n12365), .B2(n13828), .ZN(
        n12318) );
  XNOR2_X1 U14570 ( .A(n12318), .B(n12366), .ZN(n12320) );
  AOI22_X1 U14571 ( .A1(n13965), .A2(n12365), .B1(n12364), .B2(n13828), .ZN(
        n12319) );
  XNOR2_X1 U14572 ( .A(n12320), .B(n12319), .ZN(n13483) );
  NAND2_X1 U14573 ( .A1(n12320), .A2(n12319), .ZN(n12321) );
  NAND2_X1 U14574 ( .A1(n13960), .A2(n12363), .ZN(n12323) );
  NAND2_X1 U14575 ( .A1(n12365), .A2(n13583), .ZN(n12322) );
  NAND2_X1 U14576 ( .A1(n12323), .A2(n12322), .ZN(n12324) );
  XNOR2_X1 U14577 ( .A(n12324), .B(n12366), .ZN(n12325) );
  AOI22_X1 U14578 ( .A1(n13960), .A2(n12365), .B1(n12364), .B2(n13583), .ZN(
        n12326) );
  XNOR2_X1 U14579 ( .A(n12325), .B(n12326), .ZN(n13527) );
  INV_X1 U14580 ( .A(n12325), .ZN(n12327) );
  NAND2_X1 U14581 ( .A1(n12327), .A2(n12326), .ZN(n12328) );
  NAND2_X1 U14582 ( .A1(n13952), .A2(n12363), .ZN(n12330) );
  NAND2_X1 U14583 ( .A1(n12365), .A2(n13827), .ZN(n12329) );
  NAND2_X1 U14584 ( .A1(n12330), .A2(n12329), .ZN(n12331) );
  XNOR2_X1 U14585 ( .A(n12331), .B(n12366), .ZN(n12332) );
  AOI22_X1 U14586 ( .A1(n13952), .A2(n12365), .B1(n12364), .B2(n13827), .ZN(
        n12333) );
  XNOR2_X1 U14587 ( .A(n12332), .B(n12333), .ZN(n13458) );
  INV_X1 U14588 ( .A(n12332), .ZN(n12334) );
  NAND2_X1 U14589 ( .A1(n13805), .A2(n12363), .ZN(n12336) );
  NAND2_X1 U14590 ( .A1(n12365), .A2(n13779), .ZN(n12335) );
  NAND2_X1 U14591 ( .A1(n12336), .A2(n12335), .ZN(n12337) );
  XNOR2_X1 U14592 ( .A(n12337), .B(n12366), .ZN(n12338) );
  AOI22_X1 U14593 ( .A1(n13805), .A2(n12365), .B1(n12364), .B2(n13779), .ZN(
        n12339) );
  XNOR2_X1 U14594 ( .A(n12338), .B(n12339), .ZN(n13518) );
  NAND2_X1 U14595 ( .A1(n13517), .A2(n13518), .ZN(n12342) );
  INV_X1 U14596 ( .A(n12338), .ZN(n12340) );
  NAND2_X1 U14597 ( .A1(n12340), .A2(n12339), .ZN(n12341) );
  NAND2_X1 U14598 ( .A1(n12342), .A2(n12341), .ZN(n13489) );
  NAND2_X1 U14599 ( .A1(n13942), .A2(n12363), .ZN(n12344) );
  NAND2_X1 U14600 ( .A1(n12365), .A2(n13799), .ZN(n12343) );
  NAND2_X1 U14601 ( .A1(n12344), .A2(n12343), .ZN(n12345) );
  XNOR2_X1 U14602 ( .A(n12345), .B(n12366), .ZN(n12346) );
  AOI22_X1 U14603 ( .A1(n13942), .A2(n12365), .B1(n12364), .B2(n13799), .ZN(
        n12347) );
  XNOR2_X1 U14604 ( .A(n12346), .B(n12347), .ZN(n13490) );
  INV_X1 U14605 ( .A(n12346), .ZN(n12348) );
  NAND2_X1 U14606 ( .A1(n12348), .A2(n12347), .ZN(n12349) );
  NAND2_X1 U14607 ( .A1(n13562), .A2(n12363), .ZN(n12351) );
  NAND2_X1 U14608 ( .A1(n12365), .A2(n13778), .ZN(n12350) );
  NAND2_X1 U14609 ( .A1(n12351), .A2(n12350), .ZN(n12352) );
  XNOR2_X1 U14610 ( .A(n12352), .B(n12366), .ZN(n12353) );
  AOI22_X1 U14611 ( .A1(n13562), .A2(n12365), .B1(n12364), .B2(n13778), .ZN(
        n12354) );
  XNOR2_X1 U14612 ( .A(n12353), .B(n12354), .ZN(n13556) );
  INV_X1 U14613 ( .A(n12353), .ZN(n12355) );
  NAND2_X1 U14614 ( .A1(n13454), .A2(n12363), .ZN(n12358) );
  NAND2_X1 U14615 ( .A1(n12365), .A2(n13765), .ZN(n12357) );
  NAND2_X1 U14616 ( .A1(n12358), .A2(n12357), .ZN(n12359) );
  XNOR2_X1 U14617 ( .A(n12359), .B(n12366), .ZN(n12360) );
  AOI22_X1 U14618 ( .A1(n13454), .A2(n12365), .B1(n12364), .B2(n13765), .ZN(
        n12361) );
  XNOR2_X1 U14619 ( .A(n12360), .B(n12361), .ZN(n13448) );
  INV_X1 U14620 ( .A(n12360), .ZN(n12362) );
  AOI22_X1 U14621 ( .A1(n13927), .A2(n12363), .B1(n12365), .B2(n13582), .ZN(
        n12369) );
  AOI22_X1 U14622 ( .A1(n13927), .A2(n12365), .B1(n12364), .B2(n13582), .ZN(
        n12367) );
  XNOR2_X1 U14623 ( .A(n12367), .B(n12366), .ZN(n12368) );
  XOR2_X1 U14624 ( .A(n12369), .B(n12368), .Z(n12370) );
  XNOR2_X1 U14625 ( .A(n12371), .B(n12370), .ZN(n12379) );
  INV_X1 U14626 ( .A(n13748), .ZN(n12376) );
  OR2_X1 U14627 ( .A1(n12372), .A2(n13892), .ZN(n12374) );
  NAND2_X1 U14628 ( .A1(n14131), .A2(n13765), .ZN(n12373) );
  NAND2_X1 U14629 ( .A1(n12374), .A2(n12373), .ZN(n13926) );
  AOI22_X1 U14630 ( .A1(n14141), .A2(n13926), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12375) );
  OAI21_X1 U14631 ( .B1(n12376), .B2(n14146), .A(n12375), .ZN(n12377) );
  AOI21_X1 U14632 ( .B1(n13927), .B2(n14142), .A(n12377), .ZN(n12378) );
  OAI21_X1 U14633 ( .B1(n12379), .B2(n13564), .A(n12378), .ZN(P1_U3220) );
  OAI222_X1 U14634 ( .A1(n14012), .A2(n12382), .B1(n14014), .B2(n12381), .C1(
        P1_U3086), .C2(n12380), .ZN(P1_U3334) );
  XNOR2_X1 U14635 ( .A(n12781), .B(n12444), .ZN(n12441) );
  XNOR2_X1 U14636 ( .A(n12441), .B(n12536), .ZN(n12442) );
  XNOR2_X1 U14637 ( .A(n12857), .B(n12444), .ZN(n12391) );
  INV_X1 U14638 ( .A(n12391), .ZN(n12392) );
  XNOR2_X1 U14639 ( .A(n12385), .B(n12444), .ZN(n12387) );
  XNOR2_X1 U14640 ( .A(n12387), .B(n12764), .ZN(n12473) );
  NAND2_X1 U14641 ( .A1(n12474), .A2(n12473), .ZN(n12472) );
  NAND2_X1 U14642 ( .A1(n12472), .A2(n12388), .ZN(n12512) );
  XNOR2_X1 U14643 ( .A(n12774), .B(n12444), .ZN(n12389) );
  XNOR2_X1 U14644 ( .A(n12389), .B(n12543), .ZN(n12511) );
  NAND2_X1 U14645 ( .A1(n12512), .A2(n12511), .ZN(n12510) );
  NAND2_X1 U14646 ( .A1(n12510), .A2(n12390), .ZN(n12437) );
  XNOR2_X1 U14647 ( .A(n12391), .B(n12514), .ZN(n12436) );
  XNOR2_X1 U14648 ( .A(n12853), .B(n12444), .ZN(n12393) );
  XNOR2_X1 U14649 ( .A(n12393), .B(n12394), .ZN(n12495) );
  NAND2_X1 U14650 ( .A1(n12393), .A2(n12542), .ZN(n12395) );
  XNOR2_X1 U14651 ( .A(n12460), .B(n12444), .ZN(n12397) );
  XNOR2_X1 U14652 ( .A(n12397), .B(n12396), .ZN(n12457) );
  XNOR2_X1 U14653 ( .A(n12845), .B(n12444), .ZN(n12399) );
  INV_X1 U14654 ( .A(n12399), .ZN(n12400) );
  NAND2_X1 U14655 ( .A1(n7327), .A2(n12400), .ZN(n12401) );
  OAI21_X2 U14656 ( .B1(n12501), .B2(n12540), .A(n12401), .ZN(n12404) );
  XNOR2_X1 U14657 ( .A(n12842), .B(n12444), .ZN(n12402) );
  XNOR2_X1 U14658 ( .A(n12404), .B(n12402), .ZN(n12427) );
  NAND2_X1 U14659 ( .A1(n12427), .A2(n12487), .ZN(n12406) );
  INV_X1 U14660 ( .A(n12402), .ZN(n12403) );
  NAND2_X1 U14661 ( .A1(n12404), .A2(n12403), .ZN(n12405) );
  NAND2_X1 U14662 ( .A1(n12406), .A2(n12405), .ZN(n12484) );
  XNOR2_X1 U14663 ( .A(n12491), .B(n12444), .ZN(n12408) );
  XNOR2_X1 U14664 ( .A(n12408), .B(n12538), .ZN(n12486) );
  NAND2_X1 U14665 ( .A1(n12484), .A2(n12486), .ZN(n12410) );
  NAND2_X1 U14666 ( .A1(n12408), .A2(n12407), .ZN(n12409) );
  NAND2_X1 U14667 ( .A1(n12410), .A2(n12409), .ZN(n12464) );
  XNOR2_X1 U14668 ( .A(n12834), .B(n12444), .ZN(n12411) );
  XNOR2_X1 U14669 ( .A(n12411), .B(n12670), .ZN(n12465) );
  NAND2_X1 U14670 ( .A1(n12464), .A2(n12465), .ZN(n12414) );
  INV_X1 U14671 ( .A(n12411), .ZN(n12412) );
  NAND2_X1 U14672 ( .A1(n12412), .A2(n12670), .ZN(n12413) );
  NAND2_X1 U14673 ( .A1(n12414), .A2(n12413), .ZN(n12519) );
  XNOR2_X1 U14674 ( .A(n12529), .B(n12444), .ZN(n12416) );
  XNOR2_X1 U14675 ( .A(n12416), .B(n12537), .ZN(n12521) );
  NAND2_X1 U14676 ( .A1(n12519), .A2(n12521), .ZN(n12418) );
  NAND2_X1 U14677 ( .A1(n12416), .A2(n12415), .ZN(n12417) );
  XOR2_X1 U14678 ( .A(n12442), .B(n12443), .Z(n12426) );
  OR2_X1 U14679 ( .A1(n12419), .A2(n14760), .ZN(n12421) );
  NAND2_X1 U14680 ( .A1(n12537), .A2(n12763), .ZN(n12420) );
  NAND2_X1 U14681 ( .A1(n12421), .A2(n12420), .ZN(n12657) );
  INV_X1 U14682 ( .A(n12657), .ZN(n12423) );
  AOI22_X1 U14683 ( .A1(n12659), .A2(n12523), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12422) );
  OAI21_X1 U14684 ( .B1(n12423), .B2(n12503), .A(n12422), .ZN(n12424) );
  AOI21_X1 U14685 ( .B1(n12781), .B2(n12528), .A(n12424), .ZN(n12425) );
  OAI21_X1 U14686 ( .B1(n12426), .B2(n12531), .A(n12425), .ZN(P3_U3154) );
  XNOR2_X1 U14687 ( .A(n12427), .B(n12539), .ZN(n12434) );
  NOR2_X1 U14688 ( .A1(n12500), .A2(n14762), .ZN(n12428) );
  AOI21_X1 U14689 ( .B1(n12538), .B2(n12765), .A(n12428), .ZN(n12707) );
  NAND2_X1 U14690 ( .A1(P3_U3151), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n12430)
         );
  NAND2_X1 U14691 ( .A1(n12523), .A2(n12712), .ZN(n12429) );
  OAI211_X1 U14692 ( .C1(n12707), .C2(n12503), .A(n12430), .B(n12429), .ZN(
        n12431) );
  AOI21_X1 U14693 ( .B1(n12432), .B2(n12528), .A(n12431), .ZN(n12433) );
  OAI21_X1 U14694 ( .B1(n12434), .B2(n12531), .A(n12433), .ZN(P3_U3156) );
  OAI211_X1 U14695 ( .C1(n12437), .C2(n12436), .A(n12435), .B(n12509), .ZN(
        n12440) );
  AOI22_X1 U14696 ( .A1(n12543), .A2(n12763), .B1(n12765), .B2(n12542), .ZN(
        n12750) );
  NAND2_X1 U14697 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12626)
         );
  OAI21_X1 U14698 ( .B1(n12750), .B2(n12503), .A(n12626), .ZN(n12438) );
  AOI21_X1 U14699 ( .B1(n12754), .B2(n12523), .A(n12438), .ZN(n12439) );
  OAI211_X1 U14700 ( .C1(n12518), .C2(n12857), .A(n12440), .B(n12439), .ZN(
        P3_U3159) );
  AOI22_X1 U14701 ( .A1(n12443), .A2(n12442), .B1(n12671), .B2(n12441), .ZN(
        n12447) );
  XNOR2_X1 U14702 ( .A(n12445), .B(n12444), .ZN(n12446) );
  XNOR2_X1 U14703 ( .A(n12447), .B(n12446), .ZN(n12455) );
  INV_X1 U14704 ( .A(n12448), .ZN(n12648) );
  OAI22_X1 U14705 ( .A1(n12648), .A2(n12450), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12449), .ZN(n12453) );
  OAI22_X1 U14706 ( .A1(n12451), .A2(n12526), .B1(n12671), .B2(n12475), .ZN(
        n12452) );
  AOI211_X1 U14707 ( .C1(n12652), .C2(n12528), .A(n12453), .B(n12452), .ZN(
        n12454) );
  OAI21_X1 U14708 ( .B1(n12455), .B2(n12531), .A(n12454), .ZN(P3_U3160) );
  AOI21_X1 U14709 ( .B1(n12457), .B2(n12456), .A(n6581), .ZN(n12463) );
  AOI22_X1 U14710 ( .A1(n12540), .A2(n12765), .B1(n12763), .B2(n12542), .ZN(
        n12728) );
  OAI22_X1 U14711 ( .A1(n12728), .A2(n12503), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12458), .ZN(n12459) );
  AOI21_X1 U14712 ( .B1(n12732), .B2(n12523), .A(n12459), .ZN(n12462) );
  NAND2_X1 U14713 ( .A1(n12460), .A2(n12528), .ZN(n12461) );
  OAI211_X1 U14714 ( .C1(n12463), .C2(n12531), .A(n12462), .B(n12461), .ZN(
        P3_U3163) );
  XOR2_X1 U14715 ( .A(n12465), .B(n12464), .Z(n12471) );
  AND2_X1 U14716 ( .A1(n12538), .A2(n12763), .ZN(n12466) );
  AOI21_X1 U14717 ( .B1(n12537), .B2(n12765), .A(n12466), .ZN(n12684) );
  AOI22_X1 U14718 ( .A1(n12689), .A2(n12523), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12467) );
  OAI21_X1 U14719 ( .B1(n12684), .B2(n12503), .A(n12467), .ZN(n12468) );
  AOI21_X1 U14720 ( .B1(n12469), .B2(n12528), .A(n12468), .ZN(n12470) );
  OAI21_X1 U14721 ( .B1(n12471), .B2(n12531), .A(n12470), .ZN(P3_U3165) );
  OAI211_X1 U14722 ( .C1(n12474), .C2(n12473), .A(n12472), .B(n12509), .ZN(
        n12483) );
  NOR2_X1 U14723 ( .A1(n12476), .A2(n12475), .ZN(n12480) );
  OAI22_X1 U14724 ( .A1(n12478), .A2(n12526), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12477), .ZN(n12479) );
  AOI211_X1 U14725 ( .C1(n12481), .C2(n12523), .A(n12480), .B(n12479), .ZN(
        n12482) );
  OAI211_X1 U14726 ( .C1(n12866), .C2(n12518), .A(n12483), .B(n12482), .ZN(
        P3_U3168) );
  XOR2_X1 U14727 ( .A(n12486), .B(n12485), .Z(n12493) );
  NOR2_X1 U14728 ( .A1(n12487), .A2(n14762), .ZN(n12488) );
  AOI21_X1 U14729 ( .B1(n7178), .B2(n12765), .A(n12488), .ZN(n12698) );
  AOI22_X1 U14730 ( .A1(n12702), .A2(n12523), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12489) );
  OAI21_X1 U14731 ( .B1(n12698), .B2(n12503), .A(n12489), .ZN(n12490) );
  AOI21_X1 U14732 ( .B1(n12491), .B2(n12528), .A(n12490), .ZN(n12492) );
  OAI21_X1 U14733 ( .B1(n12493), .B2(n12531), .A(n12492), .ZN(P3_U3169) );
  OAI211_X1 U14734 ( .C1(n12496), .C2(n12495), .A(n12494), .B(n12509), .ZN(
        n12499) );
  AOI22_X1 U14735 ( .A1(n12766), .A2(n12763), .B1(n12541), .B2(n12765), .ZN(
        n12740) );
  OAI22_X1 U14736 ( .A1(n12740), .A2(n12503), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14920), .ZN(n12497) );
  AOI21_X1 U14737 ( .B1(n12744), .B2(n12523), .A(n12497), .ZN(n12498) );
  OAI211_X1 U14738 ( .C1(n12853), .C2(n12518), .A(n12499), .B(n12498), .ZN(
        P3_U3173) );
  XNOR2_X1 U14739 ( .A(n12501), .B(n12500), .ZN(n12508) );
  AOI22_X1 U14740 ( .A1(n12539), .A2(n12765), .B1(n12763), .B2(n12541), .ZN(
        n12718) );
  INV_X1 U14741 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n12502) );
  OAI22_X1 U14742 ( .A1(n12718), .A2(n12503), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12502), .ZN(n12504) );
  AOI21_X1 U14743 ( .B1(n12722), .B2(n12523), .A(n12504), .ZN(n12507) );
  NAND2_X1 U14744 ( .A1(n12505), .A2(n12528), .ZN(n12506) );
  OAI211_X1 U14745 ( .C1(n12508), .C2(n12531), .A(n12507), .B(n12506), .ZN(
        P3_U3175) );
  INV_X1 U14746 ( .A(n12774), .ZN(n12861) );
  OAI211_X1 U14747 ( .C1(n12512), .C2(n12511), .A(n12510), .B(n12509), .ZN(
        n12517) );
  NAND2_X1 U14748 ( .A1(n12764), .A2(n12522), .ZN(n12513) );
  NAND2_X1 U14749 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12590)
         );
  OAI211_X1 U14750 ( .C1(n12514), .C2(n12526), .A(n12513), .B(n12590), .ZN(
        n12515) );
  AOI21_X1 U14751 ( .B1(n12769), .B2(n12523), .A(n12515), .ZN(n12516) );
  OAI211_X1 U14752 ( .C1(n12861), .C2(n12518), .A(n12517), .B(n12516), .ZN(
        P3_U3178) );
  XOR2_X1 U14753 ( .A(n12521), .B(n12520), .Z(n12532) );
  AOI22_X1 U14754 ( .A1(n7178), .A2(n12522), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12525) );
  NAND2_X1 U14755 ( .A1(n12675), .A2(n12523), .ZN(n12524) );
  OAI211_X1 U14756 ( .C1(n12671), .C2(n12526), .A(n12525), .B(n12524), .ZN(
        n12527) );
  AOI21_X1 U14757 ( .B1(n12529), .B2(n12528), .A(n12527), .ZN(n12530) );
  OAI21_X1 U14758 ( .B1(n12532), .B2(n12531), .A(n12530), .ZN(P3_U3180) );
  MUX2_X1 U14759 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12533), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14760 ( .A(n12534), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12552), .Z(
        P3_U3521) );
  MUX2_X1 U14761 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12535), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14762 ( .A(n12536), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12552), .Z(
        P3_U3518) );
  MUX2_X1 U14763 ( .A(n12537), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12552), .Z(
        P3_U3517) );
  MUX2_X1 U14764 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n7178), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14765 ( .A(n12538), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12552), .Z(
        P3_U3515) );
  MUX2_X1 U14766 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12539), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14767 ( .A(n12540), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12552), .Z(
        P3_U3513) );
  MUX2_X1 U14768 ( .A(n12541), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12552), .Z(
        P3_U3512) );
  MUX2_X1 U14769 ( .A(n12542), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12552), .Z(
        P3_U3511) );
  MUX2_X1 U14770 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12766), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14771 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12543), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14772 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12764), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14773 ( .A(n12544), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12552), .Z(
        P3_U3507) );
  MUX2_X1 U14774 ( .A(n12545), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12552), .Z(
        P3_U3505) );
  MUX2_X1 U14775 ( .A(n12546), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12552), .Z(
        P3_U3504) );
  MUX2_X1 U14776 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12547), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14777 ( .A(n12548), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12552), .Z(
        P3_U3502) );
  MUX2_X1 U14778 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12549), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14779 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12550), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14780 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12551), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14781 ( .A(n12553), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12552), .Z(
        P3_U3498) );
  MUX2_X1 U14782 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12554), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14783 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12555), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14784 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12556), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14785 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n10201), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14786 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12557), .S(P3_U3897), .Z(
        P3_U3492) );
  AOI21_X2 U14787 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n12561), .A(n12558), 
        .ZN(n12604) );
  XNOR2_X1 U14788 ( .A(n12604), .B(n12605), .ZN(n12559) );
  AOI21_X1 U14789 ( .B1(n12560), .B2(n12559), .A(n12606), .ZN(n12582) );
  NAND2_X1 U14790 ( .A1(n12561), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12566) );
  NAND2_X1 U14791 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12563), .ZN(n12594) );
  OAI21_X1 U14792 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12563), .A(n12594), 
        .ZN(n12580) );
  NOR2_X1 U14793 ( .A1(n12565), .A2(n12564), .ZN(n12568) );
  INV_X1 U14794 ( .A(n12566), .ZN(n12567) );
  MUX2_X1 U14795 ( .A(n12568), .B(n12567), .S(n12073), .Z(n12569) );
  XNOR2_X1 U14796 ( .A(n12571), .B(n12593), .ZN(n12573) );
  MUX2_X1 U14797 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12073), .Z(n12572) );
  NOR2_X1 U14798 ( .A1(n12573), .A2(n12572), .ZN(n12583) );
  AOI21_X1 U14799 ( .B1(n12573), .B2(n12572), .A(n12583), .ZN(n12578) );
  AND2_X1 U14800 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12576) );
  NOR2_X1 U14801 ( .A1(n14727), .A2(n12574), .ZN(n12575) );
  AOI211_X1 U14802 ( .C1(n14718), .C2(n12605), .A(n12576), .B(n12575), .ZN(
        n12577) );
  OAI21_X1 U14803 ( .B1(n12578), .B2(n14709), .A(n12577), .ZN(n12579) );
  AOI21_X1 U14804 ( .B1(n14746), .B2(n12580), .A(n12579), .ZN(n12581) );
  OAI21_X1 U14805 ( .B1(n12582), .B2(n14750), .A(n12581), .ZN(P3_U3197) );
  MUX2_X1 U14806 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12073), .Z(n12589) );
  MUX2_X1 U14807 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12073), .Z(n12587) );
  AOI21_X1 U14808 ( .B1(n12584), .B2(n12605), .A(n12583), .ZN(n14059) );
  MUX2_X1 U14809 ( .A(n12585), .B(n12591), .S(n12073), .Z(n12586) );
  NOR2_X1 U14810 ( .A1(n12586), .A2(n14054), .ZN(n14055) );
  NAND2_X1 U14811 ( .A1(n12586), .A2(n14054), .ZN(n14056) );
  OAI21_X1 U14812 ( .B1(n14059), .B2(n14055), .A(n14056), .ZN(n14075) );
  XNOR2_X1 U14813 ( .A(n12587), .B(n14025), .ZN(n14076) );
  NOR2_X1 U14814 ( .A1(n14075), .A2(n14076), .ZN(n14074) );
  AOI21_X1 U14815 ( .B1(n12589), .B2(n12588), .A(n12627), .ZN(n12617) );
  INV_X1 U14816 ( .A(n14041), .ZN(n12628) );
  OAI21_X1 U14817 ( .B1(n14727), .B2(n9487), .A(n12590), .ZN(n12603) );
  NAND2_X1 U14818 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12609), .ZN(n12596) );
  AOI22_X1 U14819 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12609), .B1(n14054), 
        .B2(n12591), .ZN(n14062) );
  NAND2_X1 U14820 ( .A1(n12593), .A2(n12592), .ZN(n12595) );
  NAND2_X1 U14821 ( .A1(n12595), .A2(n12594), .ZN(n14061) );
  NAND2_X1 U14822 ( .A1(n14062), .A2(n14061), .ZN(n14060) );
  NAND2_X1 U14823 ( .A1(n12596), .A2(n14060), .ZN(n12597) );
  XNOR2_X1 U14824 ( .A(n14071), .B(n12597), .ZN(n14073) );
  NAND2_X1 U14825 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14073), .ZN(n14072) );
  NAND2_X1 U14826 ( .A1(n12597), .A2(n14025), .ZN(n12598) );
  XNOR2_X1 U14827 ( .A(n14041), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n12599) );
  INV_X1 U14828 ( .A(n12622), .ZN(n12601) );
  NAND3_X1 U14829 ( .A1(n14072), .A2(n12599), .A3(n12598), .ZN(n12600) );
  INV_X1 U14830 ( .A(n14746), .ZN(n14607) );
  AOI21_X1 U14831 ( .B1(n12601), .B2(n12600), .A(n14607), .ZN(n12602) );
  AOI211_X1 U14832 ( .C1(n14718), .C2(n12628), .A(n12603), .B(n12602), .ZN(
        n12616) );
  NOR2_X1 U14833 ( .A1(n12605), .A2(n12604), .ZN(n12607) );
  NAND2_X1 U14834 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12609), .ZN(n12608) );
  OAI21_X1 U14835 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n12609), .A(n12608), 
        .ZN(n14065) );
  OR2_X2 U14836 ( .A1(n14081), .A2(n14082), .ZN(n14079) );
  OR2_X1 U14837 ( .A1(n12610), .A2(n14071), .ZN(n12613) );
  NAND2_X1 U14838 ( .A1(n14041), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12618) );
  OR2_X1 U14839 ( .A1(n14041), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12611) );
  NAND2_X1 U14840 ( .A1(n12618), .A2(n12611), .ZN(n12612) );
  AOI21_X1 U14841 ( .B1(n14079), .B2(n12613), .A(n12612), .ZN(n12620) );
  AND3_X1 U14842 ( .A1(n14079), .A2(n12613), .A3(n12612), .ZN(n12614) );
  OAI21_X1 U14843 ( .B1(n12620), .B2(n12614), .A(n14080), .ZN(n12615) );
  OAI211_X1 U14844 ( .C1(n12617), .C2(n14709), .A(n12616), .B(n12615), .ZN(
        P3_U3200) );
  INV_X1 U14845 ( .A(n12618), .ZN(n12619) );
  NOR2_X1 U14846 ( .A1(n12620), .A2(n12619), .ZN(n12621) );
  XNOR2_X1 U14847 ( .A(n12623), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12630) );
  XNOR2_X1 U14848 ( .A(n12621), .B(n12630), .ZN(n12636) );
  XNOR2_X1 U14849 ( .A(n12623), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12629) );
  INV_X1 U14850 ( .A(n12629), .ZN(n12624) );
  NAND2_X1 U14851 ( .A1(n14743), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12625) );
  OAI211_X1 U14852 ( .C1(n14740), .C2(n12105), .A(n12626), .B(n12625), .ZN(
        n12634) );
  MUX2_X1 U14853 ( .A(n12630), .B(n12629), .S(n12073), .Z(n12631) );
  XNOR2_X1 U14854 ( .A(n12632), .B(n12631), .ZN(n12633) );
  OAI21_X1 U14855 ( .B1(n12636), .B2(n14750), .A(n12635), .ZN(P3_U3201) );
  NAND2_X1 U14856 ( .A1(n12637), .A2(n12755), .ZN(n12641) );
  INV_X1 U14857 ( .A(n12638), .ZN(n12639) );
  AOI21_X1 U14858 ( .B1(n12641), .B2(n14088), .A(n14772), .ZN(n12646) );
  AOI21_X1 U14859 ( .B1(n14772), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12646), 
        .ZN(n12642) );
  OAI21_X1 U14860 ( .B1(n12643), .B2(n12757), .A(n12642), .ZN(P3_U3202) );
  OAI22_X1 U14861 ( .A1(n12644), .A2(n14770), .B1(n12757), .B2(n14091), .ZN(
        n12645) );
  OR2_X1 U14862 ( .A1(n12646), .A2(n12645), .ZN(P3_U3203) );
  OAI22_X1 U14863 ( .A1(n12648), .A2(n14755), .B1(n14770), .B2(n12647), .ZN(
        n12651) );
  NOR2_X1 U14864 ( .A1(n12649), .A2(n12663), .ZN(n12650) );
  AOI211_X1 U14865 ( .C1(n12773), .C2(n12652), .A(n12651), .B(n12650), .ZN(
        n12653) );
  OAI21_X1 U14866 ( .B1(n12654), .B2(n14772), .A(n12653), .ZN(P3_U3205) );
  OAI21_X1 U14867 ( .B1(n12656), .B2(n8646), .A(n12655), .ZN(n12658) );
  AOI21_X1 U14868 ( .B1(n12658), .B2(n12768), .A(n12657), .ZN(n12783) );
  INV_X1 U14869 ( .A(n12659), .ZN(n12661) );
  OAI22_X1 U14870 ( .A1(n12661), .A2(n14755), .B1(n14770), .B2(n12660), .ZN(
        n12665) );
  XNOR2_X1 U14871 ( .A(n12662), .B(n8646), .ZN(n12784) );
  NOR2_X1 U14872 ( .A1(n12784), .A2(n12663), .ZN(n12664) );
  AOI211_X1 U14873 ( .C1(n12773), .C2(n12781), .A(n12665), .B(n12664), .ZN(
        n12666) );
  OAI21_X1 U14874 ( .B1(n12783), .B2(n14772), .A(n12666), .ZN(P3_U3206) );
  XOR2_X1 U14875 ( .A(n12667), .B(n12669), .Z(n12674) );
  XNOR2_X1 U14876 ( .A(n12668), .B(n12669), .ZN(n12786) );
  OAI22_X1 U14877 ( .A1(n12671), .A2(n14760), .B1(n12670), .B2(n14762), .ZN(
        n12672) );
  AOI21_X1 U14878 ( .B1(n12786), .B2(n14805), .A(n12672), .ZN(n12673) );
  OAI21_X1 U14879 ( .B1(n12674), .B2(n14767), .A(n12673), .ZN(n12785) );
  INV_X1 U14880 ( .A(n12785), .ZN(n12680) );
  AOI22_X1 U14881 ( .A1(n12675), .A2(n12755), .B1(n14772), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12676) );
  OAI21_X1 U14882 ( .B1(n12831), .B2(n12757), .A(n12676), .ZN(n12677) );
  AOI21_X1 U14883 ( .B1(n12786), .B2(n12678), .A(n12677), .ZN(n12679) );
  OAI21_X1 U14884 ( .B1(n12680), .B2(n14772), .A(n12679), .ZN(P3_U3207) );
  OAI211_X1 U14885 ( .C1(n12683), .C2(n12682), .A(n12681), .B(n12768), .ZN(
        n12685) );
  NAND2_X1 U14886 ( .A1(n12685), .A2(n12684), .ZN(n12789) );
  INV_X1 U14887 ( .A(n12789), .ZN(n12693) );
  OAI21_X1 U14888 ( .B1(n12688), .B2(n12687), .A(n12686), .ZN(n12790) );
  AOI22_X1 U14889 ( .A1(n12689), .A2(n12755), .B1(n14772), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12690) );
  OAI21_X1 U14890 ( .B1(n12834), .B2(n12757), .A(n12690), .ZN(n12691) );
  AOI21_X1 U14891 ( .B1(n12790), .B2(n12778), .A(n12691), .ZN(n12692) );
  OAI21_X1 U14892 ( .B1(n12693), .B2(n14772), .A(n12692), .ZN(P3_U3208) );
  NAND2_X1 U14893 ( .A1(n12695), .A2(n12694), .ZN(n12697) );
  OAI211_X1 U14894 ( .C1(n12708), .C2(n12697), .A(n12696), .B(n12768), .ZN(
        n12699) );
  NAND2_X1 U14895 ( .A1(n12699), .A2(n12698), .ZN(n12793) );
  INV_X1 U14896 ( .A(n12793), .ZN(n12706) );
  XNOR2_X1 U14897 ( .A(n12700), .B(n12701), .ZN(n12794) );
  AOI22_X1 U14898 ( .A1(n12702), .A2(n12755), .B1(n14772), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12703) );
  OAI21_X1 U14899 ( .B1(n12838), .B2(n12757), .A(n12703), .ZN(n12704) );
  AOI21_X1 U14900 ( .B1(n12794), .B2(n12778), .A(n12704), .ZN(n12705) );
  OAI21_X1 U14901 ( .B1(n12706), .B2(n14772), .A(n12705), .ZN(P3_U3209) );
  OAI21_X1 U14902 ( .B1(n6515), .B2(n12710), .A(n12768), .ZN(n12709) );
  OAI21_X1 U14903 ( .B1(n12709), .B2(n12708), .A(n12707), .ZN(n12797) );
  INV_X1 U14904 ( .A(n12797), .ZN(n12716) );
  XNOR2_X1 U14905 ( .A(n12711), .B(n12710), .ZN(n12798) );
  AOI22_X1 U14906 ( .A1(n14772), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n12755), 
        .B2(n12712), .ZN(n12713) );
  OAI21_X1 U14907 ( .B1(n12842), .B2(n12757), .A(n12713), .ZN(n12714) );
  AOI21_X1 U14908 ( .B1(n12798), .B2(n12778), .A(n12714), .ZN(n12715) );
  OAI21_X1 U14909 ( .B1(n12716), .B2(n14772), .A(n12715), .ZN(P3_U3210) );
  XNOR2_X1 U14910 ( .A(n12717), .B(n12721), .ZN(n12719) );
  OAI21_X1 U14911 ( .B1(n12719), .B2(n14767), .A(n12718), .ZN(n12801) );
  INV_X1 U14912 ( .A(n12801), .ZN(n12726) );
  XNOR2_X1 U14913 ( .A(n12720), .B(n12721), .ZN(n12802) );
  AOI22_X1 U14914 ( .A1(n14772), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n12755), 
        .B2(n12722), .ZN(n12723) );
  OAI21_X1 U14915 ( .B1(n12845), .B2(n12757), .A(n12723), .ZN(n12724) );
  AOI21_X1 U14916 ( .B1(n12802), .B2(n12778), .A(n12724), .ZN(n12725) );
  OAI21_X1 U14917 ( .B1(n12726), .B2(n14772), .A(n12725), .ZN(P3_U3211) );
  XOR2_X1 U14918 ( .A(n12727), .B(n12730), .Z(n12729) );
  OAI21_X1 U14919 ( .B1(n12729), .B2(n14767), .A(n12728), .ZN(n12805) );
  INV_X1 U14920 ( .A(n12805), .ZN(n12736) );
  XOR2_X1 U14921 ( .A(n12731), .B(n12730), .Z(n12806) );
  AOI22_X1 U14922 ( .A1(n14772), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n12755), 
        .B2(n12732), .ZN(n12733) );
  OAI21_X1 U14923 ( .B1(n12849), .B2(n12757), .A(n12733), .ZN(n12734) );
  AOI21_X1 U14924 ( .B1(n12806), .B2(n12778), .A(n12734), .ZN(n12735) );
  OAI21_X1 U14925 ( .B1(n12736), .B2(n14772), .A(n12735), .ZN(P3_U3212) );
  OAI211_X1 U14926 ( .C1(n12739), .C2(n12738), .A(n12737), .B(n12768), .ZN(
        n12741) );
  NAND2_X1 U14927 ( .A1(n12741), .A2(n12740), .ZN(n12809) );
  INV_X1 U14928 ( .A(n12809), .ZN(n12748) );
  XNOR2_X1 U14929 ( .A(n12743), .B(n12742), .ZN(n12810) );
  AOI22_X1 U14930 ( .A1(n14772), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n12755), 
        .B2(n12744), .ZN(n12745) );
  OAI21_X1 U14931 ( .B1(n12853), .B2(n12757), .A(n12745), .ZN(n12746) );
  AOI21_X1 U14932 ( .B1(n12810), .B2(n12778), .A(n12746), .ZN(n12747) );
  OAI21_X1 U14933 ( .B1(n12748), .B2(n14772), .A(n12747), .ZN(P3_U3213) );
  XNOR2_X1 U14934 ( .A(n12749), .B(n12752), .ZN(n12751) );
  OAI21_X1 U14935 ( .B1(n12751), .B2(n14767), .A(n12750), .ZN(n12813) );
  INV_X1 U14936 ( .A(n12813), .ZN(n12760) );
  XOR2_X1 U14937 ( .A(n12753), .B(n12752), .Z(n12814) );
  AOI22_X1 U14938 ( .A1(n14772), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n12755), 
        .B2(n12754), .ZN(n12756) );
  OAI21_X1 U14939 ( .B1(n12857), .B2(n12757), .A(n12756), .ZN(n12758) );
  AOI21_X1 U14940 ( .B1(n12814), .B2(n12778), .A(n12758), .ZN(n12759) );
  OAI21_X1 U14941 ( .B1(n12760), .B2(n14772), .A(n12759), .ZN(P3_U3214) );
  OAI21_X1 U14942 ( .B1(n12762), .B2(n12777), .A(n12761), .ZN(n12767) );
  AOI222_X1 U14943 ( .A1(n12768), .A2(n12767), .B1(n12766), .B2(n12765), .C1(
        n12764), .C2(n12763), .ZN(n12819) );
  INV_X1 U14944 ( .A(n12769), .ZN(n12770) );
  OAI22_X1 U14945 ( .A1(n14770), .A2(n12771), .B1(n12770), .B2(n14755), .ZN(
        n12772) );
  AOI21_X1 U14946 ( .B1(n12774), .B2(n12773), .A(n12772), .ZN(n12780) );
  NAND2_X1 U14947 ( .A1(n12776), .A2(n12777), .ZN(n12817) );
  NAND3_X1 U14948 ( .A1(n12775), .A2(n12817), .A3(n12778), .ZN(n12779) );
  OAI211_X1 U14949 ( .C1(n12819), .C2(n14772), .A(n12780), .B(n12779), .ZN(
        P3_U3215) );
  NAND2_X1 U14950 ( .A1(n12781), .A2(n14812), .ZN(n12782) );
  OAI211_X1 U14951 ( .C1(n14828), .C2(n12784), .A(n12783), .B(n12782), .ZN(
        n12827) );
  MUX2_X1 U14952 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n12827), .S(n14846), .Z(
        P3_U3486) );
  INV_X1 U14953 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12787) );
  INV_X1 U14954 ( .A(n14821), .ZN(n14780) );
  AOI21_X1 U14955 ( .B1(n14780), .B2(n12786), .A(n12785), .ZN(n12828) );
  MUX2_X1 U14956 ( .A(n12787), .B(n12828), .S(n14846), .Z(n12788) );
  OAI21_X1 U14957 ( .B1(n12831), .B2(n12826), .A(n12788), .ZN(P3_U3485) );
  INV_X1 U14958 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12791) );
  AOI21_X1 U14959 ( .B1(n14106), .B2(n12790), .A(n12789), .ZN(n12832) );
  MUX2_X1 U14960 ( .A(n12791), .B(n12832), .S(n14846), .Z(n12792) );
  OAI21_X1 U14961 ( .B1(n12834), .B2(n12826), .A(n12792), .ZN(P3_U3484) );
  INV_X1 U14962 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12795) );
  AOI21_X1 U14963 ( .B1(n12794), .B2(n14106), .A(n12793), .ZN(n12835) );
  MUX2_X1 U14964 ( .A(n12795), .B(n12835), .S(n14846), .Z(n12796) );
  OAI21_X1 U14965 ( .B1(n12838), .B2(n12826), .A(n12796), .ZN(P3_U3483) );
  INV_X1 U14966 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12799) );
  AOI21_X1 U14967 ( .B1(n12798), .B2(n14106), .A(n12797), .ZN(n12839) );
  MUX2_X1 U14968 ( .A(n12799), .B(n12839), .S(n14846), .Z(n12800) );
  OAI21_X1 U14969 ( .B1(n12842), .B2(n12826), .A(n12800), .ZN(P3_U3482) );
  INV_X1 U14970 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12803) );
  AOI21_X1 U14971 ( .B1(n12802), .B2(n14106), .A(n12801), .ZN(n12843) );
  MUX2_X1 U14972 ( .A(n12803), .B(n12843), .S(n14846), .Z(n12804) );
  OAI21_X1 U14973 ( .B1(n12845), .B2(n12826), .A(n12804), .ZN(P3_U3481) );
  AOI21_X1 U14974 ( .B1(n12806), .B2(n14106), .A(n12805), .ZN(n12846) );
  MUX2_X1 U14975 ( .A(n12807), .B(n12846), .S(n14846), .Z(n12808) );
  OAI21_X1 U14976 ( .B1(n12849), .B2(n12826), .A(n12808), .ZN(P3_U3480) );
  INV_X1 U14977 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12811) );
  AOI21_X1 U14978 ( .B1(n12810), .B2(n14106), .A(n12809), .ZN(n12850) );
  MUX2_X1 U14979 ( .A(n12811), .B(n12850), .S(n14846), .Z(n12812) );
  OAI21_X1 U14980 ( .B1(n12853), .B2(n12826), .A(n12812), .ZN(P3_U3479) );
  INV_X1 U14981 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12815) );
  AOI21_X1 U14982 ( .B1(n12814), .B2(n14106), .A(n12813), .ZN(n12854) );
  MUX2_X1 U14983 ( .A(n12815), .B(n12854), .S(n14846), .Z(n12816) );
  OAI21_X1 U14984 ( .B1(n12826), .B2(n12857), .A(n12816), .ZN(P3_U3478) );
  INV_X1 U14985 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12820) );
  NAND3_X1 U14986 ( .A1(n12775), .A2(n14106), .A3(n12817), .ZN(n12818) );
  AND2_X1 U14987 ( .A1(n12819), .A2(n12818), .ZN(n12858) );
  MUX2_X1 U14988 ( .A(n12820), .B(n12858), .S(n14846), .Z(n12821) );
  OAI21_X1 U14989 ( .B1(n12861), .B2(n12826), .A(n12821), .ZN(P3_U3477) );
  INV_X1 U14990 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12824) );
  AOI21_X1 U14991 ( .B1(n12823), .B2(n14106), .A(n12822), .ZN(n12862) );
  MUX2_X1 U14992 ( .A(n12824), .B(n12862), .S(n14846), .Z(n12825) );
  OAI21_X1 U14993 ( .B1(n12866), .B2(n12826), .A(n12825), .ZN(P3_U3476) );
  MUX2_X1 U14994 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n12827), .S(n14833), .Z(
        P3_U3454) );
  INV_X1 U14995 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12829) );
  MUX2_X1 U14996 ( .A(n12829), .B(n12828), .S(n14833), .Z(n12830) );
  OAI21_X1 U14997 ( .B1(n12831), .B2(n12865), .A(n12830), .ZN(P3_U3453) );
  MUX2_X1 U14998 ( .A(n14849), .B(n12832), .S(n14833), .Z(n12833) );
  OAI21_X1 U14999 ( .B1(n12834), .B2(n12865), .A(n12833), .ZN(P3_U3452) );
  INV_X1 U15000 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12836) );
  MUX2_X1 U15001 ( .A(n12836), .B(n12835), .S(n14833), .Z(n12837) );
  OAI21_X1 U15002 ( .B1(n12838), .B2(n12865), .A(n12837), .ZN(P3_U3451) );
  INV_X1 U15003 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12840) );
  MUX2_X1 U15004 ( .A(n12840), .B(n12839), .S(n14833), .Z(n12841) );
  OAI21_X1 U15005 ( .B1(n12842), .B2(n12865), .A(n12841), .ZN(P3_U3450) );
  INV_X1 U15006 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n14893) );
  MUX2_X1 U15007 ( .A(n14893), .B(n12843), .S(n14833), .Z(n12844) );
  OAI21_X1 U15008 ( .B1(n12845), .B2(n12865), .A(n12844), .ZN(P3_U3449) );
  INV_X1 U15009 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12847) );
  MUX2_X1 U15010 ( .A(n12847), .B(n12846), .S(n14833), .Z(n12848) );
  OAI21_X1 U15011 ( .B1(n12849), .B2(n12865), .A(n12848), .ZN(P3_U3448) );
  INV_X1 U15012 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12851) );
  MUX2_X1 U15013 ( .A(n12851), .B(n12850), .S(n14833), .Z(n12852) );
  OAI21_X1 U15014 ( .B1(n12853), .B2(n12865), .A(n12852), .ZN(P3_U3447) );
  INV_X1 U15015 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12855) );
  MUX2_X1 U15016 ( .A(n12855), .B(n12854), .S(n14833), .Z(n12856) );
  OAI21_X1 U15017 ( .B1(n12865), .B2(n12857), .A(n12856), .ZN(P3_U3446) );
  INV_X1 U15018 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12859) );
  MUX2_X1 U15019 ( .A(n12859), .B(n12858), .S(n14833), .Z(n12860) );
  OAI21_X1 U15020 ( .B1(n12861), .B2(n12865), .A(n12860), .ZN(P3_U3444) );
  INV_X1 U15021 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12863) );
  MUX2_X1 U15022 ( .A(n12863), .B(n12862), .S(n14833), .Z(n12864) );
  OAI21_X1 U15023 ( .B1(n12866), .B2(n12865), .A(n12864), .ZN(P3_U3441) );
  NAND2_X1 U15024 ( .A1(n12867), .A2(n14038), .ZN(n12871) );
  INV_X1 U15025 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n12869) );
  NAND4_X1 U15026 ( .A1(n12868), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .A4(n12869), .ZN(n12870) );
  OAI211_X1 U15027 ( .C1(n12872), .C2(n12874), .A(n12871), .B(n12870), .ZN(
        P3_U3264) );
  INV_X1 U15028 ( .A(n12873), .ZN(n12876) );
  OAI222_X1 U15029 ( .A1(P3_U3151), .A2(n12877), .B1(n12880), .B2(n12876), 
        .C1(n12875), .C2(n12874), .ZN(P3_U3266) );
  INV_X1 U15030 ( .A(n12878), .ZN(n12879) );
  XNOR2_X1 U15031 ( .A(n13338), .B(n12948), .ZN(n12910) );
  INV_X1 U15032 ( .A(n12910), .ZN(n12912) );
  NAND2_X1 U15033 ( .A1(n10256), .A2(n13052), .ZN(n12911) );
  INV_X1 U15034 ( .A(n12881), .ZN(n12882) );
  NAND2_X1 U15035 ( .A1(n12883), .A2(n12882), .ZN(n12884) );
  XNOR2_X1 U15036 ( .A(n13369), .B(n12917), .ZN(n12887) );
  NAND2_X1 U15037 ( .A1(n13057), .A2(n6458), .ZN(n12888) );
  XNOR2_X1 U15038 ( .A(n12887), .B(n12888), .ZN(n13024) );
  INV_X1 U15039 ( .A(n13024), .ZN(n12886) );
  INV_X1 U15040 ( .A(n12887), .ZN(n12890) );
  INV_X1 U15041 ( .A(n12888), .ZN(n12889) );
  NAND2_X1 U15042 ( .A1(n12890), .A2(n12889), .ZN(n12891) );
  NAND2_X1 U15043 ( .A1(n13026), .A2(n12891), .ZN(n12936) );
  XNOR2_X1 U15044 ( .A(n13365), .B(n12917), .ZN(n12892) );
  NAND2_X1 U15045 ( .A1(n13056), .A2(n6458), .ZN(n12893) );
  NAND2_X1 U15046 ( .A1(n12892), .A2(n12893), .ZN(n12935) );
  INV_X1 U15047 ( .A(n12892), .ZN(n12895) );
  INV_X1 U15048 ( .A(n12893), .ZN(n12894) );
  NAND2_X1 U15049 ( .A1(n12895), .A2(n12894), .ZN(n12934) );
  XNOR2_X1 U15050 ( .A(n13359), .B(n12917), .ZN(n12896) );
  NAND2_X1 U15051 ( .A1(n13055), .A2(n10256), .ZN(n12897) );
  NAND2_X1 U15052 ( .A1(n12896), .A2(n12897), .ZN(n12901) );
  INV_X1 U15053 ( .A(n12896), .ZN(n12899) );
  INV_X1 U15054 ( .A(n12897), .ZN(n12898) );
  NAND2_X1 U15055 ( .A1(n12899), .A2(n12898), .ZN(n12900) );
  NAND2_X1 U15056 ( .A1(n12901), .A2(n12900), .ZN(n12994) );
  XNOR2_X1 U15057 ( .A(n13354), .B(n12917), .ZN(n12902) );
  NAND2_X1 U15058 ( .A1(n13054), .A2(n10256), .ZN(n12903) );
  XNOR2_X1 U15059 ( .A(n12902), .B(n12903), .ZN(n12958) );
  XNOR2_X1 U15060 ( .A(n13349), .B(n12917), .ZN(n13008) );
  NAND2_X1 U15061 ( .A1(n13012), .A2(n10256), .ZN(n13010) );
  INV_X1 U15062 ( .A(n12902), .ZN(n12905) );
  INV_X1 U15063 ( .A(n12903), .ZN(n12904) );
  NAND2_X1 U15064 ( .A1(n12905), .A2(n12904), .ZN(n13005) );
  OAI21_X1 U15065 ( .B1(n13008), .B2(n13010), .A(n13005), .ZN(n12908) );
  INV_X1 U15066 ( .A(n13010), .ZN(n12907) );
  INV_X1 U15067 ( .A(n13008), .ZN(n12906) );
  XNOR2_X1 U15068 ( .A(n12910), .B(n12911), .ZN(n12984) );
  XNOR2_X1 U15069 ( .A(n13167), .B(n12948), .ZN(n12914) );
  NAND2_X1 U15070 ( .A1(n13051), .A2(n10256), .ZN(n12913) );
  XNOR2_X1 U15071 ( .A(n12914), .B(n12913), .ZN(n12965) );
  INV_X1 U15072 ( .A(n12913), .ZN(n12915) );
  AND2_X1 U15073 ( .A1(n13050), .A2(n10256), .ZN(n12919) );
  XNOR2_X1 U15074 ( .A(n13326), .B(n12917), .ZN(n12918) );
  NOR2_X1 U15075 ( .A1(n12918), .A2(n12919), .ZN(n12920) );
  AOI21_X1 U15076 ( .B1(n12919), .B2(n12918), .A(n12920), .ZN(n13033) );
  XNOR2_X1 U15077 ( .A(n13128), .B(n12948), .ZN(n12944) );
  NAND2_X1 U15078 ( .A1(n13049), .A2(n10256), .ZN(n12943) );
  XNOR2_X1 U15079 ( .A(n12944), .B(n12943), .ZN(n12945) );
  XNOR2_X1 U15080 ( .A(n12946), .B(n12945), .ZN(n12926) );
  OAI22_X1 U15081 ( .A1(n12922), .A2(n12997), .B1(n12968), .B2(n12995), .ZN(
        n13126) );
  AOI22_X1 U15082 ( .A1(n12999), .A2(n13126), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12923) );
  OAI21_X1 U15083 ( .B1(n13015), .B2(n13133), .A(n12923), .ZN(n12924) );
  AOI21_X1 U15084 ( .B1(n8135), .B2(n6418), .A(n12924), .ZN(n12925) );
  OAI21_X1 U15085 ( .B1(n12926), .B2(n13023), .A(n12925), .ZN(P2_U3186) );
  OAI22_X1 U15086 ( .A1(n12928), .A2(n12995), .B1(n12927), .B2(n12997), .ZN(
        n13190) );
  AOI22_X1 U15087 ( .A1(n13190), .A2(n12999), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12929) );
  OAI21_X1 U15088 ( .B1(n13197), .B2(n13015), .A(n12929), .ZN(n12930) );
  AOI21_X1 U15089 ( .B1(n13344), .B2(n6418), .A(n12930), .ZN(n12933) );
  NAND3_X1 U15090 ( .A1(n12931), .A2(n13013), .A3(n13053), .ZN(n12932) );
  OAI211_X1 U15091 ( .C1(n6716), .C2(n13023), .A(n12933), .B(n12932), .ZN(
        P2_U3188) );
  NAND2_X1 U15092 ( .A1(n12935), .A2(n12934), .ZN(n12937) );
  XOR2_X1 U15093 ( .A(n12937), .B(n12936), .Z(n12942) );
  AND2_X1 U15094 ( .A1(n13057), .A2(n13038), .ZN(n12938) );
  AOI21_X1 U15095 ( .B1(n13055), .B2(n13037), .A(n12938), .ZN(n13255) );
  NAND2_X1 U15096 ( .A1(n13042), .A2(n13260), .ZN(n12939) );
  NAND2_X1 U15097 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13095)
         );
  OAI211_X1 U15098 ( .C1(n13255), .C2(n13040), .A(n12939), .B(n13095), .ZN(
        n12940) );
  AOI21_X1 U15099 ( .B1(n13365), .B2(n6418), .A(n12940), .ZN(n12941) );
  OAI21_X1 U15100 ( .B1(n12942), .B2(n13023), .A(n12941), .ZN(P2_U3191) );
  NAND2_X1 U15101 ( .A1(n13048), .A2(n10256), .ZN(n12947) );
  XOR2_X1 U15102 ( .A(n12948), .B(n12947), .Z(n12949) );
  XNOR2_X1 U15103 ( .A(n13118), .B(n12949), .ZN(n12950) );
  XNOR2_X1 U15104 ( .A(n12951), .B(n12950), .ZN(n12957) );
  OAI22_X1 U15105 ( .A1(n12953), .A2(n12997), .B1(n12952), .B2(n12995), .ZN(
        n13111) );
  AOI22_X1 U15106 ( .A1(n12999), .A2(n13111), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12954) );
  OAI21_X1 U15107 ( .B1(n13015), .B2(n13114), .A(n12954), .ZN(n12955) );
  AOI21_X1 U15108 ( .B1(n13315), .B2(n6418), .A(n12955), .ZN(n12956) );
  OAI21_X1 U15109 ( .B1(n12957), .B2(n13023), .A(n12956), .ZN(P2_U3192) );
  XNOR2_X1 U15110 ( .A(n12959), .B(n12958), .ZN(n12964) );
  AOI22_X1 U15111 ( .A1(n13012), .A2(n13037), .B1(n13038), .B2(n13055), .ZN(
        n13219) );
  OAI22_X1 U15112 ( .A1(n13219), .A2(n13040), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12960), .ZN(n12962) );
  NOR2_X1 U15113 ( .A1(n13230), .A2(n13045), .ZN(n12961) );
  AOI211_X1 U15114 ( .C1(n13042), .C2(n13227), .A(n12962), .B(n12961), .ZN(
        n12963) );
  OAI21_X1 U15115 ( .B1(n12964), .B2(n13023), .A(n12963), .ZN(P2_U3195) );
  XNOR2_X1 U15116 ( .A(n12966), .B(n12965), .ZN(n12972) );
  NAND2_X1 U15117 ( .A1(n13038), .A2(n13052), .ZN(n12967) );
  OAI21_X1 U15118 ( .B1(n12968), .B2(n12997), .A(n12967), .ZN(n13158) );
  AOI22_X1 U15119 ( .A1(n12999), .A2(n13158), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12969) );
  OAI21_X1 U15120 ( .B1(n13015), .B2(n13165), .A(n12969), .ZN(n12970) );
  AOI21_X1 U15121 ( .B1(n13167), .B2(n6418), .A(n12970), .ZN(n12971) );
  OAI21_X1 U15122 ( .B1(n12972), .B2(n13023), .A(n12971), .ZN(P2_U3197) );
  INV_X1 U15123 ( .A(n11977), .ZN(n12973) );
  AOI21_X1 U15124 ( .B1(n12975), .B2(n12974), .A(n12973), .ZN(n12982) );
  NAND2_X1 U15125 ( .A1(n12999), .A2(n12976), .ZN(n12977) );
  OAI211_X1 U15126 ( .C1(n13015), .C2(n12979), .A(n12978), .B(n12977), .ZN(
        n12980) );
  AOI21_X1 U15127 ( .B1(n13378), .B2(n6418), .A(n12980), .ZN(n12981) );
  OAI21_X1 U15128 ( .B1(n12982), .B2(n13023), .A(n12981), .ZN(P2_U3198) );
  OAI211_X1 U15129 ( .C1(n6555), .C2(n12984), .A(n12983), .B(n13035), .ZN(
        n12990) );
  OAI22_X1 U15130 ( .A1(n12986), .A2(n12995), .B1(n12985), .B2(n12997), .ZN(
        n13176) );
  AOI22_X1 U15131 ( .A1(n13176), .A2(n12999), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12987) );
  OAI21_X1 U15132 ( .B1(n13181), .B2(n13015), .A(n12987), .ZN(n12988) );
  AOI21_X1 U15133 ( .B1(n13338), .B2(n6418), .A(n12988), .ZN(n12989) );
  NAND2_X1 U15134 ( .A1(n12990), .A2(n12989), .ZN(P2_U3201) );
  INV_X1 U15135 ( .A(n12991), .ZN(n12992) );
  AOI21_X1 U15136 ( .B1(n12994), .B2(n12993), .A(n12992), .ZN(n13004) );
  OAI22_X1 U15137 ( .A1(n12998), .A2(n12997), .B1(n12996), .B2(n12995), .ZN(
        n13237) );
  AOI22_X1 U15138 ( .A1(n13237), .A2(n12999), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13000) );
  OAI21_X1 U15139 ( .B1(n13244), .B2(n13015), .A(n13000), .ZN(n13001) );
  AOI21_X1 U15140 ( .B1(n13359), .B2(n6418), .A(n13001), .ZN(n13003) );
  OAI21_X1 U15141 ( .B1(n13004), .B2(n13023), .A(n13003), .ZN(P2_U3205) );
  INV_X1 U15142 ( .A(n13005), .ZN(n13006) );
  OR2_X1 U15143 ( .A1(n13007), .A2(n13006), .ZN(n13009) );
  XNOR2_X1 U15144 ( .A(n13009), .B(n13008), .ZN(n13011) );
  NAND3_X1 U15145 ( .A1(n13011), .A2(n13035), .A3(n13010), .ZN(n13022) );
  INV_X1 U15146 ( .A(n13011), .ZN(n13014) );
  NAND3_X1 U15147 ( .A1(n13014), .A2(n13013), .A3(n13012), .ZN(n13021) );
  NOR2_X1 U15148 ( .A1(n13015), .A2(n13211), .ZN(n13019) );
  AND2_X1 U15149 ( .A1(n13054), .A2(n13038), .ZN(n13016) );
  AOI21_X1 U15150 ( .B1(n13053), .B2(n13037), .A(n13016), .ZN(n13204) );
  OAI22_X1 U15151 ( .A1(n13204), .A2(n13040), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13017), .ZN(n13018) );
  AOI211_X1 U15152 ( .C1(n13349), .C2(n6418), .A(n13019), .B(n13018), .ZN(
        n13020) );
  NAND3_X1 U15153 ( .A1(n13022), .A2(n13021), .A3(n13020), .ZN(P2_U3207) );
  AOI21_X1 U15154 ( .B1(n13025), .B2(n13024), .A(n13023), .ZN(n13027) );
  NAND2_X1 U15155 ( .A1(n13027), .A2(n13026), .ZN(n13031) );
  INV_X1 U15156 ( .A(n13028), .ZN(n13272) );
  AOI22_X1 U15157 ( .A1(n13056), .A2(n13037), .B1(n13038), .B2(n13058), .ZN(
        n13267) );
  OAI22_X1 U15158 ( .A1(n13040), .A2(n13267), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14533), .ZN(n13029) );
  AOI21_X1 U15159 ( .B1(n13272), .B2(n13042), .A(n13029), .ZN(n13030) );
  OAI211_X1 U15160 ( .C1(n13274), .C2(n13045), .A(n13031), .B(n13030), .ZN(
        P2_U3210) );
  INV_X1 U15161 ( .A(n13147), .ZN(n13043) );
  AOI22_X1 U15162 ( .A1(n13038), .A2(n13051), .B1(n13049), .B2(n13037), .ZN(
        n13141) );
  OAI22_X1 U15163 ( .A1(n13040), .A2(n13141), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13039), .ZN(n13041) );
  AOI21_X1 U15164 ( .B1(n13043), .B2(n13042), .A(n13041), .ZN(n13044) );
  MUX2_X1 U15165 ( .A(n13101), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13072), .Z(
        P2_U3562) );
  MUX2_X1 U15166 ( .A(n13046), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13072), .Z(
        P2_U3561) );
  MUX2_X1 U15167 ( .A(n13047), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13072), .Z(
        P2_U3560) );
  MUX2_X1 U15168 ( .A(n13048), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13072), .Z(
        P2_U3559) );
  MUX2_X1 U15169 ( .A(n13049), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13072), .Z(
        P2_U3558) );
  MUX2_X1 U15170 ( .A(n13050), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13072), .Z(
        P2_U3557) );
  MUX2_X1 U15171 ( .A(n13051), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13072), .Z(
        P2_U3556) );
  MUX2_X1 U15172 ( .A(n13052), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13072), .Z(
        P2_U3555) );
  MUX2_X1 U15173 ( .A(n13053), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13072), .Z(
        P2_U3554) );
  MUX2_X1 U15174 ( .A(n13054), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13072), .Z(
        P2_U3552) );
  MUX2_X1 U15175 ( .A(n13055), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13072), .Z(
        P2_U3551) );
  MUX2_X1 U15176 ( .A(n13056), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13072), .Z(
        P2_U3550) );
  MUX2_X1 U15177 ( .A(n13057), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13072), .Z(
        P2_U3549) );
  MUX2_X1 U15178 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13058), .S(P2_U3947), .Z(
        P2_U3548) );
  MUX2_X1 U15179 ( .A(n13059), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13072), .Z(
        P2_U3547) );
  MUX2_X1 U15180 ( .A(n13060), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13072), .Z(
        P2_U3546) );
  MUX2_X1 U15181 ( .A(n13061), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13072), .Z(
        P2_U3545) );
  MUX2_X1 U15182 ( .A(n13062), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13072), .Z(
        P2_U3544) );
  MUX2_X1 U15183 ( .A(n13063), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13072), .Z(
        P2_U3543) );
  MUX2_X1 U15184 ( .A(n13064), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13072), .Z(
        P2_U3542) );
  MUX2_X1 U15185 ( .A(n13065), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13072), .Z(
        P2_U3541) );
  MUX2_X1 U15186 ( .A(n13066), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13072), .Z(
        P2_U3540) );
  MUX2_X1 U15187 ( .A(n13067), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13072), .Z(
        P2_U3539) );
  MUX2_X1 U15188 ( .A(n13068), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13072), .Z(
        P2_U3538) );
  MUX2_X1 U15189 ( .A(n13069), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13072), .Z(
        P2_U3537) );
  MUX2_X1 U15190 ( .A(n13070), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13072), .Z(
        P2_U3536) );
  MUX2_X1 U15191 ( .A(n13071), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13072), .Z(
        P2_U3535) );
  MUX2_X1 U15192 ( .A(n8149), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13072), .Z(
        P2_U3534) );
  MUX2_X1 U15193 ( .A(n8146), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13072), .Z(
        P2_U3533) );
  MUX2_X1 U15194 ( .A(n8148), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13072), .Z(
        P2_U3532) );
  MUX2_X1 U15195 ( .A(n9869), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13072), .Z(
        P2_U3531) );
  NAND2_X1 U15196 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n14520), .ZN(n13077) );
  INV_X1 U15197 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13074) );
  INV_X1 U15198 ( .A(n13077), .ZN(n13073) );
  AOI21_X1 U15199 ( .B1(n13074), .B2(n13085), .A(n13073), .ZN(n14528) );
  INV_X1 U15200 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13076) );
  OAI21_X1 U15201 ( .B1(n13083), .B2(n13076), .A(n13075), .ZN(n14527) );
  NAND2_X1 U15202 ( .A1(n14528), .A2(n14527), .ZN(n14525) );
  NOR2_X1 U15203 ( .A1(n13087), .A2(n13078), .ZN(n13079) );
  XNOR2_X1 U15204 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13080), .ZN(n13091) );
  INV_X1 U15205 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13084) );
  XNOR2_X1 U15206 ( .A(n13085), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14524) );
  INV_X1 U15207 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n13082) );
  OAI21_X1 U15208 ( .B1(n13083), .B2(n13082), .A(n13081), .ZN(n14523) );
  NAND2_X1 U15209 ( .A1(n14524), .A2(n14523), .ZN(n14522) );
  OAI21_X1 U15210 ( .B1(n13085), .B2(n13084), .A(n14522), .ZN(n13086) );
  XNOR2_X1 U15211 ( .A(n14546), .B(n13086), .ZN(n14543) );
  NAND2_X1 U15212 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n14543), .ZN(n14541) );
  NAND2_X1 U15213 ( .A1(n13087), .A2(n13086), .ZN(n13088) );
  NAND2_X1 U15214 ( .A1(n14541), .A2(n13088), .ZN(n13089) );
  XOR2_X1 U15215 ( .A(n13089), .B(P2_REG1_REG_19__SCAN_IN), .Z(n13092) );
  OAI21_X1 U15216 ( .B1(n13092), .B2(n14483), .A(n14547), .ZN(n13090) );
  AOI21_X1 U15217 ( .B1(n13091), .B2(n14526), .A(n13090), .ZN(n13094) );
  NAND2_X1 U15218 ( .A1(n13107), .A2(n13308), .ZN(n13106) );
  INV_X1 U15219 ( .A(n13100), .ZN(n13102) );
  NAND2_X1 U15220 ( .A1(n13102), .A2(n13101), .ZN(n13306) );
  NOR2_X1 U15221 ( .A1(n13304), .A2(n13306), .ZN(n13109) );
  NOR2_X1 U15222 ( .A1(n13098), .A2(n13294), .ZN(n13104) );
  AOI211_X1 U15223 ( .C1(n13304), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13109), 
        .B(n13104), .ZN(n13105) );
  OAI21_X1 U15224 ( .B1(n13170), .B2(n13305), .A(n13105), .ZN(P2_U3234) );
  OAI211_X1 U15225 ( .C1(n13107), .C2(n13308), .A(n13379), .B(n13106), .ZN(
        n13307) );
  NOR2_X1 U15226 ( .A1(n13308), .A2(n13294), .ZN(n13108) );
  AOI211_X1 U15227 ( .C1(n13304), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13109), 
        .B(n13108), .ZN(n13110) );
  OAI21_X1 U15228 ( .B1(n13170), .B2(n13307), .A(n13110), .ZN(P2_U3235) );
  OR2_X1 U15229 ( .A1(n13118), .A2(n13130), .ZN(n13112) );
  AND3_X1 U15230 ( .A1(n13113), .A2(n13112), .A3(n13379), .ZN(n13314) );
  INV_X1 U15231 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13115) );
  OAI22_X1 U15232 ( .A1(n13257), .A2(n13115), .B1(n13114), .B2(n13245), .ZN(
        n13116) );
  INV_X1 U15233 ( .A(n13116), .ZN(n13117) );
  OAI21_X1 U15234 ( .B1(n13118), .B2(n13294), .A(n13117), .ZN(n13123) );
  OAI21_X1 U15235 ( .B1(n13121), .B2(n13120), .A(n13119), .ZN(n13318) );
  NOR2_X1 U15236 ( .A1(n13318), .A2(n13299), .ZN(n13122) );
  AOI211_X1 U15237 ( .C1(n13314), .C2(n13302), .A(n13123), .B(n13122), .ZN(
        n13124) );
  OAI21_X1 U15238 ( .B1(n13317), .B2(n13304), .A(n13124), .ZN(P2_U3237) );
  XNOR2_X1 U15239 ( .A(n13125), .B(n13131), .ZN(n13127) );
  AOI21_X1 U15240 ( .B1(n13127), .B2(n13284), .A(n13126), .ZN(n13324) );
  OAI21_X1 U15241 ( .B1(n13128), .B2(n13146), .A(n13379), .ZN(n13129) );
  OR2_X1 U15242 ( .A1(n13130), .A2(n13129), .ZN(n13323) );
  OR2_X1 U15243 ( .A1(n13132), .A2(n13131), .ZN(n13320) );
  NAND3_X1 U15244 ( .A1(n13320), .A2(n13319), .A3(n13232), .ZN(n13137) );
  INV_X1 U15245 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13134) );
  OAI22_X1 U15246 ( .A1(n13257), .A2(n13134), .B1(n13133), .B2(n13245), .ZN(
        n13135) );
  AOI21_X1 U15247 ( .B1(n8135), .B2(n13241), .A(n13135), .ZN(n13136) );
  OAI211_X1 U15248 ( .C1(n13323), .C2(n13170), .A(n13137), .B(n13136), .ZN(
        n13138) );
  INV_X1 U15249 ( .A(n13138), .ZN(n13139) );
  OAI21_X1 U15250 ( .B1(n13324), .B2(n13304), .A(n13139), .ZN(P2_U3238) );
  XNOR2_X1 U15251 ( .A(n13140), .B(n13143), .ZN(n13142) );
  OAI21_X1 U15252 ( .B1(n13142), .B2(n13268), .A(n13141), .ZN(n13327) );
  INV_X1 U15253 ( .A(n13327), .ZN(n13154) );
  XNOR2_X1 U15254 ( .A(n13144), .B(n13143), .ZN(n13329) );
  OAI21_X1 U15255 ( .B1(n13164), .B2(n13326), .A(n13379), .ZN(n13145) );
  OR2_X1 U15256 ( .A1(n13146), .A2(n13145), .ZN(n13325) );
  INV_X1 U15257 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13148) );
  OAI22_X1 U15258 ( .A1(n13257), .A2(n13148), .B1(n13147), .B2(n13245), .ZN(
        n13149) );
  AOI21_X1 U15259 ( .B1(n13150), .B2(n13241), .A(n13149), .ZN(n13151) );
  OAI21_X1 U15260 ( .B1(n13325), .B2(n13170), .A(n13151), .ZN(n13152) );
  AOI21_X1 U15261 ( .B1(n13329), .B2(n13232), .A(n13152), .ZN(n13153) );
  OAI21_X1 U15262 ( .B1(n13154), .B2(n13304), .A(n13153), .ZN(P2_U3239) );
  OAI21_X1 U15263 ( .B1(n13157), .B2(n13156), .A(n13155), .ZN(n13159) );
  AOI21_X1 U15264 ( .B1(n13159), .B2(n13284), .A(n13158), .ZN(n13336) );
  OAI21_X1 U15265 ( .B1(n13162), .B2(n13161), .A(n13160), .ZN(n13334) );
  OAI21_X1 U15266 ( .B1(n13179), .B2(n13332), .A(n13379), .ZN(n13163) );
  OR2_X1 U15267 ( .A1(n13164), .A2(n13163), .ZN(n13331) );
  INV_X1 U15268 ( .A(n13165), .ZN(n13166) );
  AOI22_X1 U15269 ( .A1(n13304), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n13166), 
        .B2(n13291), .ZN(n13169) );
  NAND2_X1 U15270 ( .A1(n13167), .A2(n13241), .ZN(n13168) );
  OAI211_X1 U15271 ( .C1(n13331), .C2(n13170), .A(n13169), .B(n13168), .ZN(
        n13171) );
  AOI21_X1 U15272 ( .B1(n13334), .B2(n13232), .A(n13171), .ZN(n13172) );
  OAI21_X1 U15273 ( .B1(n13336), .B2(n13304), .A(n13172), .ZN(P2_U3240) );
  XNOR2_X1 U15274 ( .A(n13173), .B(n13174), .ZN(n13178) );
  XNOR2_X1 U15275 ( .A(n13175), .B(n13174), .ZN(n13342) );
  NOR2_X1 U15276 ( .A1(n13342), .A2(n9868), .ZN(n13177) );
  AOI211_X1 U15277 ( .C1(n13178), .C2(n13284), .A(n13177), .B(n13176), .ZN(
        n13340) );
  INV_X1 U15278 ( .A(n13194), .ZN(n13180) );
  AOI211_X1 U15279 ( .C1(n13338), .C2(n13180), .A(n13289), .B(n13179), .ZN(
        n13337) );
  INV_X1 U15280 ( .A(n13181), .ZN(n13182) );
  AOI22_X1 U15281 ( .A1(n13304), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13182), 
        .B2(n13291), .ZN(n13183) );
  OAI21_X1 U15282 ( .B1(n13184), .B2(n13294), .A(n13183), .ZN(n13187) );
  NOR2_X1 U15283 ( .A1(n13342), .A2(n13185), .ZN(n13186) );
  AOI211_X1 U15284 ( .C1(n13337), .C2(n13302), .A(n13187), .B(n13186), .ZN(
        n13188) );
  OAI21_X1 U15285 ( .B1(n13340), .B2(n13304), .A(n13188), .ZN(P2_U3241) );
  XOR2_X1 U15286 ( .A(n13198), .B(n13189), .Z(n13191) );
  AOI21_X1 U15287 ( .B1(n13191), .B2(n13284), .A(n13190), .ZN(n13346) );
  NAND2_X1 U15288 ( .A1(n13344), .A2(n13207), .ZN(n13192) );
  NAND2_X1 U15289 ( .A1(n13192), .A2(n13379), .ZN(n13193) );
  NOR2_X1 U15290 ( .A1(n13194), .A2(n13193), .ZN(n13343) );
  NAND2_X1 U15291 ( .A1(n13344), .A2(n13241), .ZN(n13196) );
  NAND2_X1 U15292 ( .A1(n13304), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n13195) );
  OAI211_X1 U15293 ( .C1(n13245), .C2(n13197), .A(n13196), .B(n13195), .ZN(
        n13201) );
  XNOR2_X1 U15294 ( .A(n13199), .B(n13198), .ZN(n13347) );
  NOR2_X1 U15295 ( .A1(n13347), .A2(n13299), .ZN(n13200) );
  AOI211_X1 U15296 ( .C1(n13343), .C2(n13302), .A(n13201), .B(n13200), .ZN(
        n13202) );
  OAI21_X1 U15297 ( .B1(n13346), .B2(n13304), .A(n13202), .ZN(P2_U3242) );
  AOI211_X1 U15298 ( .C1(n13213), .C2(n13203), .A(n13268), .B(n6514), .ZN(
        n13206) );
  INV_X1 U15299 ( .A(n13204), .ZN(n13205) );
  NOR2_X1 U15300 ( .A1(n13206), .A2(n13205), .ZN(n13351) );
  AOI21_X1 U15301 ( .B1(n13349), .B2(n13226), .A(n13289), .ZN(n13208) );
  AND2_X1 U15302 ( .A1(n13208), .A2(n13207), .ZN(n13348) );
  NAND2_X1 U15303 ( .A1(n13349), .A2(n13241), .ZN(n13210) );
  NAND2_X1 U15304 ( .A1(n13304), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n13209) );
  OAI211_X1 U15305 ( .C1(n13245), .C2(n13211), .A(n13210), .B(n13209), .ZN(
        n13216) );
  OAI21_X1 U15306 ( .B1(n13214), .B2(n13213), .A(n13212), .ZN(n13352) );
  NOR2_X1 U15307 ( .A1(n13352), .A2(n13299), .ZN(n13215) );
  AOI211_X1 U15308 ( .C1(n13348), .C2(n13302), .A(n13216), .B(n13215), .ZN(
        n13217) );
  OAI21_X1 U15309 ( .B1(n13351), .B2(n13304), .A(n13217), .ZN(P2_U3243) );
  XNOR2_X1 U15310 ( .A(n13218), .B(n13222), .ZN(n13221) );
  INV_X1 U15311 ( .A(n13219), .ZN(n13220) );
  AOI21_X1 U15312 ( .B1(n13221), .B2(n13284), .A(n13220), .ZN(n13356) );
  XOR2_X1 U15313 ( .A(n13223), .B(n13222), .Z(n13357) );
  INV_X1 U15314 ( .A(n13357), .ZN(n13233) );
  AOI21_X1 U15315 ( .B1(n13354), .B2(n13239), .A(n13289), .ZN(n13225) );
  AND2_X1 U15316 ( .A1(n13226), .A2(n13225), .ZN(n13353) );
  NAND2_X1 U15317 ( .A1(n13353), .A2(n13302), .ZN(n13229) );
  AOI22_X1 U15318 ( .A1(n13304), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13227), 
        .B2(n13291), .ZN(n13228) );
  OAI211_X1 U15319 ( .C1(n13230), .C2(n13294), .A(n13229), .B(n13228), .ZN(
        n13231) );
  AOI21_X1 U15320 ( .B1(n13233), .B2(n13232), .A(n13231), .ZN(n13234) );
  OAI21_X1 U15321 ( .B1(n13356), .B2(n13304), .A(n13234), .ZN(P2_U3244) );
  XNOR2_X1 U15322 ( .A(n13236), .B(n13235), .ZN(n13238) );
  AOI21_X1 U15323 ( .B1(n13238), .B2(n13284), .A(n13237), .ZN(n13361) );
  AOI21_X1 U15324 ( .B1(n13359), .B2(n13258), .A(n13289), .ZN(n13240) );
  AND2_X1 U15325 ( .A1(n13240), .A2(n13239), .ZN(n13358) );
  NAND2_X1 U15326 ( .A1(n13359), .A2(n13241), .ZN(n13243) );
  NAND2_X1 U15327 ( .A1(n13304), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n13242) );
  OAI211_X1 U15328 ( .C1(n13245), .C2(n13244), .A(n13243), .B(n13242), .ZN(
        n13249) );
  XNOR2_X1 U15329 ( .A(n13247), .B(n13246), .ZN(n13362) );
  NOR2_X1 U15330 ( .A1(n13362), .A2(n13299), .ZN(n13248) );
  AOI211_X1 U15331 ( .C1(n13358), .C2(n13302), .A(n13249), .B(n13248), .ZN(
        n13250) );
  OAI21_X1 U15332 ( .B1(n13361), .B2(n13304), .A(n13250), .ZN(P2_U3245) );
  NAND2_X1 U15333 ( .A1(n13275), .A2(n13251), .ZN(n13252) );
  XOR2_X1 U15334 ( .A(n13254), .B(n13252), .Z(n13367) );
  XOR2_X1 U15335 ( .A(n13254), .B(n13253), .Z(n13256) );
  OAI21_X1 U15336 ( .B1(n13256), .B2(n13268), .A(n13255), .ZN(n13363) );
  NAND2_X1 U15337 ( .A1(n13363), .A2(n13257), .ZN(n13265) );
  INV_X1 U15338 ( .A(n13258), .ZN(n13259) );
  AOI211_X1 U15339 ( .C1(n13365), .C2(n13271), .A(n13289), .B(n13259), .ZN(
        n13364) );
  AOI22_X1 U15340 ( .A1(n13304), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13260), 
        .B2(n13291), .ZN(n13261) );
  OAI21_X1 U15341 ( .B1(n13262), .B2(n13294), .A(n13261), .ZN(n13263) );
  AOI21_X1 U15342 ( .B1(n13364), .B2(n13302), .A(n13263), .ZN(n13264) );
  OAI211_X1 U15343 ( .C1(n13299), .C2(n13367), .A(n13265), .B(n13264), .ZN(
        P2_U3246) );
  XNOR2_X1 U15344 ( .A(n13266), .B(n13278), .ZN(n13269) );
  OAI21_X1 U15345 ( .B1(n13269), .B2(n13268), .A(n13267), .ZN(n13270) );
  INV_X1 U15346 ( .A(n13270), .ZN(n13371) );
  AOI211_X1 U15347 ( .C1(n13369), .C2(n13287), .A(n13289), .B(n6930), .ZN(
        n13368) );
  AOI22_X1 U15348 ( .A1(n13304), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13272), 
        .B2(n13291), .ZN(n13273) );
  OAI21_X1 U15349 ( .B1(n13274), .B2(n13294), .A(n13273), .ZN(n13280) );
  INV_X1 U15350 ( .A(n13275), .ZN(n13276) );
  AOI21_X1 U15351 ( .B1(n13278), .B2(n13277), .A(n13276), .ZN(n13372) );
  NOR2_X1 U15352 ( .A1(n13372), .A2(n13299), .ZN(n13279) );
  AOI211_X1 U15353 ( .C1(n13368), .C2(n13302), .A(n13280), .B(n13279), .ZN(
        n13281) );
  OAI21_X1 U15354 ( .B1(n13304), .B2(n13371), .A(n13281), .ZN(P2_U3247) );
  XNOR2_X1 U15355 ( .A(n13282), .B(n13297), .ZN(n13285) );
  AOI21_X1 U15356 ( .B1(n13285), .B2(n13284), .A(n13283), .ZN(n13376) );
  INV_X1 U15357 ( .A(n13286), .ZN(n13290) );
  INV_X1 U15358 ( .A(n13287), .ZN(n13288) );
  AOI211_X1 U15359 ( .C1(n13374), .C2(n13290), .A(n13289), .B(n13288), .ZN(
        n13373) );
  AOI22_X1 U15360 ( .A1(n13304), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13292), 
        .B2(n13291), .ZN(n13293) );
  OAI21_X1 U15361 ( .B1(n13295), .B2(n13294), .A(n13293), .ZN(n13301) );
  OAI21_X1 U15362 ( .B1(n13298), .B2(n13297), .A(n13296), .ZN(n13377) );
  NOR2_X1 U15363 ( .A1(n13377), .A2(n13299), .ZN(n13300) );
  AOI211_X1 U15364 ( .C1(n13373), .C2(n13302), .A(n13301), .B(n13300), .ZN(
        n13303) );
  OAI21_X1 U15365 ( .B1(n13304), .B2(n13376), .A(n13303), .ZN(P2_U3248) );
  OAI211_X1 U15366 ( .C1(n13098), .C2(n14592), .A(n13305), .B(n13306), .ZN(
        n13407) );
  MUX2_X1 U15367 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13407), .S(n10988), .Z(
        P2_U3530) );
  OAI211_X1 U15368 ( .C1(n13308), .C2(n14592), .A(n13307), .B(n13306), .ZN(
        n13408) );
  MUX2_X1 U15369 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13408), .S(n10988), .Z(
        P2_U3529) );
  AOI21_X1 U15370 ( .B1(n14567), .B2(n13310), .A(n13309), .ZN(n13311) );
  MUX2_X1 U15371 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13409), .S(n10988), .Z(
        P2_U3528) );
  AOI21_X1 U15372 ( .B1(n14567), .B2(n13315), .A(n13314), .ZN(n13316) );
  MUX2_X1 U15373 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13410), .S(n10988), .Z(
        P2_U3527) );
  NAND3_X1 U15374 ( .A1(n13320), .A2(n13319), .A3(n14589), .ZN(n13322) );
  NAND2_X1 U15375 ( .A1(n8135), .A2(n14567), .ZN(n13321) );
  NAND4_X1 U15376 ( .A1(n13324), .A2(n13323), .A3(n13322), .A4(n13321), .ZN(
        n13411) );
  MUX2_X1 U15377 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13411), .S(n10988), .Z(
        P2_U3526) );
  OAI21_X1 U15378 ( .B1(n13326), .B2(n14592), .A(n13325), .ZN(n13328) );
  AOI211_X1 U15379 ( .C1(n14589), .C2(n13329), .A(n13328), .B(n13327), .ZN(
        n13330) );
  INV_X1 U15380 ( .A(n13330), .ZN(n13412) );
  MUX2_X1 U15381 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13412), .S(n10988), .Z(
        P2_U3525) );
  OAI21_X1 U15382 ( .B1(n13332), .B2(n14592), .A(n13331), .ZN(n13333) );
  AOI21_X1 U15383 ( .B1(n13334), .B2(n14589), .A(n13333), .ZN(n13335) );
  NAND2_X1 U15384 ( .A1(n13336), .A2(n13335), .ZN(n13413) );
  MUX2_X1 U15385 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13413), .S(n10988), .Z(
        P2_U3524) );
  AOI21_X1 U15386 ( .B1(n14567), .B2(n13338), .A(n13337), .ZN(n13339) );
  OAI211_X1 U15387 ( .C1(n13342), .C2(n13341), .A(n13340), .B(n13339), .ZN(
        n13414) );
  MUX2_X1 U15388 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13414), .S(n10988), .Z(
        P2_U3523) );
  AOI21_X1 U15389 ( .B1(n14567), .B2(n13344), .A(n13343), .ZN(n13345) );
  OAI211_X1 U15390 ( .C1(n14571), .C2(n13347), .A(n13346), .B(n13345), .ZN(
        n13415) );
  MUX2_X1 U15391 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13415), .S(n10988), .Z(
        P2_U3522) );
  AOI21_X1 U15392 ( .B1(n14567), .B2(n13349), .A(n13348), .ZN(n13350) );
  OAI211_X1 U15393 ( .C1(n14571), .C2(n13352), .A(n13351), .B(n13350), .ZN(
        n13416) );
  MUX2_X1 U15394 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13416), .S(n10988), .Z(
        P2_U3521) );
  AOI21_X1 U15395 ( .B1(n14567), .B2(n13354), .A(n13353), .ZN(n13355) );
  OAI211_X1 U15396 ( .C1(n14571), .C2(n13357), .A(n13356), .B(n13355), .ZN(
        n13417) );
  MUX2_X1 U15397 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13417), .S(n10988), .Z(
        P2_U3520) );
  AOI21_X1 U15398 ( .B1(n14567), .B2(n13359), .A(n13358), .ZN(n13360) );
  OAI211_X1 U15399 ( .C1(n14571), .C2(n13362), .A(n13361), .B(n13360), .ZN(
        n13418) );
  MUX2_X1 U15400 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13418), .S(n10988), .Z(
        P2_U3519) );
  AOI211_X1 U15401 ( .C1(n14567), .C2(n13365), .A(n13364), .B(n13363), .ZN(
        n13366) );
  OAI21_X1 U15402 ( .B1(n14571), .B2(n13367), .A(n13366), .ZN(n13419) );
  MUX2_X1 U15403 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13419), .S(n10988), .Z(
        P2_U3518) );
  AOI21_X1 U15404 ( .B1(n14567), .B2(n13369), .A(n13368), .ZN(n13370) );
  OAI211_X1 U15405 ( .C1(n14571), .C2(n13372), .A(n13371), .B(n13370), .ZN(
        n13420) );
  MUX2_X1 U15406 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13420), .S(n10988), .Z(
        P2_U3517) );
  AOI21_X1 U15407 ( .B1(n14567), .B2(n13374), .A(n13373), .ZN(n13375) );
  OAI211_X1 U15408 ( .C1(n14571), .C2(n13377), .A(n13376), .B(n13375), .ZN(
        n13421) );
  MUX2_X1 U15409 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13421), .S(n10988), .Z(
        P2_U3516) );
  AOI22_X1 U15410 ( .A1(n13380), .A2(n13379), .B1(n14567), .B2(n13378), .ZN(
        n13384) );
  NAND3_X1 U15411 ( .A1(n13382), .A2(n13381), .A3(n14589), .ZN(n13383) );
  NAND3_X1 U15412 ( .A1(n13385), .A2(n13384), .A3(n13383), .ZN(n13422) );
  MUX2_X1 U15413 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13422), .S(n10988), .Z(
        P2_U3515) );
  AOI21_X1 U15414 ( .B1(n14567), .B2(n13387), .A(n13386), .ZN(n13388) );
  OAI211_X1 U15415 ( .C1(n14571), .C2(n13390), .A(n13389), .B(n13388), .ZN(
        n13423) );
  MUX2_X1 U15416 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13423), .S(n10988), .Z(
        P2_U3514) );
  AOI21_X1 U15417 ( .B1(n14567), .B2(n13392), .A(n13391), .ZN(n13393) );
  OAI211_X1 U15418 ( .C1(n13395), .C2(n14571), .A(n13394), .B(n13393), .ZN(
        n13424) );
  MUX2_X1 U15419 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13424), .S(n10988), .Z(
        P2_U3513) );
  AOI211_X1 U15420 ( .C1(n14567), .C2(n13398), .A(n13397), .B(n13396), .ZN(
        n13399) );
  OAI21_X1 U15421 ( .B1(n14571), .B2(n13400), .A(n13399), .ZN(n13425) );
  MUX2_X1 U15422 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n13425), .S(n10988), .Z(
        P2_U3512) );
  AOI211_X1 U15423 ( .C1(n14567), .C2(n13403), .A(n13402), .B(n13401), .ZN(
        n13404) );
  OAI21_X1 U15424 ( .B1(n14571), .B2(n13405), .A(n13404), .ZN(n13426) );
  MUX2_X1 U15425 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n13426), .S(n10988), .Z(
        P2_U3511) );
  MUX2_X1 U15426 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n13406), .S(n10988), .Z(
        P2_U3501) );
  MUX2_X1 U15427 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13407), .S(n10992), .Z(
        P2_U3498) );
  MUX2_X1 U15428 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13408), .S(n10992), .Z(
        P2_U3497) );
  MUX2_X1 U15429 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13410), .S(n10992), .Z(
        P2_U3495) );
  MUX2_X1 U15430 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13411), .S(n10992), .Z(
        P2_U3494) );
  MUX2_X1 U15431 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13412), .S(n10992), .Z(
        P2_U3493) );
  MUX2_X1 U15432 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13413), .S(n10992), .Z(
        P2_U3492) );
  MUX2_X1 U15433 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13414), .S(n10992), .Z(
        P2_U3491) );
  MUX2_X1 U15434 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13415), .S(n10992), .Z(
        P2_U3490) );
  MUX2_X1 U15435 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13416), .S(n10992), .Z(
        P2_U3489) );
  MUX2_X1 U15436 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13417), .S(n10992), .Z(
        P2_U3488) );
  MUX2_X1 U15437 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13418), .S(n10992), .Z(
        P2_U3487) );
  MUX2_X1 U15438 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13419), .S(n10992), .Z(
        P2_U3486) );
  MUX2_X1 U15439 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13420), .S(n10992), .Z(
        P2_U3484) );
  MUX2_X1 U15440 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13421), .S(n10992), .Z(
        P2_U3481) );
  MUX2_X1 U15441 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13422), .S(n10992), .Z(
        P2_U3478) );
  MUX2_X1 U15442 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13423), .S(n10992), .Z(
        P2_U3475) );
  MUX2_X1 U15443 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13424), .S(n10992), .Z(
        P2_U3472) );
  MUX2_X1 U15444 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n13425), .S(n10992), .Z(
        P2_U3469) );
  MUX2_X1 U15445 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n13426), .S(n10992), .Z(
        P2_U3466) );
  INV_X1 U15446 ( .A(n13427), .ZN(n14002) );
  INV_X1 U15447 ( .A(n13428), .ZN(n13429) );
  NOR4_X1 U15448 ( .A1(n13429), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14924), .A4(
        P2_U3088), .ZN(n13430) );
  AOI21_X1 U15449 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n13431), .A(n13430), 
        .ZN(n13432) );
  OAI21_X1 U15450 ( .B1(n14002), .B2(n13444), .A(n13432), .ZN(P2_U3296) );
  INV_X1 U15451 ( .A(n13433), .ZN(n14006) );
  OAI222_X1 U15452 ( .A1(n13444), .A2(n14006), .B1(n13435), .B2(P2_U3088), 
        .C1(n13434), .C2(n12041), .ZN(P2_U3298) );
  NAND2_X1 U15453 ( .A1(n14008), .A2(n13436), .ZN(n13438) );
  OAI211_X1 U15454 ( .C1(n12041), .C2(n13439), .A(n13438), .B(n13437), .ZN(
        P2_U3299) );
  OAI222_X1 U15455 ( .A1(n13444), .A2(n13440), .B1(n8183), .B2(P2_U3088), .C1(
        n14882), .C2(n12041), .ZN(P2_U3300) );
  INV_X1 U15456 ( .A(n13441), .ZN(n14013) );
  OAI222_X1 U15457 ( .A1(n13444), .A2(n14013), .B1(n13443), .B2(P2_U3088), 
        .C1(n13442), .C2(n12041), .ZN(P2_U3301) );
  INV_X1 U15458 ( .A(n13445), .ZN(n13446) );
  MUX2_X1 U15459 ( .A(n13446), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U15460 ( .A(n13448), .B(n13447), .Z(n13456) );
  AOI22_X1 U15461 ( .A1(n13557), .A2(n13778), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13451) );
  NAND2_X1 U15462 ( .A1(n13576), .A2(n13449), .ZN(n13450) );
  OAI211_X1 U15463 ( .C1(n13452), .C2(n13570), .A(n13451), .B(n13450), .ZN(
        n13453) );
  AOI21_X1 U15464 ( .B1(n13454), .B2(n14142), .A(n13453), .ZN(n13455) );
  OAI21_X1 U15465 ( .B1(n13456), .B2(n13564), .A(n13455), .ZN(P1_U3214) );
  XOR2_X1 U15466 ( .A(n13458), .B(n13457), .Z(n13465) );
  NAND2_X1 U15467 ( .A1(n14292), .A2(n13779), .ZN(n13460) );
  NAND2_X1 U15468 ( .A1(n14131), .A2(n13583), .ZN(n13459) );
  AND2_X1 U15469 ( .A1(n13460), .A2(n13459), .ZN(n13953) );
  OAI22_X1 U15470 ( .A1(n13513), .A2(n13953), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13461), .ZN(n13462) );
  AOI21_X1 U15471 ( .B1(n13817), .B2(n13576), .A(n13462), .ZN(n13464) );
  NAND2_X1 U15472 ( .A1(n13952), .A2(n14142), .ZN(n13463) );
  OAI211_X1 U15473 ( .C1(n13465), .C2(n13564), .A(n13464), .B(n13463), .ZN(
        P1_U3216) );
  NAND2_X1 U15474 ( .A1(n13466), .A2(n13467), .ZN(n13472) );
  NAND2_X1 U15475 ( .A1(n13472), .A2(n13468), .ZN(n13470) );
  AOI21_X1 U15476 ( .B1(n13470), .B2(n13469), .A(n13564), .ZN(n13474) );
  NAND2_X1 U15477 ( .A1(n13472), .A2(n13471), .ZN(n13473) );
  NAND2_X1 U15478 ( .A1(n13474), .A2(n13473), .ZN(n13479) );
  NAND2_X1 U15479 ( .A1(n13557), .A2(n13875), .ZN(n13475) );
  NAND2_X1 U15480 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13730)
         );
  OAI211_X1 U15481 ( .C1(n13476), .C2(n13570), .A(n13475), .B(n13730), .ZN(
        n13477) );
  AOI21_X1 U15482 ( .B1(n13877), .B2(n13576), .A(n13477), .ZN(n13478) );
  OAI211_X1 U15483 ( .C1(n13977), .C2(n13579), .A(n13479), .B(n13478), .ZN(
        P1_U3219) );
  INV_X1 U15484 ( .A(n13480), .ZN(n13481) );
  AOI21_X1 U15485 ( .B1(n13483), .B2(n13482), .A(n13481), .ZN(n13488) );
  AOI22_X1 U15486 ( .A1(n13876), .A2(n14131), .B1(n14292), .B2(n13583), .ZN(
        n13843) );
  OAI22_X1 U15487 ( .A1(n13843), .A2(n13513), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13484), .ZN(n13485) );
  AOI21_X1 U15488 ( .B1(n13846), .B2(n13576), .A(n13485), .ZN(n13487) );
  NAND2_X1 U15489 ( .A1(n13965), .A2(n14142), .ZN(n13486) );
  OAI211_X1 U15490 ( .C1(n13488), .C2(n13564), .A(n13487), .B(n13486), .ZN(
        P1_U3223) );
  XOR2_X1 U15491 ( .A(n13490), .B(n13489), .Z(n13496) );
  AOI22_X1 U15492 ( .A1(n13557), .A2(n13779), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13492) );
  NAND2_X1 U15493 ( .A1(n13576), .A2(n13782), .ZN(n13491) );
  OAI211_X1 U15494 ( .C1(n13493), .C2(n13570), .A(n13492), .B(n13491), .ZN(
        n13494) );
  AOI21_X1 U15495 ( .B1(n13942), .B2(n14142), .A(n13494), .ZN(n13495) );
  OAI21_X1 U15496 ( .B1(n13496), .B2(n13564), .A(n13495), .ZN(P1_U3225) );
  INV_X1 U15497 ( .A(n13497), .ZN(n13498) );
  AOI21_X1 U15498 ( .B1(n13500), .B2(n13499), .A(n13498), .ZN(n13507) );
  OAI21_X1 U15499 ( .B1(n13570), .B2(n13891), .A(n13501), .ZN(n13502) );
  AOI21_X1 U15500 ( .B1(n13557), .B2(n13587), .A(n13502), .ZN(n13503) );
  OAI21_X1 U15501 ( .B1(n13504), .B2(n14146), .A(n13503), .ZN(n13505) );
  AOI21_X1 U15502 ( .B1(n14195), .B2(n14142), .A(n13505), .ZN(n13506) );
  OAI21_X1 U15503 ( .B1(n13507), .B2(n13564), .A(n13506), .ZN(P1_U3226) );
  NAND2_X1 U15504 ( .A1(n13466), .A2(n13508), .ZN(n13547) );
  OAI21_X1 U15505 ( .B1(n13508), .B2(n13466), .A(n13547), .ZN(n13509) );
  NAND2_X1 U15506 ( .A1(n13509), .A2(n14139), .ZN(n13516) );
  INV_X1 U15507 ( .A(n13510), .ZN(n14153) );
  AND2_X1 U15508 ( .A1(n14131), .A2(n13586), .ZN(n13511) );
  AOI21_X1 U15509 ( .B1(n13875), .B2(n14292), .A(n13511), .ZN(n14149) );
  OAI21_X1 U15510 ( .B1(n13513), .B2(n14149), .A(n13512), .ZN(n13514) );
  AOI21_X1 U15511 ( .B1(n14153), .B2(n13576), .A(n13514), .ZN(n13515) );
  OAI211_X1 U15512 ( .C1(n14190), .C2(n13579), .A(n13516), .B(n13515), .ZN(
        P1_U3228) );
  XOR2_X1 U15513 ( .A(n13518), .B(n13517), .Z(n13524) );
  INV_X1 U15514 ( .A(n13799), .ZN(n13521) );
  AOI22_X1 U15515 ( .A1(n13557), .A2(n13827), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13520) );
  NAND2_X1 U15516 ( .A1(n13576), .A2(n13804), .ZN(n13519) );
  OAI211_X1 U15517 ( .C1(n13521), .C2(n13570), .A(n13520), .B(n13519), .ZN(
        n13522) );
  AOI21_X1 U15518 ( .B1(n13805), .B2(n14142), .A(n13522), .ZN(n13523) );
  OAI21_X1 U15519 ( .B1(n13524), .B2(n13564), .A(n13523), .ZN(P1_U3229) );
  OAI21_X1 U15520 ( .B1(n13527), .B2(n13526), .A(n13525), .ZN(n13528) );
  NAND2_X1 U15521 ( .A1(n13528), .A2(n14139), .ZN(n13535) );
  OAI22_X1 U15522 ( .A1(n13570), .A2(n13530), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13529), .ZN(n13533) );
  NOR2_X1 U15523 ( .A1(n13572), .A2(n13531), .ZN(n13532) );
  AOI211_X1 U15524 ( .C1(n13576), .C2(n13833), .A(n13533), .B(n13532), .ZN(
        n13534) );
  OAI211_X1 U15525 ( .C1(n13579), .C2(n13835), .A(n13535), .B(n13534), .ZN(
        P1_U3235) );
  OAI21_X1 U15526 ( .B1(n13538), .B2(n13537), .A(n13536), .ZN(n13539) );
  NAND2_X1 U15527 ( .A1(n13539), .A2(n14139), .ZN(n13545) );
  AOI22_X1 U15528 ( .A1(n13541), .A2(n13596), .B1(n13540), .B2(n14142), .ZN(
        n13544) );
  AOI22_X1 U15529 ( .A1(n13557), .A2(n9761), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n13542), .ZN(n13543) );
  NAND3_X1 U15530 ( .A1(n13545), .A2(n13544), .A3(n13543), .ZN(P1_U3237) );
  NAND2_X1 U15531 ( .A1(n13547), .A2(n13546), .ZN(n13548) );
  XOR2_X1 U15532 ( .A(n13549), .B(n13548), .Z(n13554) );
  NAND2_X1 U15533 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13705)
         );
  OAI21_X1 U15534 ( .B1(n13570), .B2(n13893), .A(n13705), .ZN(n13550) );
  AOI21_X1 U15535 ( .B1(n13557), .B2(n13585), .A(n13550), .ZN(n13551) );
  OAI21_X1 U15536 ( .B1(n13903), .B2(n14146), .A(n13551), .ZN(n13552) );
  AOI21_X1 U15537 ( .B1(n14180), .B2(n14142), .A(n13552), .ZN(n13553) );
  OAI21_X1 U15538 ( .B1(n13554), .B2(n13564), .A(n13553), .ZN(P1_U3238) );
  XOR2_X1 U15539 ( .A(n13556), .B(n13555), .Z(n13565) );
  AOI22_X1 U15540 ( .A1(n13557), .A2(n13799), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13559) );
  NAND2_X1 U15541 ( .A1(n13576), .A2(n13768), .ZN(n13558) );
  OAI211_X1 U15542 ( .C1(n13560), .C2(n13570), .A(n13559), .B(n13558), .ZN(
        n13561) );
  AOI21_X1 U15543 ( .B1(n13562), .B2(n14142), .A(n13561), .ZN(n13563) );
  OAI21_X1 U15544 ( .B1(n13565), .B2(n13564), .A(n13563), .ZN(P1_U3240) );
  OAI211_X1 U15545 ( .C1(n13568), .C2(n13567), .A(n13566), .B(n14139), .ZN(
        n13578) );
  OAI22_X1 U15546 ( .A1(n13570), .A2(n13569), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14977), .ZN(n13574) );
  NOR2_X1 U15547 ( .A1(n13572), .A2(n13571), .ZN(n13573) );
  AOI211_X1 U15548 ( .C1(n13576), .C2(n13575), .A(n13574), .B(n13573), .ZN(
        n13577) );
  OAI211_X1 U15549 ( .C1(n6891), .C2(n13579), .A(n13578), .B(n13577), .ZN(
        P1_U3241) );
  MUX2_X1 U15550 ( .A(n13734), .B(P1_DATAO_REG_31__SCAN_IN), .S(n13615), .Z(
        P1_U3591) );
  MUX2_X1 U15551 ( .A(n13580), .B(P1_DATAO_REG_30__SCAN_IN), .S(n13615), .Z(
        P1_U3590) );
  MUX2_X1 U15552 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13581), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15553 ( .A(n13582), .B(P1_DATAO_REG_28__SCAN_IN), .S(n13615), .Z(
        P1_U3588) );
  MUX2_X1 U15554 ( .A(n13765), .B(P1_DATAO_REG_27__SCAN_IN), .S(n13615), .Z(
        P1_U3587) );
  MUX2_X1 U15555 ( .A(n13778), .B(P1_DATAO_REG_26__SCAN_IN), .S(n13615), .Z(
        P1_U3586) );
  MUX2_X1 U15556 ( .A(n13799), .B(P1_DATAO_REG_25__SCAN_IN), .S(n13615), .Z(
        P1_U3585) );
  MUX2_X1 U15557 ( .A(n13779), .B(P1_DATAO_REG_24__SCAN_IN), .S(n13615), .Z(
        P1_U3584) );
  MUX2_X1 U15558 ( .A(n13827), .B(P1_DATAO_REG_23__SCAN_IN), .S(n13615), .Z(
        P1_U3583) );
  MUX2_X1 U15559 ( .A(n13583), .B(P1_DATAO_REG_22__SCAN_IN), .S(n13615), .Z(
        P1_U3582) );
  MUX2_X1 U15560 ( .A(n13828), .B(P1_DATAO_REG_21__SCAN_IN), .S(n13615), .Z(
        P1_U3581) );
  MUX2_X1 U15561 ( .A(n13876), .B(P1_DATAO_REG_20__SCAN_IN), .S(n13615), .Z(
        P1_U3580) );
  MUX2_X1 U15562 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13584), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15563 ( .A(n13875), .B(P1_DATAO_REG_18__SCAN_IN), .S(n13615), .Z(
        P1_U3578) );
  MUX2_X1 U15564 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13585), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15565 ( .A(n13586), .B(P1_DATAO_REG_16__SCAN_IN), .S(n13615), .Z(
        P1_U3576) );
  MUX2_X1 U15566 ( .A(n13587), .B(P1_DATAO_REG_15__SCAN_IN), .S(n13615), .Z(
        P1_U3575) );
  MUX2_X1 U15567 ( .A(n13588), .B(P1_DATAO_REG_14__SCAN_IN), .S(n13615), .Z(
        P1_U3574) );
  MUX2_X1 U15568 ( .A(n13589), .B(P1_DATAO_REG_13__SCAN_IN), .S(n13615), .Z(
        P1_U3573) );
  MUX2_X1 U15569 ( .A(n14129), .B(P1_DATAO_REG_12__SCAN_IN), .S(n13615), .Z(
        P1_U3572) );
  MUX2_X1 U15570 ( .A(n14291), .B(P1_DATAO_REG_11__SCAN_IN), .S(n13615), .Z(
        P1_U3571) );
  MUX2_X1 U15571 ( .A(n14130), .B(P1_DATAO_REG_10__SCAN_IN), .S(n13615), .Z(
        P1_U3570) );
  MUX2_X1 U15572 ( .A(n13590), .B(P1_DATAO_REG_9__SCAN_IN), .S(n13615), .Z(
        P1_U3569) );
  MUX2_X1 U15573 ( .A(n13591), .B(P1_DATAO_REG_8__SCAN_IN), .S(n13615), .Z(
        P1_U3568) );
  MUX2_X1 U15574 ( .A(n13592), .B(P1_DATAO_REG_7__SCAN_IN), .S(n13615), .Z(
        P1_U3567) );
  MUX2_X1 U15575 ( .A(n13593), .B(P1_DATAO_REG_6__SCAN_IN), .S(n13615), .Z(
        P1_U3566) );
  MUX2_X1 U15576 ( .A(n13594), .B(P1_DATAO_REG_5__SCAN_IN), .S(n13615), .Z(
        P1_U3565) );
  MUX2_X1 U15577 ( .A(n13595), .B(P1_DATAO_REG_4__SCAN_IN), .S(n13615), .Z(
        P1_U3564) );
  MUX2_X1 U15578 ( .A(n13596), .B(P1_DATAO_REG_3__SCAN_IN), .S(n13615), .Z(
        P1_U3563) );
  MUX2_X1 U15579 ( .A(n13597), .B(P1_DATAO_REG_2__SCAN_IN), .S(n13615), .Z(
        P1_U3562) );
  MUX2_X1 U15580 ( .A(n9761), .B(P1_DATAO_REG_1__SCAN_IN), .S(n13615), .Z(
        P1_U3561) );
  MUX2_X1 U15581 ( .A(n13598), .B(P1_DATAO_REG_0__SCAN_IN), .S(n13615), .Z(
        P1_U3560) );
  OAI22_X1 U15582 ( .A1(n14278), .A2(n13600), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13599), .ZN(n13601) );
  AOI21_X1 U15583 ( .B1(n13602), .B2(n13723), .A(n13601), .ZN(n13612) );
  OAI21_X1 U15584 ( .B1(n9753), .B2(n13617), .A(n13603), .ZN(n13604) );
  NAND3_X1 U15585 ( .A1(n13726), .A2(n13628), .A3(n13604), .ZN(n13611) );
  MUX2_X1 U15586 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n13606), .S(n13605), .Z(
        n13607) );
  NAND2_X1 U15587 ( .A1(n13607), .A2(n13614), .ZN(n13608) );
  NAND3_X1 U15588 ( .A1(n13725), .A2(n13609), .A3(n13608), .ZN(n13610) );
  NAND3_X1 U15589 ( .A1(n13612), .A2(n13611), .A3(n13610), .ZN(P1_U3244) );
  MUX2_X1 U15590 ( .A(n13614), .B(n13613), .S(n8847), .Z(n13619) );
  AOI21_X1 U15591 ( .B1(n13617), .B2(n13616), .A(n13615), .ZN(n13618) );
  OAI21_X1 U15592 ( .B1(n13619), .B2(n14009), .A(n13618), .ZN(n13651) );
  AOI22_X1 U15593 ( .A1(n13708), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n13633) );
  INV_X1 U15594 ( .A(n13620), .ZN(n13622) );
  XNOR2_X1 U15595 ( .A(n13622), .B(n13621), .ZN(n13624) );
  AOI22_X1 U15596 ( .A1(n13725), .A2(n13624), .B1(n13723), .B2(n13623), .ZN(
        n13632) );
  INV_X1 U15597 ( .A(n13625), .ZN(n13630) );
  NAND3_X1 U15598 ( .A1(n13628), .A2(n13627), .A3(n13626), .ZN(n13629) );
  NAND3_X1 U15599 ( .A1(n13726), .A2(n13630), .A3(n13629), .ZN(n13631) );
  NAND4_X1 U15600 ( .A1(n13651), .A2(n13633), .A3(n13632), .A4(n13631), .ZN(
        P1_U3245) );
  NAND2_X1 U15601 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n13708), .ZN(n13650) );
  AND3_X1 U15602 ( .A1(n13636), .A2(n13635), .A3(n13634), .ZN(n13637) );
  NOR3_X1 U15603 ( .A1(n14272), .A2(n13638), .A3(n13637), .ZN(n13648) );
  OAI21_X1 U15604 ( .B1(n14274), .B2(n13640), .A(n13639), .ZN(n13647) );
  INV_X1 U15605 ( .A(n13663), .ZN(n13645) );
  NOR3_X1 U15606 ( .A1(n13643), .A2(n13642), .A3(n13641), .ZN(n13644) );
  NOR3_X1 U15607 ( .A1(n14270), .A2(n13645), .A3(n13644), .ZN(n13646) );
  NOR3_X1 U15608 ( .A1(n13648), .A2(n13647), .A3(n13646), .ZN(n13649) );
  NAND3_X1 U15609 ( .A1(n13651), .A2(n13650), .A3(n13649), .ZN(P1_U3247) );
  OAI21_X1 U15610 ( .B1(n14278), .B2(n13653), .A(n13652), .ZN(n13654) );
  AOI21_X1 U15611 ( .B1(n13655), .B2(n13723), .A(n13654), .ZN(n13668) );
  OAI21_X1 U15612 ( .B1(n13658), .B2(n13657), .A(n13656), .ZN(n13659) );
  NAND2_X1 U15613 ( .A1(n13726), .A2(n13659), .ZN(n13667) );
  INV_X1 U15614 ( .A(n13660), .ZN(n13665) );
  NAND3_X1 U15615 ( .A1(n13663), .A2(n13662), .A3(n13661), .ZN(n13664) );
  NAND3_X1 U15616 ( .A1(n13725), .A2(n13665), .A3(n13664), .ZN(n13666) );
  NAND3_X1 U15617 ( .A1(n13668), .A2(n13667), .A3(n13666), .ZN(P1_U3248) );
  OAI21_X1 U15618 ( .B1(n13670), .B2(n13669), .A(n13685), .ZN(n13671) );
  NAND2_X1 U15619 ( .A1(n13671), .A2(n13726), .ZN(n13682) );
  INV_X1 U15620 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n13672) );
  NAND2_X1 U15621 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14143)
         );
  OAI21_X1 U15622 ( .B1(n14278), .B2(n13672), .A(n14143), .ZN(n13673) );
  AOI21_X1 U15623 ( .B1(n13674), .B2(n13723), .A(n13673), .ZN(n13681) );
  OR3_X1 U15624 ( .A1(n13677), .A2(n13676), .A3(n13675), .ZN(n13678) );
  NAND3_X1 U15625 ( .A1(n13679), .A2(n13725), .A3(n13678), .ZN(n13680) );
  NAND3_X1 U15626 ( .A1(n13682), .A2(n13681), .A3(n13680), .ZN(P1_U3254) );
  AND3_X1 U15627 ( .A1(n13685), .A2(n13684), .A3(n13683), .ZN(n13686) );
  OAI21_X1 U15628 ( .B1(n13687), .B2(n13686), .A(n13726), .ZN(n13698) );
  NOR2_X1 U15629 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13688), .ZN(n13689) );
  AOI21_X1 U15630 ( .B1(n13708), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n13689), 
        .ZN(n13697) );
  AOI21_X1 U15631 ( .B1(n13692), .B2(n13691), .A(n13690), .ZN(n13693) );
  OR2_X1 U15632 ( .A1(n13693), .A2(n14270), .ZN(n13696) );
  NAND2_X1 U15633 ( .A1(n13723), .A2(n13694), .ZN(n13695) );
  NAND4_X1 U15634 ( .A1(n13698), .A2(n13697), .A3(n13696), .A4(n13695), .ZN(
        P1_U3255) );
  NAND2_X1 U15635 ( .A1(n13700), .A2(n13699), .ZN(n13718) );
  XNOR2_X1 U15636 ( .A(n13718), .B(n13711), .ZN(n13716) );
  XNOR2_X1 U15637 ( .A(n13716), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n13710) );
  INV_X1 U15638 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14193) );
  XNOR2_X1 U15639 ( .A(n13712), .B(n13711), .ZN(n13703) );
  NAND2_X1 U15640 ( .A1(n13703), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n13714) );
  OAI211_X1 U15641 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n13703), .A(n13726), 
        .B(n13714), .ZN(n13704) );
  NAND2_X1 U15642 ( .A1(n13705), .A2(n13704), .ZN(n13707) );
  NOR2_X1 U15643 ( .A1(n14274), .A2(n13711), .ZN(n13706) );
  AOI211_X1 U15644 ( .C1(n13708), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n13707), 
        .B(n13706), .ZN(n13709) );
  OAI21_X1 U15645 ( .B1(n13710), .B2(n14270), .A(n13709), .ZN(P1_U3261) );
  INV_X1 U15646 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n14851) );
  INV_X1 U15647 ( .A(n13711), .ZN(n13717) );
  NAND2_X1 U15648 ( .A1(n13712), .A2(n13717), .ZN(n13713) );
  NAND2_X1 U15649 ( .A1(n13714), .A2(n13713), .ZN(n13715) );
  NAND2_X1 U15650 ( .A1(n13716), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n13720) );
  NAND2_X1 U15651 ( .A1(n13718), .A2(n13717), .ZN(n13719) );
  NAND2_X1 U15652 ( .A1(n13720), .A2(n13719), .ZN(n13721) );
  XOR2_X1 U15653 ( .A(n13721), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13724) );
  NOR2_X1 U15654 ( .A1(n13724), .A2(n14270), .ZN(n13722) );
  AOI211_X1 U15655 ( .C1(n6607), .C2(n13726), .A(n13723), .B(n13722), .ZN(
        n13729) );
  AOI22_X1 U15656 ( .A1(n13727), .A2(n13726), .B1(n13725), .B2(n13724), .ZN(
        n13728) );
  MUX2_X1 U15657 ( .A(n13729), .B(n13728), .S(n10556), .Z(n13731) );
  OAI211_X1 U15658 ( .C1(n14851), .C2(n14278), .A(n13731), .B(n13730), .ZN(
        P1_U3262) );
  NAND2_X1 U15659 ( .A1(n13739), .A2(n13915), .ZN(n13733) );
  NAND2_X1 U15660 ( .A1(n13735), .A2(n13734), .ZN(n13913) );
  NOR2_X1 U15661 ( .A1(n13880), .A2(n13913), .ZN(n13742) );
  AOI21_X1 U15662 ( .B1(n13880), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13742), 
        .ZN(n13737) );
  NAND2_X1 U15663 ( .A1(n13732), .A2(n14306), .ZN(n13736) );
  OAI211_X1 U15664 ( .C1(n13912), .C2(n13907), .A(n13737), .B(n13736), .ZN(
        P1_U3263) );
  XNOR2_X1 U15665 ( .A(n13739), .B(n13738), .ZN(n13740) );
  NAND2_X1 U15666 ( .A1(n13740), .A2(n14310), .ZN(n13914) );
  NOR2_X1 U15667 ( .A1(n13915), .A2(n13883), .ZN(n13741) );
  AOI211_X1 U15668 ( .C1(n13880), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13742), 
        .B(n13741), .ZN(n13743) );
  OAI21_X1 U15669 ( .B1(n14160), .B2(n13914), .A(n13743), .ZN(P1_U3264) );
  XNOR2_X1 U15670 ( .A(n13744), .B(n13746), .ZN(n13924) );
  OAI21_X1 U15671 ( .B1(n13747), .B2(n13746), .A(n13745), .ZN(n13929) );
  INV_X1 U15672 ( .A(n13926), .ZN(n13751) );
  NAND2_X1 U15673 ( .A1(n14284), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n13750) );
  NAND2_X1 U15674 ( .A1(n14285), .A2(n13748), .ZN(n13749) );
  OAI211_X1 U15675 ( .C1(n14318), .C2(n13751), .A(n13750), .B(n13749), .ZN(
        n13752) );
  AOI21_X1 U15676 ( .B1(n13927), .B2(n14306), .A(n13752), .ZN(n13757) );
  AOI21_X1 U15677 ( .B1(n13927), .B2(n13753), .A(n14182), .ZN(n13755) );
  NAND2_X1 U15678 ( .A1(n13925), .A2(n14314), .ZN(n13756) );
  OAI211_X1 U15679 ( .C1(n13929), .C2(n13887), .A(n13757), .B(n13756), .ZN(
        n13758) );
  AOI21_X1 U15680 ( .B1(n13885), .B2(n13924), .A(n13758), .ZN(n13759) );
  INV_X1 U15681 ( .A(n13759), .ZN(P1_U3265) );
  XNOR2_X1 U15682 ( .A(n13761), .B(n13760), .ZN(n13940) );
  OAI21_X1 U15683 ( .B1(n13763), .B2(n13762), .A(n12043), .ZN(n13938) );
  OAI211_X1 U15684 ( .C1(n13936), .C2(n13781), .A(n14310), .B(n13764), .ZN(
        n13935) );
  NAND2_X1 U15685 ( .A1(n14292), .A2(n13765), .ZN(n13767) );
  NAND2_X1 U15686 ( .A1(n14131), .A2(n13799), .ZN(n13766) );
  AND2_X1 U15687 ( .A1(n13767), .A2(n13766), .ZN(n13934) );
  INV_X1 U15688 ( .A(n13768), .ZN(n13769) );
  OAI22_X1 U15689 ( .A1(n13880), .A2(n13934), .B1(n13769), .B2(n14302), .ZN(
        n13771) );
  NOR2_X1 U15690 ( .A1(n13936), .A2(n13883), .ZN(n13770) );
  AOI211_X1 U15691 ( .C1(n13880), .C2(P1_REG2_REG_26__SCAN_IN), .A(n13771), 
        .B(n13770), .ZN(n13772) );
  OAI21_X1 U15692 ( .B1(n14160), .B2(n13935), .A(n13772), .ZN(n13773) );
  AOI21_X1 U15693 ( .B1(n13938), .B2(n13885), .A(n13773), .ZN(n13774) );
  OAI21_X1 U15694 ( .B1(n13887), .B2(n13940), .A(n13774), .ZN(P1_U3267) );
  AND2_X1 U15695 ( .A1(n13798), .A2(n13775), .ZN(n13777) );
  OAI21_X1 U15696 ( .B1(n13777), .B2(n13785), .A(n13776), .ZN(n13780) );
  AOI222_X1 U15697 ( .A1(n14353), .A2(n13780), .B1(n13779), .B2(n14131), .C1(
        n13778), .C2(n14292), .ZN(n13944) );
  AOI211_X1 U15698 ( .C1(n13942), .C2(n6487), .A(n14182), .B(n13781), .ZN(
        n13941) );
  AOI22_X1 U15699 ( .A1(n14284), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n13782), 
        .B2(n14285), .ZN(n13783) );
  OAI21_X1 U15700 ( .B1(n13784), .B2(n13883), .A(n13783), .ZN(n13790) );
  NAND2_X1 U15701 ( .A1(n13786), .A2(n13785), .ZN(n13787) );
  NAND2_X1 U15702 ( .A1(n13788), .A2(n13787), .ZN(n13945) );
  NOR2_X1 U15703 ( .A1(n13945), .A2(n13887), .ZN(n13789) );
  AOI211_X1 U15704 ( .C1(n13941), .C2(n14314), .A(n13790), .B(n13789), .ZN(
        n13791) );
  OAI21_X1 U15705 ( .B1(n13944), .B2(n14284), .A(n13791), .ZN(P1_U3268) );
  XNOR2_X1 U15706 ( .A(n13792), .B(n13793), .ZN(n13794) );
  NAND2_X1 U15707 ( .A1(n13794), .A2(n14375), .ZN(n13802) );
  NAND2_X1 U15708 ( .A1(n13796), .A2(n13795), .ZN(n13797) );
  NAND3_X1 U15709 ( .A1(n13798), .A2(n14353), .A3(n13797), .ZN(n13801) );
  AOI22_X1 U15710 ( .A1(n14292), .A2(n13799), .B1(n14131), .B2(n13827), .ZN(
        n13800) );
  NAND3_X1 U15711 ( .A1(n13802), .A2(n13801), .A3(n13800), .ZN(n13949) );
  AOI21_X1 U15712 ( .B1(n13816), .B2(n13805), .A(n14182), .ZN(n13803) );
  NAND2_X1 U15713 ( .A1(n13803), .A2(n6487), .ZN(n13946) );
  AOI22_X1 U15714 ( .A1(n14284), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n13804), 
        .B2(n14285), .ZN(n13807) );
  NAND2_X1 U15715 ( .A1(n13805), .A2(n14306), .ZN(n13806) );
  OAI211_X1 U15716 ( .C1(n13946), .C2(n14160), .A(n13807), .B(n13806), .ZN(
        n13808) );
  AOI21_X1 U15717 ( .B1(n13949), .B2(n14303), .A(n13808), .ZN(n13809) );
  INV_X1 U15718 ( .A(n13809), .ZN(P1_U3269) );
  XNOR2_X1 U15719 ( .A(n13811), .B(n13813), .ZN(n13958) );
  OAI21_X1 U15720 ( .B1(n13814), .B2(n13813), .A(n13812), .ZN(n13956) );
  NAND2_X1 U15721 ( .A1(n13831), .A2(n13952), .ZN(n13815) );
  NAND3_X1 U15722 ( .A1(n13816), .A2(n14310), .A3(n13815), .ZN(n13954) );
  INV_X1 U15723 ( .A(n13817), .ZN(n13818) );
  OAI21_X1 U15724 ( .B1(n14302), .B2(n13818), .A(n13953), .ZN(n13819) );
  INV_X1 U15725 ( .A(n13819), .ZN(n13821) );
  NAND2_X1 U15726 ( .A1(n14284), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n13820) );
  OAI21_X1 U15727 ( .B1(n14318), .B2(n13821), .A(n13820), .ZN(n13822) );
  AOI21_X1 U15728 ( .B1(n13952), .B2(n14306), .A(n13822), .ZN(n13823) );
  OAI21_X1 U15729 ( .B1(n13954), .B2(n14160), .A(n13823), .ZN(n13824) );
  AOI21_X1 U15730 ( .B1(n13956), .B2(n13885), .A(n13824), .ZN(n13825) );
  OAI21_X1 U15731 ( .B1(n13887), .B2(n13958), .A(n13825), .ZN(P1_U3270) );
  XNOR2_X1 U15732 ( .A(n13826), .B(n13837), .ZN(n13829) );
  AOI222_X1 U15733 ( .A1(n14353), .A2(n13829), .B1(n13828), .B2(n14131), .C1(
        n13827), .C2(n14292), .ZN(n13962) );
  INV_X1 U15734 ( .A(n13831), .ZN(n13832) );
  AOI211_X1 U15735 ( .C1(n13960), .C2(n6888), .A(n14182), .B(n13832), .ZN(
        n13959) );
  AOI22_X1 U15736 ( .A1(n14284), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n13833), 
        .B2(n14285), .ZN(n13834) );
  OAI21_X1 U15737 ( .B1(n13835), .B2(n13883), .A(n13834), .ZN(n13839) );
  XOR2_X1 U15738 ( .A(n13836), .B(n13837), .Z(n13963) );
  NOR2_X1 U15739 ( .A1(n13963), .A2(n13887), .ZN(n13838) );
  AOI211_X1 U15740 ( .C1(n13959), .C2(n14314), .A(n13839), .B(n13838), .ZN(
        n13840) );
  OAI21_X1 U15741 ( .B1(n13880), .B2(n13962), .A(n13840), .ZN(P1_U3271) );
  XNOR2_X1 U15742 ( .A(n13841), .B(n13842), .ZN(n13845) );
  INV_X1 U15743 ( .A(n13843), .ZN(n13844) );
  AOI21_X1 U15744 ( .B1(n13845), .B2(n14353), .A(n13844), .ZN(n13967) );
  AOI211_X1 U15745 ( .C1(n13965), .C2(n13860), .A(n14182), .B(n13830), .ZN(
        n13964) );
  INV_X1 U15746 ( .A(n13965), .ZN(n13848) );
  AOI22_X1 U15747 ( .A1(n14284), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n13846), 
        .B2(n14285), .ZN(n13847) );
  OAI21_X1 U15748 ( .B1(n13848), .B2(n13883), .A(n13847), .ZN(n13852) );
  AOI21_X1 U15749 ( .B1(n13850), .B2(n13849), .A(n6516), .ZN(n13968) );
  NOR2_X1 U15750 ( .A1(n13968), .A2(n13887), .ZN(n13851) );
  AOI211_X1 U15751 ( .C1(n13964), .C2(n14314), .A(n13852), .B(n13851), .ZN(
        n13853) );
  OAI21_X1 U15752 ( .B1(n13880), .B2(n13967), .A(n13853), .ZN(P1_U3272) );
  OAI21_X1 U15753 ( .B1(n13855), .B2(n13859), .A(n13854), .ZN(n13975) );
  INV_X1 U15754 ( .A(n13856), .ZN(n13857) );
  AOI21_X1 U15755 ( .B1(n13859), .B2(n13858), .A(n13857), .ZN(n13973) );
  NAND2_X1 U15756 ( .A1(n13973), .A2(n14315), .ZN(n13867) );
  OAI211_X1 U15757 ( .C1(n13971), .C2(n13873), .A(n14310), .B(n13860), .ZN(
        n13970) );
  INV_X1 U15758 ( .A(n13970), .ZN(n13865) );
  OAI22_X1 U15759 ( .A1(n13969), .A2(n14284), .B1(n13861), .B2(n14302), .ZN(
        n13862) );
  AOI21_X1 U15760 ( .B1(P1_REG2_REG_20__SCAN_IN), .B2(n14284), .A(n13862), 
        .ZN(n13863) );
  OAI21_X1 U15761 ( .B1(n13971), .B2(n13883), .A(n13863), .ZN(n13864) );
  AOI21_X1 U15762 ( .B1(n13865), .B2(n14314), .A(n13864), .ZN(n13866) );
  OAI211_X1 U15763 ( .C1(n13975), .C2(n13868), .A(n13867), .B(n13866), .ZN(
        P1_U3273) );
  XNOR2_X1 U15764 ( .A(n13869), .B(n13871), .ZN(n13982) );
  OAI21_X1 U15765 ( .B1(n13872), .B2(n13871), .A(n13870), .ZN(n13980) );
  AOI211_X1 U15766 ( .C1(n13874), .C2(n13902), .A(n14182), .B(n13873), .ZN(
        n13979) );
  NAND2_X1 U15767 ( .A1(n13979), .A2(n14314), .ZN(n13882) );
  AOI22_X1 U15768 ( .A1(n13876), .A2(n14292), .B1(n14131), .B2(n13875), .ZN(
        n13976) );
  INV_X1 U15769 ( .A(n13877), .ZN(n13878) );
  OAI22_X1 U15770 ( .A1(n13976), .A2(n14284), .B1(n13878), .B2(n14302), .ZN(
        n13879) );
  AOI21_X1 U15771 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(n13880), .A(n13879), 
        .ZN(n13881) );
  OAI211_X1 U15772 ( .C1(n13977), .C2(n13883), .A(n13882), .B(n13881), .ZN(
        n13884) );
  AOI21_X1 U15773 ( .B1(n13980), .B2(n13885), .A(n13884), .ZN(n13886) );
  OAI21_X1 U15774 ( .B1(n13982), .B2(n13887), .A(n13886), .ZN(P1_U3274) );
  XNOR2_X1 U15775 ( .A(n13888), .B(n11847), .ZN(n13889) );
  NAND2_X1 U15776 ( .A1(n13889), .A2(n14353), .ZN(n13896) );
  OAI22_X1 U15777 ( .A1(n13893), .A2(n13892), .B1(n13891), .B2(n13890), .ZN(
        n13894) );
  INV_X1 U15778 ( .A(n13894), .ZN(n13895) );
  NAND2_X1 U15779 ( .A1(n13896), .A2(n13895), .ZN(n14186) );
  INV_X1 U15780 ( .A(n14186), .ZN(n13910) );
  NAND2_X1 U15781 ( .A1(n13898), .A2(n13897), .ZN(n13899) );
  NAND2_X1 U15782 ( .A1(n13900), .A2(n13899), .ZN(n14179) );
  NAND2_X1 U15783 ( .A1(n14158), .A2(n14180), .ZN(n13901) );
  NAND2_X1 U15784 ( .A1(n13902), .A2(n13901), .ZN(n14183) );
  INV_X1 U15785 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n13904) );
  OAI22_X1 U15786 ( .A1(n14303), .A2(n13904), .B1(n13903), .B2(n14302), .ZN(
        n13905) );
  AOI21_X1 U15787 ( .B1(n14180), .B2(n14306), .A(n13905), .ZN(n13906) );
  OAI21_X1 U15788 ( .B1(n14183), .B2(n13907), .A(n13906), .ZN(n13908) );
  AOI21_X1 U15789 ( .B1(n14179), .B2(n14315), .A(n13908), .ZN(n13909) );
  OAI21_X1 U15790 ( .B1(n13910), .B2(n14284), .A(n13909), .ZN(P1_U3275) );
  NAND2_X1 U15791 ( .A1(n13732), .A2(n14345), .ZN(n13911) );
  OAI211_X1 U15792 ( .C1(n13912), .C2(n14182), .A(n13911), .B(n13913), .ZN(
        n13983) );
  MUX2_X1 U15793 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n13983), .S(n14391), .Z(
        P1_U3559) );
  OAI211_X1 U15794 ( .C1(n13915), .C2(n14371), .A(n13914), .B(n13913), .ZN(
        n13984) );
  MUX2_X1 U15795 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n13984), .S(n14391), .Z(
        P1_U3558) );
  OAI211_X1 U15796 ( .C1(n13919), .C2(n14371), .A(n13918), .B(n13917), .ZN(
        n13920) );
  OAI211_X1 U15797 ( .C1(n13923), .C2(n14349), .A(n13922), .B(n7357), .ZN(
        n13985) );
  MUX2_X1 U15798 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n13985), .S(n14391), .Z(
        P1_U3557) );
  NAND2_X1 U15799 ( .A1(n13924), .A2(n14353), .ZN(n13928) );
  MUX2_X1 U15800 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n13986), .S(n14391), .Z(
        P1_U3556) );
  NAND2_X1 U15801 ( .A1(n13933), .A2(n13932), .ZN(n13987) );
  MUX2_X1 U15802 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n13987), .S(n14391), .Z(
        P1_U3555) );
  OAI211_X1 U15803 ( .C1(n13936), .C2(n14371), .A(n13935), .B(n13934), .ZN(
        n13937) );
  AOI21_X1 U15804 ( .B1(n13938), .B2(n14353), .A(n13937), .ZN(n13939) );
  OAI21_X1 U15805 ( .B1(n14349), .B2(n13940), .A(n13939), .ZN(n13988) );
  MUX2_X1 U15806 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n13988), .S(n14391), .Z(
        P1_U3554) );
  AOI21_X1 U15807 ( .B1(n14345), .B2(n13942), .A(n13941), .ZN(n13943) );
  OAI211_X1 U15808 ( .C1(n14349), .C2(n13945), .A(n13944), .B(n13943), .ZN(
        n13989) );
  MUX2_X1 U15809 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n13989), .S(n14391), .Z(
        P1_U3553) );
  OAI21_X1 U15810 ( .B1(n13947), .B2(n14371), .A(n13946), .ZN(n13948) );
  NOR2_X1 U15811 ( .A1(n13949), .A2(n13948), .ZN(n13990) );
  INV_X1 U15812 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n13950) );
  MUX2_X1 U15813 ( .A(n13990), .B(n13950), .S(n14388), .Z(n13951) );
  INV_X1 U15814 ( .A(n13951), .ZN(P1_U3552) );
  OAI211_X1 U15815 ( .C1(n6884), .C2(n14371), .A(n13954), .B(n13953), .ZN(
        n13955) );
  AOI21_X1 U15816 ( .B1(n13956), .B2(n14353), .A(n13955), .ZN(n13957) );
  OAI21_X1 U15817 ( .B1(n14349), .B2(n13958), .A(n13957), .ZN(n13993) );
  MUX2_X1 U15818 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n13993), .S(n14391), .Z(
        P1_U3551) );
  AOI21_X1 U15819 ( .B1(n14345), .B2(n13960), .A(n13959), .ZN(n13961) );
  OAI211_X1 U15820 ( .C1(n13963), .C2(n14349), .A(n13962), .B(n13961), .ZN(
        n13994) );
  MUX2_X1 U15821 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n13994), .S(n14391), .Z(
        P1_U3550) );
  AOI21_X1 U15822 ( .B1(n14345), .B2(n13965), .A(n13964), .ZN(n13966) );
  OAI211_X1 U15823 ( .C1(n13968), .C2(n14349), .A(n13967), .B(n13966), .ZN(
        n13995) );
  MUX2_X1 U15824 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n13995), .S(n14391), .Z(
        P1_U3549) );
  OAI211_X1 U15825 ( .C1(n13971), .C2(n14371), .A(n13970), .B(n13969), .ZN(
        n13972) );
  AOI21_X1 U15826 ( .B1(n13973), .B2(n14375), .A(n13972), .ZN(n13974) );
  OAI21_X1 U15827 ( .B1(n14357), .B2(n13975), .A(n13974), .ZN(n13996) );
  MUX2_X1 U15828 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n13996), .S(n14391), .Z(
        P1_U3548) );
  OAI21_X1 U15829 ( .B1(n13977), .B2(n14371), .A(n13976), .ZN(n13978) );
  AOI211_X1 U15830 ( .C1(n13980), .C2(n14353), .A(n13979), .B(n13978), .ZN(
        n13981) );
  OAI21_X1 U15831 ( .B1(n13982), .B2(n14349), .A(n13981), .ZN(n13997) );
  MUX2_X1 U15832 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n13997), .S(n14391), .Z(
        P1_U3547) );
  MUX2_X1 U15833 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n13983), .S(n14378), .Z(
        P1_U3527) );
  MUX2_X1 U15834 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n13984), .S(n14378), .Z(
        P1_U3526) );
  MUX2_X1 U15835 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n13985), .S(n14378), .Z(
        P1_U3525) );
  MUX2_X1 U15836 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n13986), .S(n14378), .Z(
        P1_U3524) );
  MUX2_X1 U15837 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n13987), .S(n14378), .Z(
        P1_U3523) );
  MUX2_X1 U15838 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n13988), .S(n14378), .Z(
        P1_U3522) );
  MUX2_X1 U15839 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n13989), .S(n14378), .Z(
        P1_U3521) );
  INV_X1 U15840 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n13991) );
  MUX2_X1 U15841 ( .A(n13991), .B(n13990), .S(n14378), .Z(n13992) );
  INV_X1 U15842 ( .A(n13992), .ZN(P1_U3520) );
  MUX2_X1 U15843 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n13993), .S(n14378), .Z(
        P1_U3519) );
  MUX2_X1 U15844 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n13994), .S(n14378), .Z(
        P1_U3518) );
  MUX2_X1 U15845 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n13995), .S(n14378), .Z(
        P1_U3517) );
  MUX2_X1 U15846 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n13996), .S(n14378), .Z(
        P1_U3516) );
  MUX2_X1 U15847 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n13997), .S(n14378), .Z(
        P1_U3515) );
  INV_X1 U15848 ( .A(n8776), .ZN(n13998) );
  NOR4_X1 U15849 ( .A1(n13998), .A2(P1_IR_REG_30__SCAN_IN), .A3(n6613), .A4(
        P1_U3086), .ZN(n13999) );
  AOI21_X1 U15850 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n14000), .A(n13999), 
        .ZN(n14001) );
  OAI21_X1 U15851 ( .B1(n14002), .B2(n14014), .A(n14001), .ZN(P1_U3324) );
  OAI222_X1 U15852 ( .A1(n14012), .A2(n14879), .B1(n14014), .B2(n14004), .C1(
        n14003), .C2(P1_U3086), .ZN(P1_U3325) );
  OAI222_X1 U15853 ( .A1(n14012), .A2(n14007), .B1(n14014), .B2(n14006), .C1(
        n14005), .C2(P1_U3086), .ZN(P1_U3326) );
  INV_X1 U15854 ( .A(n14008), .ZN(n14010) );
  OAI222_X1 U15855 ( .A1(n14012), .A2(n14011), .B1(n14014), .B2(n14010), .C1(
        P1_U3086), .C2(n14009), .ZN(P1_U3327) );
  OAI222_X1 U15856 ( .A1(n14015), .A2(P1_U3086), .B1(n14014), .B2(n14013), 
        .C1(n6674), .C2(n14012), .ZN(P1_U3329) );
  MUX2_X1 U15857 ( .A(n14017), .B(n14016), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U15858 ( .A(n14018), .ZN(n14019) );
  MUX2_X1 U15859 ( .A(n14019), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U15860 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14020), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U15861 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14021) );
  OAI21_X1 U15862 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14021), 
        .ZN(U28) );
  AOI21_X1 U15863 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14022) );
  OAI21_X1 U15864 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14022), 
        .ZN(U29) );
  AOI22_X1 U15865 ( .A1(n14023), .A2(n14038), .B1(SI_17_), .B2(n14037), .ZN(
        n14024) );
  OAI21_X1 U15866 ( .B1(P3_U3151), .B2(n14025), .A(n14024), .ZN(P3_U3278) );
  AOI21_X1 U15867 ( .B1(n14028), .B2(n14027), .A(n14026), .ZN(n14029) );
  XOR2_X1 U15868 ( .A(n14029), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  INV_X1 U15869 ( .A(n14030), .ZN(n14031) );
  AOI22_X1 U15870 ( .A1(n14031), .A2(n14038), .B1(SI_10_), .B2(n14037), .ZN(
        n14032) );
  OAI21_X1 U15871 ( .B1(P3_U3151), .B2(n14033), .A(n14032), .ZN(P3_U3285) );
  XOR2_X1 U15872 ( .A(n14035), .B(n14034), .Z(SUB_1596_U57) );
  XNOR2_X1 U15873 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14036), .ZN(SUB_1596_U55)
         );
  AOI22_X1 U15874 ( .A1(n14039), .A2(n14038), .B1(SI_18_), .B2(n14037), .ZN(
        n14040) );
  OAI21_X1 U15875 ( .B1(P3_U3151), .B2(n14041), .A(n14040), .ZN(P3_U3277) );
  XOR2_X1 U15876 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14043), .Z(SUB_1596_U54) );
  OAI21_X1 U15877 ( .B1(n14046), .B2(n14045), .A(n14044), .ZN(n14048) );
  XOR2_X1 U15878 ( .A(n14048), .B(n14047), .Z(SUB_1596_U70) );
  OAI21_X1 U15879 ( .B1(n14051), .B2(n14050), .A(n14049), .ZN(n14053) );
  XOR2_X1 U15880 ( .A(n14053), .B(n14052), .Z(SUB_1596_U63) );
  AOI22_X1 U15881 ( .A1(n14718), .A2(n14054), .B1(n14743), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n14070) );
  INV_X1 U15882 ( .A(n14055), .ZN(n14057) );
  NAND2_X1 U15883 ( .A1(n14057), .A2(n14056), .ZN(n14058) );
  XNOR2_X1 U15884 ( .A(n14059), .B(n14058), .ZN(n14064) );
  OAI21_X1 U15885 ( .B1(n14062), .B2(n14061), .A(n14060), .ZN(n14063) );
  AOI22_X1 U15886 ( .A1(n14064), .A2(n14735), .B1(n14746), .B2(n14063), .ZN(
        n14069) );
  NAND2_X1 U15887 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n14068)
         );
  OAI221_X1 U15888 ( .B1(n14066), .B2(n6565), .C1(n14066), .C2(n14065), .A(
        n14080), .ZN(n14067) );
  NAND4_X1 U15889 ( .A1(n14070), .A2(n14069), .A3(n14068), .A4(n14067), .ZN(
        P3_U3198) );
  AOI22_X1 U15890 ( .A1(n14718), .A2(n14071), .B1(n14743), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14087) );
  OAI21_X1 U15891 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n14073), .A(n14072), 
        .ZN(n14078) );
  AOI211_X1 U15892 ( .C1(n14076), .C2(n14075), .A(n14709), .B(n14074), .ZN(
        n14077) );
  AOI21_X1 U15893 ( .B1(n14746), .B2(n14078), .A(n14077), .ZN(n14086) );
  NAND2_X1 U15894 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_U3151), .ZN(n14085)
         );
  OAI221_X1 U15895 ( .B1(n14083), .B2(n14082), .C1(n14083), .C2(n14081), .A(
        n14080), .ZN(n14084) );
  NAND4_X1 U15896 ( .A1(n14087), .A2(n14086), .A3(n14085), .A4(n14084), .ZN(
        P3_U3199) );
  AOI21_X1 U15897 ( .B1(n14089), .B2(n14812), .A(n14092), .ZN(n14112) );
  INV_X1 U15898 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14090) );
  AOI22_X1 U15899 ( .A1(n14846), .A2(n14112), .B1(n14090), .B2(n14844), .ZN(
        P3_U3490) );
  INV_X1 U15900 ( .A(n14091), .ZN(n14093) );
  AOI21_X1 U15901 ( .B1(n14812), .B2(n14093), .A(n14092), .ZN(n14113) );
  INV_X1 U15902 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14094) );
  AOI22_X1 U15903 ( .A1(n14846), .A2(n14113), .B1(n14094), .B2(n14844), .ZN(
        P3_U3489) );
  OAI22_X1 U15904 ( .A1(n14096), .A2(n14828), .B1(n14827), .B2(n14095), .ZN(
        n14097) );
  NOR2_X1 U15905 ( .A1(n14098), .A2(n14097), .ZN(n14115) );
  INV_X1 U15906 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14099) );
  AOI22_X1 U15907 ( .A1(n14846), .A2(n14115), .B1(n14099), .B2(n14844), .ZN(
        P3_U3472) );
  OAI22_X1 U15908 ( .A1(n14101), .A2(n14828), .B1(n14100), .B2(n14827), .ZN(
        n14102) );
  NOR2_X1 U15909 ( .A1(n14103), .A2(n14102), .ZN(n14117) );
  AOI22_X1 U15910 ( .A1(n14846), .A2(n14117), .B1(n14104), .B2(n14844), .ZN(
        P3_U3471) );
  AOI22_X1 U15911 ( .A1(n14107), .A2(n14106), .B1(n14812), .B2(n14105), .ZN(
        n14108) );
  AND2_X1 U15912 ( .A1(n14109), .A2(n14108), .ZN(n14119) );
  INV_X1 U15913 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14110) );
  AOI22_X1 U15914 ( .A1(n14846), .A2(n14119), .B1(n14110), .B2(n14844), .ZN(
        P3_U3470) );
  INV_X1 U15915 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14111) );
  AOI22_X1 U15916 ( .A1(n14833), .A2(n14112), .B1(n14111), .B2(n14832), .ZN(
        P3_U3458) );
  INV_X1 U15917 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14968) );
  AOI22_X1 U15918 ( .A1(n14833), .A2(n14113), .B1(n14968), .B2(n14832), .ZN(
        P3_U3457) );
  INV_X1 U15919 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14114) );
  AOI22_X1 U15920 ( .A1(n14833), .A2(n14115), .B1(n14114), .B2(n14832), .ZN(
        P3_U3429) );
  INV_X1 U15921 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14116) );
  AOI22_X1 U15922 ( .A1(n14833), .A2(n14117), .B1(n14116), .B2(n14832), .ZN(
        P3_U3426) );
  INV_X1 U15923 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14118) );
  AOI22_X1 U15924 ( .A1(n14833), .A2(n14119), .B1(n14118), .B2(n14832), .ZN(
        P3_U3423) );
  AND2_X1 U15925 ( .A1(n14121), .A2(n14120), .ZN(n14124) );
  OAI21_X1 U15926 ( .B1(n14124), .B2(n14123), .A(n14122), .ZN(n14125) );
  AOI222_X1 U15927 ( .A1(n14142), .A2(n14210), .B1(n14209), .B2(n14141), .C1(
        n14125), .C2(n14139), .ZN(n14127) );
  OAI211_X1 U15928 ( .C1(n14146), .C2(n14128), .A(n14127), .B(n14126), .ZN(
        P1_U3215) );
  NAND2_X1 U15929 ( .A1(n14292), .A2(n14129), .ZN(n14133) );
  NAND2_X1 U15930 ( .A1(n14131), .A2(n14130), .ZN(n14132) );
  NAND2_X1 U15931 ( .A1(n14133), .A2(n14132), .ZN(n14166) );
  AND2_X1 U15932 ( .A1(n14135), .A2(n14134), .ZN(n14138) );
  OAI21_X1 U15933 ( .B1(n14138), .B2(n14137), .A(n14136), .ZN(n14140) );
  AOI222_X1 U15934 ( .A1(n14142), .A2(n14172), .B1(n14166), .B2(n14141), .C1(
        n14140), .C2(n14139), .ZN(n14144) );
  OAI211_X1 U15935 ( .C1(n14146), .C2(n14145), .A(n14144), .B(n14143), .ZN(
        P1_U3236) );
  AOI21_X1 U15936 ( .B1(n14148), .B2(n14147), .A(n14357), .ZN(n14152) );
  INV_X1 U15937 ( .A(n14149), .ZN(n14150) );
  AOI21_X1 U15938 ( .B1(n14152), .B2(n14151), .A(n14150), .ZN(n14189) );
  AOI222_X1 U15939 ( .A1(n14154), .A2(n14306), .B1(P1_REG2_REG_17__SCAN_IN), 
        .B2(n14284), .C1(n14285), .C2(n14153), .ZN(n14163) );
  NAND2_X1 U15940 ( .A1(n14156), .A2(n14155), .ZN(n14157) );
  AND2_X1 U15941 ( .A1(n7361), .A2(n14157), .ZN(n14192) );
  OAI211_X1 U15942 ( .C1(n14159), .C2(n14190), .A(n14310), .B(n14158), .ZN(
        n14188) );
  NOR2_X1 U15943 ( .A1(n14188), .A2(n14160), .ZN(n14161) );
  AOI21_X1 U15944 ( .B1(n14192), .B2(n14315), .A(n14161), .ZN(n14162) );
  OAI211_X1 U15945 ( .C1(n14318), .C2(n14189), .A(n14163), .B(n14162), .ZN(
        P1_U3276) );
  INV_X1 U15946 ( .A(n14164), .ZN(n14165) );
  AOI21_X1 U15947 ( .B1(n14165), .B2(n14171), .A(n14357), .ZN(n14168) );
  AOI21_X1 U15948 ( .B1(n14168), .B2(n14167), .A(n14166), .ZN(n14224) );
  AOI222_X1 U15949 ( .A1(n14172), .A2(n14306), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n14284), .C1(n14285), .C2(n14169), .ZN(n14178) );
  XNOR2_X1 U15950 ( .A(n14170), .B(n14171), .ZN(n14227) );
  INV_X1 U15951 ( .A(n14172), .ZN(n14225) );
  INV_X1 U15952 ( .A(n14173), .ZN(n14175) );
  OAI211_X1 U15953 ( .C1(n14225), .C2(n14175), .A(n14310), .B(n14174), .ZN(
        n14223) );
  INV_X1 U15954 ( .A(n14223), .ZN(n14176) );
  AOI22_X1 U15955 ( .A1(n14227), .A2(n14315), .B1(n14314), .B2(n14176), .ZN(
        n14177) );
  OAI211_X1 U15956 ( .C1(n14318), .C2(n14224), .A(n14178), .B(n14177), .ZN(
        P1_U3282) );
  AND2_X1 U15957 ( .A1(n14179), .A2(n14375), .ZN(n14185) );
  INV_X1 U15958 ( .A(n14180), .ZN(n14181) );
  OAI22_X1 U15959 ( .A1(n14183), .A2(n14182), .B1(n14181), .B2(n14371), .ZN(
        n14184) );
  NOR3_X1 U15960 ( .A1(n14186), .A2(n14185), .A3(n14184), .ZN(n14230) );
  INV_X1 U15961 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14187) );
  AOI22_X1 U15962 ( .A1(n14391), .A2(n14230), .B1(n14187), .B2(n14388), .ZN(
        P1_U3546) );
  OAI211_X1 U15963 ( .C1(n14190), .C2(n14371), .A(n14189), .B(n14188), .ZN(
        n14191) );
  AOI21_X1 U15964 ( .B1(n14375), .B2(n14192), .A(n14191), .ZN(n14232) );
  AOI22_X1 U15965 ( .A1(n14391), .A2(n14232), .B1(n14193), .B2(n14388), .ZN(
        P1_U3545) );
  AND2_X1 U15966 ( .A1(n14194), .A2(n14375), .ZN(n14199) );
  INV_X1 U15967 ( .A(n14195), .ZN(n14197) );
  OAI21_X1 U15968 ( .B1(n14197), .B2(n14371), .A(n14196), .ZN(n14198) );
  NOR3_X1 U15969 ( .A1(n14200), .A2(n14199), .A3(n14198), .ZN(n14234) );
  AOI22_X1 U15970 ( .A1(n14391), .A2(n14234), .B1(n14201), .B2(n14388), .ZN(
        P1_U3544) );
  AND2_X1 U15971 ( .A1(n14202), .A2(n14375), .ZN(n14205) );
  OAI21_X1 U15972 ( .B1(n6891), .B2(n14371), .A(n14203), .ZN(n14204) );
  NOR3_X1 U15973 ( .A1(n14206), .A2(n14205), .A3(n14204), .ZN(n14236) );
  INV_X1 U15974 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14207) );
  AOI22_X1 U15975 ( .A1(n14391), .A2(n14236), .B1(n14207), .B2(n14388), .ZN(
        P1_U3543) );
  AOI211_X1 U15976 ( .C1(n14345), .C2(n14210), .A(n14209), .B(n14208), .ZN(
        n14213) );
  NAND3_X1 U15977 ( .A1(n11546), .A2(n14211), .A3(n14375), .ZN(n14212) );
  OAI211_X1 U15978 ( .C1(n14357), .C2(n14214), .A(n14213), .B(n14212), .ZN(
        n14215) );
  INV_X1 U15979 ( .A(n14215), .ZN(n14238) );
  AOI22_X1 U15980 ( .A1(n14391), .A2(n14238), .B1(n14216), .B2(n14388), .ZN(
        P1_U3542) );
  NOR2_X1 U15981 ( .A1(n14217), .A2(n14349), .ZN(n14221) );
  OAI21_X1 U15982 ( .B1(n14219), .B2(n14371), .A(n14218), .ZN(n14220) );
  NOR3_X1 U15983 ( .A1(n14222), .A2(n14221), .A3(n14220), .ZN(n14240) );
  AOI22_X1 U15984 ( .A1(n14391), .A2(n14240), .B1(n10382), .B2(n14388), .ZN(
        P1_U3541) );
  OAI211_X1 U15985 ( .C1(n14225), .C2(n14371), .A(n14224), .B(n14223), .ZN(
        n14226) );
  AOI21_X1 U15986 ( .B1(n14375), .B2(n14227), .A(n14226), .ZN(n14242) );
  AOI22_X1 U15987 ( .A1(n14391), .A2(n14242), .B1(n14228), .B2(n14388), .ZN(
        P1_U3539) );
  INV_X1 U15988 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n14229) );
  AOI22_X1 U15989 ( .A1(n14378), .A2(n14230), .B1(n14229), .B2(n14376), .ZN(
        P1_U3513) );
  INV_X1 U15990 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14231) );
  AOI22_X1 U15991 ( .A1(n14378), .A2(n14232), .B1(n14231), .B2(n14376), .ZN(
        P1_U3510) );
  INV_X1 U15992 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14233) );
  AOI22_X1 U15993 ( .A1(n14378), .A2(n14234), .B1(n14233), .B2(n14376), .ZN(
        P1_U3507) );
  INV_X1 U15994 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14235) );
  AOI22_X1 U15995 ( .A1(n14378), .A2(n14236), .B1(n14235), .B2(n14376), .ZN(
        P1_U3504) );
  INV_X1 U15996 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14237) );
  AOI22_X1 U15997 ( .A1(n14378), .A2(n14238), .B1(n14237), .B2(n14376), .ZN(
        P1_U3501) );
  INV_X1 U15998 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14239) );
  AOI22_X1 U15999 ( .A1(n14378), .A2(n14240), .B1(n14239), .B2(n14376), .ZN(
        P1_U3498) );
  INV_X1 U16000 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14241) );
  AOI22_X1 U16001 ( .A1(n14378), .A2(n14242), .B1(n14241), .B2(n14376), .ZN(
        P1_U3492) );
  AOI21_X1 U16002 ( .B1(n14245), .B2(n14244), .A(n14243), .ZN(n14246) );
  XOR2_X1 U16003 ( .A(n14246), .B(P2_ADDR_REG_11__SCAN_IN), .Z(SUB_1596_U69)
         );
  OAI21_X1 U16004 ( .B1(n14248), .B2(n6592), .A(n14247), .ZN(n14249) );
  XOR2_X1 U16005 ( .A(n14249), .B(n14498), .Z(SUB_1596_U68) );
  OAI21_X1 U16006 ( .B1(n14252), .B2(n14251), .A(n14250), .ZN(n14254) );
  XOR2_X1 U16007 ( .A(n14254), .B(n14253), .Z(SUB_1596_U67) );
  AOI21_X1 U16008 ( .B1(n14257), .B2(n14256), .A(n14255), .ZN(n14258) );
  XOR2_X1 U16009 ( .A(n14258), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  NOR2_X1 U16010 ( .A1(n14260), .A2(n14259), .ZN(n14261) );
  XOR2_X1 U16011 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14261), .Z(SUB_1596_U65)
         );
  NOR2_X1 U16012 ( .A1(n14263), .A2(n14262), .ZN(n14264) );
  XOR2_X1 U16013 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14264), .Z(SUB_1596_U64)
         );
  AOI21_X1 U16014 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n14266), .A(n14265), 
        .ZN(n14271) );
  AOI21_X1 U16015 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14268), .A(n14267), 
        .ZN(n14269) );
  OAI222_X1 U16016 ( .A1(n14274), .A2(n14273), .B1(n14272), .B2(n14271), .C1(
        n14270), .C2(n14269), .ZN(n14275) );
  INV_X1 U16017 ( .A(n14275), .ZN(n14277) );
  NAND2_X1 U16018 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14276)
         );
  OAI211_X1 U16019 ( .C1(n14279), .C2(n14278), .A(n14277), .B(n14276), .ZN(
        P1_U3258) );
  AOI21_X1 U16020 ( .B1(n14280), .B2(n14289), .A(n14357), .ZN(n14283) );
  AOI21_X1 U16021 ( .B1(n14283), .B2(n14282), .A(n14281), .ZN(n14370) );
  AOI222_X1 U16022 ( .A1(n14287), .A2(n14306), .B1(n14286), .B2(n14285), .C1(
        P1_REG2_REG_10__SCAN_IN), .C2(n14284), .ZN(n14296) );
  XNOR2_X1 U16023 ( .A(n14288), .B(n14289), .ZN(n14374) );
  XNOR2_X1 U16024 ( .A(n14372), .B(n14290), .ZN(n14293) );
  AOI22_X1 U16025 ( .A1(n14293), .A2(n14310), .B1(n14292), .B2(n14291), .ZN(
        n14369) );
  INV_X1 U16026 ( .A(n14369), .ZN(n14294) );
  AOI22_X1 U16027 ( .A1(n14374), .A2(n14315), .B1(n14314), .B2(n14294), .ZN(
        n14295) );
  OAI211_X1 U16028 ( .C1(n14318), .C2(n14370), .A(n14296), .B(n14295), .ZN(
        P1_U3283) );
  XNOR2_X1 U16029 ( .A(n14297), .B(n14298), .ZN(n14301) );
  INV_X1 U16030 ( .A(n14299), .ZN(n14300) );
  AOI21_X1 U16031 ( .B1(n14301), .B2(n14353), .A(n14300), .ZN(n14329) );
  OAI22_X1 U16032 ( .A1(n14303), .A2(n9606), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n14302), .ZN(n14304) );
  AOI21_X1 U16033 ( .B1(n14306), .B2(n14305), .A(n14304), .ZN(n14317) );
  XNOR2_X1 U16034 ( .A(n14307), .B(n14308), .ZN(n14332) );
  INV_X1 U16035 ( .A(n14309), .ZN(n14311) );
  OAI211_X1 U16036 ( .C1(n14328), .C2(n14312), .A(n14311), .B(n14310), .ZN(
        n14327) );
  INV_X1 U16037 ( .A(n14327), .ZN(n14313) );
  AOI22_X1 U16038 ( .A1(n14332), .A2(n14315), .B1(n14314), .B2(n14313), .ZN(
        n14316) );
  OAI211_X1 U16039 ( .C1(n14318), .C2(n14329), .A(n14317), .B(n14316), .ZN(
        P1_U3290) );
  AND2_X1 U16040 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14320), .ZN(P1_U3294) );
  AND2_X1 U16041 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14320), .ZN(P1_U3295) );
  AND2_X1 U16042 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14320), .ZN(P1_U3296) );
  AND2_X1 U16043 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14320), .ZN(P1_U3297) );
  AND2_X1 U16044 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14320), .ZN(P1_U3298) );
  AND2_X1 U16045 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14320), .ZN(P1_U3299) );
  AND2_X1 U16046 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14320), .ZN(P1_U3300) );
  AND2_X1 U16047 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14320), .ZN(P1_U3301) );
  AND2_X1 U16048 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14320), .ZN(P1_U3302) );
  AND2_X1 U16049 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14320), .ZN(P1_U3303) );
  AND2_X1 U16050 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14320), .ZN(P1_U3304) );
  AND2_X1 U16051 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14320), .ZN(P1_U3305) );
  AND2_X1 U16052 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14320), .ZN(P1_U3306) );
  INV_X1 U16053 ( .A(n14320), .ZN(n14319) );
  INV_X1 U16054 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n14950) );
  NOR2_X1 U16055 ( .A1(n14319), .A2(n14950), .ZN(P1_U3307) );
  AND2_X1 U16056 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14320), .ZN(P1_U3308) );
  AND2_X1 U16057 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14320), .ZN(P1_U3309) );
  AND2_X1 U16058 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14320), .ZN(P1_U3310) );
  AND2_X1 U16059 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14320), .ZN(P1_U3311) );
  INV_X1 U16060 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n14869) );
  NOR2_X1 U16061 ( .A1(n14319), .A2(n14869), .ZN(P1_U3312) );
  INV_X1 U16062 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n14866) );
  NOR2_X1 U16063 ( .A1(n14319), .A2(n14866), .ZN(P1_U3313) );
  AND2_X1 U16064 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14320), .ZN(P1_U3314) );
  AND2_X1 U16065 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14320), .ZN(P1_U3315) );
  AND2_X1 U16066 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14320), .ZN(P1_U3316) );
  AND2_X1 U16067 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14320), .ZN(P1_U3317) );
  AND2_X1 U16068 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14320), .ZN(P1_U3318) );
  AND2_X1 U16069 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14320), .ZN(P1_U3319) );
  AND2_X1 U16070 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14320), .ZN(P1_U3320) );
  AND2_X1 U16071 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14320), .ZN(P1_U3321) );
  AND2_X1 U16072 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14320), .ZN(P1_U3322) );
  AND2_X1 U16073 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14320), .ZN(P1_U3323) );
  OAI21_X1 U16074 ( .B1(n14322), .B2(n14371), .A(n14321), .ZN(n14324) );
  AOI211_X1 U16075 ( .C1(n14375), .C2(n14325), .A(n14324), .B(n14323), .ZN(
        n14380) );
  INV_X1 U16076 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14326) );
  AOI22_X1 U16077 ( .A1(n14378), .A2(n14380), .B1(n14326), .B2(n14376), .ZN(
        P1_U3462) );
  OAI21_X1 U16078 ( .B1(n14328), .B2(n14371), .A(n14327), .ZN(n14331) );
  INV_X1 U16079 ( .A(n14329), .ZN(n14330) );
  AOI211_X1 U16080 ( .C1(n14375), .C2(n14332), .A(n14331), .B(n14330), .ZN(
        n14381) );
  INV_X1 U16081 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14333) );
  AOI22_X1 U16082 ( .A1(n14378), .A2(n14381), .B1(n14333), .B2(n14376), .ZN(
        P1_U3468) );
  NAND2_X1 U16083 ( .A1(n14334), .A2(n14375), .ZN(n14339) );
  NAND2_X1 U16084 ( .A1(n14335), .A2(n14345), .ZN(n14336) );
  NAND4_X1 U16085 ( .A1(n14339), .A2(n14338), .A3(n14337), .A4(n14336), .ZN(
        n14340) );
  AOI21_X1 U16086 ( .B1(n14353), .B2(n14341), .A(n14340), .ZN(n14382) );
  INV_X1 U16087 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14342) );
  AOI22_X1 U16088 ( .A1(n14378), .A2(n14382), .B1(n14342), .B2(n14376), .ZN(
        P1_U3471) );
  INV_X1 U16089 ( .A(n14343), .ZN(n14344) );
  AOI21_X1 U16090 ( .B1(n14346), .B2(n14345), .A(n14344), .ZN(n14348) );
  OAI211_X1 U16091 ( .C1(n14350), .C2(n14349), .A(n14348), .B(n14347), .ZN(
        n14351) );
  AOI21_X1 U16092 ( .B1(n14353), .B2(n14352), .A(n14351), .ZN(n14384) );
  INV_X1 U16093 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14354) );
  AOI22_X1 U16094 ( .A1(n14378), .A2(n14384), .B1(n14354), .B2(n14376), .ZN(
        P1_U3477) );
  OAI211_X1 U16095 ( .C1(n6881), .C2(n14371), .A(n14356), .B(n14355), .ZN(
        n14360) );
  NOR2_X1 U16096 ( .A1(n14358), .A2(n14357), .ZN(n14359) );
  AOI211_X1 U16097 ( .C1(n14375), .C2(n14361), .A(n14360), .B(n14359), .ZN(
        n14386) );
  INV_X1 U16098 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14362) );
  AOI22_X1 U16099 ( .A1(n14378), .A2(n14386), .B1(n14362), .B2(n14376), .ZN(
        P1_U3480) );
  OAI21_X1 U16100 ( .B1(n14364), .B2(n14371), .A(n14363), .ZN(n14366) );
  AOI211_X1 U16101 ( .C1(n14375), .C2(n14367), .A(n14366), .B(n14365), .ZN(
        n14387) );
  INV_X1 U16102 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14368) );
  AOI22_X1 U16103 ( .A1(n14378), .A2(n14387), .B1(n14368), .B2(n14376), .ZN(
        P1_U3483) );
  OAI211_X1 U16104 ( .C1(n14372), .C2(n14371), .A(n14370), .B(n14369), .ZN(
        n14373) );
  AOI21_X1 U16105 ( .B1(n14375), .B2(n14374), .A(n14373), .ZN(n14390) );
  INV_X1 U16106 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14377) );
  AOI22_X1 U16107 ( .A1(n14378), .A2(n14390), .B1(n14377), .B2(n14376), .ZN(
        P1_U3489) );
  AOI22_X1 U16108 ( .A1(n14391), .A2(n14380), .B1(n14379), .B2(n14388), .ZN(
        P1_U3529) );
  AOI22_X1 U16109 ( .A1(n14391), .A2(n14381), .B1(n9595), .B2(n14388), .ZN(
        P1_U3531) );
  AOI22_X1 U16110 ( .A1(n14391), .A2(n14382), .B1(n14877), .B2(n14388), .ZN(
        P1_U3532) );
  AOI22_X1 U16111 ( .A1(n14391), .A2(n14384), .B1(n14383), .B2(n14388), .ZN(
        P1_U3534) );
  AOI22_X1 U16112 ( .A1(n14391), .A2(n14386), .B1(n14385), .B2(n14388), .ZN(
        P1_U3535) );
  AOI22_X1 U16113 ( .A1(n14391), .A2(n14387), .B1(n9593), .B2(n14388), .ZN(
        P1_U3536) );
  AOI22_X1 U16114 ( .A1(n14391), .A2(n14390), .B1(n14389), .B2(n14388), .ZN(
        P1_U3538) );
  NOR2_X1 U16115 ( .A1(n14540), .A2(P2_U3947), .ZN(P2_U3087) );
  NAND2_X1 U16116 ( .A1(n14392), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14467) );
  NAND2_X1 U16117 ( .A1(P2_U3088), .A2(n14393), .ZN(n14394) );
  OAI211_X1 U16118 ( .C1(n14395), .C2(P2_U3088), .A(n14467), .B(n14394), .ZN(
        n14407) );
  OAI21_X1 U16119 ( .B1(n14398), .B2(n14397), .A(n14396), .ZN(n14399) );
  NAND3_X1 U16120 ( .A1(n14542), .A2(n14400), .A3(n14399), .ZN(n14406) );
  AOI21_X1 U16121 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(P2_REG2_REG_0__SCAN_IN), 
        .A(n14401), .ZN(n14402) );
  OR3_X1 U16122 ( .A1(n14536), .A2(n14403), .A3(n14402), .ZN(n14405) );
  NAND2_X1 U16123 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14540), .ZN(n14404) );
  NAND4_X1 U16124 ( .A1(n14407), .A2(n14406), .A3(n14405), .A4(n14404), .ZN(
        P2_U3215) );
  NAND2_X1 U16125 ( .A1(P2_U3088), .A2(n14408), .ZN(n14409) );
  OAI211_X1 U16126 ( .C1(n14411), .C2(P2_U3088), .A(n14467), .B(n14409), .ZN(
        n14422) );
  XOR2_X1 U16127 ( .A(n14413), .B(n14412), .Z(n14414) );
  NAND2_X1 U16128 ( .A1(n14542), .A2(n14414), .ZN(n14421) );
  AOI211_X1 U16129 ( .C1(n14417), .C2(n14416), .A(n14415), .B(n14536), .ZN(
        n14418) );
  INV_X1 U16130 ( .A(n14418), .ZN(n14420) );
  NAND2_X1 U16131 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(n14540), .ZN(n14419) );
  NAND4_X1 U16132 ( .A1(n14422), .A2(n14421), .A3(n14420), .A4(n14419), .ZN(
        P2_U3216) );
  INV_X1 U16133 ( .A(n14423), .ZN(n14424) );
  OAI21_X1 U16134 ( .B1(n14547), .B2(n14425), .A(n14424), .ZN(n14426) );
  AOI21_X1 U16135 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n14540), .A(n14426), .ZN(
        n14436) );
  AOI211_X1 U16136 ( .C1(n14429), .C2(n14428), .A(n14427), .B(n14536), .ZN(
        n14430) );
  INV_X1 U16137 ( .A(n14430), .ZN(n14435) );
  OAI211_X1 U16138 ( .C1(n14433), .C2(n14432), .A(n14542), .B(n14431), .ZN(
        n14434) );
  NAND3_X1 U16139 ( .A1(n14436), .A2(n14435), .A3(n14434), .ZN(P2_U3217) );
  INV_X1 U16140 ( .A(n14437), .ZN(n14439) );
  NAND2_X1 U16141 ( .A1(n14540), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n14438) );
  OAI211_X1 U16142 ( .C1(n14547), .C2(n14440), .A(n14439), .B(n14438), .ZN(
        n14441) );
  INV_X1 U16143 ( .A(n14441), .ZN(n14450) );
  AOI211_X1 U16144 ( .C1(n6601), .C2(n14443), .A(n14536), .B(n14442), .ZN(
        n14444) );
  INV_X1 U16145 ( .A(n14444), .ZN(n14449) );
  OAI211_X1 U16146 ( .C1(n14447), .C2(n14446), .A(n14542), .B(n14445), .ZN(
        n14448) );
  NAND3_X1 U16147 ( .A1(n14450), .A2(n14449), .A3(n14448), .ZN(P2_U3221) );
  NAND2_X1 U16148 ( .A1(n14451), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14452) );
  OAI211_X1 U16149 ( .C1(P2_STATE_REG_SCAN_IN), .C2(P2_REG3_REG_8__SCAN_IN), 
        .A(n14467), .B(n14452), .ZN(n14464) );
  INV_X1 U16150 ( .A(n14453), .ZN(n14454) );
  OAI211_X1 U16151 ( .C1(n14456), .C2(n14455), .A(n14542), .B(n14454), .ZN(
        n14463) );
  AOI211_X1 U16152 ( .C1(n14459), .C2(n14458), .A(n14536), .B(n14457), .ZN(
        n14460) );
  INV_X1 U16153 ( .A(n14460), .ZN(n14462) );
  NAND2_X1 U16154 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n14540), .ZN(n14461) );
  NAND4_X1 U16155 ( .A1(n14464), .A2(n14463), .A3(n14462), .A4(n14461), .ZN(
        P2_U3222) );
  NAND2_X1 U16156 ( .A1(n14465), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14466) );
  OAI211_X1 U16157 ( .C1(P2_STATE_REG_SCAN_IN), .C2(P2_REG3_REG_10__SCAN_IN), 
        .A(n14467), .B(n14466), .ZN(n14478) );
  OAI211_X1 U16158 ( .C1(n14470), .C2(n14469), .A(n14468), .B(n14542), .ZN(
        n14477) );
  NAND2_X1 U16159 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n14540), .ZN(n14476) );
  AOI211_X1 U16160 ( .C1(n14473), .C2(n14472), .A(n14536), .B(n14471), .ZN(
        n14474) );
  INV_X1 U16161 ( .A(n14474), .ZN(n14475) );
  NAND4_X1 U16162 ( .A1(n14478), .A2(n14477), .A3(n14476), .A4(n14475), .ZN(
        P2_U3224) );
  INV_X1 U16163 ( .A(n14479), .ZN(n14485) );
  OAI21_X1 U16164 ( .B1(n14482), .B2(n14481), .A(n14480), .ZN(n14484) );
  AOI21_X1 U16165 ( .B1(n14485), .B2(n14484), .A(n14483), .ZN(n14493) );
  INV_X1 U16166 ( .A(n14486), .ZN(n14491) );
  NAND3_X1 U16167 ( .A1(n14489), .A2(n14488), .A3(n14487), .ZN(n14490) );
  AOI21_X1 U16168 ( .B1(n14491), .B2(n14490), .A(n14536), .ZN(n14492) );
  AOI211_X1 U16169 ( .C1(n14521), .C2(n14494), .A(n14493), .B(n14492), .ZN(
        n14496) );
  NAND2_X1 U16170 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14495)
         );
  OAI211_X1 U16171 ( .C1(n14498), .C2(n14497), .A(n14496), .B(n14495), .ZN(
        P2_U3226) );
  NAND2_X1 U16172 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n14503)
         );
  OAI211_X1 U16173 ( .C1(n14501), .C2(n14500), .A(n14499), .B(n14526), .ZN(
        n14502) );
  NAND2_X1 U16174 ( .A1(n14503), .A2(n14502), .ZN(n14504) );
  AOI21_X1 U16175 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(n14540), .A(n14504), 
        .ZN(n14509) );
  OAI211_X1 U16176 ( .C1(n14507), .C2(n14506), .A(n14505), .B(n14542), .ZN(
        n14508) );
  OAI211_X1 U16177 ( .C1(n14547), .C2(n14510), .A(n14509), .B(n14508), .ZN(
        P2_U3227) );
  AOI22_X1 U16178 ( .A1(n14540), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14519) );
  NAND2_X1 U16179 ( .A1(n14521), .A2(n14511), .ZN(n14518) );
  OAI211_X1 U16180 ( .C1(n14513), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14526), 
        .B(n14512), .ZN(n14517) );
  OAI211_X1 U16181 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n14515), .A(n14542), 
        .B(n14514), .ZN(n14516) );
  NAND4_X1 U16182 ( .A1(n14519), .A2(n14518), .A3(n14517), .A4(n14516), .ZN(
        P2_U3229) );
  AOI22_X1 U16183 ( .A1(n14540), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3088), .ZN(n14532) );
  NAND2_X1 U16184 ( .A1(n14521), .A2(n14520), .ZN(n14531) );
  OAI211_X1 U16185 ( .C1(n14524), .C2(n14523), .A(n14542), .B(n14522), .ZN(
        n14530) );
  OAI211_X1 U16186 ( .C1(n14528), .C2(n14527), .A(n14526), .B(n14525), .ZN(
        n14529) );
  NAND4_X1 U16187 ( .A1(n14532), .A2(n14531), .A3(n14530), .A4(n14529), .ZN(
        P2_U3231) );
  NOR2_X1 U16188 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14533), .ZN(n14539) );
  AOI21_X1 U16189 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n14535), .A(n14534), 
        .ZN(n14537) );
  NOR2_X1 U16190 ( .A1(n14537), .A2(n14536), .ZN(n14538) );
  AOI211_X1 U16191 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n14540), .A(n14539), 
        .B(n14538), .ZN(n14545) );
  OAI211_X1 U16192 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n14543), .A(n14542), 
        .B(n14541), .ZN(n14544) );
  OAI211_X1 U16193 ( .C1(n14547), .C2(n14546), .A(n14545), .B(n14544), .ZN(
        P2_U3232) );
  AND2_X1 U16194 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14550), .ZN(P2_U3266) );
  AND2_X1 U16195 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14550), .ZN(P2_U3267) );
  AND2_X1 U16196 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14550), .ZN(P2_U3268) );
  AND2_X1 U16197 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14550), .ZN(P2_U3269) );
  AND2_X1 U16198 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14550), .ZN(P2_U3270) );
  AND2_X1 U16199 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14550), .ZN(P2_U3271) );
  AND2_X1 U16200 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14550), .ZN(P2_U3272) );
  AND2_X1 U16201 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14550), .ZN(P2_U3273) );
  AND2_X1 U16202 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14550), .ZN(P2_U3274) );
  AND2_X1 U16203 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14550), .ZN(P2_U3275) );
  AND2_X1 U16204 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14550), .ZN(P2_U3276) );
  AND2_X1 U16205 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14550), .ZN(P2_U3277) );
  AND2_X1 U16206 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14550), .ZN(P2_U3278) );
  AND2_X1 U16207 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14550), .ZN(P2_U3279) );
  AND2_X1 U16208 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14550), .ZN(P2_U3280) );
  AND2_X1 U16209 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14550), .ZN(P2_U3281) );
  AND2_X1 U16210 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14550), .ZN(P2_U3282) );
  AND2_X1 U16211 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14550), .ZN(P2_U3283) );
  AND2_X1 U16212 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14550), .ZN(P2_U3284) );
  AND2_X1 U16213 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14550), .ZN(P2_U3285) );
  INV_X1 U16214 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n14855) );
  NOR2_X1 U16215 ( .A1(n14549), .A2(n14855), .ZN(P2_U3286) );
  AND2_X1 U16216 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14550), .ZN(P2_U3287) );
  AND2_X1 U16217 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14550), .ZN(P2_U3288) );
  AND2_X1 U16218 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14550), .ZN(P2_U3289) );
  AND2_X1 U16219 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14550), .ZN(P2_U3290) );
  AND2_X1 U16220 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14550), .ZN(P2_U3291) );
  AND2_X1 U16221 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14550), .ZN(P2_U3292) );
  AND2_X1 U16222 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14550), .ZN(P2_U3293) );
  AND2_X1 U16223 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14550), .ZN(P2_U3294) );
  AND2_X1 U16224 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14550), .ZN(P2_U3295) );
  OAI21_X1 U16225 ( .B1(n14556), .B2(n14552), .A(n14551), .ZN(P2_U3416) );
  AOI22_X1 U16226 ( .A1(n14556), .A2(n14555), .B1(n14554), .B2(n14553), .ZN(
        P2_U3417) );
  INV_X1 U16227 ( .A(n14557), .ZN(n14563) );
  INV_X1 U16228 ( .A(n14558), .ZN(n14559) );
  OAI211_X1 U16229 ( .C1(n14561), .C2(n14592), .A(n14560), .B(n14559), .ZN(
        n14562) );
  AOI21_X1 U16230 ( .B1(n14589), .B2(n14563), .A(n14562), .ZN(n14599) );
  INV_X1 U16231 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14564) );
  AOI22_X1 U16232 ( .A1(n10992), .A2(n14599), .B1(n14564), .B2(n14597), .ZN(
        P2_U3439) );
  AOI21_X1 U16233 ( .B1(n14567), .B2(n14566), .A(n14565), .ZN(n14569) );
  OAI211_X1 U16234 ( .C1(n14571), .C2(n14570), .A(n14569), .B(n14568), .ZN(
        n14572) );
  INV_X1 U16235 ( .A(n14572), .ZN(n14600) );
  INV_X1 U16236 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14573) );
  AOI22_X1 U16237 ( .A1(n10992), .A2(n14600), .B1(n14573), .B2(n14597), .ZN(
        P2_U3442) );
  INV_X1 U16238 ( .A(n14574), .ZN(n14579) );
  OAI21_X1 U16239 ( .B1(n14576), .B2(n14592), .A(n14575), .ZN(n14578) );
  AOI211_X1 U16240 ( .C1(n14580), .C2(n14579), .A(n14578), .B(n14577), .ZN(
        n14601) );
  INV_X1 U16241 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n14581) );
  AOI22_X1 U16242 ( .A1(n10992), .A2(n14601), .B1(n14581), .B2(n14597), .ZN(
        P2_U3448) );
  OAI21_X1 U16243 ( .B1(n14583), .B2(n14592), .A(n14582), .ZN(n14586) );
  INV_X1 U16244 ( .A(n14584), .ZN(n14585) );
  AOI211_X1 U16245 ( .C1(n14587), .C2(n14589), .A(n14586), .B(n14585), .ZN(
        n14602) );
  INV_X1 U16246 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n14588) );
  AOI22_X1 U16247 ( .A1(n10992), .A2(n14602), .B1(n14588), .B2(n14597), .ZN(
        P2_U3451) );
  AND2_X1 U16248 ( .A1(n14590), .A2(n14589), .ZN(n14595) );
  OAI21_X1 U16249 ( .B1(n14593), .B2(n14592), .A(n14591), .ZN(n14594) );
  NOR3_X1 U16250 ( .A1(n14596), .A2(n14595), .A3(n14594), .ZN(n14604) );
  INV_X1 U16251 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14598) );
  AOI22_X1 U16252 ( .A1(n10992), .A2(n14604), .B1(n14598), .B2(n14597), .ZN(
        P2_U3463) );
  AOI22_X1 U16253 ( .A1(n10988), .A2(n14599), .B1(n9645), .B2(n14603), .ZN(
        P2_U3502) );
  AOI22_X1 U16254 ( .A1(n10988), .A2(n14600), .B1(n9658), .B2(n14603), .ZN(
        P2_U3503) );
  AOI22_X1 U16255 ( .A1(n10988), .A2(n14601), .B1(n9675), .B2(n14603), .ZN(
        P2_U3505) );
  AOI22_X1 U16256 ( .A1(n10988), .A2(n14602), .B1(n9950), .B2(n14603), .ZN(
        P2_U3506) );
  AOI22_X1 U16257 ( .A1(n10988), .A2(n14604), .B1(n10431), .B2(n14603), .ZN(
        P2_U3510) );
  NOR2_X1 U16258 ( .A1(P3_U3897), .A2(n14743), .ZN(P3_U3150) );
  MUX2_X1 U16259 ( .A(n14605), .B(n10309), .S(n12073), .Z(n14606) );
  NAND3_X1 U16260 ( .A1(n14607), .A2(n14750), .A3(n14709), .ZN(n14608) );
  OAI21_X1 U16261 ( .B1(n14610), .B2(n14609), .A(n14608), .ZN(n14612) );
  OAI211_X1 U16262 ( .C1(n14613), .C2(n14727), .A(n14612), .B(n14611), .ZN(
        P3_U3182) );
  AOI21_X1 U16263 ( .B1(n14615), .B2(n10595), .A(n14614), .ZN(n14620) );
  OAI21_X1 U16264 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(n14617), .A(n14616), .ZN(
        n14618) );
  NAND2_X1 U16265 ( .A1(n14746), .A2(n14618), .ZN(n14619) );
  OAI21_X1 U16266 ( .B1(n14620), .B2(n14750), .A(n14619), .ZN(n14626) );
  OR3_X1 U16267 ( .A1(n14623), .A2(n14622), .A3(n14621), .ZN(n14624) );
  AOI21_X1 U16268 ( .B1(n14642), .B2(n14624), .A(n14709), .ZN(n14625) );
  AOI211_X1 U16269 ( .C1(n14718), .C2(n14627), .A(n14626), .B(n14625), .ZN(
        n14629) );
  NAND2_X1 U16270 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_U3151), .ZN(n14628) );
  OAI211_X1 U16271 ( .C1(n9384), .C2(n14727), .A(n14629), .B(n14628), .ZN(
        P3_U3185) );
  INV_X1 U16272 ( .A(n14630), .ZN(n14631) );
  AOI21_X1 U16273 ( .B1(n14633), .B2(n14632), .A(n14631), .ZN(n14639) );
  OAI21_X1 U16274 ( .B1(n14636), .B2(n14635), .A(n14634), .ZN(n14637) );
  NAND2_X1 U16275 ( .A1(n14746), .A2(n14637), .ZN(n14638) );
  OAI21_X1 U16276 ( .B1(n14639), .B2(n14750), .A(n14638), .ZN(n14646) );
  INV_X1 U16277 ( .A(n14655), .ZN(n14644) );
  NAND3_X1 U16278 ( .A1(n14642), .A2(n14641), .A3(n14640), .ZN(n14643) );
  AOI21_X1 U16279 ( .B1(n14644), .B2(n14643), .A(n14709), .ZN(n14645) );
  AOI211_X1 U16280 ( .C1(n14718), .C2(n14647), .A(n14646), .B(n14645), .ZN(
        n14649) );
  NAND2_X1 U16281 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n14648) );
  OAI211_X1 U16282 ( .C1(n14650), .C2(n14727), .A(n14649), .B(n14648), .ZN(
        P3_U3186) );
  AOI21_X1 U16283 ( .B1(n14652), .B2(n10720), .A(n14651), .ZN(n14664) );
  INV_X1 U16284 ( .A(n14679), .ZN(n14657) );
  NOR3_X1 U16285 ( .A1(n14655), .A2(n14654), .A3(n14653), .ZN(n14656) );
  OAI21_X1 U16286 ( .B1(n14657), .B2(n14656), .A(n14735), .ZN(n14663) );
  OAI21_X1 U16287 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n14659), .A(n14658), .ZN(
        n14660) );
  AOI22_X1 U16288 ( .A1(n14718), .A2(n14661), .B1(n14746), .B2(n14660), .ZN(
        n14662) );
  OAI211_X1 U16289 ( .C1(n14664), .C2(n14750), .A(n14663), .B(n14662), .ZN(
        n14665) );
  INV_X1 U16290 ( .A(n14665), .ZN(n14667) );
  NAND2_X1 U16291 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(P3_U3151), .ZN(n14666) );
  OAI211_X1 U16292 ( .C1(n14668), .C2(n14727), .A(n14667), .B(n14666), .ZN(
        P3_U3187) );
  AOI21_X1 U16293 ( .B1(n14670), .B2(n14669), .A(n6597), .ZN(n14676) );
  OAI21_X1 U16294 ( .B1(n14673), .B2(n14672), .A(n14671), .ZN(n14674) );
  NAND2_X1 U16295 ( .A1(n14746), .A2(n14674), .ZN(n14675) );
  OAI21_X1 U16296 ( .B1(n14676), .B2(n14750), .A(n14675), .ZN(n14683) );
  INV_X1 U16297 ( .A(n14693), .ZN(n14681) );
  NAND3_X1 U16298 ( .A1(n14679), .A2(n14678), .A3(n14677), .ZN(n14680) );
  AOI21_X1 U16299 ( .B1(n14681), .B2(n14680), .A(n14709), .ZN(n14682) );
  AOI211_X1 U16300 ( .C1(n14718), .C2(n14684), .A(n14683), .B(n14682), .ZN(
        n14686) );
  NAND2_X1 U16301 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n14685) );
  OAI211_X1 U16302 ( .C1(n14687), .C2(n14727), .A(n14686), .B(n14685), .ZN(
        P3_U3188) );
  AOI21_X1 U16303 ( .B1(n10612), .B2(n14689), .A(n14688), .ZN(n14705) );
  INV_X1 U16304 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n14690) );
  NOR2_X1 U16305 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14690), .ZN(n14699) );
  INV_X1 U16306 ( .A(n14708), .ZN(n14695) );
  NOR3_X1 U16307 ( .A1(n14693), .A2(n14692), .A3(n14691), .ZN(n14694) );
  OAI21_X1 U16308 ( .B1(n14695), .B2(n14694), .A(n14735), .ZN(n14696) );
  OAI21_X1 U16309 ( .B1(n14740), .B2(n14697), .A(n14696), .ZN(n14698) );
  AOI211_X1 U16310 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n14743), .A(n14699), .B(
        n14698), .ZN(n14704) );
  OAI21_X1 U16311 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n14701), .A(n14700), .ZN(
        n14702) );
  NAND2_X1 U16312 ( .A1(n14702), .A2(n14746), .ZN(n14703) );
  OAI211_X1 U16313 ( .C1(n14705), .C2(n14750), .A(n14704), .B(n14703), .ZN(
        P3_U3189) );
  INV_X1 U16314 ( .A(n14734), .ZN(n14711) );
  NAND3_X1 U16315 ( .A1(n14708), .A2(n14707), .A3(n14706), .ZN(n14710) );
  AOI21_X1 U16316 ( .B1(n14711), .B2(n14710), .A(n14709), .ZN(n14724) );
  AOI21_X1 U16317 ( .B1(n14714), .B2(n14713), .A(n14712), .ZN(n14722) );
  OAI21_X1 U16318 ( .B1(n14717), .B2(n14716), .A(n14715), .ZN(n14720) );
  AOI22_X1 U16319 ( .A1(n14720), .A2(n14746), .B1(n14719), .B2(n14718), .ZN(
        n14721) );
  OAI21_X1 U16320 ( .B1(n14722), .B2(n14750), .A(n14721), .ZN(n14723) );
  NOR2_X1 U16321 ( .A1(n14724), .A2(n14723), .ZN(n14726) );
  OAI211_X1 U16322 ( .C1(n14728), .C2(n14727), .A(n14726), .B(n14725), .ZN(
        P3_U3190) );
  AOI21_X1 U16323 ( .B1(n10624), .B2(n14730), .A(n14729), .ZN(n14751) );
  INV_X1 U16324 ( .A(n14731), .ZN(n14737) );
  NOR3_X1 U16325 ( .A1(n14734), .A2(n14733), .A3(n14732), .ZN(n14736) );
  OAI21_X1 U16326 ( .B1(n14737), .B2(n14736), .A(n14735), .ZN(n14738) );
  OAI21_X1 U16327 ( .B1(n14740), .B2(n14739), .A(n14738), .ZN(n14741) );
  AOI211_X1 U16328 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n14743), .A(n14742), .B(
        n14741), .ZN(n14749) );
  OAI21_X1 U16329 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n14745), .A(n14744), .ZN(
        n14747) );
  NAND2_X1 U16330 ( .A1(n14747), .A2(n14746), .ZN(n14748) );
  OAI211_X1 U16331 ( .C1(n14751), .C2(n14750), .A(n14749), .B(n14748), .ZN(
        P3_U3191) );
  OAI21_X1 U16332 ( .B1(n14753), .B2(n14758), .A(n14752), .ZN(n14779) );
  NOR2_X1 U16333 ( .A1(n14754), .A2(n14827), .ZN(n14778) );
  INV_X1 U16334 ( .A(n14778), .ZN(n14757) );
  OAI22_X1 U16335 ( .A1(n14757), .A2(n14756), .B1(n10077), .B2(n14755), .ZN(
        n14768) );
  XNOR2_X1 U16336 ( .A(n14759), .B(n14758), .ZN(n14766) );
  OAI22_X1 U16337 ( .A1(n14763), .A2(n14762), .B1(n14761), .B2(n14760), .ZN(
        n14764) );
  AOI21_X1 U16338 ( .B1(n14779), .B2(n14805), .A(n14764), .ZN(n14765) );
  OAI21_X1 U16339 ( .B1(n14767), .B2(n14766), .A(n14765), .ZN(n14777) );
  AOI211_X1 U16340 ( .C1(n14769), .C2(n14779), .A(n14768), .B(n14777), .ZN(
        n14771) );
  AOI22_X1 U16341 ( .A1(n14772), .A2(n10333), .B1(n14771), .B2(n14770), .ZN(
        P3_U3231) );
  AOI211_X1 U16342 ( .C1(n14780), .C2(n14775), .A(n14774), .B(n14773), .ZN(
        n14834) );
  AOI22_X1 U16343 ( .A1(n14833), .A2(n14834), .B1(n14776), .B2(n14832), .ZN(
        P3_U3393) );
  AOI211_X1 U16344 ( .C1(n14780), .C2(n14779), .A(n14778), .B(n14777), .ZN(
        n14836) );
  INV_X1 U16345 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n14781) );
  AOI22_X1 U16346 ( .A1(n14833), .A2(n14836), .B1(n14781), .B2(n14832), .ZN(
        P3_U3396) );
  OAI22_X1 U16347 ( .A1(n14783), .A2(n14821), .B1(n14827), .B2(n14782), .ZN(
        n14784) );
  NOR2_X1 U16348 ( .A1(n14785), .A2(n14784), .ZN(n14837) );
  AOI22_X1 U16349 ( .A1(n14833), .A2(n14837), .B1(n14786), .B2(n14832), .ZN(
        P3_U3399) );
  AOI21_X1 U16350 ( .B1(n14808), .B2(n14821), .A(n14787), .ZN(n14790) );
  INV_X1 U16351 ( .A(n14788), .ZN(n14789) );
  AOI211_X1 U16352 ( .C1(n14812), .C2(n14791), .A(n14790), .B(n14789), .ZN(
        n14838) );
  INV_X1 U16353 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n14792) );
  AOI22_X1 U16354 ( .A1(n14833), .A2(n14838), .B1(n14792), .B2(n14832), .ZN(
        P3_U3402) );
  INV_X1 U16355 ( .A(n14793), .ZN(n14797) );
  OAI22_X1 U16356 ( .A1(n14795), .A2(n14828), .B1(n14827), .B2(n14794), .ZN(
        n14796) );
  NOR2_X1 U16357 ( .A1(n14797), .A2(n14796), .ZN(n14839) );
  INV_X1 U16358 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n14798) );
  AOI22_X1 U16359 ( .A1(n14833), .A2(n14839), .B1(n14798), .B2(n14832), .ZN(
        P3_U3405) );
  INV_X1 U16360 ( .A(n14800), .ZN(n14804) );
  OAI22_X1 U16361 ( .A1(n14800), .A2(n14821), .B1(n14799), .B2(n14827), .ZN(
        n14803) );
  INV_X1 U16362 ( .A(n14801), .ZN(n14802) );
  AOI211_X1 U16363 ( .C1(n14805), .C2(n14804), .A(n14803), .B(n14802), .ZN(
        n14840) );
  INV_X1 U16364 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n14806) );
  AOI22_X1 U16365 ( .A1(n14833), .A2(n14840), .B1(n14806), .B2(n14832), .ZN(
        P3_U3408) );
  AOI21_X1 U16366 ( .B1(n14808), .B2(n14821), .A(n14807), .ZN(n14809) );
  AOI211_X1 U16367 ( .C1(n14812), .C2(n14811), .A(n14810), .B(n14809), .ZN(
        n14841) );
  INV_X1 U16368 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n14813) );
  AOI22_X1 U16369 ( .A1(n14833), .A2(n14841), .B1(n14813), .B2(n14832), .ZN(
        P3_U3411) );
  INV_X1 U16370 ( .A(n14814), .ZN(n14816) );
  OAI22_X1 U16371 ( .A1(n14816), .A2(n14821), .B1(n14815), .B2(n14827), .ZN(
        n14817) );
  NOR2_X1 U16372 ( .A1(n14818), .A2(n14817), .ZN(n14842) );
  INV_X1 U16373 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n14819) );
  AOI22_X1 U16374 ( .A1(n14833), .A2(n14842), .B1(n14819), .B2(n14832), .ZN(
        P3_U3414) );
  OAI22_X1 U16375 ( .A1(n14822), .A2(n14821), .B1(n14827), .B2(n14820), .ZN(
        n14823) );
  NOR2_X1 U16376 ( .A1(n14824), .A2(n14823), .ZN(n14843) );
  INV_X1 U16377 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n14825) );
  AOI22_X1 U16378 ( .A1(n14833), .A2(n14843), .B1(n14825), .B2(n14832), .ZN(
        P3_U3417) );
  OAI22_X1 U16379 ( .A1(n14829), .A2(n14828), .B1(n14827), .B2(n14826), .ZN(
        n14830) );
  NOR2_X1 U16380 ( .A1(n14831), .A2(n14830), .ZN(n14845) );
  INV_X1 U16381 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n14976) );
  AOI22_X1 U16382 ( .A1(n14833), .A2(n14845), .B1(n14976), .B2(n14832), .ZN(
        P3_U3420) );
  AOI22_X1 U16383 ( .A1(n14846), .A2(n14834), .B1(n8328), .B2(n14844), .ZN(
        P3_U3460) );
  AOI22_X1 U16384 ( .A1(n14846), .A2(n14836), .B1(n14835), .B2(n14844), .ZN(
        P3_U3461) );
  AOI22_X1 U16385 ( .A1(n14846), .A2(n14837), .B1(n10594), .B2(n14844), .ZN(
        P3_U3462) );
  AOI22_X1 U16386 ( .A1(n14846), .A2(n14838), .B1(n10640), .B2(n14844), .ZN(
        P3_U3463) );
  AOI22_X1 U16387 ( .A1(n14846), .A2(n14839), .B1(n10603), .B2(n14844), .ZN(
        P3_U3464) );
  AOI22_X1 U16388 ( .A1(n14846), .A2(n14840), .B1(n10638), .B2(n14844), .ZN(
        P3_U3465) );
  AOI22_X1 U16389 ( .A1(n14846), .A2(n14841), .B1(n10611), .B2(n14844), .ZN(
        P3_U3466) );
  AOI22_X1 U16390 ( .A1(n14846), .A2(n14842), .B1(n10617), .B2(n14844), .ZN(
        P3_U3467) );
  AOI22_X1 U16391 ( .A1(n14846), .A2(n14843), .B1(n10623), .B2(n14844), .ZN(
        P3_U3468) );
  AOI22_X1 U16392 ( .A1(n14846), .A2(n14845), .B1(n10657), .B2(n14844), .ZN(
        P3_U3469) );
  INV_X1 U16393 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n14848) );
  AOI22_X1 U16394 ( .A1(n14849), .A2(keyinput51), .B1(keyinput40), .B2(n14848), 
        .ZN(n14847) );
  OAI221_X1 U16395 ( .B1(n14849), .B2(keyinput51), .C1(n14848), .C2(keyinput40), .A(n14847), .ZN(n14861) );
  AOI22_X1 U16396 ( .A1(n14852), .A2(keyinput23), .B1(n14851), .B2(keyinput14), 
        .ZN(n14850) );
  OAI221_X1 U16397 ( .B1(n14852), .B2(keyinput23), .C1(n14851), .C2(keyinput14), .A(n14850), .ZN(n14860) );
  AOI22_X1 U16398 ( .A1(n14855), .A2(keyinput60), .B1(keyinput1), .B2(n14854), 
        .ZN(n14853) );
  OAI221_X1 U16399 ( .B1(n14855), .B2(keyinput60), .C1(n14854), .C2(keyinput1), 
        .A(n14853), .ZN(n14859) );
  XNOR2_X1 U16400 ( .A(P1_REG3_REG_25__SCAN_IN), .B(keyinput30), .ZN(n14857)
         );
  XNOR2_X1 U16401 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput9), .ZN(n14856) );
  NAND2_X1 U16402 ( .A1(n14857), .A2(n14856), .ZN(n14858) );
  NOR4_X1 U16403 ( .A1(n14861), .A2(n14860), .A3(n14859), .A4(n14858), .ZN(
        n14905) );
  INV_X1 U16404 ( .A(SI_28_), .ZN(n14863) );
  AOI22_X1 U16405 ( .A1(n14864), .A2(keyinput46), .B1(keyinput56), .B2(n14863), 
        .ZN(n14862) );
  OAI221_X1 U16406 ( .B1(n14864), .B2(keyinput46), .C1(n14863), .C2(keyinput56), .A(n14862), .ZN(n14875) );
  AOI22_X1 U16407 ( .A1(n14867), .A2(keyinput19), .B1(keyinput20), .B2(n14866), 
        .ZN(n14865) );
  OAI221_X1 U16408 ( .B1(n14867), .B2(keyinput19), .C1(n14866), .C2(keyinput20), .A(n14865), .ZN(n14874) );
  AOI22_X1 U16409 ( .A1(n14869), .A2(keyinput32), .B1(n14968), .B2(keyinput31), 
        .ZN(n14868) );
  OAI221_X1 U16410 ( .B1(n14869), .B2(keyinput32), .C1(n14968), .C2(keyinput31), .A(n14868), .ZN(n14873) );
  XNOR2_X1 U16411 ( .A(P3_REG1_REG_16__SCAN_IN), .B(keyinput47), .ZN(n14871)
         );
  XNOR2_X1 U16412 ( .A(P3_IR_REG_6__SCAN_IN), .B(keyinput57), .ZN(n14870) );
  NAND2_X1 U16413 ( .A1(n14871), .A2(n14870), .ZN(n14872) );
  NOR4_X1 U16414 ( .A1(n14875), .A2(n14874), .A3(n14873), .A4(n14872), .ZN(
        n14904) );
  AOI22_X1 U16415 ( .A1(n8628), .A2(keyinput53), .B1(keyinput55), .B2(n14877), 
        .ZN(n14876) );
  OAI221_X1 U16416 ( .B1(n8628), .B2(keyinput53), .C1(n14877), .C2(keyinput55), 
        .A(n14876), .ZN(n14889) );
  AOI22_X1 U16417 ( .A1(n14880), .A2(keyinput49), .B1(n14879), .B2(keyinput52), 
        .ZN(n14878) );
  OAI221_X1 U16418 ( .B1(n14880), .B2(keyinput49), .C1(n14879), .C2(keyinput52), .A(n14878), .ZN(n14888) );
  AOI22_X1 U16419 ( .A1(n14883), .A2(keyinput7), .B1(n14882), .B2(keyinput38), 
        .ZN(n14881) );
  OAI221_X1 U16420 ( .B1(n14883), .B2(keyinput7), .C1(n14882), .C2(keyinput38), 
        .A(n14881), .ZN(n14887) );
  XNOR2_X1 U16421 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput41), .ZN(n14885) );
  XNOR2_X1 U16422 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput35), .ZN(n14884) );
  NAND2_X1 U16423 ( .A1(n14885), .A2(n14884), .ZN(n14886) );
  NOR4_X1 U16424 ( .A1(n14889), .A2(n14888), .A3(n14887), .A4(n14886), .ZN(
        n14903) );
  AOI22_X1 U16425 ( .A1(n12458), .A2(keyinput6), .B1(keyinput28), .B2(n14891), 
        .ZN(n14890) );
  OAI221_X1 U16426 ( .B1(n12458), .B2(keyinput6), .C1(n14891), .C2(keyinput28), 
        .A(n14890), .ZN(n14901) );
  AOI22_X1 U16427 ( .A1(n9611), .A2(keyinput43), .B1(n14893), .B2(keyinput12), 
        .ZN(n14892) );
  OAI221_X1 U16428 ( .B1(n9611), .B2(keyinput43), .C1(n14893), .C2(keyinput12), 
        .A(n14892), .ZN(n14900) );
  XNOR2_X1 U16429 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput11), .ZN(n14896)
         );
  XNOR2_X1 U16430 ( .A(P1_REG2_REG_2__SCAN_IN), .B(keyinput42), .ZN(n14895) );
  XNOR2_X1 U16431 ( .A(P2_IR_REG_0__SCAN_IN), .B(keyinput25), .ZN(n14894) );
  NAND3_X1 U16432 ( .A1(n14896), .A2(n14895), .A3(n14894), .ZN(n14899) );
  XNOR2_X1 U16433 ( .A(n14897), .B(keyinput59), .ZN(n14898) );
  NOR4_X1 U16434 ( .A1(n14901), .A2(n14900), .A3(n14899), .A4(n14898), .ZN(
        n14902) );
  NAND4_X1 U16435 ( .A1(n14905), .A2(n14904), .A3(n14903), .A4(n14902), .ZN(
        n14964) );
  INV_X1 U16436 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14907) );
  AOI22_X1 U16437 ( .A1(n14907), .A2(keyinput45), .B1(n9720), .B2(keyinput39), 
        .ZN(n14906) );
  OAI221_X1 U16438 ( .B1(n14907), .B2(keyinput45), .C1(n9720), .C2(keyinput39), 
        .A(n14906), .ZN(n14918) );
  INV_X1 U16439 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14909) );
  AOI22_X1 U16440 ( .A1(n10623), .A2(keyinput21), .B1(keyinput33), .B2(n14909), 
        .ZN(n14908) );
  OAI221_X1 U16441 ( .B1(n10623), .B2(keyinput21), .C1(n14909), .C2(keyinput33), .A(n14908), .ZN(n14917) );
  AOI22_X1 U16442 ( .A1(n14912), .A2(keyinput48), .B1(keyinput58), .B2(n14911), 
        .ZN(n14910) );
  OAI221_X1 U16443 ( .B1(n14912), .B2(keyinput48), .C1(n14911), .C2(keyinput58), .A(n14910), .ZN(n14916) );
  XNOR2_X1 U16444 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput8), .ZN(n14914)
         );
  XNOR2_X1 U16445 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput18), .ZN(n14913) );
  NAND2_X1 U16446 ( .A1(n14914), .A2(n14913), .ZN(n14915) );
  NOR4_X1 U16447 ( .A1(n14918), .A2(n14917), .A3(n14916), .A4(n14915), .ZN(
        n14962) );
  AOI22_X1 U16448 ( .A1(n14920), .A2(keyinput37), .B1(keyinput5), .B2(n10929), 
        .ZN(n14919) );
  OAI221_X1 U16449 ( .B1(n14920), .B2(keyinput37), .C1(n10929), .C2(keyinput5), 
        .A(n14919), .ZN(n14933) );
  AOI22_X1 U16450 ( .A1(n14922), .A2(keyinput22), .B1(n14977), .B2(keyinput61), 
        .ZN(n14921) );
  OAI221_X1 U16451 ( .B1(n14922), .B2(keyinput22), .C1(n14977), .C2(keyinput61), .A(n14921), .ZN(n14927) );
  XNOR2_X1 U16452 ( .A(n14923), .B(keyinput3), .ZN(n14926) );
  XNOR2_X1 U16453 ( .A(n14924), .B(keyinput13), .ZN(n14925) );
  OR3_X1 U16454 ( .A1(n14927), .A2(n14926), .A3(n14925), .ZN(n14932) );
  AOI22_X1 U16455 ( .A1(n14930), .A2(keyinput24), .B1(n14929), .B2(keyinput62), 
        .ZN(n14928) );
  OAI221_X1 U16456 ( .B1(n14930), .B2(keyinput24), .C1(n14929), .C2(keyinput62), .A(n14928), .ZN(n14931) );
  NOR3_X1 U16457 ( .A1(n14933), .A2(n14932), .A3(n14931), .ZN(n14961) );
  AOI22_X1 U16458 ( .A1(n7745), .A2(keyinput63), .B1(keyinput34), .B2(n14935), 
        .ZN(n14934) );
  OAI221_X1 U16459 ( .B1(n7745), .B2(keyinput63), .C1(n14935), .C2(keyinput34), 
        .A(n14934), .ZN(n14945) );
  AOI22_X1 U16460 ( .A1(n14938), .A2(keyinput4), .B1(n14937), .B2(keyinput15), 
        .ZN(n14936) );
  OAI221_X1 U16461 ( .B1(n14938), .B2(keyinput4), .C1(n14937), .C2(keyinput15), 
        .A(n14936), .ZN(n14944) );
  XOR2_X1 U16462 ( .A(n14976), .B(keyinput36), .Z(n14942) );
  XNOR2_X1 U16463 ( .A(P1_REG1_REG_30__SCAN_IN), .B(keyinput54), .ZN(n14941)
         );
  XNOR2_X1 U16464 ( .A(P3_IR_REG_4__SCAN_IN), .B(keyinput26), .ZN(n14940) );
  XNOR2_X1 U16465 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput17), .ZN(n14939) );
  NAND4_X1 U16466 ( .A1(n14942), .A2(n14941), .A3(n14940), .A4(n14939), .ZN(
        n14943) );
  NOR3_X1 U16467 ( .A1(n14945), .A2(n14944), .A3(n14943), .ZN(n14960) );
  AOI22_X1 U16468 ( .A1(n14948), .A2(keyinput29), .B1(keyinput27), .B2(n14947), 
        .ZN(n14946) );
  OAI221_X1 U16469 ( .B1(n14948), .B2(keyinput29), .C1(n14947), .C2(keyinput27), .A(n14946), .ZN(n14958) );
  AOI22_X1 U16470 ( .A1(n14950), .A2(keyinput50), .B1(n8558), .B2(keyinput16), 
        .ZN(n14949) );
  OAI221_X1 U16471 ( .B1(n14950), .B2(keyinput50), .C1(n8558), .C2(keyinput16), 
        .A(n14949), .ZN(n14957) );
  XNOR2_X1 U16472 ( .A(P3_REG1_REG_15__SCAN_IN), .B(keyinput2), .ZN(n14953) );
  XNOR2_X1 U16473 ( .A(SI_1_), .B(keyinput10), .ZN(n14952) );
  XNOR2_X1 U16474 ( .A(P3_IR_REG_20__SCAN_IN), .B(keyinput44), .ZN(n14951) );
  NAND3_X1 U16475 ( .A1(n14953), .A2(n14952), .A3(n14951), .ZN(n14956) );
  XNOR2_X1 U16476 ( .A(n14954), .B(keyinput0), .ZN(n14955) );
  NOR4_X1 U16477 ( .A1(n14958), .A2(n14957), .A3(n14956), .A4(n14955), .ZN(
        n14959) );
  NAND4_X1 U16478 ( .A1(n14962), .A2(n14961), .A3(n14960), .A4(n14959), .ZN(
        n14963) );
  NOR2_X1 U16479 ( .A1(n14964), .A2(n14963), .ZN(n14967) );
  NAND2_X1 U16480 ( .A1(n14965), .A2(P3_D_REG_20__SCAN_IN), .ZN(n14966) );
  XNOR2_X1 U16481 ( .A(n14967), .B(n14966), .ZN(n14994) );
  NOR4_X1 U16482 ( .A1(SI_12_), .A2(P3_REG3_REG_21__SCAN_IN), .A3(
        P3_REG2_REG_20__SCAN_IN), .A4(n14968), .ZN(n14992) );
  NAND4_X1 U16483 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P3_REG0_REG_25__SCAN_IN), 
        .A3(P3_DATAO_REG_0__SCAN_IN), .A4(P3_DATAO_REG_4__SCAN_IN), .ZN(n14971) );
  NAND4_X1 U16484 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_DATAO_REG_6__SCAN_IN), 
        .A3(P2_REG0_REG_14__SCAN_IN), .A4(P3_DATAO_REG_15__SCAN_IN), .ZN(
        n14970) );
  NAND4_X1 U16485 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_REG2_REG_21__SCAN_IN), .A4(P1_REG2_REG_8__SCAN_IN), .ZN(n14969) );
  NOR3_X1 U16486 ( .A1(n14971), .A2(n14970), .A3(n14969), .ZN(n14991) );
  NAND4_X1 U16487 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(P1_REG0_REG_0__SCAN_IN), 
        .A3(P1_REG1_REG_4__SCAN_IN), .A4(P3_ADDR_REG_13__SCAN_IN), .ZN(n14975)
         );
  NAND4_X1 U16488 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(P2_REG0_REG_17__SCAN_IN), .A3(P3_REG0_REG_22__SCAN_IN), .A4(P2_DATAO_REG_30__SCAN_IN), .ZN(n14974) );
  NAND4_X1 U16489 ( .A1(P3_REG3_REG_20__SCAN_IN), .A2(P3_REG2_REG_26__SCAN_IN), 
        .A3(P3_REG1_REG_16__SCAN_IN), .A4(SI_30_), .ZN(n14973) );
  NAND4_X1 U16490 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_DATAO_REG_23__SCAN_IN), .A3(SI_1_), .A4(P1_ADDR_REG_16__SCAN_IN), .ZN(n14972) );
  NOR4_X1 U16491 ( .A1(n14975), .A2(n14974), .A3(n14973), .A4(n14972), .ZN(
        n14990) );
  NAND3_X1 U16492 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), 
        .A3(P3_IR_REG_4__SCAN_IN), .ZN(n14988) );
  NAND4_X1 U16493 ( .A1(n14977), .A2(n14976), .A3(n10929), .A4(n10623), .ZN(
        n14979) );
  NOR4_X1 U16494 ( .A1(n14979), .A2(n14978), .A3(P2_IR_REG_25__SCAN_IN), .A4(
        P1_REG3_REG_25__SCAN_IN), .ZN(n14981) );
  NAND4_X1 U16495 ( .A1(n14981), .A2(n14980), .A3(P3_ADDR_REG_2__SCAN_IN), 
        .A4(P1_ADDR_REG_2__SCAN_IN), .ZN(n14987) );
  NOR4_X1 U16496 ( .A1(P2_REG1_REG_25__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(P2_REG1_REG_31__SCAN_IN), .A4(P1_REG1_REG_30__SCAN_IN), .ZN(n14985) );
  NOR4_X1 U16497 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .A3(
        P1_REG2_REG_22__SCAN_IN), .A4(P1_REG2_REG_20__SCAN_IN), .ZN(n14984) );
  NOR4_X1 U16498 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(P2_REG2_REG_15__SCAN_IN), 
        .A3(P3_REG3_REG_13__SCAN_IN), .A4(P1_IR_REG_18__SCAN_IN), .ZN(n14983)
         );
  NOR4_X1 U16499 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(P2_DATAO_REG_14__SCAN_IN), .A3(SI_28_), .A4(P3_REG1_REG_15__SCAN_IN), .ZN(n14982) );
  NAND4_X1 U16500 ( .A1(n14985), .A2(n14984), .A3(n14983), .A4(n14982), .ZN(
        n14986) );
  NOR4_X1 U16501 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(n14988), .A3(n14987), 
        .A4(n14986), .ZN(n14989) );
  NAND4_X1 U16502 ( .A1(n14992), .A2(n14991), .A3(n14990), .A4(n14989), .ZN(
        n14993) );
  XNOR2_X1 U16503 ( .A(n14994), .B(n14993), .ZN(P3_U3245) );
  XOR2_X1 U16504 ( .A(n14996), .B(n14995), .Z(SUB_1596_U59) );
  XNOR2_X1 U16505 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n14997), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16506 ( .B1(n14999), .B2(n14998), .A(n15008), .ZN(SUB_1596_U53) );
  XOR2_X1 U16507 ( .A(n15000), .B(n15001), .Z(SUB_1596_U56) );
  OAI21_X1 U16508 ( .B1(n15004), .B2(n15003), .A(n15002), .ZN(n15006) );
  XOR2_X1 U16509 ( .A(n15006), .B(n15005), .Z(SUB_1596_U60) );
  XOR2_X1 U16510 ( .A(n15008), .B(n15007), .Z(SUB_1596_U5) );
  CLKBUF_X1 U7174 ( .A(n8888), .Z(n6464) );
  CLKBUF_X1 U7196 ( .A(n10256), .Z(n6458) );
  NAND2_X1 U7200 ( .A1(n11020), .A2(n8812), .ZN(n9747) );
  CLKBUF_X1 U7205 ( .A(n7508), .Z(n8077) );
  CLKBUF_X1 U7229 ( .A(n8889), .Z(n9266) );
  NAND2_X1 U7472 ( .A1(n6463), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8834) );
  CLKBUF_X1 U7490 ( .A(n8681), .Z(n12073) );
endmodule

